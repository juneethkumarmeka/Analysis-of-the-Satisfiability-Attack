module basic_1000_10000_1500_5_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_96,In_136);
nand U1 (N_1,In_356,In_348);
or U2 (N_2,In_627,In_359);
nand U3 (N_3,In_671,In_503);
nor U4 (N_4,In_786,In_816);
nor U5 (N_5,In_443,In_183);
or U6 (N_6,In_631,In_640);
or U7 (N_7,In_154,In_63);
nor U8 (N_8,In_692,In_150);
and U9 (N_9,In_804,In_181);
or U10 (N_10,In_938,In_794);
nand U11 (N_11,In_702,In_590);
nand U12 (N_12,In_821,In_15);
or U13 (N_13,In_713,In_43);
xnor U14 (N_14,In_543,In_198);
nor U15 (N_15,In_20,In_781);
or U16 (N_16,In_965,In_628);
nand U17 (N_17,In_836,In_859);
nor U18 (N_18,In_410,In_295);
or U19 (N_19,In_604,In_187);
and U20 (N_20,In_813,In_822);
nor U21 (N_21,In_315,In_351);
nand U22 (N_22,In_635,In_677);
nor U23 (N_23,In_742,In_500);
and U24 (N_24,In_478,In_833);
and U25 (N_25,In_828,In_439);
xor U26 (N_26,In_101,In_600);
or U27 (N_27,In_976,In_773);
and U28 (N_28,In_842,In_846);
xor U29 (N_29,In_762,In_966);
nor U30 (N_30,In_64,In_58);
nand U31 (N_31,In_511,In_621);
xnor U32 (N_32,In_643,In_213);
or U33 (N_33,In_681,In_520);
or U34 (N_34,In_361,In_927);
nand U35 (N_35,In_583,In_219);
nand U36 (N_36,In_358,In_548);
or U37 (N_37,In_386,In_745);
nand U38 (N_38,In_584,In_115);
nor U39 (N_39,In_116,In_112);
or U40 (N_40,In_273,In_454);
nor U41 (N_41,In_592,In_790);
or U42 (N_42,In_59,In_51);
nand U43 (N_43,In_678,In_298);
nand U44 (N_44,In_419,In_75);
or U45 (N_45,In_201,In_263);
xor U46 (N_46,In_484,In_951);
nand U47 (N_47,In_283,In_151);
nand U48 (N_48,In_143,In_759);
nand U49 (N_49,In_166,In_429);
xor U50 (N_50,In_542,In_318);
or U51 (N_51,In_84,In_504);
nor U52 (N_52,In_885,In_236);
or U53 (N_53,In_598,In_614);
and U54 (N_54,In_26,In_83);
and U55 (N_55,In_801,In_480);
nand U56 (N_56,In_698,In_563);
or U57 (N_57,In_290,In_721);
and U58 (N_58,In_778,In_936);
nor U59 (N_59,In_831,In_928);
or U60 (N_60,In_495,In_460);
nor U61 (N_61,In_407,In_765);
xnor U62 (N_62,In_264,In_321);
nor U63 (N_63,In_505,In_550);
nand U64 (N_64,In_714,In_62);
and U65 (N_65,In_941,In_696);
or U66 (N_66,In_887,In_568);
nand U67 (N_67,In_73,In_239);
nor U68 (N_68,In_602,In_779);
nor U69 (N_69,In_313,In_577);
nor U70 (N_70,In_400,In_871);
nor U71 (N_71,In_14,In_8);
and U72 (N_72,In_82,In_684);
nand U73 (N_73,In_658,In_570);
or U74 (N_74,In_618,In_567);
nand U75 (N_75,In_29,In_695);
nand U76 (N_76,In_109,In_922);
xor U77 (N_77,In_444,In_19);
or U78 (N_78,In_16,In_872);
and U79 (N_79,In_986,In_483);
and U80 (N_80,In_10,In_297);
or U81 (N_81,In_482,In_332);
xor U82 (N_82,In_134,In_86);
nand U83 (N_83,In_106,In_881);
nand U84 (N_84,In_336,In_795);
or U85 (N_85,In_225,In_608);
and U86 (N_86,In_565,In_724);
nand U87 (N_87,In_597,In_237);
nor U88 (N_88,In_895,In_921);
or U89 (N_89,In_329,In_796);
and U90 (N_90,In_57,In_975);
nand U91 (N_91,In_42,In_240);
nor U92 (N_92,In_850,In_47);
or U93 (N_93,In_133,In_432);
or U94 (N_94,In_957,In_2);
xor U95 (N_95,In_860,In_797);
and U96 (N_96,In_540,In_962);
nor U97 (N_97,In_380,In_78);
and U98 (N_98,In_653,In_485);
nand U99 (N_99,In_716,In_494);
and U100 (N_100,In_224,In_369);
nor U101 (N_101,In_427,In_272);
nor U102 (N_102,In_748,In_507);
nand U103 (N_103,In_424,In_413);
and U104 (N_104,In_431,In_411);
and U105 (N_105,In_149,In_210);
or U106 (N_106,In_280,In_931);
and U107 (N_107,In_254,In_23);
nor U108 (N_108,In_949,In_360);
or U109 (N_109,In_586,In_102);
xor U110 (N_110,In_525,In_223);
nand U111 (N_111,In_164,In_591);
nand U112 (N_112,In_277,In_925);
nor U113 (N_113,In_655,In_377);
nor U114 (N_114,In_71,In_649);
or U115 (N_115,In_516,In_746);
nor U116 (N_116,In_910,In_868);
or U117 (N_117,In_858,In_362);
xnor U118 (N_118,In_368,In_49);
nand U119 (N_119,In_776,In_126);
or U120 (N_120,In_719,In_30);
nor U121 (N_121,In_193,In_509);
nor U122 (N_122,In_670,In_123);
nand U123 (N_123,In_118,In_693);
and U124 (N_124,In_666,In_50);
and U125 (N_125,In_566,In_445);
nand U126 (N_126,In_481,In_961);
or U127 (N_127,In_825,In_387);
or U128 (N_128,In_757,In_248);
or U129 (N_129,In_120,In_398);
nor U130 (N_130,In_302,In_569);
nand U131 (N_131,In_863,In_37);
and U132 (N_132,In_36,In_955);
and U133 (N_133,In_967,In_611);
and U134 (N_134,In_146,In_447);
nand U135 (N_135,In_416,In_383);
or U136 (N_136,In_463,In_688);
nand U137 (N_137,In_807,In_984);
nand U138 (N_138,In_200,In_382);
and U139 (N_139,In_905,In_171);
nand U140 (N_140,In_709,In_390);
nor U141 (N_141,In_541,In_969);
xnor U142 (N_142,In_366,In_624);
and U143 (N_143,In_685,In_492);
and U144 (N_144,In_153,In_190);
nor U145 (N_145,In_355,In_903);
nor U146 (N_146,In_580,In_581);
nand U147 (N_147,In_531,In_189);
or U148 (N_148,In_403,In_593);
or U149 (N_149,In_772,In_227);
nor U150 (N_150,In_266,In_393);
nand U151 (N_151,In_241,In_970);
or U152 (N_152,In_184,In_983);
nor U153 (N_153,In_426,In_912);
nor U154 (N_154,In_891,In_341);
nand U155 (N_155,In_551,In_324);
or U156 (N_156,In_855,In_683);
nand U157 (N_157,In_79,In_766);
and U158 (N_158,In_256,In_125);
and U159 (N_159,In_18,In_522);
and U160 (N_160,In_616,In_527);
nand U161 (N_161,In_459,In_956);
xor U162 (N_162,In_60,In_838);
and U163 (N_163,In_320,In_869);
and U164 (N_164,In_353,In_67);
and U165 (N_165,In_165,In_27);
nor U166 (N_166,In_251,In_980);
and U167 (N_167,In_350,In_305);
or U168 (N_168,In_376,In_72);
nor U169 (N_169,In_619,In_453);
nand U170 (N_170,In_303,In_992);
nor U171 (N_171,In_758,In_650);
nor U172 (N_172,In_562,In_769);
nor U173 (N_173,In_942,In_7);
nor U174 (N_174,In_747,In_207);
or U175 (N_175,In_767,In_926);
xor U176 (N_176,In_206,In_395);
nor U177 (N_177,In_379,In_438);
and U178 (N_178,In_898,In_310);
nand U179 (N_179,In_645,In_648);
and U180 (N_180,In_734,In_117);
nor U181 (N_181,In_723,In_943);
nand U182 (N_182,In_873,In_622);
nand U183 (N_183,In_717,In_634);
nor U184 (N_184,In_587,In_609);
or U185 (N_185,In_397,In_736);
xor U186 (N_186,In_66,In_322);
or U187 (N_187,In_365,In_446);
or U188 (N_188,In_840,In_196);
and U189 (N_189,In_557,In_857);
or U190 (N_190,In_108,In_394);
and U191 (N_191,In_344,In_185);
or U192 (N_192,In_124,In_462);
and U193 (N_193,In_718,In_279);
nand U194 (N_194,In_406,In_740);
nor U195 (N_195,In_521,In_890);
nand U196 (N_196,In_245,In_632);
nand U197 (N_197,In_589,In_792);
or U198 (N_198,In_706,In_339);
or U199 (N_199,In_437,In_89);
and U200 (N_200,In_363,In_560);
or U201 (N_201,In_372,In_595);
or U202 (N_202,In_107,In_261);
xor U203 (N_203,In_103,In_973);
and U204 (N_204,In_11,In_182);
nor U205 (N_205,In_232,In_700);
nor U206 (N_206,In_725,In_515);
and U207 (N_207,In_325,In_971);
nor U208 (N_208,In_764,In_893);
or U209 (N_209,In_793,In_889);
or U210 (N_210,In_605,In_642);
or U211 (N_211,In_334,In_506);
nand U212 (N_212,In_135,In_412);
nand U213 (N_213,In_585,In_289);
or U214 (N_214,In_866,In_301);
and U215 (N_215,In_238,In_988);
or U216 (N_216,In_474,In_498);
xor U217 (N_217,In_247,In_343);
nand U218 (N_218,In_24,In_493);
and U219 (N_219,In_275,In_985);
and U220 (N_220,In_31,In_708);
nor U221 (N_221,In_991,In_944);
or U222 (N_222,In_654,In_497);
and U223 (N_223,In_217,In_571);
and U224 (N_224,In_138,In_537);
nand U225 (N_225,In_442,In_286);
and U226 (N_226,In_130,In_630);
nor U227 (N_227,In_612,In_647);
nand U228 (N_228,In_327,In_851);
or U229 (N_229,In_421,In_730);
and U230 (N_230,In_113,In_197);
nand U231 (N_231,In_33,In_676);
xnor U232 (N_232,In_897,In_751);
or U233 (N_233,In_701,In_791);
or U234 (N_234,In_916,In_911);
and U235 (N_235,In_270,In_775);
and U236 (N_236,In_704,In_954);
or U237 (N_237,In_374,In_787);
nand U238 (N_238,In_697,In_782);
or U239 (N_239,In_156,In_999);
or U240 (N_240,In_902,In_385);
nand U241 (N_241,In_203,In_798);
xor U242 (N_242,In_259,In_430);
xor U243 (N_243,In_579,In_732);
and U244 (N_244,In_77,In_906);
nor U245 (N_245,In_572,In_220);
nand U246 (N_246,In_300,In_715);
xnor U247 (N_247,In_409,In_180);
and U248 (N_248,In_545,In_691);
and U249 (N_249,In_996,In_744);
nor U250 (N_250,In_13,In_475);
nand U251 (N_251,In_434,In_425);
xor U252 (N_252,In_104,In_880);
nor U253 (N_253,In_333,In_523);
or U254 (N_254,In_547,In_907);
nor U255 (N_255,In_464,In_417);
or U256 (N_256,In_168,In_282);
nor U257 (N_257,In_933,In_534);
and U258 (N_258,In_28,In_338);
and U259 (N_259,In_526,In_188);
nor U260 (N_260,In_221,In_594);
nor U261 (N_261,In_761,In_141);
and U262 (N_262,In_755,In_712);
or U263 (N_263,In_981,In_337);
or U264 (N_264,In_667,In_760);
xnor U265 (N_265,In_0,In_235);
and U266 (N_266,In_230,In_352);
nor U267 (N_267,In_867,In_899);
nor U268 (N_268,In_304,In_639);
nand U269 (N_269,In_137,In_435);
nor U270 (N_270,In_95,In_741);
or U271 (N_271,In_849,In_119);
nand U272 (N_272,In_939,In_780);
nand U273 (N_273,In_163,In_122);
or U274 (N_274,In_870,In_389);
xor U275 (N_275,In_864,In_328);
nand U276 (N_276,In_306,In_226);
and U277 (N_277,In_690,In_392);
or U278 (N_278,In_588,In_530);
xnor U279 (N_279,In_662,In_707);
xor U280 (N_280,In_179,In_12);
or U281 (N_281,In_646,In_285);
nor U282 (N_282,In_265,In_162);
and U283 (N_283,In_257,In_599);
or U284 (N_284,In_573,In_293);
nand U285 (N_285,In_783,In_874);
or U286 (N_286,In_110,In_705);
nand U287 (N_287,In_276,In_896);
nand U288 (N_288,In_620,In_105);
and U289 (N_289,In_205,In_802);
or U290 (N_290,In_830,In_74);
and U291 (N_291,In_111,In_799);
or U292 (N_292,In_405,In_178);
nor U293 (N_293,In_148,In_308);
nand U294 (N_294,In_252,In_924);
nand U295 (N_295,In_128,In_55);
and U296 (N_296,In_937,In_458);
nand U297 (N_297,In_669,In_391);
or U298 (N_298,In_753,In_161);
and U299 (N_299,In_211,In_820);
nor U300 (N_300,In_307,In_656);
and U301 (N_301,In_402,In_703);
and U302 (N_302,In_218,In_519);
and U303 (N_303,In_625,In_686);
and U304 (N_304,In_808,In_953);
or U305 (N_305,In_750,In_711);
nor U306 (N_306,In_340,In_56);
and U307 (N_307,In_553,In_346);
xnor U308 (N_308,In_81,In_659);
and U309 (N_309,In_139,In_488);
and U310 (N_310,In_54,In_158);
and U311 (N_311,In_843,In_948);
and U312 (N_312,In_22,In_132);
nor U313 (N_313,In_192,In_209);
and U314 (N_314,In_839,In_617);
nand U315 (N_315,In_997,In_452);
nor U316 (N_316,In_652,In_884);
and U317 (N_317,In_644,In_559);
nand U318 (N_318,In_533,In_449);
and U319 (N_319,In_255,In_32);
nand U320 (N_320,In_763,In_291);
nand U321 (N_321,In_817,In_878);
or U322 (N_322,In_316,In_578);
nor U323 (N_323,In_502,In_835);
nand U324 (N_324,In_477,In_722);
nand U325 (N_325,In_909,In_811);
nor U326 (N_326,In_513,In_147);
xnor U327 (N_327,In_172,In_5);
and U328 (N_328,In_53,In_809);
nand U329 (N_329,In_408,In_675);
nor U330 (N_330,In_660,In_114);
or U331 (N_331,In_420,In_803);
xnor U332 (N_332,In_784,In_246);
nor U333 (N_333,In_877,In_278);
or U334 (N_334,In_876,In_919);
and U335 (N_335,In_623,In_915);
nor U336 (N_336,In_680,In_940);
nor U337 (N_337,In_456,In_470);
nand U338 (N_338,In_155,In_471);
nand U339 (N_339,In_490,In_977);
nand U340 (N_340,In_689,In_287);
or U341 (N_341,In_865,In_127);
nand U342 (N_342,In_731,In_45);
nor U343 (N_343,In_665,In_556);
or U344 (N_344,In_90,In_97);
or U345 (N_345,In_242,In_963);
nor U346 (N_346,In_294,In_544);
or U347 (N_347,In_38,In_388);
xnor U348 (N_348,In_231,In_202);
and U349 (N_349,In_234,In_25);
or U350 (N_350,In_229,In_214);
xor U351 (N_351,In_668,In_68);
and U352 (N_352,In_735,In_455);
nand U353 (N_353,In_538,In_574);
nand U354 (N_354,In_433,In_892);
nor U355 (N_355,In_404,In_879);
or U356 (N_356,In_737,In_837);
nor U357 (N_357,In_342,In_990);
nand U358 (N_358,In_661,In_958);
xnor U359 (N_359,In_422,In_862);
xnor U360 (N_360,In_535,In_549);
nand U361 (N_361,In_87,In_823);
xnor U362 (N_362,In_262,In_140);
and U363 (N_363,In_41,In_467);
or U364 (N_364,In_486,In_726);
nor U365 (N_365,In_673,In_886);
and U366 (N_366,In_311,In_9);
and U367 (N_367,In_749,In_694);
and U368 (N_368,In_17,In_528);
and U369 (N_369,In_35,In_65);
nand U370 (N_370,In_99,In_901);
nor U371 (N_371,In_52,In_768);
and U372 (N_372,In_743,In_228);
xor U373 (N_373,In_271,In_98);
nor U374 (N_374,In_908,In_536);
nand U375 (N_375,In_894,In_177);
and U376 (N_376,In_727,In_524);
nor U377 (N_377,In_260,In_312);
xnor U378 (N_378,In_810,In_682);
or U379 (N_379,In_175,In_436);
nand U380 (N_380,In_46,In_85);
nand U381 (N_381,In_978,In_93);
or U382 (N_382,In_679,In_819);
nand U383 (N_383,In_317,In_174);
nor U384 (N_384,In_848,In_80);
and U385 (N_385,In_469,In_479);
nor U386 (N_386,In_882,In_558);
xor U387 (N_387,In_674,In_529);
and U388 (N_388,In_4,In_968);
nand U389 (N_389,In_552,In_167);
nand U390 (N_390,In_964,In_752);
and U391 (N_391,In_267,In_354);
or U392 (N_392,In_687,In_274);
and U393 (N_393,In_800,In_331);
nor U394 (N_394,In_243,In_194);
or U395 (N_395,In_699,In_48);
nand U396 (N_396,In_76,In_142);
nor U397 (N_397,In_347,In_204);
or U398 (N_398,In_518,In_465);
nor U399 (N_399,In_423,In_345);
xnor U400 (N_400,In_920,In_129);
nor U401 (N_401,In_918,In_199);
or U402 (N_402,In_222,In_473);
and U403 (N_403,In_284,In_844);
or U404 (N_404,In_468,In_440);
nand U405 (N_405,In_827,In_92);
nor U406 (N_406,In_629,In_253);
nand U407 (N_407,In_250,In_900);
or U408 (N_408,In_487,In_607);
nor U409 (N_409,In_771,In_215);
nand U410 (N_410,In_466,In_789);
or U411 (N_411,In_296,In_3);
nor U412 (N_412,In_861,In_805);
or U413 (N_413,In_613,In_637);
xor U414 (N_414,In_34,In_364);
nor U415 (N_415,In_972,In_945);
nor U416 (N_416,In_774,In_754);
nand U417 (N_417,In_987,In_738);
or U418 (N_418,In_657,In_923);
and U419 (N_419,In_917,In_994);
nand U420 (N_420,In_501,In_314);
xnor U421 (N_421,In_615,In_672);
nand U422 (N_422,In_989,In_852);
and U423 (N_423,In_788,In_216);
nand U424 (N_424,In_739,In_729);
or U425 (N_425,In_349,In_309);
nand U426 (N_426,In_856,In_960);
or U427 (N_427,In_476,In_499);
and U428 (N_428,In_875,In_319);
xor U429 (N_429,In_145,In_539);
or U430 (N_430,In_288,In_100);
nor U431 (N_431,In_244,In_44);
xnor U432 (N_432,In_384,In_375);
or U433 (N_433,In_636,In_664);
and U434 (N_434,In_157,In_663);
or U435 (N_435,In_854,In_281);
nand U436 (N_436,In_806,In_371);
nand U437 (N_437,In_935,In_575);
nor U438 (N_438,In_576,In_512);
xnor U439 (N_439,In_829,In_292);
nor U440 (N_440,In_606,In_212);
nor U441 (N_441,In_441,In_88);
nand U442 (N_442,In_159,In_651);
or U443 (N_443,In_70,In_934);
and U444 (N_444,In_176,In_929);
xnor U445 (N_445,In_638,In_152);
nand U446 (N_446,In_582,In_950);
nor U447 (N_447,In_94,In_489);
and U448 (N_448,In_418,In_510);
or U449 (N_449,In_546,In_845);
nor U450 (N_450,In_258,In_461);
nand U451 (N_451,In_39,In_564);
and U452 (N_452,In_191,In_428);
xnor U453 (N_453,In_169,In_834);
nor U454 (N_454,In_914,In_982);
nand U455 (N_455,In_832,In_888);
xor U456 (N_456,In_532,In_335);
and U457 (N_457,In_777,In_373);
nand U458 (N_458,In_69,In_952);
nand U459 (N_459,In_414,In_491);
and U460 (N_460,In_979,In_208);
or U461 (N_461,In_610,In_299);
and U462 (N_462,In_993,In_974);
nor U463 (N_463,In_728,In_61);
or U464 (N_464,In_841,In_415);
or U465 (N_465,In_249,In_448);
xnor U466 (N_466,In_173,In_818);
xor U467 (N_467,In_186,In_160);
nor U468 (N_468,In_195,In_770);
nor U469 (N_469,In_998,In_517);
nand U470 (N_470,In_472,In_814);
nor U471 (N_471,In_6,In_170);
nand U472 (N_472,In_959,In_330);
or U473 (N_473,In_378,In_946);
and U474 (N_474,In_268,In_457);
nand U475 (N_475,In_144,In_450);
and U476 (N_476,In_561,In_733);
nand U477 (N_477,In_932,In_323);
or U478 (N_478,In_596,In_451);
or U479 (N_479,In_269,In_554);
nand U480 (N_480,In_370,In_396);
and U481 (N_481,In_720,In_947);
nor U482 (N_482,In_904,In_853);
nor U483 (N_483,In_367,In_21);
nand U484 (N_484,In_785,In_1);
nand U485 (N_485,In_633,In_812);
nor U486 (N_486,In_824,In_381);
and U487 (N_487,In_756,In_326);
and U488 (N_488,In_847,In_496);
nand U489 (N_489,In_40,In_913);
nor U490 (N_490,In_995,In_121);
or U491 (N_491,In_131,In_508);
or U492 (N_492,In_815,In_401);
nand U493 (N_493,In_555,In_357);
xnor U494 (N_494,In_930,In_710);
nor U495 (N_495,In_601,In_91);
xor U496 (N_496,In_399,In_883);
and U497 (N_497,In_514,In_826);
nand U498 (N_498,In_603,In_626);
and U499 (N_499,In_641,In_233);
nor U500 (N_500,In_822,In_452);
nor U501 (N_501,In_935,In_836);
or U502 (N_502,In_881,In_698);
xnor U503 (N_503,In_315,In_470);
or U504 (N_504,In_617,In_54);
xnor U505 (N_505,In_282,In_467);
or U506 (N_506,In_889,In_204);
or U507 (N_507,In_70,In_152);
or U508 (N_508,In_502,In_687);
nor U509 (N_509,In_522,In_991);
xnor U510 (N_510,In_228,In_13);
nand U511 (N_511,In_314,In_573);
and U512 (N_512,In_276,In_157);
or U513 (N_513,In_3,In_79);
and U514 (N_514,In_999,In_434);
nand U515 (N_515,In_544,In_85);
nor U516 (N_516,In_625,In_243);
xnor U517 (N_517,In_262,In_938);
nor U518 (N_518,In_731,In_421);
or U519 (N_519,In_555,In_967);
nor U520 (N_520,In_689,In_29);
nor U521 (N_521,In_964,In_652);
or U522 (N_522,In_184,In_24);
and U523 (N_523,In_752,In_856);
or U524 (N_524,In_119,In_405);
xor U525 (N_525,In_375,In_257);
or U526 (N_526,In_256,In_468);
xnor U527 (N_527,In_556,In_153);
nand U528 (N_528,In_704,In_829);
or U529 (N_529,In_164,In_470);
and U530 (N_530,In_826,In_326);
and U531 (N_531,In_940,In_731);
nor U532 (N_532,In_195,In_640);
and U533 (N_533,In_466,In_439);
nor U534 (N_534,In_766,In_694);
nor U535 (N_535,In_657,In_173);
nor U536 (N_536,In_891,In_552);
or U537 (N_537,In_849,In_779);
nand U538 (N_538,In_871,In_861);
and U539 (N_539,In_785,In_766);
and U540 (N_540,In_435,In_449);
or U541 (N_541,In_749,In_673);
nor U542 (N_542,In_831,In_472);
xor U543 (N_543,In_412,In_69);
and U544 (N_544,In_15,In_407);
xnor U545 (N_545,In_221,In_737);
and U546 (N_546,In_722,In_70);
nor U547 (N_547,In_801,In_0);
or U548 (N_548,In_443,In_518);
nor U549 (N_549,In_804,In_543);
nand U550 (N_550,In_376,In_508);
nand U551 (N_551,In_472,In_118);
and U552 (N_552,In_962,In_133);
xnor U553 (N_553,In_477,In_621);
xor U554 (N_554,In_194,In_691);
nor U555 (N_555,In_374,In_942);
nor U556 (N_556,In_172,In_904);
nor U557 (N_557,In_709,In_821);
nor U558 (N_558,In_13,In_281);
nor U559 (N_559,In_571,In_544);
or U560 (N_560,In_320,In_564);
or U561 (N_561,In_830,In_991);
or U562 (N_562,In_743,In_991);
and U563 (N_563,In_892,In_620);
or U564 (N_564,In_438,In_203);
or U565 (N_565,In_105,In_802);
or U566 (N_566,In_759,In_949);
nor U567 (N_567,In_992,In_372);
and U568 (N_568,In_418,In_635);
nor U569 (N_569,In_908,In_520);
and U570 (N_570,In_516,In_585);
and U571 (N_571,In_72,In_215);
nand U572 (N_572,In_334,In_499);
and U573 (N_573,In_645,In_845);
nor U574 (N_574,In_276,In_72);
nand U575 (N_575,In_551,In_51);
or U576 (N_576,In_33,In_392);
nand U577 (N_577,In_623,In_675);
nand U578 (N_578,In_966,In_697);
nand U579 (N_579,In_471,In_465);
and U580 (N_580,In_778,In_980);
and U581 (N_581,In_590,In_386);
nor U582 (N_582,In_492,In_328);
nand U583 (N_583,In_567,In_486);
and U584 (N_584,In_571,In_188);
xor U585 (N_585,In_611,In_813);
or U586 (N_586,In_830,In_547);
nor U587 (N_587,In_123,In_612);
or U588 (N_588,In_7,In_780);
and U589 (N_589,In_41,In_2);
or U590 (N_590,In_993,In_125);
and U591 (N_591,In_173,In_700);
xor U592 (N_592,In_396,In_604);
nor U593 (N_593,In_253,In_381);
or U594 (N_594,In_625,In_942);
nor U595 (N_595,In_539,In_552);
nor U596 (N_596,In_522,In_699);
nor U597 (N_597,In_631,In_579);
and U598 (N_598,In_296,In_575);
nand U599 (N_599,In_571,In_122);
nor U600 (N_600,In_817,In_193);
xor U601 (N_601,In_168,In_612);
nand U602 (N_602,In_776,In_273);
or U603 (N_603,In_430,In_517);
nand U604 (N_604,In_750,In_402);
nor U605 (N_605,In_880,In_855);
and U606 (N_606,In_599,In_291);
or U607 (N_607,In_687,In_542);
or U608 (N_608,In_109,In_788);
or U609 (N_609,In_401,In_603);
nor U610 (N_610,In_393,In_250);
or U611 (N_611,In_651,In_101);
or U612 (N_612,In_975,In_519);
and U613 (N_613,In_139,In_936);
or U614 (N_614,In_50,In_428);
nand U615 (N_615,In_697,In_990);
and U616 (N_616,In_808,In_309);
and U617 (N_617,In_701,In_960);
and U618 (N_618,In_373,In_599);
and U619 (N_619,In_444,In_979);
nand U620 (N_620,In_515,In_795);
nand U621 (N_621,In_837,In_42);
nor U622 (N_622,In_486,In_796);
xnor U623 (N_623,In_884,In_902);
nand U624 (N_624,In_492,In_86);
nor U625 (N_625,In_275,In_763);
or U626 (N_626,In_464,In_213);
nand U627 (N_627,In_563,In_839);
and U628 (N_628,In_350,In_69);
nand U629 (N_629,In_12,In_579);
or U630 (N_630,In_902,In_589);
or U631 (N_631,In_950,In_328);
nand U632 (N_632,In_396,In_930);
nand U633 (N_633,In_765,In_12);
or U634 (N_634,In_350,In_121);
nand U635 (N_635,In_397,In_962);
nand U636 (N_636,In_754,In_532);
nor U637 (N_637,In_474,In_791);
or U638 (N_638,In_794,In_728);
nand U639 (N_639,In_120,In_905);
or U640 (N_640,In_299,In_791);
nor U641 (N_641,In_831,In_200);
nor U642 (N_642,In_4,In_222);
xor U643 (N_643,In_433,In_114);
nor U644 (N_644,In_301,In_231);
or U645 (N_645,In_560,In_427);
nand U646 (N_646,In_982,In_918);
or U647 (N_647,In_356,In_756);
or U648 (N_648,In_26,In_256);
nor U649 (N_649,In_134,In_21);
nor U650 (N_650,In_87,In_706);
or U651 (N_651,In_83,In_175);
nor U652 (N_652,In_323,In_711);
nand U653 (N_653,In_754,In_428);
nand U654 (N_654,In_304,In_928);
nor U655 (N_655,In_168,In_100);
and U656 (N_656,In_262,In_948);
nor U657 (N_657,In_57,In_450);
or U658 (N_658,In_426,In_693);
or U659 (N_659,In_698,In_906);
xnor U660 (N_660,In_733,In_531);
or U661 (N_661,In_26,In_422);
and U662 (N_662,In_550,In_161);
or U663 (N_663,In_193,In_927);
nor U664 (N_664,In_454,In_114);
and U665 (N_665,In_741,In_571);
or U666 (N_666,In_303,In_127);
or U667 (N_667,In_278,In_741);
and U668 (N_668,In_637,In_559);
nand U669 (N_669,In_65,In_49);
nand U670 (N_670,In_302,In_581);
nand U671 (N_671,In_981,In_298);
nand U672 (N_672,In_235,In_923);
or U673 (N_673,In_160,In_543);
nor U674 (N_674,In_137,In_887);
and U675 (N_675,In_291,In_623);
nand U676 (N_676,In_428,In_874);
nand U677 (N_677,In_351,In_391);
nand U678 (N_678,In_105,In_386);
or U679 (N_679,In_395,In_207);
nor U680 (N_680,In_716,In_261);
or U681 (N_681,In_248,In_29);
nand U682 (N_682,In_160,In_240);
and U683 (N_683,In_564,In_701);
and U684 (N_684,In_535,In_203);
nor U685 (N_685,In_392,In_914);
and U686 (N_686,In_551,In_760);
nor U687 (N_687,In_694,In_286);
xnor U688 (N_688,In_458,In_214);
and U689 (N_689,In_718,In_469);
and U690 (N_690,In_496,In_105);
or U691 (N_691,In_991,In_291);
nor U692 (N_692,In_382,In_800);
and U693 (N_693,In_225,In_851);
xor U694 (N_694,In_424,In_852);
and U695 (N_695,In_62,In_378);
nor U696 (N_696,In_938,In_909);
nor U697 (N_697,In_299,In_278);
nand U698 (N_698,In_365,In_828);
nor U699 (N_699,In_125,In_649);
nand U700 (N_700,In_829,In_388);
xor U701 (N_701,In_469,In_797);
nand U702 (N_702,In_992,In_831);
and U703 (N_703,In_112,In_299);
or U704 (N_704,In_278,In_404);
nand U705 (N_705,In_118,In_218);
or U706 (N_706,In_467,In_455);
and U707 (N_707,In_38,In_592);
nand U708 (N_708,In_867,In_370);
nor U709 (N_709,In_368,In_524);
and U710 (N_710,In_977,In_894);
nor U711 (N_711,In_331,In_960);
nor U712 (N_712,In_974,In_150);
nand U713 (N_713,In_191,In_822);
xnor U714 (N_714,In_843,In_730);
or U715 (N_715,In_859,In_402);
and U716 (N_716,In_593,In_860);
nand U717 (N_717,In_548,In_728);
and U718 (N_718,In_60,In_246);
or U719 (N_719,In_584,In_225);
nor U720 (N_720,In_416,In_518);
and U721 (N_721,In_207,In_642);
or U722 (N_722,In_540,In_965);
xnor U723 (N_723,In_931,In_75);
or U724 (N_724,In_870,In_129);
and U725 (N_725,In_719,In_991);
and U726 (N_726,In_946,In_288);
or U727 (N_727,In_294,In_145);
and U728 (N_728,In_513,In_851);
and U729 (N_729,In_199,In_336);
xnor U730 (N_730,In_726,In_388);
and U731 (N_731,In_454,In_427);
nor U732 (N_732,In_168,In_576);
or U733 (N_733,In_5,In_938);
xor U734 (N_734,In_444,In_514);
or U735 (N_735,In_666,In_191);
and U736 (N_736,In_405,In_97);
or U737 (N_737,In_619,In_488);
or U738 (N_738,In_108,In_889);
nand U739 (N_739,In_799,In_672);
and U740 (N_740,In_451,In_522);
or U741 (N_741,In_887,In_451);
or U742 (N_742,In_980,In_348);
and U743 (N_743,In_582,In_238);
and U744 (N_744,In_976,In_162);
nor U745 (N_745,In_94,In_979);
nand U746 (N_746,In_524,In_567);
and U747 (N_747,In_427,In_622);
and U748 (N_748,In_366,In_122);
and U749 (N_749,In_553,In_126);
xor U750 (N_750,In_940,In_869);
or U751 (N_751,In_104,In_508);
or U752 (N_752,In_308,In_609);
nor U753 (N_753,In_522,In_701);
and U754 (N_754,In_299,In_442);
nand U755 (N_755,In_147,In_38);
nand U756 (N_756,In_69,In_234);
or U757 (N_757,In_352,In_278);
or U758 (N_758,In_122,In_499);
or U759 (N_759,In_586,In_831);
xor U760 (N_760,In_721,In_494);
nor U761 (N_761,In_64,In_554);
nand U762 (N_762,In_968,In_462);
xor U763 (N_763,In_365,In_58);
and U764 (N_764,In_787,In_137);
and U765 (N_765,In_186,In_122);
xor U766 (N_766,In_348,In_157);
nand U767 (N_767,In_591,In_71);
or U768 (N_768,In_468,In_765);
nand U769 (N_769,In_362,In_377);
nand U770 (N_770,In_326,In_187);
nand U771 (N_771,In_522,In_439);
and U772 (N_772,In_642,In_191);
or U773 (N_773,In_206,In_948);
nor U774 (N_774,In_713,In_868);
nor U775 (N_775,In_304,In_982);
and U776 (N_776,In_853,In_940);
and U777 (N_777,In_436,In_154);
or U778 (N_778,In_397,In_668);
nand U779 (N_779,In_233,In_80);
and U780 (N_780,In_862,In_975);
nand U781 (N_781,In_633,In_146);
and U782 (N_782,In_935,In_959);
and U783 (N_783,In_893,In_577);
and U784 (N_784,In_516,In_664);
nand U785 (N_785,In_414,In_709);
xor U786 (N_786,In_147,In_39);
nand U787 (N_787,In_765,In_672);
nand U788 (N_788,In_145,In_547);
or U789 (N_789,In_524,In_589);
or U790 (N_790,In_770,In_404);
nor U791 (N_791,In_180,In_96);
nor U792 (N_792,In_52,In_38);
nand U793 (N_793,In_605,In_499);
and U794 (N_794,In_743,In_92);
nand U795 (N_795,In_72,In_805);
nand U796 (N_796,In_2,In_146);
nand U797 (N_797,In_14,In_95);
nor U798 (N_798,In_701,In_559);
xor U799 (N_799,In_756,In_137);
and U800 (N_800,In_904,In_430);
and U801 (N_801,In_115,In_632);
nand U802 (N_802,In_496,In_936);
nand U803 (N_803,In_273,In_942);
nor U804 (N_804,In_297,In_336);
or U805 (N_805,In_89,In_988);
and U806 (N_806,In_415,In_124);
and U807 (N_807,In_479,In_415);
nand U808 (N_808,In_56,In_148);
and U809 (N_809,In_924,In_637);
nand U810 (N_810,In_906,In_556);
xor U811 (N_811,In_453,In_296);
nor U812 (N_812,In_181,In_922);
or U813 (N_813,In_411,In_911);
or U814 (N_814,In_81,In_571);
nand U815 (N_815,In_653,In_208);
or U816 (N_816,In_53,In_40);
nand U817 (N_817,In_431,In_867);
or U818 (N_818,In_723,In_445);
and U819 (N_819,In_960,In_542);
nor U820 (N_820,In_933,In_23);
or U821 (N_821,In_799,In_452);
nand U822 (N_822,In_828,In_616);
xor U823 (N_823,In_813,In_591);
nand U824 (N_824,In_272,In_34);
nor U825 (N_825,In_141,In_33);
nand U826 (N_826,In_804,In_601);
or U827 (N_827,In_249,In_327);
nor U828 (N_828,In_813,In_485);
nand U829 (N_829,In_800,In_129);
nand U830 (N_830,In_575,In_420);
and U831 (N_831,In_876,In_638);
xnor U832 (N_832,In_488,In_646);
and U833 (N_833,In_168,In_87);
nand U834 (N_834,In_765,In_944);
and U835 (N_835,In_419,In_318);
and U836 (N_836,In_87,In_44);
nand U837 (N_837,In_269,In_916);
or U838 (N_838,In_926,In_181);
or U839 (N_839,In_758,In_392);
and U840 (N_840,In_163,In_731);
or U841 (N_841,In_337,In_940);
or U842 (N_842,In_328,In_938);
xnor U843 (N_843,In_250,In_627);
nor U844 (N_844,In_27,In_21);
nor U845 (N_845,In_51,In_345);
nor U846 (N_846,In_635,In_931);
nor U847 (N_847,In_36,In_948);
xor U848 (N_848,In_142,In_267);
nand U849 (N_849,In_208,In_256);
nor U850 (N_850,In_774,In_629);
nand U851 (N_851,In_131,In_201);
and U852 (N_852,In_309,In_668);
nand U853 (N_853,In_193,In_139);
nand U854 (N_854,In_858,In_161);
or U855 (N_855,In_519,In_302);
or U856 (N_856,In_420,In_819);
or U857 (N_857,In_2,In_209);
or U858 (N_858,In_963,In_104);
nand U859 (N_859,In_426,In_973);
nor U860 (N_860,In_659,In_646);
nor U861 (N_861,In_543,In_98);
nor U862 (N_862,In_793,In_581);
nand U863 (N_863,In_3,In_960);
or U864 (N_864,In_536,In_871);
nand U865 (N_865,In_536,In_307);
or U866 (N_866,In_375,In_288);
and U867 (N_867,In_453,In_682);
or U868 (N_868,In_84,In_701);
or U869 (N_869,In_792,In_465);
nor U870 (N_870,In_871,In_478);
or U871 (N_871,In_157,In_45);
nor U872 (N_872,In_893,In_807);
xor U873 (N_873,In_443,In_945);
and U874 (N_874,In_348,In_50);
nor U875 (N_875,In_689,In_632);
nand U876 (N_876,In_641,In_982);
and U877 (N_877,In_177,In_721);
nor U878 (N_878,In_774,In_684);
nand U879 (N_879,In_218,In_946);
nor U880 (N_880,In_748,In_125);
xnor U881 (N_881,In_659,In_380);
or U882 (N_882,In_212,In_944);
or U883 (N_883,In_610,In_653);
nor U884 (N_884,In_667,In_525);
and U885 (N_885,In_843,In_779);
nor U886 (N_886,In_95,In_861);
and U887 (N_887,In_784,In_391);
xor U888 (N_888,In_598,In_987);
or U889 (N_889,In_412,In_263);
nand U890 (N_890,In_964,In_537);
and U891 (N_891,In_901,In_868);
or U892 (N_892,In_251,In_272);
nand U893 (N_893,In_484,In_84);
or U894 (N_894,In_813,In_511);
or U895 (N_895,In_169,In_870);
or U896 (N_896,In_669,In_594);
nand U897 (N_897,In_242,In_142);
or U898 (N_898,In_623,In_790);
nor U899 (N_899,In_578,In_52);
nand U900 (N_900,In_589,In_302);
nand U901 (N_901,In_364,In_293);
nand U902 (N_902,In_421,In_52);
nand U903 (N_903,In_516,In_23);
nand U904 (N_904,In_412,In_390);
or U905 (N_905,In_143,In_283);
nor U906 (N_906,In_19,In_364);
and U907 (N_907,In_991,In_119);
or U908 (N_908,In_728,In_667);
xor U909 (N_909,In_129,In_931);
and U910 (N_910,In_911,In_259);
or U911 (N_911,In_14,In_435);
or U912 (N_912,In_737,In_129);
and U913 (N_913,In_823,In_610);
or U914 (N_914,In_986,In_997);
nor U915 (N_915,In_267,In_211);
xor U916 (N_916,In_797,In_137);
nand U917 (N_917,In_407,In_604);
nor U918 (N_918,In_551,In_910);
nor U919 (N_919,In_428,In_152);
nand U920 (N_920,In_214,In_946);
and U921 (N_921,In_759,In_247);
or U922 (N_922,In_394,In_797);
nor U923 (N_923,In_440,In_603);
nor U924 (N_924,In_439,In_699);
nand U925 (N_925,In_654,In_883);
or U926 (N_926,In_482,In_437);
and U927 (N_927,In_817,In_655);
nand U928 (N_928,In_871,In_406);
and U929 (N_929,In_75,In_216);
nor U930 (N_930,In_811,In_457);
xor U931 (N_931,In_596,In_628);
nor U932 (N_932,In_611,In_224);
or U933 (N_933,In_229,In_604);
nor U934 (N_934,In_972,In_561);
nand U935 (N_935,In_429,In_184);
and U936 (N_936,In_708,In_694);
and U937 (N_937,In_579,In_422);
or U938 (N_938,In_31,In_421);
and U939 (N_939,In_621,In_575);
and U940 (N_940,In_152,In_846);
xnor U941 (N_941,In_187,In_106);
nand U942 (N_942,In_132,In_663);
xor U943 (N_943,In_127,In_486);
nor U944 (N_944,In_607,In_476);
nor U945 (N_945,In_161,In_650);
and U946 (N_946,In_50,In_576);
nor U947 (N_947,In_733,In_730);
or U948 (N_948,In_306,In_707);
or U949 (N_949,In_864,In_452);
nor U950 (N_950,In_713,In_895);
and U951 (N_951,In_819,In_942);
nor U952 (N_952,In_701,In_235);
nor U953 (N_953,In_333,In_235);
nand U954 (N_954,In_104,In_725);
nand U955 (N_955,In_885,In_168);
nor U956 (N_956,In_87,In_306);
nor U957 (N_957,In_419,In_927);
nand U958 (N_958,In_97,In_863);
xor U959 (N_959,In_160,In_455);
nand U960 (N_960,In_416,In_935);
nand U961 (N_961,In_782,In_14);
or U962 (N_962,In_310,In_612);
nand U963 (N_963,In_40,In_673);
nand U964 (N_964,In_453,In_132);
nand U965 (N_965,In_222,In_48);
nor U966 (N_966,In_332,In_991);
nor U967 (N_967,In_603,In_808);
and U968 (N_968,In_509,In_841);
and U969 (N_969,In_685,In_772);
nor U970 (N_970,In_851,In_96);
or U971 (N_971,In_562,In_341);
nor U972 (N_972,In_187,In_69);
nor U973 (N_973,In_970,In_223);
nor U974 (N_974,In_639,In_670);
nand U975 (N_975,In_828,In_950);
nand U976 (N_976,In_16,In_262);
and U977 (N_977,In_403,In_345);
xor U978 (N_978,In_898,In_756);
nor U979 (N_979,In_434,In_180);
and U980 (N_980,In_924,In_430);
or U981 (N_981,In_340,In_285);
nand U982 (N_982,In_29,In_691);
nor U983 (N_983,In_419,In_657);
and U984 (N_984,In_321,In_760);
xor U985 (N_985,In_380,In_487);
or U986 (N_986,In_123,In_80);
nand U987 (N_987,In_143,In_507);
xnor U988 (N_988,In_215,In_25);
nand U989 (N_989,In_925,In_664);
or U990 (N_990,In_415,In_271);
or U991 (N_991,In_340,In_359);
and U992 (N_992,In_918,In_680);
and U993 (N_993,In_943,In_812);
nor U994 (N_994,In_164,In_285);
and U995 (N_995,In_49,In_475);
and U996 (N_996,In_81,In_333);
and U997 (N_997,In_184,In_303);
nand U998 (N_998,In_886,In_930);
or U999 (N_999,In_377,In_242);
nor U1000 (N_1000,In_607,In_46);
or U1001 (N_1001,In_669,In_554);
or U1002 (N_1002,In_827,In_223);
nor U1003 (N_1003,In_8,In_977);
nand U1004 (N_1004,In_368,In_162);
nor U1005 (N_1005,In_780,In_302);
nor U1006 (N_1006,In_142,In_16);
and U1007 (N_1007,In_146,In_893);
nand U1008 (N_1008,In_980,In_123);
and U1009 (N_1009,In_390,In_371);
nor U1010 (N_1010,In_532,In_686);
xor U1011 (N_1011,In_36,In_309);
nand U1012 (N_1012,In_890,In_354);
and U1013 (N_1013,In_50,In_836);
nand U1014 (N_1014,In_371,In_73);
nor U1015 (N_1015,In_630,In_308);
or U1016 (N_1016,In_115,In_751);
or U1017 (N_1017,In_359,In_750);
and U1018 (N_1018,In_477,In_555);
or U1019 (N_1019,In_315,In_827);
nor U1020 (N_1020,In_1,In_709);
nor U1021 (N_1021,In_617,In_528);
or U1022 (N_1022,In_726,In_178);
nor U1023 (N_1023,In_966,In_329);
nor U1024 (N_1024,In_314,In_417);
nor U1025 (N_1025,In_278,In_128);
and U1026 (N_1026,In_556,In_233);
nor U1027 (N_1027,In_671,In_728);
nand U1028 (N_1028,In_361,In_918);
and U1029 (N_1029,In_948,In_551);
nand U1030 (N_1030,In_657,In_193);
or U1031 (N_1031,In_702,In_352);
nor U1032 (N_1032,In_382,In_120);
nand U1033 (N_1033,In_24,In_92);
xor U1034 (N_1034,In_765,In_285);
nand U1035 (N_1035,In_752,In_523);
nor U1036 (N_1036,In_401,In_318);
or U1037 (N_1037,In_558,In_297);
and U1038 (N_1038,In_555,In_204);
nor U1039 (N_1039,In_908,In_930);
nor U1040 (N_1040,In_179,In_403);
nor U1041 (N_1041,In_666,In_845);
nor U1042 (N_1042,In_428,In_263);
and U1043 (N_1043,In_224,In_686);
nand U1044 (N_1044,In_787,In_897);
and U1045 (N_1045,In_340,In_379);
nor U1046 (N_1046,In_59,In_831);
xor U1047 (N_1047,In_661,In_77);
and U1048 (N_1048,In_794,In_38);
nor U1049 (N_1049,In_421,In_906);
nor U1050 (N_1050,In_977,In_979);
or U1051 (N_1051,In_952,In_388);
or U1052 (N_1052,In_834,In_143);
nand U1053 (N_1053,In_993,In_199);
nand U1054 (N_1054,In_319,In_713);
xnor U1055 (N_1055,In_714,In_265);
nor U1056 (N_1056,In_41,In_639);
and U1057 (N_1057,In_431,In_465);
and U1058 (N_1058,In_105,In_773);
or U1059 (N_1059,In_385,In_324);
or U1060 (N_1060,In_569,In_800);
and U1061 (N_1061,In_173,In_806);
or U1062 (N_1062,In_297,In_857);
nand U1063 (N_1063,In_383,In_920);
or U1064 (N_1064,In_667,In_369);
and U1065 (N_1065,In_936,In_177);
nor U1066 (N_1066,In_596,In_321);
and U1067 (N_1067,In_610,In_283);
nor U1068 (N_1068,In_889,In_881);
or U1069 (N_1069,In_666,In_585);
nand U1070 (N_1070,In_503,In_967);
and U1071 (N_1071,In_894,In_812);
xor U1072 (N_1072,In_846,In_367);
nor U1073 (N_1073,In_800,In_441);
nor U1074 (N_1074,In_686,In_883);
nand U1075 (N_1075,In_90,In_743);
xor U1076 (N_1076,In_675,In_79);
nand U1077 (N_1077,In_366,In_881);
nand U1078 (N_1078,In_899,In_194);
xnor U1079 (N_1079,In_922,In_667);
and U1080 (N_1080,In_252,In_334);
xor U1081 (N_1081,In_939,In_709);
nand U1082 (N_1082,In_425,In_985);
nor U1083 (N_1083,In_983,In_385);
or U1084 (N_1084,In_177,In_80);
nor U1085 (N_1085,In_185,In_663);
nand U1086 (N_1086,In_84,In_990);
or U1087 (N_1087,In_41,In_14);
and U1088 (N_1088,In_830,In_580);
or U1089 (N_1089,In_188,In_285);
or U1090 (N_1090,In_177,In_904);
or U1091 (N_1091,In_421,In_771);
or U1092 (N_1092,In_391,In_751);
nand U1093 (N_1093,In_895,In_863);
nand U1094 (N_1094,In_858,In_619);
nand U1095 (N_1095,In_24,In_869);
or U1096 (N_1096,In_288,In_666);
nor U1097 (N_1097,In_641,In_723);
nor U1098 (N_1098,In_631,In_14);
and U1099 (N_1099,In_335,In_541);
or U1100 (N_1100,In_753,In_929);
and U1101 (N_1101,In_917,In_566);
or U1102 (N_1102,In_333,In_60);
nor U1103 (N_1103,In_284,In_888);
nor U1104 (N_1104,In_381,In_548);
and U1105 (N_1105,In_820,In_240);
and U1106 (N_1106,In_333,In_992);
or U1107 (N_1107,In_923,In_468);
nor U1108 (N_1108,In_758,In_221);
or U1109 (N_1109,In_792,In_964);
or U1110 (N_1110,In_221,In_36);
xnor U1111 (N_1111,In_720,In_582);
or U1112 (N_1112,In_80,In_905);
xor U1113 (N_1113,In_52,In_536);
xor U1114 (N_1114,In_230,In_583);
or U1115 (N_1115,In_189,In_977);
or U1116 (N_1116,In_686,In_80);
and U1117 (N_1117,In_764,In_372);
or U1118 (N_1118,In_576,In_675);
nor U1119 (N_1119,In_839,In_700);
or U1120 (N_1120,In_930,In_95);
nand U1121 (N_1121,In_930,In_354);
nand U1122 (N_1122,In_521,In_284);
nor U1123 (N_1123,In_424,In_57);
or U1124 (N_1124,In_416,In_144);
nor U1125 (N_1125,In_987,In_796);
and U1126 (N_1126,In_867,In_166);
or U1127 (N_1127,In_729,In_776);
nand U1128 (N_1128,In_292,In_181);
nand U1129 (N_1129,In_445,In_766);
xnor U1130 (N_1130,In_709,In_3);
nor U1131 (N_1131,In_414,In_201);
or U1132 (N_1132,In_911,In_733);
nor U1133 (N_1133,In_572,In_274);
nand U1134 (N_1134,In_811,In_660);
nor U1135 (N_1135,In_336,In_782);
and U1136 (N_1136,In_304,In_369);
nand U1137 (N_1137,In_860,In_6);
nor U1138 (N_1138,In_943,In_45);
nand U1139 (N_1139,In_965,In_844);
nand U1140 (N_1140,In_100,In_844);
and U1141 (N_1141,In_774,In_640);
xor U1142 (N_1142,In_658,In_150);
xor U1143 (N_1143,In_420,In_407);
or U1144 (N_1144,In_882,In_775);
or U1145 (N_1145,In_712,In_444);
or U1146 (N_1146,In_584,In_524);
nor U1147 (N_1147,In_111,In_926);
or U1148 (N_1148,In_266,In_180);
nor U1149 (N_1149,In_548,In_925);
nor U1150 (N_1150,In_220,In_517);
nand U1151 (N_1151,In_72,In_606);
and U1152 (N_1152,In_111,In_919);
nand U1153 (N_1153,In_636,In_253);
or U1154 (N_1154,In_253,In_430);
or U1155 (N_1155,In_386,In_371);
nand U1156 (N_1156,In_758,In_969);
or U1157 (N_1157,In_922,In_281);
and U1158 (N_1158,In_846,In_626);
and U1159 (N_1159,In_776,In_257);
or U1160 (N_1160,In_478,In_124);
or U1161 (N_1161,In_24,In_32);
nand U1162 (N_1162,In_909,In_131);
or U1163 (N_1163,In_420,In_396);
nand U1164 (N_1164,In_461,In_111);
and U1165 (N_1165,In_319,In_819);
nand U1166 (N_1166,In_451,In_802);
nor U1167 (N_1167,In_115,In_68);
and U1168 (N_1168,In_589,In_629);
nand U1169 (N_1169,In_542,In_372);
nand U1170 (N_1170,In_698,In_271);
nor U1171 (N_1171,In_659,In_135);
or U1172 (N_1172,In_863,In_30);
or U1173 (N_1173,In_348,In_323);
or U1174 (N_1174,In_300,In_678);
nand U1175 (N_1175,In_576,In_292);
nor U1176 (N_1176,In_565,In_481);
xnor U1177 (N_1177,In_559,In_787);
xnor U1178 (N_1178,In_499,In_330);
or U1179 (N_1179,In_959,In_340);
nor U1180 (N_1180,In_123,In_405);
and U1181 (N_1181,In_950,In_663);
or U1182 (N_1182,In_427,In_930);
and U1183 (N_1183,In_914,In_252);
nand U1184 (N_1184,In_768,In_767);
nor U1185 (N_1185,In_66,In_96);
and U1186 (N_1186,In_231,In_282);
nand U1187 (N_1187,In_861,In_18);
or U1188 (N_1188,In_38,In_30);
nor U1189 (N_1189,In_179,In_411);
nor U1190 (N_1190,In_336,In_107);
nand U1191 (N_1191,In_825,In_434);
or U1192 (N_1192,In_175,In_96);
or U1193 (N_1193,In_202,In_461);
or U1194 (N_1194,In_321,In_211);
nand U1195 (N_1195,In_86,In_263);
nand U1196 (N_1196,In_407,In_882);
and U1197 (N_1197,In_281,In_126);
nor U1198 (N_1198,In_832,In_643);
nand U1199 (N_1199,In_474,In_311);
nand U1200 (N_1200,In_650,In_726);
nand U1201 (N_1201,In_227,In_412);
or U1202 (N_1202,In_230,In_559);
nor U1203 (N_1203,In_466,In_760);
and U1204 (N_1204,In_132,In_558);
or U1205 (N_1205,In_400,In_298);
and U1206 (N_1206,In_237,In_670);
and U1207 (N_1207,In_418,In_284);
nor U1208 (N_1208,In_707,In_920);
or U1209 (N_1209,In_644,In_388);
nor U1210 (N_1210,In_216,In_871);
nand U1211 (N_1211,In_799,In_581);
nor U1212 (N_1212,In_351,In_398);
and U1213 (N_1213,In_866,In_901);
nor U1214 (N_1214,In_686,In_808);
nand U1215 (N_1215,In_988,In_342);
nor U1216 (N_1216,In_947,In_569);
nand U1217 (N_1217,In_315,In_247);
and U1218 (N_1218,In_99,In_198);
nor U1219 (N_1219,In_113,In_517);
nor U1220 (N_1220,In_489,In_906);
and U1221 (N_1221,In_404,In_453);
or U1222 (N_1222,In_894,In_317);
or U1223 (N_1223,In_530,In_804);
and U1224 (N_1224,In_785,In_264);
nand U1225 (N_1225,In_996,In_831);
and U1226 (N_1226,In_15,In_535);
nand U1227 (N_1227,In_847,In_594);
or U1228 (N_1228,In_17,In_307);
xnor U1229 (N_1229,In_771,In_611);
or U1230 (N_1230,In_617,In_277);
nor U1231 (N_1231,In_449,In_748);
nand U1232 (N_1232,In_953,In_49);
xor U1233 (N_1233,In_628,In_394);
or U1234 (N_1234,In_494,In_796);
and U1235 (N_1235,In_913,In_496);
nor U1236 (N_1236,In_494,In_167);
nand U1237 (N_1237,In_411,In_652);
or U1238 (N_1238,In_844,In_661);
or U1239 (N_1239,In_870,In_416);
or U1240 (N_1240,In_373,In_213);
nor U1241 (N_1241,In_292,In_749);
and U1242 (N_1242,In_870,In_922);
and U1243 (N_1243,In_209,In_213);
xnor U1244 (N_1244,In_574,In_440);
nand U1245 (N_1245,In_392,In_908);
or U1246 (N_1246,In_831,In_552);
nor U1247 (N_1247,In_354,In_831);
nor U1248 (N_1248,In_60,In_887);
nor U1249 (N_1249,In_60,In_444);
nand U1250 (N_1250,In_13,In_625);
or U1251 (N_1251,In_303,In_741);
nand U1252 (N_1252,In_359,In_885);
nand U1253 (N_1253,In_442,In_65);
nand U1254 (N_1254,In_139,In_951);
and U1255 (N_1255,In_776,In_921);
nor U1256 (N_1256,In_436,In_89);
nor U1257 (N_1257,In_127,In_22);
or U1258 (N_1258,In_451,In_740);
and U1259 (N_1259,In_632,In_301);
and U1260 (N_1260,In_240,In_180);
xnor U1261 (N_1261,In_934,In_708);
nor U1262 (N_1262,In_799,In_258);
nor U1263 (N_1263,In_897,In_738);
xnor U1264 (N_1264,In_491,In_958);
nand U1265 (N_1265,In_832,In_894);
or U1266 (N_1266,In_240,In_762);
and U1267 (N_1267,In_889,In_734);
xnor U1268 (N_1268,In_549,In_252);
nand U1269 (N_1269,In_100,In_251);
nand U1270 (N_1270,In_659,In_297);
nand U1271 (N_1271,In_746,In_65);
or U1272 (N_1272,In_698,In_488);
nand U1273 (N_1273,In_292,In_324);
nand U1274 (N_1274,In_199,In_521);
nor U1275 (N_1275,In_777,In_543);
and U1276 (N_1276,In_924,In_932);
nand U1277 (N_1277,In_51,In_701);
nor U1278 (N_1278,In_161,In_528);
nand U1279 (N_1279,In_310,In_144);
nand U1280 (N_1280,In_926,In_594);
xor U1281 (N_1281,In_509,In_383);
or U1282 (N_1282,In_689,In_999);
nor U1283 (N_1283,In_186,In_832);
xnor U1284 (N_1284,In_395,In_438);
nor U1285 (N_1285,In_954,In_409);
and U1286 (N_1286,In_47,In_962);
and U1287 (N_1287,In_485,In_175);
and U1288 (N_1288,In_148,In_292);
and U1289 (N_1289,In_400,In_203);
xor U1290 (N_1290,In_896,In_778);
xor U1291 (N_1291,In_759,In_589);
or U1292 (N_1292,In_628,In_959);
nand U1293 (N_1293,In_709,In_416);
nor U1294 (N_1294,In_620,In_455);
nor U1295 (N_1295,In_191,In_820);
nor U1296 (N_1296,In_384,In_843);
or U1297 (N_1297,In_334,In_323);
xnor U1298 (N_1298,In_520,In_323);
or U1299 (N_1299,In_585,In_228);
nand U1300 (N_1300,In_726,In_679);
nor U1301 (N_1301,In_913,In_994);
nor U1302 (N_1302,In_192,In_494);
and U1303 (N_1303,In_106,In_55);
nor U1304 (N_1304,In_2,In_344);
nor U1305 (N_1305,In_580,In_871);
or U1306 (N_1306,In_975,In_11);
xnor U1307 (N_1307,In_906,In_175);
xor U1308 (N_1308,In_481,In_372);
nand U1309 (N_1309,In_971,In_669);
nor U1310 (N_1310,In_58,In_393);
nand U1311 (N_1311,In_226,In_976);
nand U1312 (N_1312,In_974,In_548);
nor U1313 (N_1313,In_223,In_557);
or U1314 (N_1314,In_808,In_81);
nand U1315 (N_1315,In_698,In_229);
nand U1316 (N_1316,In_117,In_400);
nand U1317 (N_1317,In_357,In_874);
nand U1318 (N_1318,In_154,In_628);
or U1319 (N_1319,In_841,In_73);
nor U1320 (N_1320,In_905,In_50);
or U1321 (N_1321,In_247,In_930);
and U1322 (N_1322,In_149,In_322);
or U1323 (N_1323,In_126,In_835);
nor U1324 (N_1324,In_104,In_288);
and U1325 (N_1325,In_270,In_609);
nor U1326 (N_1326,In_585,In_397);
nand U1327 (N_1327,In_918,In_365);
xor U1328 (N_1328,In_867,In_411);
or U1329 (N_1329,In_215,In_475);
or U1330 (N_1330,In_343,In_136);
and U1331 (N_1331,In_123,In_42);
nor U1332 (N_1332,In_185,In_75);
xor U1333 (N_1333,In_502,In_454);
xor U1334 (N_1334,In_707,In_17);
xor U1335 (N_1335,In_147,In_391);
or U1336 (N_1336,In_797,In_416);
nor U1337 (N_1337,In_837,In_118);
nor U1338 (N_1338,In_554,In_498);
and U1339 (N_1339,In_903,In_562);
or U1340 (N_1340,In_960,In_176);
nor U1341 (N_1341,In_713,In_726);
nor U1342 (N_1342,In_82,In_286);
nor U1343 (N_1343,In_187,In_660);
nor U1344 (N_1344,In_58,In_144);
and U1345 (N_1345,In_165,In_571);
xor U1346 (N_1346,In_919,In_510);
or U1347 (N_1347,In_214,In_503);
and U1348 (N_1348,In_884,In_464);
nand U1349 (N_1349,In_588,In_323);
nand U1350 (N_1350,In_576,In_596);
xor U1351 (N_1351,In_74,In_965);
nor U1352 (N_1352,In_610,In_379);
nand U1353 (N_1353,In_566,In_456);
nand U1354 (N_1354,In_380,In_439);
or U1355 (N_1355,In_642,In_308);
and U1356 (N_1356,In_404,In_33);
or U1357 (N_1357,In_49,In_592);
or U1358 (N_1358,In_354,In_936);
nor U1359 (N_1359,In_604,In_203);
nand U1360 (N_1360,In_479,In_754);
or U1361 (N_1361,In_326,In_764);
and U1362 (N_1362,In_399,In_603);
and U1363 (N_1363,In_989,In_224);
and U1364 (N_1364,In_118,In_263);
or U1365 (N_1365,In_294,In_864);
and U1366 (N_1366,In_888,In_613);
nor U1367 (N_1367,In_177,In_734);
nand U1368 (N_1368,In_694,In_248);
nor U1369 (N_1369,In_628,In_962);
or U1370 (N_1370,In_614,In_714);
nand U1371 (N_1371,In_609,In_176);
xnor U1372 (N_1372,In_398,In_313);
nand U1373 (N_1373,In_915,In_871);
nor U1374 (N_1374,In_32,In_860);
nor U1375 (N_1375,In_349,In_449);
and U1376 (N_1376,In_723,In_376);
or U1377 (N_1377,In_3,In_434);
or U1378 (N_1378,In_846,In_711);
or U1379 (N_1379,In_327,In_446);
xor U1380 (N_1380,In_971,In_874);
nand U1381 (N_1381,In_548,In_705);
or U1382 (N_1382,In_293,In_677);
or U1383 (N_1383,In_564,In_727);
and U1384 (N_1384,In_743,In_16);
or U1385 (N_1385,In_306,In_951);
and U1386 (N_1386,In_772,In_458);
or U1387 (N_1387,In_107,In_449);
nand U1388 (N_1388,In_263,In_215);
nand U1389 (N_1389,In_856,In_81);
nor U1390 (N_1390,In_289,In_618);
nand U1391 (N_1391,In_116,In_852);
nand U1392 (N_1392,In_733,In_810);
nand U1393 (N_1393,In_447,In_840);
or U1394 (N_1394,In_213,In_608);
nand U1395 (N_1395,In_127,In_650);
and U1396 (N_1396,In_398,In_519);
nor U1397 (N_1397,In_889,In_495);
or U1398 (N_1398,In_288,In_292);
nand U1399 (N_1399,In_908,In_977);
nand U1400 (N_1400,In_101,In_639);
nand U1401 (N_1401,In_804,In_36);
nand U1402 (N_1402,In_559,In_37);
and U1403 (N_1403,In_768,In_569);
nand U1404 (N_1404,In_904,In_97);
or U1405 (N_1405,In_626,In_374);
nand U1406 (N_1406,In_347,In_61);
and U1407 (N_1407,In_46,In_58);
nor U1408 (N_1408,In_12,In_702);
nor U1409 (N_1409,In_782,In_395);
nand U1410 (N_1410,In_865,In_41);
or U1411 (N_1411,In_304,In_151);
nand U1412 (N_1412,In_659,In_514);
or U1413 (N_1413,In_32,In_627);
nand U1414 (N_1414,In_244,In_594);
and U1415 (N_1415,In_604,In_924);
xnor U1416 (N_1416,In_77,In_365);
or U1417 (N_1417,In_727,In_718);
nand U1418 (N_1418,In_768,In_378);
and U1419 (N_1419,In_570,In_169);
or U1420 (N_1420,In_319,In_761);
and U1421 (N_1421,In_803,In_890);
nor U1422 (N_1422,In_378,In_762);
or U1423 (N_1423,In_833,In_558);
nand U1424 (N_1424,In_996,In_779);
nand U1425 (N_1425,In_525,In_951);
xnor U1426 (N_1426,In_81,In_559);
or U1427 (N_1427,In_222,In_118);
and U1428 (N_1428,In_106,In_821);
or U1429 (N_1429,In_206,In_581);
xor U1430 (N_1430,In_814,In_595);
or U1431 (N_1431,In_110,In_835);
nand U1432 (N_1432,In_310,In_782);
nor U1433 (N_1433,In_152,In_375);
or U1434 (N_1434,In_821,In_990);
or U1435 (N_1435,In_379,In_523);
and U1436 (N_1436,In_89,In_381);
nand U1437 (N_1437,In_929,In_764);
xnor U1438 (N_1438,In_277,In_228);
nor U1439 (N_1439,In_144,In_299);
nor U1440 (N_1440,In_634,In_815);
nand U1441 (N_1441,In_437,In_654);
nand U1442 (N_1442,In_144,In_828);
and U1443 (N_1443,In_366,In_353);
nand U1444 (N_1444,In_857,In_241);
nand U1445 (N_1445,In_252,In_555);
nand U1446 (N_1446,In_164,In_486);
or U1447 (N_1447,In_947,In_101);
or U1448 (N_1448,In_835,In_924);
or U1449 (N_1449,In_948,In_530);
nor U1450 (N_1450,In_856,In_157);
nand U1451 (N_1451,In_904,In_579);
or U1452 (N_1452,In_904,In_441);
xnor U1453 (N_1453,In_311,In_1);
nor U1454 (N_1454,In_123,In_325);
or U1455 (N_1455,In_334,In_983);
xor U1456 (N_1456,In_887,In_40);
or U1457 (N_1457,In_141,In_71);
or U1458 (N_1458,In_67,In_909);
nor U1459 (N_1459,In_23,In_470);
nor U1460 (N_1460,In_856,In_20);
nand U1461 (N_1461,In_575,In_118);
nor U1462 (N_1462,In_550,In_365);
nand U1463 (N_1463,In_763,In_534);
nor U1464 (N_1464,In_587,In_351);
nor U1465 (N_1465,In_184,In_759);
nand U1466 (N_1466,In_544,In_586);
nor U1467 (N_1467,In_960,In_955);
nand U1468 (N_1468,In_328,In_860);
or U1469 (N_1469,In_702,In_28);
and U1470 (N_1470,In_755,In_496);
nand U1471 (N_1471,In_423,In_134);
nor U1472 (N_1472,In_853,In_711);
nor U1473 (N_1473,In_272,In_253);
xnor U1474 (N_1474,In_497,In_500);
or U1475 (N_1475,In_87,In_536);
nand U1476 (N_1476,In_397,In_574);
or U1477 (N_1477,In_871,In_668);
nor U1478 (N_1478,In_16,In_249);
nor U1479 (N_1479,In_472,In_743);
nor U1480 (N_1480,In_121,In_222);
and U1481 (N_1481,In_379,In_853);
or U1482 (N_1482,In_15,In_115);
and U1483 (N_1483,In_603,In_965);
xnor U1484 (N_1484,In_251,In_71);
or U1485 (N_1485,In_154,In_432);
and U1486 (N_1486,In_332,In_894);
nor U1487 (N_1487,In_64,In_300);
and U1488 (N_1488,In_671,In_373);
and U1489 (N_1489,In_891,In_926);
and U1490 (N_1490,In_269,In_206);
and U1491 (N_1491,In_894,In_346);
nand U1492 (N_1492,In_442,In_585);
nor U1493 (N_1493,In_821,In_532);
nor U1494 (N_1494,In_77,In_923);
nor U1495 (N_1495,In_465,In_648);
or U1496 (N_1496,In_398,In_908);
nor U1497 (N_1497,In_784,In_320);
xnor U1498 (N_1498,In_944,In_767);
xor U1499 (N_1499,In_869,In_453);
nor U1500 (N_1500,In_377,In_6);
nor U1501 (N_1501,In_754,In_587);
nand U1502 (N_1502,In_229,In_179);
and U1503 (N_1503,In_968,In_350);
nor U1504 (N_1504,In_212,In_983);
nand U1505 (N_1505,In_973,In_137);
nor U1506 (N_1506,In_385,In_798);
nor U1507 (N_1507,In_639,In_235);
and U1508 (N_1508,In_596,In_4);
or U1509 (N_1509,In_927,In_698);
or U1510 (N_1510,In_837,In_30);
and U1511 (N_1511,In_365,In_800);
or U1512 (N_1512,In_136,In_418);
xnor U1513 (N_1513,In_9,In_983);
and U1514 (N_1514,In_944,In_213);
nor U1515 (N_1515,In_168,In_53);
nand U1516 (N_1516,In_320,In_309);
or U1517 (N_1517,In_160,In_316);
or U1518 (N_1518,In_124,In_953);
xor U1519 (N_1519,In_763,In_357);
nand U1520 (N_1520,In_432,In_61);
or U1521 (N_1521,In_841,In_83);
nand U1522 (N_1522,In_372,In_472);
or U1523 (N_1523,In_94,In_717);
or U1524 (N_1524,In_988,In_577);
xor U1525 (N_1525,In_256,In_887);
or U1526 (N_1526,In_909,In_831);
nor U1527 (N_1527,In_63,In_704);
or U1528 (N_1528,In_502,In_414);
or U1529 (N_1529,In_557,In_388);
nand U1530 (N_1530,In_859,In_297);
and U1531 (N_1531,In_58,In_243);
nor U1532 (N_1532,In_538,In_196);
and U1533 (N_1533,In_701,In_696);
and U1534 (N_1534,In_666,In_636);
nor U1535 (N_1535,In_692,In_19);
and U1536 (N_1536,In_340,In_914);
and U1537 (N_1537,In_287,In_148);
nor U1538 (N_1538,In_635,In_291);
nor U1539 (N_1539,In_102,In_366);
xnor U1540 (N_1540,In_574,In_502);
nand U1541 (N_1541,In_498,In_61);
nor U1542 (N_1542,In_289,In_919);
and U1543 (N_1543,In_940,In_126);
and U1544 (N_1544,In_370,In_919);
nor U1545 (N_1545,In_477,In_757);
nor U1546 (N_1546,In_446,In_673);
nor U1547 (N_1547,In_18,In_392);
nor U1548 (N_1548,In_772,In_690);
or U1549 (N_1549,In_699,In_579);
and U1550 (N_1550,In_985,In_104);
or U1551 (N_1551,In_17,In_148);
and U1552 (N_1552,In_25,In_575);
or U1553 (N_1553,In_92,In_226);
or U1554 (N_1554,In_339,In_4);
nor U1555 (N_1555,In_679,In_882);
and U1556 (N_1556,In_800,In_706);
nor U1557 (N_1557,In_910,In_90);
nand U1558 (N_1558,In_392,In_580);
nand U1559 (N_1559,In_794,In_165);
or U1560 (N_1560,In_829,In_837);
nor U1561 (N_1561,In_470,In_61);
nor U1562 (N_1562,In_919,In_444);
nand U1563 (N_1563,In_541,In_58);
nand U1564 (N_1564,In_205,In_433);
or U1565 (N_1565,In_162,In_61);
or U1566 (N_1566,In_727,In_455);
nand U1567 (N_1567,In_137,In_774);
nor U1568 (N_1568,In_574,In_48);
nor U1569 (N_1569,In_423,In_999);
nor U1570 (N_1570,In_512,In_244);
and U1571 (N_1571,In_694,In_340);
and U1572 (N_1572,In_771,In_557);
and U1573 (N_1573,In_770,In_566);
xor U1574 (N_1574,In_575,In_17);
nand U1575 (N_1575,In_469,In_674);
and U1576 (N_1576,In_895,In_876);
xor U1577 (N_1577,In_540,In_83);
xor U1578 (N_1578,In_768,In_225);
nand U1579 (N_1579,In_685,In_736);
and U1580 (N_1580,In_864,In_868);
nor U1581 (N_1581,In_829,In_880);
xnor U1582 (N_1582,In_482,In_407);
or U1583 (N_1583,In_574,In_343);
nor U1584 (N_1584,In_797,In_142);
nor U1585 (N_1585,In_682,In_972);
and U1586 (N_1586,In_948,In_194);
and U1587 (N_1587,In_858,In_696);
nor U1588 (N_1588,In_26,In_623);
and U1589 (N_1589,In_370,In_123);
and U1590 (N_1590,In_397,In_476);
xnor U1591 (N_1591,In_758,In_155);
and U1592 (N_1592,In_400,In_738);
or U1593 (N_1593,In_491,In_663);
nand U1594 (N_1594,In_543,In_754);
nor U1595 (N_1595,In_838,In_785);
nor U1596 (N_1596,In_877,In_151);
nor U1597 (N_1597,In_6,In_757);
nor U1598 (N_1598,In_367,In_343);
or U1599 (N_1599,In_718,In_519);
nor U1600 (N_1600,In_688,In_448);
nand U1601 (N_1601,In_563,In_318);
and U1602 (N_1602,In_390,In_719);
nor U1603 (N_1603,In_89,In_210);
nor U1604 (N_1604,In_390,In_990);
and U1605 (N_1605,In_802,In_537);
xor U1606 (N_1606,In_422,In_115);
nor U1607 (N_1607,In_621,In_922);
nand U1608 (N_1608,In_276,In_639);
nand U1609 (N_1609,In_853,In_190);
nor U1610 (N_1610,In_249,In_858);
nor U1611 (N_1611,In_293,In_814);
and U1612 (N_1612,In_358,In_799);
or U1613 (N_1613,In_719,In_173);
and U1614 (N_1614,In_430,In_437);
nand U1615 (N_1615,In_704,In_160);
nand U1616 (N_1616,In_829,In_332);
or U1617 (N_1617,In_914,In_588);
nand U1618 (N_1618,In_566,In_354);
nor U1619 (N_1619,In_722,In_456);
and U1620 (N_1620,In_18,In_667);
xnor U1621 (N_1621,In_50,In_102);
or U1622 (N_1622,In_206,In_662);
or U1623 (N_1623,In_144,In_327);
and U1624 (N_1624,In_14,In_750);
nor U1625 (N_1625,In_427,In_523);
or U1626 (N_1626,In_307,In_649);
or U1627 (N_1627,In_159,In_149);
nand U1628 (N_1628,In_725,In_994);
nand U1629 (N_1629,In_719,In_336);
and U1630 (N_1630,In_148,In_591);
nor U1631 (N_1631,In_122,In_825);
nor U1632 (N_1632,In_574,In_638);
or U1633 (N_1633,In_71,In_222);
nand U1634 (N_1634,In_752,In_765);
and U1635 (N_1635,In_422,In_804);
nor U1636 (N_1636,In_144,In_40);
nand U1637 (N_1637,In_831,In_485);
and U1638 (N_1638,In_851,In_280);
and U1639 (N_1639,In_43,In_410);
or U1640 (N_1640,In_148,In_422);
nor U1641 (N_1641,In_18,In_42);
xor U1642 (N_1642,In_354,In_857);
nand U1643 (N_1643,In_979,In_108);
and U1644 (N_1644,In_498,In_672);
and U1645 (N_1645,In_953,In_637);
and U1646 (N_1646,In_307,In_340);
xnor U1647 (N_1647,In_322,In_355);
nand U1648 (N_1648,In_984,In_628);
or U1649 (N_1649,In_663,In_617);
nor U1650 (N_1650,In_382,In_429);
xnor U1651 (N_1651,In_750,In_388);
nor U1652 (N_1652,In_835,In_139);
and U1653 (N_1653,In_734,In_124);
nand U1654 (N_1654,In_207,In_618);
nor U1655 (N_1655,In_994,In_387);
or U1656 (N_1656,In_532,In_956);
and U1657 (N_1657,In_134,In_695);
nor U1658 (N_1658,In_690,In_991);
nor U1659 (N_1659,In_929,In_727);
nor U1660 (N_1660,In_322,In_415);
xor U1661 (N_1661,In_375,In_468);
nand U1662 (N_1662,In_708,In_732);
and U1663 (N_1663,In_901,In_766);
and U1664 (N_1664,In_972,In_833);
nor U1665 (N_1665,In_635,In_229);
and U1666 (N_1666,In_100,In_741);
xor U1667 (N_1667,In_419,In_418);
and U1668 (N_1668,In_375,In_44);
and U1669 (N_1669,In_755,In_100);
nand U1670 (N_1670,In_578,In_628);
xor U1671 (N_1671,In_187,In_194);
nand U1672 (N_1672,In_782,In_778);
xor U1673 (N_1673,In_151,In_963);
or U1674 (N_1674,In_722,In_953);
and U1675 (N_1675,In_139,In_599);
or U1676 (N_1676,In_930,In_731);
nor U1677 (N_1677,In_504,In_27);
or U1678 (N_1678,In_72,In_229);
or U1679 (N_1679,In_458,In_310);
and U1680 (N_1680,In_817,In_213);
nand U1681 (N_1681,In_889,In_234);
nor U1682 (N_1682,In_71,In_142);
xnor U1683 (N_1683,In_495,In_247);
nor U1684 (N_1684,In_238,In_400);
nand U1685 (N_1685,In_354,In_316);
or U1686 (N_1686,In_209,In_784);
nor U1687 (N_1687,In_977,In_509);
nand U1688 (N_1688,In_16,In_730);
or U1689 (N_1689,In_528,In_252);
nor U1690 (N_1690,In_785,In_671);
nor U1691 (N_1691,In_124,In_107);
or U1692 (N_1692,In_769,In_775);
nand U1693 (N_1693,In_143,In_287);
or U1694 (N_1694,In_366,In_478);
nor U1695 (N_1695,In_562,In_155);
nor U1696 (N_1696,In_444,In_462);
xor U1697 (N_1697,In_458,In_558);
xor U1698 (N_1698,In_123,In_359);
and U1699 (N_1699,In_502,In_136);
or U1700 (N_1700,In_975,In_522);
or U1701 (N_1701,In_87,In_896);
and U1702 (N_1702,In_9,In_91);
nor U1703 (N_1703,In_634,In_207);
nor U1704 (N_1704,In_736,In_477);
or U1705 (N_1705,In_81,In_60);
and U1706 (N_1706,In_409,In_512);
nand U1707 (N_1707,In_474,In_145);
nand U1708 (N_1708,In_494,In_918);
and U1709 (N_1709,In_797,In_431);
or U1710 (N_1710,In_415,In_237);
nand U1711 (N_1711,In_220,In_970);
or U1712 (N_1712,In_446,In_1);
nand U1713 (N_1713,In_574,In_446);
xor U1714 (N_1714,In_771,In_418);
nand U1715 (N_1715,In_979,In_594);
nor U1716 (N_1716,In_884,In_868);
xnor U1717 (N_1717,In_11,In_322);
nor U1718 (N_1718,In_490,In_313);
nand U1719 (N_1719,In_316,In_667);
or U1720 (N_1720,In_657,In_127);
and U1721 (N_1721,In_906,In_50);
or U1722 (N_1722,In_406,In_719);
xnor U1723 (N_1723,In_89,In_284);
nand U1724 (N_1724,In_790,In_344);
nand U1725 (N_1725,In_976,In_214);
nand U1726 (N_1726,In_912,In_45);
or U1727 (N_1727,In_627,In_892);
and U1728 (N_1728,In_483,In_882);
nor U1729 (N_1729,In_762,In_2);
nand U1730 (N_1730,In_151,In_878);
nor U1731 (N_1731,In_721,In_813);
xnor U1732 (N_1732,In_133,In_913);
or U1733 (N_1733,In_12,In_978);
or U1734 (N_1734,In_642,In_222);
and U1735 (N_1735,In_429,In_570);
nand U1736 (N_1736,In_918,In_610);
nor U1737 (N_1737,In_890,In_624);
nor U1738 (N_1738,In_702,In_998);
xor U1739 (N_1739,In_46,In_336);
nor U1740 (N_1740,In_264,In_809);
and U1741 (N_1741,In_886,In_676);
and U1742 (N_1742,In_171,In_177);
nand U1743 (N_1743,In_848,In_633);
nand U1744 (N_1744,In_458,In_978);
and U1745 (N_1745,In_730,In_142);
xnor U1746 (N_1746,In_752,In_40);
nor U1747 (N_1747,In_335,In_798);
and U1748 (N_1748,In_975,In_595);
and U1749 (N_1749,In_927,In_529);
xnor U1750 (N_1750,In_810,In_447);
and U1751 (N_1751,In_638,In_530);
or U1752 (N_1752,In_808,In_76);
nand U1753 (N_1753,In_484,In_783);
or U1754 (N_1754,In_188,In_278);
xnor U1755 (N_1755,In_716,In_190);
xor U1756 (N_1756,In_938,In_153);
or U1757 (N_1757,In_571,In_275);
nor U1758 (N_1758,In_453,In_370);
or U1759 (N_1759,In_892,In_736);
nor U1760 (N_1760,In_720,In_268);
nand U1761 (N_1761,In_298,In_213);
xor U1762 (N_1762,In_496,In_910);
xor U1763 (N_1763,In_764,In_930);
xnor U1764 (N_1764,In_773,In_400);
and U1765 (N_1765,In_700,In_207);
xnor U1766 (N_1766,In_706,In_700);
or U1767 (N_1767,In_958,In_778);
or U1768 (N_1768,In_395,In_420);
or U1769 (N_1769,In_202,In_765);
and U1770 (N_1770,In_337,In_605);
or U1771 (N_1771,In_724,In_102);
nand U1772 (N_1772,In_569,In_108);
or U1773 (N_1773,In_609,In_435);
or U1774 (N_1774,In_594,In_639);
or U1775 (N_1775,In_845,In_758);
nand U1776 (N_1776,In_603,In_373);
or U1777 (N_1777,In_291,In_590);
or U1778 (N_1778,In_713,In_984);
nor U1779 (N_1779,In_977,In_852);
xor U1780 (N_1780,In_243,In_235);
or U1781 (N_1781,In_748,In_372);
and U1782 (N_1782,In_346,In_973);
and U1783 (N_1783,In_343,In_940);
or U1784 (N_1784,In_297,In_998);
and U1785 (N_1785,In_614,In_276);
or U1786 (N_1786,In_465,In_135);
nand U1787 (N_1787,In_115,In_719);
nand U1788 (N_1788,In_367,In_271);
or U1789 (N_1789,In_582,In_829);
xnor U1790 (N_1790,In_434,In_473);
and U1791 (N_1791,In_275,In_890);
and U1792 (N_1792,In_166,In_287);
nand U1793 (N_1793,In_1,In_857);
nand U1794 (N_1794,In_866,In_213);
and U1795 (N_1795,In_723,In_922);
or U1796 (N_1796,In_225,In_394);
nand U1797 (N_1797,In_992,In_473);
or U1798 (N_1798,In_821,In_772);
and U1799 (N_1799,In_915,In_948);
nor U1800 (N_1800,In_626,In_582);
and U1801 (N_1801,In_492,In_773);
nand U1802 (N_1802,In_217,In_307);
or U1803 (N_1803,In_306,In_114);
and U1804 (N_1804,In_534,In_743);
and U1805 (N_1805,In_6,In_379);
nor U1806 (N_1806,In_21,In_69);
or U1807 (N_1807,In_491,In_920);
or U1808 (N_1808,In_353,In_999);
or U1809 (N_1809,In_435,In_822);
nor U1810 (N_1810,In_996,In_507);
and U1811 (N_1811,In_191,In_523);
or U1812 (N_1812,In_103,In_500);
nor U1813 (N_1813,In_662,In_635);
nand U1814 (N_1814,In_881,In_361);
nand U1815 (N_1815,In_267,In_758);
or U1816 (N_1816,In_220,In_876);
xnor U1817 (N_1817,In_443,In_355);
nor U1818 (N_1818,In_179,In_27);
nor U1819 (N_1819,In_395,In_618);
and U1820 (N_1820,In_54,In_693);
and U1821 (N_1821,In_660,In_828);
nand U1822 (N_1822,In_886,In_154);
and U1823 (N_1823,In_636,In_426);
nor U1824 (N_1824,In_13,In_589);
or U1825 (N_1825,In_662,In_875);
nand U1826 (N_1826,In_819,In_145);
nor U1827 (N_1827,In_578,In_305);
nor U1828 (N_1828,In_914,In_114);
and U1829 (N_1829,In_619,In_378);
nand U1830 (N_1830,In_530,In_45);
nor U1831 (N_1831,In_594,In_800);
xnor U1832 (N_1832,In_612,In_768);
and U1833 (N_1833,In_817,In_31);
nor U1834 (N_1834,In_333,In_821);
or U1835 (N_1835,In_63,In_285);
or U1836 (N_1836,In_847,In_73);
nor U1837 (N_1837,In_388,In_443);
and U1838 (N_1838,In_246,In_38);
and U1839 (N_1839,In_337,In_705);
nor U1840 (N_1840,In_412,In_168);
and U1841 (N_1841,In_505,In_951);
and U1842 (N_1842,In_377,In_611);
nand U1843 (N_1843,In_398,In_181);
or U1844 (N_1844,In_987,In_233);
and U1845 (N_1845,In_165,In_196);
nor U1846 (N_1846,In_825,In_995);
and U1847 (N_1847,In_370,In_823);
nor U1848 (N_1848,In_14,In_372);
or U1849 (N_1849,In_42,In_396);
xor U1850 (N_1850,In_473,In_190);
nand U1851 (N_1851,In_801,In_78);
and U1852 (N_1852,In_650,In_101);
nand U1853 (N_1853,In_596,In_34);
nand U1854 (N_1854,In_987,In_194);
nand U1855 (N_1855,In_653,In_206);
nand U1856 (N_1856,In_365,In_761);
and U1857 (N_1857,In_857,In_928);
or U1858 (N_1858,In_904,In_9);
and U1859 (N_1859,In_908,In_976);
nand U1860 (N_1860,In_236,In_7);
and U1861 (N_1861,In_527,In_740);
nand U1862 (N_1862,In_468,In_982);
and U1863 (N_1863,In_105,In_444);
nor U1864 (N_1864,In_968,In_481);
and U1865 (N_1865,In_195,In_737);
xor U1866 (N_1866,In_462,In_530);
nor U1867 (N_1867,In_24,In_788);
and U1868 (N_1868,In_364,In_600);
nor U1869 (N_1869,In_794,In_452);
or U1870 (N_1870,In_475,In_914);
and U1871 (N_1871,In_725,In_133);
and U1872 (N_1872,In_579,In_135);
nand U1873 (N_1873,In_38,In_942);
or U1874 (N_1874,In_461,In_917);
nor U1875 (N_1875,In_600,In_951);
nor U1876 (N_1876,In_985,In_630);
nand U1877 (N_1877,In_386,In_379);
nand U1878 (N_1878,In_282,In_512);
or U1879 (N_1879,In_644,In_565);
xnor U1880 (N_1880,In_945,In_885);
xor U1881 (N_1881,In_331,In_141);
nor U1882 (N_1882,In_873,In_547);
or U1883 (N_1883,In_578,In_323);
and U1884 (N_1884,In_238,In_780);
nand U1885 (N_1885,In_735,In_913);
nand U1886 (N_1886,In_690,In_519);
nor U1887 (N_1887,In_272,In_441);
nand U1888 (N_1888,In_681,In_713);
nor U1889 (N_1889,In_900,In_500);
and U1890 (N_1890,In_493,In_996);
nor U1891 (N_1891,In_738,In_417);
and U1892 (N_1892,In_757,In_692);
nor U1893 (N_1893,In_694,In_618);
nor U1894 (N_1894,In_4,In_7);
and U1895 (N_1895,In_329,In_88);
and U1896 (N_1896,In_412,In_376);
and U1897 (N_1897,In_676,In_416);
nand U1898 (N_1898,In_431,In_589);
or U1899 (N_1899,In_975,In_278);
or U1900 (N_1900,In_783,In_656);
nor U1901 (N_1901,In_360,In_317);
nand U1902 (N_1902,In_798,In_673);
or U1903 (N_1903,In_281,In_135);
nand U1904 (N_1904,In_69,In_0);
xnor U1905 (N_1905,In_509,In_541);
xor U1906 (N_1906,In_338,In_352);
and U1907 (N_1907,In_235,In_668);
nor U1908 (N_1908,In_189,In_615);
nor U1909 (N_1909,In_642,In_67);
nor U1910 (N_1910,In_718,In_984);
or U1911 (N_1911,In_464,In_712);
xor U1912 (N_1912,In_957,In_384);
or U1913 (N_1913,In_944,In_246);
and U1914 (N_1914,In_195,In_430);
nand U1915 (N_1915,In_189,In_983);
nor U1916 (N_1916,In_231,In_30);
nor U1917 (N_1917,In_416,In_487);
nand U1918 (N_1918,In_125,In_807);
and U1919 (N_1919,In_109,In_87);
nor U1920 (N_1920,In_822,In_715);
or U1921 (N_1921,In_955,In_525);
nor U1922 (N_1922,In_644,In_682);
and U1923 (N_1923,In_417,In_246);
nand U1924 (N_1924,In_851,In_793);
xor U1925 (N_1925,In_69,In_317);
nand U1926 (N_1926,In_77,In_951);
and U1927 (N_1927,In_347,In_230);
nand U1928 (N_1928,In_669,In_320);
or U1929 (N_1929,In_980,In_371);
nand U1930 (N_1930,In_722,In_878);
xor U1931 (N_1931,In_693,In_115);
nand U1932 (N_1932,In_334,In_3);
nand U1933 (N_1933,In_981,In_197);
or U1934 (N_1934,In_897,In_343);
and U1935 (N_1935,In_357,In_200);
and U1936 (N_1936,In_160,In_561);
and U1937 (N_1937,In_446,In_731);
nand U1938 (N_1938,In_493,In_3);
nand U1939 (N_1939,In_627,In_46);
and U1940 (N_1940,In_646,In_554);
and U1941 (N_1941,In_544,In_315);
nor U1942 (N_1942,In_388,In_768);
xnor U1943 (N_1943,In_381,In_187);
xor U1944 (N_1944,In_421,In_218);
nor U1945 (N_1945,In_695,In_657);
or U1946 (N_1946,In_350,In_578);
nand U1947 (N_1947,In_97,In_893);
nor U1948 (N_1948,In_577,In_247);
xnor U1949 (N_1949,In_232,In_29);
or U1950 (N_1950,In_129,In_947);
and U1951 (N_1951,In_502,In_512);
nor U1952 (N_1952,In_855,In_927);
or U1953 (N_1953,In_773,In_379);
nand U1954 (N_1954,In_230,In_55);
and U1955 (N_1955,In_681,In_123);
xnor U1956 (N_1956,In_858,In_770);
nand U1957 (N_1957,In_3,In_219);
and U1958 (N_1958,In_352,In_642);
nand U1959 (N_1959,In_16,In_170);
or U1960 (N_1960,In_623,In_936);
nor U1961 (N_1961,In_588,In_675);
nand U1962 (N_1962,In_175,In_596);
nand U1963 (N_1963,In_547,In_118);
xnor U1964 (N_1964,In_28,In_320);
nor U1965 (N_1965,In_438,In_905);
and U1966 (N_1966,In_531,In_680);
nand U1967 (N_1967,In_865,In_298);
or U1968 (N_1968,In_723,In_456);
nand U1969 (N_1969,In_720,In_342);
and U1970 (N_1970,In_286,In_693);
nand U1971 (N_1971,In_239,In_727);
and U1972 (N_1972,In_838,In_892);
nand U1973 (N_1973,In_307,In_838);
nor U1974 (N_1974,In_990,In_603);
nor U1975 (N_1975,In_321,In_756);
and U1976 (N_1976,In_910,In_702);
nor U1977 (N_1977,In_550,In_813);
or U1978 (N_1978,In_820,In_142);
nand U1979 (N_1979,In_362,In_394);
and U1980 (N_1980,In_10,In_861);
nor U1981 (N_1981,In_798,In_54);
nor U1982 (N_1982,In_547,In_121);
nor U1983 (N_1983,In_425,In_186);
nand U1984 (N_1984,In_197,In_61);
nand U1985 (N_1985,In_529,In_231);
and U1986 (N_1986,In_408,In_225);
xnor U1987 (N_1987,In_131,In_928);
and U1988 (N_1988,In_787,In_482);
nor U1989 (N_1989,In_206,In_684);
and U1990 (N_1990,In_45,In_625);
nand U1991 (N_1991,In_215,In_212);
or U1992 (N_1992,In_162,In_638);
nand U1993 (N_1993,In_345,In_100);
nand U1994 (N_1994,In_439,In_879);
or U1995 (N_1995,In_384,In_879);
and U1996 (N_1996,In_120,In_906);
or U1997 (N_1997,In_244,In_353);
nor U1998 (N_1998,In_89,In_863);
and U1999 (N_1999,In_106,In_530);
or U2000 (N_2000,N_1713,N_1504);
and U2001 (N_2001,N_827,N_1279);
and U2002 (N_2002,N_1829,N_689);
or U2003 (N_2003,N_243,N_106);
and U2004 (N_2004,N_1082,N_622);
nor U2005 (N_2005,N_1882,N_438);
xor U2006 (N_2006,N_444,N_339);
nor U2007 (N_2007,N_298,N_529);
xnor U2008 (N_2008,N_1622,N_601);
nand U2009 (N_2009,N_749,N_98);
and U2010 (N_2010,N_960,N_1406);
and U2011 (N_2011,N_489,N_319);
nand U2012 (N_2012,N_1246,N_1844);
nor U2013 (N_2013,N_1086,N_901);
nor U2014 (N_2014,N_338,N_214);
nor U2015 (N_2015,N_1800,N_1206);
and U2016 (N_2016,N_1,N_647);
or U2017 (N_2017,N_1377,N_379);
nor U2018 (N_2018,N_442,N_40);
and U2019 (N_2019,N_1820,N_1684);
nor U2020 (N_2020,N_1876,N_684);
xor U2021 (N_2021,N_1105,N_371);
or U2022 (N_2022,N_1679,N_457);
nand U2023 (N_2023,N_1245,N_724);
xor U2024 (N_2024,N_383,N_1848);
or U2025 (N_2025,N_65,N_1013);
nor U2026 (N_2026,N_971,N_1049);
nand U2027 (N_2027,N_1831,N_552);
or U2028 (N_2028,N_172,N_1262);
xor U2029 (N_2029,N_1032,N_779);
nor U2030 (N_2030,N_540,N_992);
nand U2031 (N_2031,N_1296,N_546);
nand U2032 (N_2032,N_735,N_13);
nor U2033 (N_2033,N_1811,N_197);
or U2034 (N_2034,N_1554,N_490);
nor U2035 (N_2035,N_1107,N_357);
nor U2036 (N_2036,N_195,N_1425);
or U2037 (N_2037,N_1147,N_1538);
or U2038 (N_2038,N_634,N_664);
nand U2039 (N_2039,N_328,N_1637);
and U2040 (N_2040,N_1416,N_1052);
xor U2041 (N_2041,N_1773,N_691);
and U2042 (N_2042,N_80,N_1438);
and U2043 (N_2043,N_1790,N_556);
and U2044 (N_2044,N_361,N_880);
and U2045 (N_2045,N_1115,N_750);
and U2046 (N_2046,N_1039,N_574);
or U2047 (N_2047,N_1874,N_1353);
xnor U2048 (N_2048,N_22,N_103);
nand U2049 (N_2049,N_1348,N_238);
or U2050 (N_2050,N_612,N_538);
nor U2051 (N_2051,N_717,N_991);
and U2052 (N_2052,N_1969,N_1217);
and U2053 (N_2053,N_1960,N_1824);
and U2054 (N_2054,N_1682,N_1788);
nor U2055 (N_2055,N_1362,N_1744);
nand U2056 (N_2056,N_1900,N_839);
nand U2057 (N_2057,N_842,N_1833);
and U2058 (N_2058,N_900,N_948);
and U2059 (N_2059,N_1952,N_87);
nand U2060 (N_2060,N_993,N_626);
nor U2061 (N_2061,N_1826,N_168);
nor U2062 (N_2062,N_795,N_1500);
and U2063 (N_2063,N_1026,N_1321);
nor U2064 (N_2064,N_882,N_1255);
nand U2065 (N_2065,N_26,N_32);
nor U2066 (N_2066,N_644,N_787);
nand U2067 (N_2067,N_281,N_973);
or U2068 (N_2068,N_49,N_280);
or U2069 (N_2069,N_1204,N_136);
nor U2070 (N_2070,N_317,N_216);
or U2071 (N_2071,N_1989,N_1997);
xor U2072 (N_2072,N_11,N_362);
nand U2073 (N_2073,N_1358,N_142);
and U2074 (N_2074,N_1176,N_236);
nor U2075 (N_2075,N_1926,N_380);
and U2076 (N_2076,N_1391,N_47);
nor U2077 (N_2077,N_1257,N_1949);
or U2078 (N_2078,N_957,N_50);
or U2079 (N_2079,N_259,N_1536);
or U2080 (N_2080,N_1539,N_1595);
nand U2081 (N_2081,N_1529,N_311);
or U2082 (N_2082,N_858,N_92);
or U2083 (N_2083,N_1813,N_1040);
and U2084 (N_2084,N_1808,N_744);
nand U2085 (N_2085,N_819,N_600);
nand U2086 (N_2086,N_997,N_781);
nor U2087 (N_2087,N_1047,N_832);
nand U2088 (N_2088,N_1227,N_1398);
nor U2089 (N_2089,N_1108,N_1664);
nand U2090 (N_2090,N_531,N_1226);
nand U2091 (N_2091,N_1635,N_1301);
nor U2092 (N_2092,N_113,N_389);
xnor U2093 (N_2093,N_462,N_1063);
nor U2094 (N_2094,N_1494,N_1476);
and U2095 (N_2095,N_1940,N_1372);
or U2096 (N_2096,N_1755,N_336);
or U2097 (N_2097,N_1902,N_310);
nand U2098 (N_2098,N_1386,N_1668);
and U2099 (N_2099,N_85,N_1719);
or U2100 (N_2100,N_599,N_1266);
and U2101 (N_2101,N_866,N_474);
and U2102 (N_2102,N_1916,N_1838);
xor U2103 (N_2103,N_613,N_1235);
nor U2104 (N_2104,N_1832,N_188);
and U2105 (N_2105,N_479,N_1191);
nand U2106 (N_2106,N_385,N_1944);
nor U2107 (N_2107,N_30,N_590);
and U2108 (N_2108,N_814,N_1648);
nand U2109 (N_2109,N_1390,N_390);
nor U2110 (N_2110,N_1317,N_895);
or U2111 (N_2111,N_554,N_1341);
and U2112 (N_2112,N_321,N_520);
xnor U2113 (N_2113,N_1122,N_1613);
xor U2114 (N_2114,N_1547,N_1769);
and U2115 (N_2115,N_1067,N_1927);
nor U2116 (N_2116,N_1911,N_181);
or U2117 (N_2117,N_915,N_1712);
and U2118 (N_2118,N_1413,N_1694);
nor U2119 (N_2119,N_308,N_1139);
or U2120 (N_2120,N_1966,N_756);
or U2121 (N_2121,N_294,N_1670);
or U2122 (N_2122,N_187,N_1929);
nand U2123 (N_2123,N_1971,N_471);
and U2124 (N_2124,N_192,N_1625);
and U2125 (N_2125,N_1205,N_1777);
nand U2126 (N_2126,N_482,N_1253);
and U2127 (N_2127,N_983,N_721);
or U2128 (N_2128,N_715,N_1477);
and U2129 (N_2129,N_1920,N_1064);
or U2130 (N_2130,N_1646,N_1890);
nor U2131 (N_2131,N_1609,N_1304);
nand U2132 (N_2132,N_1465,N_667);
or U2133 (N_2133,N_1580,N_630);
xnor U2134 (N_2134,N_1877,N_517);
nand U2135 (N_2135,N_1794,N_1376);
or U2136 (N_2136,N_653,N_513);
nor U2137 (N_2137,N_1387,N_1905);
or U2138 (N_2138,N_1671,N_898);
xnor U2139 (N_2139,N_674,N_844);
nand U2140 (N_2140,N_229,N_1633);
xnor U2141 (N_2141,N_67,N_293);
or U2142 (N_2142,N_1522,N_1355);
nor U2143 (N_2143,N_1350,N_1138);
or U2144 (N_2144,N_343,N_1014);
or U2145 (N_2145,N_1160,N_1976);
nor U2146 (N_2146,N_285,N_36);
nand U2147 (N_2147,N_1731,N_60);
or U2148 (N_2148,N_949,N_1910);
xnor U2149 (N_2149,N_1612,N_1443);
or U2150 (N_2150,N_0,N_473);
or U2151 (N_2151,N_1149,N_758);
nor U2152 (N_2152,N_1497,N_864);
or U2153 (N_2153,N_1843,N_890);
and U2154 (N_2154,N_1142,N_1543);
nand U2155 (N_2155,N_1202,N_421);
nor U2156 (N_2156,N_1421,N_1903);
or U2157 (N_2157,N_1154,N_1324);
xor U2158 (N_2158,N_1623,N_495);
and U2159 (N_2159,N_189,N_359);
xor U2160 (N_2160,N_1468,N_486);
nor U2161 (N_2161,N_1825,N_1922);
nand U2162 (N_2162,N_853,N_1275);
or U2163 (N_2163,N_884,N_675);
and U2164 (N_2164,N_1061,N_706);
nor U2165 (N_2165,N_584,N_1992);
xor U2166 (N_2166,N_1724,N_369);
or U2167 (N_2167,N_1875,N_1434);
or U2168 (N_2168,N_1248,N_1865);
nand U2169 (N_2169,N_276,N_961);
and U2170 (N_2170,N_1325,N_428);
nand U2171 (N_2171,N_1918,N_1948);
and U2172 (N_2172,N_8,N_146);
nor U2173 (N_2173,N_1837,N_782);
nor U2174 (N_2174,N_1774,N_697);
or U2175 (N_2175,N_1519,N_1126);
or U2176 (N_2176,N_157,N_1467);
xnor U2177 (N_2177,N_131,N_1162);
xnor U2178 (N_2178,N_1159,N_1548);
nor U2179 (N_2179,N_1290,N_345);
or U2180 (N_2180,N_166,N_1370);
nand U2181 (N_2181,N_857,N_397);
nor U2182 (N_2182,N_1357,N_151);
xor U2183 (N_2183,N_23,N_760);
or U2184 (N_2184,N_335,N_1688);
or U2185 (N_2185,N_1658,N_1365);
nor U2186 (N_2186,N_593,N_1056);
nand U2187 (N_2187,N_247,N_176);
or U2188 (N_2188,N_788,N_1183);
nand U2189 (N_2189,N_594,N_564);
nand U2190 (N_2190,N_855,N_1037);
nand U2191 (N_2191,N_1925,N_1216);
nor U2192 (N_2192,N_1165,N_1931);
nor U2193 (N_2193,N_841,N_1342);
or U2194 (N_2194,N_823,N_1509);
and U2195 (N_2195,N_954,N_456);
xor U2196 (N_2196,N_963,N_776);
or U2197 (N_2197,N_1456,N_826);
and U2198 (N_2198,N_804,N_1155);
nand U2199 (N_2199,N_1270,N_76);
xnor U2200 (N_2200,N_499,N_1512);
and U2201 (N_2201,N_1496,N_1428);
and U2202 (N_2202,N_1379,N_1146);
or U2203 (N_2203,N_685,N_21);
xnor U2204 (N_2204,N_731,N_1964);
nor U2205 (N_2205,N_532,N_1051);
nand U2206 (N_2206,N_1222,N_1295);
nand U2207 (N_2207,N_303,N_1400);
nand U2208 (N_2208,N_1551,N_1999);
nand U2209 (N_2209,N_666,N_1515);
or U2210 (N_2210,N_1733,N_548);
nor U2211 (N_2211,N_116,N_1187);
or U2212 (N_2212,N_1531,N_962);
nor U2213 (N_2213,N_1896,N_173);
or U2214 (N_2214,N_1153,N_1054);
nand U2215 (N_2215,N_1401,N_559);
or U2216 (N_2216,N_1656,N_929);
nand U2217 (N_2217,N_77,N_676);
and U2218 (N_2218,N_1285,N_465);
and U2219 (N_2219,N_1289,N_54);
and U2220 (N_2220,N_1395,N_563);
nand U2221 (N_2221,N_791,N_1532);
nor U2222 (N_2222,N_1935,N_1835);
nand U2223 (N_2223,N_1396,N_1088);
xor U2224 (N_2224,N_182,N_652);
and U2225 (N_2225,N_1269,N_299);
nor U2226 (N_2226,N_1722,N_344);
and U2227 (N_2227,N_1647,N_1236);
nand U2228 (N_2228,N_346,N_854);
nand U2229 (N_2229,N_598,N_154);
and U2230 (N_2230,N_266,N_933);
nand U2231 (N_2231,N_38,N_39);
and U2232 (N_2232,N_196,N_1294);
nand U2233 (N_2233,N_29,N_978);
nor U2234 (N_2234,N_153,N_932);
or U2235 (N_2235,N_1585,N_950);
nand U2236 (N_2236,N_1281,N_719);
xnor U2237 (N_2237,N_683,N_1354);
and U2238 (N_2238,N_1287,N_1839);
nor U2239 (N_2239,N_1576,N_1019);
and U2240 (N_2240,N_774,N_1924);
and U2241 (N_2241,N_789,N_1140);
xnor U2242 (N_2242,N_1091,N_887);
or U2243 (N_2243,N_292,N_497);
or U2244 (N_2244,N_99,N_631);
and U2245 (N_2245,N_1450,N_922);
nor U2246 (N_2246,N_734,N_277);
or U2247 (N_2247,N_1797,N_1862);
and U2248 (N_2248,N_1177,N_119);
nor U2249 (N_2249,N_1901,N_752);
nand U2250 (N_2250,N_665,N_1074);
xor U2251 (N_2251,N_1592,N_1097);
nor U2252 (N_2252,N_230,N_1821);
nand U2253 (N_2253,N_466,N_1846);
nor U2254 (N_2254,N_935,N_73);
xnor U2255 (N_2255,N_1895,N_184);
nor U2256 (N_2256,N_432,N_1461);
or U2257 (N_2257,N_728,N_242);
nor U2258 (N_2258,N_940,N_1619);
nor U2259 (N_2259,N_422,N_1475);
and U2260 (N_2260,N_149,N_1845);
nor U2261 (N_2261,N_1933,N_1489);
and U2262 (N_2262,N_278,N_1527);
and U2263 (N_2263,N_1566,N_1863);
xnor U2264 (N_2264,N_1402,N_365);
xor U2265 (N_2265,N_477,N_1076);
xnor U2266 (N_2266,N_1417,N_312);
and U2267 (N_2267,N_1158,N_318);
or U2268 (N_2268,N_1906,N_4);
nor U2269 (N_2269,N_250,N_1690);
xnor U2270 (N_2270,N_565,N_470);
or U2271 (N_2271,N_817,N_919);
and U2272 (N_2272,N_904,N_530);
and U2273 (N_2273,N_833,N_831);
and U2274 (N_2274,N_1508,N_1442);
nand U2275 (N_2275,N_307,N_1705);
and U2276 (N_2276,N_183,N_282);
nand U2277 (N_2277,N_633,N_1388);
or U2278 (N_2278,N_628,N_623);
nor U2279 (N_2279,N_1089,N_9);
nor U2280 (N_2280,N_1469,N_28);
nor U2281 (N_2281,N_1320,N_219);
nand U2282 (N_2282,N_1597,N_353);
and U2283 (N_2283,N_768,N_999);
or U2284 (N_2284,N_1666,N_1312);
nand U2285 (N_2285,N_1203,N_1283);
and U2286 (N_2286,N_1150,N_1079);
or U2287 (N_2287,N_51,N_1984);
nor U2288 (N_2288,N_1336,N_1516);
nand U2289 (N_2289,N_109,N_191);
nand U2290 (N_2290,N_1137,N_803);
nor U2291 (N_2291,N_1830,N_1384);
and U2292 (N_2292,N_410,N_1492);
nand U2293 (N_2293,N_257,N_1611);
nand U2294 (N_2294,N_287,N_1621);
nand U2295 (N_2295,N_1759,N_1535);
nor U2296 (N_2296,N_402,N_970);
nand U2297 (N_2297,N_1698,N_1540);
nand U2298 (N_2298,N_398,N_1654);
and U2299 (N_2299,N_678,N_1747);
or U2300 (N_2300,N_1963,N_1899);
or U2301 (N_2301,N_97,N_1286);
nand U2302 (N_2302,N_780,N_239);
nor U2303 (N_2303,N_1786,N_20);
nand U2304 (N_2304,N_133,N_1783);
and U2305 (N_2305,N_1776,N_96);
nor U2306 (N_2306,N_582,N_431);
nor U2307 (N_2307,N_1271,N_821);
nand U2308 (N_2308,N_766,N_1048);
nor U2309 (N_2309,N_1373,N_1375);
nand U2310 (N_2310,N_834,N_771);
nor U2311 (N_2311,N_1965,N_1866);
nor U2312 (N_2312,N_1602,N_1528);
nor U2313 (N_2313,N_1907,N_792);
or U2314 (N_2314,N_6,N_1228);
nor U2315 (N_2315,N_1163,N_974);
nor U2316 (N_2316,N_323,N_1382);
nand U2317 (N_2317,N_512,N_1130);
xor U2318 (N_2318,N_1513,N_914);
nor U2319 (N_2319,N_1432,N_1795);
and U2320 (N_2320,N_611,N_1859);
and U2321 (N_2321,N_562,N_148);
nor U2322 (N_2322,N_943,N_128);
or U2323 (N_2323,N_897,N_972);
and U2324 (N_2324,N_1912,N_1559);
or U2325 (N_2325,N_1305,N_454);
or U2326 (N_2326,N_135,N_1209);
nand U2327 (N_2327,N_1335,N_55);
nor U2328 (N_2328,N_1756,N_1366);
xor U2329 (N_2329,N_1463,N_129);
and U2330 (N_2330,N_170,N_604);
and U2331 (N_2331,N_372,N_1403);
or U2332 (N_2332,N_205,N_1575);
and U2333 (N_2333,N_1171,N_227);
nor U2334 (N_2334,N_291,N_426);
nor U2335 (N_2335,N_485,N_688);
and U2336 (N_2336,N_235,N_883);
and U2337 (N_2337,N_1001,N_1181);
and U2338 (N_2338,N_1590,N_56);
and U2339 (N_2339,N_1752,N_1853);
and U2340 (N_2340,N_423,N_1282);
nor U2341 (N_2341,N_1814,N_1237);
nor U2342 (N_2342,N_1740,N_93);
nor U2343 (N_2343,N_1292,N_968);
nand U2344 (N_2344,N_829,N_34);
nand U2345 (N_2345,N_1143,N_1243);
and U2346 (N_2346,N_1251,N_1729);
nor U2347 (N_2347,N_1414,N_1716);
and U2348 (N_2348,N_414,N_1995);
xnor U2349 (N_2349,N_207,N_1121);
nor U2350 (N_2350,N_1980,N_325);
and U2351 (N_2351,N_1632,N_1184);
nor U2352 (N_2352,N_411,N_94);
xnor U2353 (N_2353,N_1600,N_1210);
or U2354 (N_2354,N_386,N_288);
and U2355 (N_2355,N_902,N_406);
or U2356 (N_2356,N_1749,N_487);
or U2357 (N_2357,N_702,N_670);
and U2358 (N_2358,N_1042,N_1423);
or U2359 (N_2359,N_1479,N_1120);
nand U2360 (N_2360,N_1193,N_468);
and U2361 (N_2361,N_270,N_262);
and U2362 (N_2362,N_429,N_916);
and U2363 (N_2363,N_1148,N_873);
or U2364 (N_2364,N_677,N_1787);
and U2365 (N_2365,N_987,N_1474);
or U2366 (N_2366,N_1264,N_300);
or U2367 (N_2367,N_1033,N_545);
nand U2368 (N_2368,N_1858,N_742);
nand U2369 (N_2369,N_1340,N_164);
nand U2370 (N_2370,N_705,N_316);
nor U2371 (N_2371,N_1558,N_18);
nand U2372 (N_2372,N_1693,N_891);
nand U2373 (N_2373,N_502,N_1060);
or U2374 (N_2374,N_927,N_413);
xnor U2375 (N_2375,N_1480,N_1706);
nor U2376 (N_2376,N_1062,N_1691);
nand U2377 (N_2377,N_1288,N_1016);
and U2378 (N_2378,N_1537,N_1923);
or U2379 (N_2379,N_867,N_1069);
and U2380 (N_2380,N_1584,N_437);
nor U2381 (N_2381,N_1485,N_1420);
or U2382 (N_2382,N_1802,N_695);
nor U2383 (N_2383,N_476,N_1318);
and U2384 (N_2384,N_865,N_1332);
and U2385 (N_2385,N_1472,N_1238);
nor U2386 (N_2386,N_784,N_522);
nand U2387 (N_2387,N_1892,N_521);
nor U2388 (N_2388,N_1887,N_1211);
xnor U2389 (N_2389,N_859,N_1109);
nand U2390 (N_2390,N_366,N_580);
or U2391 (N_2391,N_1125,N_1990);
nor U2392 (N_2392,N_1102,N_1798);
and U2393 (N_2393,N_730,N_107);
nor U2394 (N_2394,N_260,N_447);
nand U2395 (N_2395,N_1113,N_1715);
and U2396 (N_2396,N_1669,N_272);
nor U2397 (N_2397,N_591,N_820);
or U2398 (N_2398,N_1847,N_1252);
or U2399 (N_2399,N_740,N_986);
or U2400 (N_2400,N_669,N_1856);
and U2401 (N_2401,N_483,N_926);
and U2402 (N_2402,N_578,N_917);
or U2403 (N_2403,N_171,N_57);
nor U2404 (N_2404,N_1702,N_152);
or U2405 (N_2405,N_863,N_1819);
nor U2406 (N_2406,N_395,N_799);
and U2407 (N_2407,N_1928,N_741);
xor U2408 (N_2408,N_1128,N_1307);
and U2409 (N_2409,N_1780,N_313);
xnor U2410 (N_2410,N_906,N_1779);
nand U2411 (N_2411,N_1807,N_1179);
and U2412 (N_2412,N_1058,N_1589);
nand U2413 (N_2413,N_672,N_718);
nor U2414 (N_2414,N_605,N_409);
or U2415 (N_2415,N_387,N_165);
nand U2416 (N_2416,N_1725,N_211);
or U2417 (N_2417,N_969,N_1166);
nand U2418 (N_2418,N_1711,N_1028);
nor U2419 (N_2419,N_137,N_608);
or U2420 (N_2420,N_232,N_838);
nand U2421 (N_2421,N_1586,N_656);
and U2422 (N_2422,N_707,N_1570);
or U2423 (N_2423,N_416,N_1483);
or U2424 (N_2424,N_894,N_114);
xor U2425 (N_2425,N_1359,N_64);
and U2426 (N_2426,N_1758,N_1015);
and U2427 (N_2427,N_1653,N_461);
and U2428 (N_2428,N_244,N_1630);
and U2429 (N_2429,N_169,N_1327);
nand U2430 (N_2430,N_813,N_896);
nand U2431 (N_2431,N_903,N_1517);
nand U2432 (N_2432,N_1643,N_1329);
nor U2433 (N_2433,N_384,N_1598);
or U2434 (N_2434,N_751,N_786);
and U2435 (N_2435,N_733,N_271);
nand U2436 (N_2436,N_710,N_433);
nand U2437 (N_2437,N_44,N_246);
nand U2438 (N_2438,N_1974,N_1549);
or U2439 (N_2439,N_279,N_1970);
and U2440 (N_2440,N_1736,N_263);
and U2441 (N_2441,N_1449,N_1717);
xnor U2442 (N_2442,N_446,N_206);
nor U2443 (N_2443,N_1784,N_1453);
or U2444 (N_2444,N_654,N_1884);
and U2445 (N_2445,N_1618,N_1010);
or U2446 (N_2446,N_441,N_1778);
nor U2447 (N_2447,N_807,N_1718);
or U2448 (N_2448,N_1129,N_1898);
xnor U2449 (N_2449,N_571,N_856);
nor U2450 (N_2450,N_660,N_7);
nor U2451 (N_2451,N_645,N_746);
nor U2452 (N_2452,N_158,N_908);
xor U2453 (N_2453,N_31,N_905);
nand U2454 (N_2454,N_1822,N_1869);
or U2455 (N_2455,N_680,N_1651);
nand U2456 (N_2456,N_1021,N_575);
and U2457 (N_2457,N_333,N_340);
or U2458 (N_2458,N_16,N_286);
and U2459 (N_2459,N_1313,N_351);
nor U2460 (N_2460,N_1167,N_445);
or U2461 (N_2461,N_852,N_375);
and U2462 (N_2462,N_690,N_687);
nand U2463 (N_2463,N_967,N_1094);
or U2464 (N_2464,N_1904,N_1663);
nand U2465 (N_2465,N_1297,N_1460);
and U2466 (N_2466,N_331,N_585);
nor U2467 (N_2467,N_794,N_1065);
or U2468 (N_2468,N_1840,N_408);
or U2469 (N_2469,N_1135,N_475);
nand U2470 (N_2470,N_1857,N_1930);
nor U2471 (N_2471,N_1757,N_394);
nand U2472 (N_2472,N_812,N_70);
or U2473 (N_2473,N_1145,N_1770);
nor U2474 (N_2474,N_725,N_958);
nor U2475 (N_2475,N_1104,N_268);
xnor U2476 (N_2476,N_1309,N_1868);
xor U2477 (N_2477,N_1962,N_1045);
and U2478 (N_2478,N_505,N_1696);
nand U2479 (N_2479,N_1550,N_1615);
and U2480 (N_2480,N_1057,N_1511);
or U2481 (N_2481,N_1681,N_37);
or U2482 (N_2482,N_1767,N_1272);
or U2483 (N_2483,N_840,N_557);
nor U2484 (N_2484,N_790,N_1680);
and U2485 (N_2485,N_500,N_696);
or U2486 (N_2486,N_1631,N_527);
or U2487 (N_2487,N_990,N_88);
and U2488 (N_2488,N_1441,N_956);
or U2489 (N_2489,N_418,N_248);
nand U2490 (N_2490,N_1175,N_1771);
nand U2491 (N_2491,N_1888,N_1331);
nand U2492 (N_2492,N_1405,N_1993);
or U2493 (N_2493,N_1178,N_1569);
or U2494 (N_2494,N_1118,N_1096);
and U2495 (N_2495,N_147,N_747);
xnor U2496 (N_2496,N_928,N_1053);
nand U2497 (N_2497,N_1945,N_753);
nand U2498 (N_2498,N_1050,N_739);
and U2499 (N_2499,N_1445,N_1567);
and U2500 (N_2500,N_1604,N_1114);
and U2501 (N_2501,N_1553,N_45);
nor U2502 (N_2502,N_156,N_452);
nand U2503 (N_2503,N_415,N_1151);
nor U2504 (N_2504,N_1972,N_764);
nand U2505 (N_2505,N_976,N_1430);
and U2506 (N_2506,N_651,N_25);
nor U2507 (N_2507,N_649,N_1867);
nor U2508 (N_2508,N_877,N_767);
and U2509 (N_2509,N_1982,N_965);
and U2510 (N_2510,N_1347,N_1748);
or U2511 (N_2511,N_1950,N_1009);
nor U2512 (N_2512,N_519,N_568);
and U2513 (N_2513,N_322,N_805);
xnor U2514 (N_2514,N_1132,N_1035);
or U2515 (N_2515,N_1284,N_139);
and U2516 (N_2516,N_71,N_995);
and U2517 (N_2517,N_692,N_118);
nor U2518 (N_2518,N_1214,N_193);
and U2519 (N_2519,N_638,N_809);
nand U2520 (N_2520,N_1170,N_694);
and U2521 (N_2521,N_876,N_449);
and U2522 (N_2522,N_679,N_459);
nor U2523 (N_2523,N_1180,N_1190);
nor U2524 (N_2524,N_130,N_1871);
xnor U2525 (N_2525,N_837,N_1103);
xor U2526 (N_2526,N_1897,N_1173);
nand U2527 (N_2527,N_1338,N_1626);
and U2528 (N_2528,N_140,N_1182);
nor U2529 (N_2529,N_33,N_727);
xnor U2530 (N_2530,N_925,N_435);
and U2531 (N_2531,N_1909,N_1499);
or U2532 (N_2532,N_1404,N_1957);
nor U2533 (N_2533,N_1380,N_348);
nor U2534 (N_2534,N_378,N_1804);
nor U2535 (N_2535,N_52,N_618);
xor U2536 (N_2536,N_736,N_1815);
or U2537 (N_2537,N_1746,N_1624);
or U2538 (N_2538,N_576,N_3);
nand U2539 (N_2539,N_231,N_1407);
xor U2540 (N_2540,N_1578,N_283);
xnor U2541 (N_2541,N_185,N_1003);
or U2542 (N_2542,N_1524,N_306);
nand U2543 (N_2543,N_1025,N_1431);
or U2544 (N_2544,N_566,N_1605);
and U2545 (N_2545,N_100,N_1345);
nor U2546 (N_2546,N_1389,N_493);
and U2547 (N_2547,N_1136,N_228);
nor U2548 (N_2548,N_1127,N_309);
and U2549 (N_2549,N_1302,N_1339);
or U2550 (N_2550,N_1034,N_918);
and U2551 (N_2551,N_104,N_1055);
nand U2552 (N_2552,N_1941,N_1201);
xor U2553 (N_2553,N_1185,N_1991);
nand U2554 (N_2554,N_614,N_434);
or U2555 (N_2555,N_24,N_1775);
nor U2556 (N_2556,N_1244,N_1603);
nor U2557 (N_2557,N_427,N_1659);
or U2558 (N_2558,N_1849,N_941);
and U2559 (N_2559,N_1583,N_132);
or U2560 (N_2560,N_587,N_1344);
or U2561 (N_2561,N_417,N_204);
nand U2562 (N_2562,N_1484,N_69);
nor U2563 (N_2563,N_1973,N_975);
or U2564 (N_2564,N_722,N_729);
or U2565 (N_2565,N_1818,N_1687);
nand U2566 (N_2566,N_201,N_1555);
nor U2567 (N_2567,N_1828,N_1000);
or U2568 (N_2568,N_828,N_655);
and U2569 (N_2569,N_240,N_1953);
or U2570 (N_2570,N_923,N_610);
nor U2571 (N_2571,N_1274,N_1561);
xnor U2572 (N_2572,N_759,N_1872);
or U2573 (N_2573,N_996,N_407);
nor U2574 (N_2574,N_48,N_1683);
nand U2575 (N_2575,N_1572,N_1674);
or U2576 (N_2576,N_1212,N_1573);
or U2577 (N_2577,N_1634,N_1542);
or U2578 (N_2578,N_472,N_1218);
nor U2579 (N_2579,N_507,N_274);
nand U2580 (N_2580,N_1249,N_953);
nor U2581 (N_2581,N_783,N_985);
nor U2582 (N_2582,N_297,N_1447);
nor U2583 (N_2583,N_1914,N_624);
and U2584 (N_2584,N_515,N_1311);
or U2585 (N_2585,N_913,N_215);
and U2586 (N_2586,N_1409,N_1782);
and U2587 (N_2587,N_1188,N_1268);
nand U2588 (N_2588,N_650,N_1368);
nand U2589 (N_2589,N_573,N_329);
nand U2590 (N_2590,N_1593,N_775);
nand U2591 (N_2591,N_455,N_980);
or U2592 (N_2592,N_82,N_1221);
or U2593 (N_2593,N_1667,N_284);
or U2594 (N_2594,N_134,N_1254);
and U2595 (N_2595,N_1709,N_1994);
nand U2596 (N_2596,N_704,N_955);
and U2597 (N_2597,N_525,N_615);
nand U2598 (N_2598,N_1408,N_1608);
and U2599 (N_2599,N_1571,N_1772);
nor U2600 (N_2600,N_1161,N_1277);
xnor U2601 (N_2601,N_1071,N_412);
and U2602 (N_2602,N_469,N_1697);
nor U2603 (N_2603,N_1451,N_1908);
and U2604 (N_2604,N_808,N_275);
or U2605 (N_2605,N_1046,N_716);
nor U2606 (N_2606,N_663,N_982);
or U2607 (N_2607,N_258,N_1700);
or U2608 (N_2608,N_1977,N_1351);
or U2609 (N_2609,N_1002,N_1454);
xor U2610 (N_2610,N_1699,N_1444);
nand U2611 (N_2611,N_712,N_400);
and U2612 (N_2612,N_824,N_1364);
nor U2613 (N_2613,N_1473,N_1587);
and U2614 (N_2614,N_15,N_1599);
nand U2615 (N_2615,N_757,N_399);
nor U2616 (N_2616,N_851,N_1328);
and U2617 (N_2617,N_661,N_251);
nor U2618 (N_2618,N_1303,N_1098);
nand U2619 (N_2619,N_930,N_163);
nand U2620 (N_2620,N_1233,N_1958);
xnor U2621 (N_2621,N_911,N_269);
or U2622 (N_2622,N_162,N_1164);
or U2623 (N_2623,N_440,N_988);
nor U2624 (N_2624,N_347,N_754);
nand U2625 (N_2625,N_818,N_535);
or U2626 (N_2626,N_203,N_1806);
and U2627 (N_2627,N_161,N_893);
xor U2628 (N_2628,N_1738,N_659);
xnor U2629 (N_2629,N_1707,N_1737);
nor U2630 (N_2630,N_1534,N_1959);
nand U2631 (N_2631,N_1419,N_1298);
and U2632 (N_2632,N_1861,N_770);
nand U2633 (N_2633,N_356,N_625);
nor U2634 (N_2634,N_1751,N_453);
xor U2635 (N_2635,N_822,N_1250);
or U2636 (N_2636,N_1685,N_1085);
nand U2637 (N_2637,N_1665,N_337);
nor U2638 (N_2638,N_91,N_304);
or U2639 (N_2639,N_503,N_516);
nor U2640 (N_2640,N_984,N_1415);
nand U2641 (N_2641,N_1703,N_1842);
nor U2642 (N_2642,N_295,N_265);
and U2643 (N_2643,N_1817,N_1988);
nor U2644 (N_2644,N_430,N_84);
nor U2645 (N_2645,N_326,N_1493);
or U2646 (N_2646,N_424,N_778);
or U2647 (N_2647,N_374,N_518);
nor U2648 (N_2648,N_843,N_1672);
nand U2649 (N_2649,N_194,N_81);
nand U2650 (N_2650,N_62,N_658);
or U2651 (N_2651,N_1657,N_2);
or U2652 (N_2652,N_221,N_1750);
nand U2653 (N_2653,N_296,N_732);
and U2654 (N_2654,N_1306,N_74);
or U2655 (N_2655,N_1308,N_41);
nand U2656 (N_2656,N_1981,N_46);
nand U2657 (N_2657,N_726,N_1642);
nor U2658 (N_2658,N_1333,N_42);
or U2659 (N_2659,N_27,N_713);
xor U2660 (N_2660,N_1381,N_1893);
and U2661 (N_2661,N_755,N_1087);
or U2662 (N_2662,N_451,N_1083);
nand U2663 (N_2663,N_561,N_1640);
or U2664 (N_2664,N_79,N_1721);
nand U2665 (N_2665,N_1110,N_1258);
nand U2666 (N_2666,N_354,N_534);
xnor U2667 (N_2667,N_112,N_1645);
or U2668 (N_2668,N_945,N_889);
or U2669 (N_2669,N_1394,N_800);
nand U2670 (N_2670,N_220,N_1796);
or U2671 (N_2671,N_1080,N_1730);
and U2672 (N_2672,N_101,N_1809);
xor U2673 (N_2673,N_1426,N_392);
nand U2674 (N_2674,N_1481,N_1701);
xor U2675 (N_2675,N_1610,N_1393);
nor U2676 (N_2676,N_606,N_17);
nand U2677 (N_2677,N_762,N_1502);
and U2678 (N_2678,N_1215,N_1987);
nand U2679 (N_2679,N_1661,N_1946);
and U2680 (N_2680,N_592,N_1792);
and U2681 (N_2681,N_539,N_1111);
nor U2682 (N_2682,N_1310,N_1436);
nand U2683 (N_2683,N_1189,N_942);
nand U2684 (N_2684,N_1636,N_254);
nor U2685 (N_2685,N_1004,N_682);
nor U2686 (N_2686,N_1186,N_1660);
or U2687 (N_2687,N_86,N_1041);
nor U2688 (N_2688,N_1915,N_1932);
xor U2689 (N_2689,N_233,N_1360);
nor U2690 (N_2690,N_218,N_1199);
nand U2691 (N_2691,N_302,N_1066);
xor U2692 (N_2692,N_1936,N_1956);
nand U2693 (N_2693,N_419,N_1985);
or U2694 (N_2694,N_881,N_1781);
nand U2695 (N_2695,N_1678,N_542);
xnor U2696 (N_2696,N_1141,N_180);
and U2697 (N_2697,N_1791,N_509);
and U2698 (N_2698,N_481,N_869);
nand U2699 (N_2699,N_989,N_1803);
nor U2700 (N_2700,N_102,N_1172);
nand U2701 (N_2701,N_443,N_492);
nor U2702 (N_2702,N_1392,N_1334);
or U2703 (N_2703,N_1727,N_1739);
or U2704 (N_2704,N_1299,N_920);
nor U2705 (N_2705,N_586,N_570);
nand U2706 (N_2706,N_671,N_1582);
nor U2707 (N_2707,N_952,N_391);
and U2708 (N_2708,N_875,N_1954);
and U2709 (N_2709,N_588,N_1518);
nor U2710 (N_2710,N_1156,N_1563);
and U2711 (N_2711,N_1322,N_1005);
nand U2712 (N_2712,N_1852,N_305);
and U2713 (N_2713,N_748,N_301);
or U2714 (N_2714,N_314,N_1482);
nor U2715 (N_2715,N_1533,N_811);
or U2716 (N_2716,N_1323,N_124);
or U2717 (N_2717,N_1734,N_708);
nor U2718 (N_2718,N_105,N_998);
and U2719 (N_2719,N_944,N_643);
or U2720 (N_2720,N_404,N_1260);
nand U2721 (N_2721,N_1077,N_1273);
and U2722 (N_2722,N_1397,N_200);
nor U2723 (N_2723,N_1031,N_450);
nand U2724 (N_2724,N_1836,N_635);
nor U2725 (N_2725,N_797,N_1092);
nor U2726 (N_2726,N_324,N_777);
and U2727 (N_2727,N_868,N_1652);
and U2728 (N_2728,N_1568,N_1213);
nand U2729 (N_2729,N_1975,N_699);
nand U2730 (N_2730,N_59,N_743);
or U2731 (N_2731,N_508,N_108);
and U2732 (N_2732,N_1446,N_662);
nor U2733 (N_2733,N_175,N_938);
or U2734 (N_2734,N_1793,N_1878);
nand U2735 (N_2735,N_1894,N_514);
or U2736 (N_2736,N_681,N_1938);
and U2737 (N_2737,N_1628,N_1240);
or U2738 (N_2738,N_673,N_639);
nand U2739 (N_2739,N_1072,N_1850);
and U2740 (N_2740,N_1823,N_765);
nand U2741 (N_2741,N_1921,N_349);
nor U2742 (N_2742,N_801,N_937);
nor U2743 (N_2743,N_1766,N_334);
nand U2744 (N_2744,N_376,N_1459);
or U2745 (N_2745,N_1591,N_701);
or U2746 (N_2746,N_75,N_1131);
or U2747 (N_2747,N_150,N_543);
nor U2748 (N_2748,N_947,N_393);
or U2749 (N_2749,N_127,N_1361);
and U2750 (N_2750,N_1805,N_547);
nor U2751 (N_2751,N_836,N_138);
nand U2752 (N_2752,N_1917,N_830);
xnor U2753 (N_2753,N_208,N_1448);
nor U2754 (N_2754,N_1947,N_959);
nor U2755 (N_2755,N_934,N_111);
xor U2756 (N_2756,N_1714,N_1399);
or U2757 (N_2757,N_1708,N_1986);
nor U2758 (N_2758,N_1157,N_315);
or U2759 (N_2759,N_1093,N_1789);
or U2760 (N_2760,N_1356,N_1073);
nor U2761 (N_2761,N_1996,N_1557);
nand U2762 (N_2762,N_467,N_1106);
nor U2763 (N_2763,N_847,N_1761);
nor U2764 (N_2764,N_1265,N_1655);
xor U2765 (N_2765,N_377,N_510);
nand U2766 (N_2766,N_1594,N_264);
nand U2767 (N_2767,N_737,N_533);
or U2768 (N_2768,N_1225,N_621);
nor U2769 (N_2769,N_1799,N_793);
or U2770 (N_2770,N_703,N_981);
nand U2771 (N_2771,N_506,N_700);
and U2772 (N_2772,N_373,N_892);
nand U2773 (N_2773,N_921,N_1649);
nor U2774 (N_2774,N_1207,N_1564);
or U2775 (N_2775,N_1196,N_253);
nor U2776 (N_2776,N_448,N_1030);
and U2777 (N_2777,N_252,N_498);
nor U2778 (N_2778,N_1510,N_1641);
or U2779 (N_2779,N_342,N_174);
and U2780 (N_2780,N_1084,N_222);
and U2781 (N_2781,N_1319,N_849);
or U2782 (N_2782,N_1020,N_720);
or U2783 (N_2783,N_1124,N_523);
nor U2784 (N_2784,N_241,N_964);
and U2785 (N_2785,N_155,N_1764);
nor U2786 (N_2786,N_609,N_1224);
or U2787 (N_2787,N_1293,N_460);
xnor U2788 (N_2788,N_43,N_810);
nor U2789 (N_2789,N_355,N_1870);
nor U2790 (N_2790,N_484,N_1673);
nand U2791 (N_2791,N_1486,N_1259);
and U2792 (N_2792,N_90,N_1961);
or U2793 (N_2793,N_1300,N_1810);
and U2794 (N_2794,N_1951,N_10);
and U2795 (N_2795,N_686,N_907);
nand U2796 (N_2796,N_117,N_1247);
xor U2797 (N_2797,N_536,N_1735);
and U2798 (N_2798,N_1239,N_496);
or U2799 (N_2799,N_1367,N_363);
and U2800 (N_2800,N_1464,N_179);
nor U2801 (N_2801,N_1078,N_1505);
nor U2802 (N_2802,N_35,N_491);
or U2803 (N_2803,N_577,N_1337);
nor U2804 (N_2804,N_1556,N_1011);
and U2805 (N_2805,N_1801,N_931);
and U2806 (N_2806,N_1710,N_1488);
nor U2807 (N_2807,N_723,N_367);
or U2808 (N_2808,N_549,N_761);
nand U2809 (N_2809,N_115,N_1195);
or U2810 (N_2810,N_141,N_579);
or U2811 (N_2811,N_143,N_648);
nor U2812 (N_2812,N_1369,N_632);
nor U2813 (N_2813,N_1741,N_1627);
nand U2814 (N_2814,N_1998,N_1059);
nand U2815 (N_2815,N_1745,N_464);
nand U2816 (N_2816,N_558,N_745);
and U2817 (N_2817,N_1241,N_1577);
or U2818 (N_2818,N_364,N_1068);
and U2819 (N_2819,N_850,N_1763);
nand U2820 (N_2820,N_210,N_544);
or U2821 (N_2821,N_1760,N_1023);
and U2822 (N_2822,N_126,N_273);
nand U2823 (N_2823,N_939,N_1470);
and U2824 (N_2824,N_121,N_1346);
nor U2825 (N_2825,N_89,N_159);
and U2826 (N_2826,N_217,N_224);
and U2827 (N_2827,N_1885,N_202);
and U2828 (N_2828,N_1081,N_785);
xor U2829 (N_2829,N_946,N_504);
nand U2830 (N_2830,N_1440,N_1455);
nor U2831 (N_2831,N_1101,N_1411);
and U2832 (N_2832,N_1913,N_1427);
xnor U2833 (N_2833,N_1276,N_698);
and U2834 (N_2834,N_245,N_802);
nand U2835 (N_2835,N_1937,N_1458);
and U2836 (N_2836,N_886,N_1732);
xor U2837 (N_2837,N_1044,N_1650);
xnor U2838 (N_2838,N_1070,N_1943);
nand U2839 (N_2839,N_1754,N_1374);
and U2840 (N_2840,N_1939,N_350);
xnor U2841 (N_2841,N_555,N_125);
nor U2842 (N_2842,N_1919,N_1644);
xor U2843 (N_2843,N_1133,N_1457);
nor U2844 (N_2844,N_1881,N_885);
and U2845 (N_2845,N_368,N_1100);
or U2846 (N_2846,N_1006,N_1968);
nand U2847 (N_2847,N_1422,N_668);
nand U2848 (N_2848,N_871,N_213);
nand U2849 (N_2849,N_403,N_816);
and U2850 (N_2850,N_420,N_1854);
or U2851 (N_2851,N_1720,N_186);
and U2852 (N_2852,N_846,N_888);
or U2853 (N_2853,N_1507,N_581);
nand U2854 (N_2854,N_1352,N_1197);
and U2855 (N_2855,N_237,N_225);
nand U2856 (N_2856,N_223,N_58);
and U2857 (N_2857,N_1620,N_1579);
nand U2858 (N_2858,N_61,N_560);
nand U2859 (N_2859,N_501,N_290);
nand U2860 (N_2860,N_370,N_190);
nand U2861 (N_2861,N_1704,N_637);
nor U2862 (N_2862,N_66,N_1326);
nand U2863 (N_2863,N_1278,N_773);
and U2864 (N_2864,N_327,N_1967);
or U2865 (N_2865,N_1231,N_1418);
nand U2866 (N_2866,N_1541,N_879);
or U2867 (N_2867,N_63,N_178);
and U2868 (N_2868,N_1024,N_1152);
nor U2869 (N_2869,N_226,N_234);
and U2870 (N_2870,N_714,N_458);
nor U2871 (N_2871,N_899,N_1841);
xnor U2872 (N_2872,N_1768,N_396);
and U2873 (N_2873,N_249,N_1038);
xor U2874 (N_2874,N_1638,N_1574);
nand U2875 (N_2875,N_68,N_1242);
nand U2876 (N_2876,N_1234,N_1523);
and U2877 (N_2877,N_480,N_1560);
nor U2878 (N_2878,N_405,N_1614);
and U2879 (N_2879,N_488,N_1229);
nor U2880 (N_2880,N_1545,N_1728);
nand U2881 (N_2881,N_1424,N_1330);
nand U2882 (N_2882,N_436,N_1383);
nand U2883 (N_2883,N_1753,N_1686);
nand U2884 (N_2884,N_1429,N_1812);
nor U2885 (N_2885,N_401,N_541);
and U2886 (N_2886,N_167,N_1267);
and U2887 (N_2887,N_861,N_620);
nand U2888 (N_2888,N_636,N_1466);
nor U2889 (N_2889,N_1099,N_1018);
or U2890 (N_2890,N_1639,N_1263);
and U2891 (N_2891,N_352,N_641);
nor U2892 (N_2892,N_1501,N_909);
or U2893 (N_2893,N_1546,N_553);
nand U2894 (N_2894,N_1873,N_1601);
or U2895 (N_2895,N_874,N_511);
nand U2896 (N_2896,N_526,N_1834);
and U2897 (N_2897,N_709,N_1552);
and U2898 (N_2898,N_439,N_1291);
and U2899 (N_2899,N_110,N_1617);
xnor U2900 (N_2900,N_198,N_1315);
and U2901 (N_2901,N_255,N_1983);
nand U2902 (N_2902,N_616,N_738);
nor U2903 (N_2903,N_1029,N_1208);
and U2904 (N_2904,N_1889,N_936);
and U2905 (N_2905,N_551,N_1008);
nand U2906 (N_2906,N_1675,N_603);
and U2907 (N_2907,N_994,N_1860);
nand U2908 (N_2908,N_1280,N_72);
nor U2909 (N_2909,N_1256,N_1891);
xnor U2910 (N_2910,N_123,N_825);
or U2911 (N_2911,N_341,N_267);
or U2912 (N_2912,N_910,N_1816);
and U2913 (N_2913,N_1978,N_796);
or U2914 (N_2914,N_5,N_1588);
nand U2915 (N_2915,N_1506,N_1435);
nor U2916 (N_2916,N_711,N_979);
xnor U2917 (N_2917,N_872,N_627);
and U2918 (N_2918,N_1629,N_1827);
or U2919 (N_2919,N_572,N_912);
nor U2920 (N_2920,N_1194,N_1134);
and U2921 (N_2921,N_860,N_878);
xnor U2922 (N_2922,N_1471,N_1514);
nand U2923 (N_2923,N_617,N_569);
nor U2924 (N_2924,N_1119,N_1075);
nand U2925 (N_2925,N_494,N_589);
nand U2926 (N_2926,N_1462,N_1363);
nand U2927 (N_2927,N_1232,N_1371);
and U2928 (N_2928,N_1879,N_1934);
nor U2929 (N_2929,N_1036,N_1864);
nand U2930 (N_2930,N_1223,N_1230);
nor U2931 (N_2931,N_19,N_640);
and U2932 (N_2932,N_567,N_596);
and U2933 (N_2933,N_358,N_1433);
and U2934 (N_2934,N_388,N_53);
or U2935 (N_2935,N_1762,N_78);
or U2936 (N_2936,N_763,N_1692);
or U2937 (N_2937,N_862,N_1095);
or U2938 (N_2938,N_1520,N_1012);
and U2939 (N_2939,N_657,N_1314);
nand U2940 (N_2940,N_83,N_1676);
or U2941 (N_2941,N_1198,N_951);
nand U2942 (N_2942,N_602,N_1412);
nand U2943 (N_2943,N_320,N_381);
or U2944 (N_2944,N_642,N_1495);
and U2945 (N_2945,N_261,N_870);
nand U2946 (N_2946,N_1955,N_95);
or U2947 (N_2947,N_209,N_1785);
nor U2948 (N_2948,N_1662,N_1530);
or U2949 (N_2949,N_122,N_1880);
or U2950 (N_2950,N_1192,N_1979);
nor U2951 (N_2951,N_382,N_1007);
nor U2952 (N_2952,N_1316,N_528);
nor U2953 (N_2953,N_769,N_1117);
nand U2954 (N_2954,N_1349,N_1168);
and U2955 (N_2955,N_160,N_1378);
nor U2956 (N_2956,N_629,N_1478);
xnor U2957 (N_2957,N_360,N_177);
nor U2958 (N_2958,N_1219,N_1112);
nor U2959 (N_2959,N_1606,N_1726);
nand U2960 (N_2960,N_1743,N_256);
or U2961 (N_2961,N_1544,N_597);
nand U2962 (N_2962,N_845,N_1503);
and U2963 (N_2963,N_1452,N_537);
nor U2964 (N_2964,N_199,N_1677);
xor U2965 (N_2965,N_1521,N_1581);
or U2966 (N_2966,N_1562,N_1200);
nor U2967 (N_2967,N_1043,N_1491);
or U2968 (N_2968,N_835,N_1439);
nand U2969 (N_2969,N_1490,N_1017);
or U2970 (N_2970,N_289,N_607);
nor U2971 (N_2971,N_966,N_1526);
or U2972 (N_2972,N_120,N_1742);
nor U2973 (N_2973,N_1410,N_1607);
nand U2974 (N_2974,N_646,N_145);
nor U2975 (N_2975,N_1144,N_212);
or U2976 (N_2976,N_1027,N_1723);
and U2977 (N_2977,N_1886,N_1689);
or U2978 (N_2978,N_1123,N_1090);
xor U2979 (N_2979,N_550,N_524);
nand U2980 (N_2980,N_1942,N_848);
nor U2981 (N_2981,N_330,N_14);
xnor U2982 (N_2982,N_1174,N_1565);
nor U2983 (N_2983,N_595,N_425);
nor U2984 (N_2984,N_1498,N_12);
xor U2985 (N_2985,N_1487,N_332);
or U2986 (N_2986,N_1437,N_1261);
nand U2987 (N_2987,N_1385,N_806);
xnor U2988 (N_2988,N_977,N_1116);
and U2989 (N_2989,N_924,N_1883);
nor U2990 (N_2990,N_1765,N_772);
or U2991 (N_2991,N_583,N_619);
or U2992 (N_2992,N_693,N_798);
and U2993 (N_2993,N_478,N_1220);
and U2994 (N_2994,N_1525,N_1343);
and U2995 (N_2995,N_1169,N_1695);
or U2996 (N_2996,N_463,N_1596);
nand U2997 (N_2997,N_1851,N_1616);
xor U2998 (N_2998,N_144,N_1855);
nor U2999 (N_2999,N_1022,N_815);
nand U3000 (N_3000,N_788,N_1189);
and U3001 (N_3001,N_1232,N_799);
and U3002 (N_3002,N_1511,N_1109);
and U3003 (N_3003,N_111,N_998);
nand U3004 (N_3004,N_1483,N_422);
nor U3005 (N_3005,N_1064,N_294);
or U3006 (N_3006,N_379,N_1125);
nand U3007 (N_3007,N_399,N_900);
or U3008 (N_3008,N_233,N_1743);
and U3009 (N_3009,N_1969,N_221);
xnor U3010 (N_3010,N_1914,N_770);
nor U3011 (N_3011,N_607,N_153);
nor U3012 (N_3012,N_1055,N_518);
and U3013 (N_3013,N_1584,N_1490);
nor U3014 (N_3014,N_1610,N_1203);
xor U3015 (N_3015,N_621,N_1206);
nor U3016 (N_3016,N_293,N_321);
or U3017 (N_3017,N_1468,N_1933);
xnor U3018 (N_3018,N_1259,N_1122);
nor U3019 (N_3019,N_978,N_621);
nand U3020 (N_3020,N_1598,N_1697);
and U3021 (N_3021,N_1528,N_353);
or U3022 (N_3022,N_1913,N_1530);
or U3023 (N_3023,N_19,N_1981);
or U3024 (N_3024,N_1074,N_828);
nand U3025 (N_3025,N_1293,N_752);
and U3026 (N_3026,N_1118,N_1966);
or U3027 (N_3027,N_1086,N_403);
and U3028 (N_3028,N_158,N_996);
xor U3029 (N_3029,N_1011,N_847);
and U3030 (N_3030,N_142,N_82);
or U3031 (N_3031,N_1049,N_888);
and U3032 (N_3032,N_1878,N_567);
nand U3033 (N_3033,N_1334,N_832);
and U3034 (N_3034,N_469,N_228);
and U3035 (N_3035,N_1899,N_1569);
nand U3036 (N_3036,N_1776,N_802);
nand U3037 (N_3037,N_754,N_1674);
or U3038 (N_3038,N_1720,N_798);
and U3039 (N_3039,N_1261,N_1940);
or U3040 (N_3040,N_585,N_985);
nor U3041 (N_3041,N_1203,N_346);
xor U3042 (N_3042,N_1689,N_1656);
nand U3043 (N_3043,N_1334,N_1824);
and U3044 (N_3044,N_919,N_899);
and U3045 (N_3045,N_1303,N_26);
and U3046 (N_3046,N_1561,N_1910);
or U3047 (N_3047,N_596,N_172);
nor U3048 (N_3048,N_781,N_1043);
nor U3049 (N_3049,N_1275,N_1559);
and U3050 (N_3050,N_466,N_660);
and U3051 (N_3051,N_992,N_1029);
or U3052 (N_3052,N_297,N_788);
nand U3053 (N_3053,N_1565,N_1512);
nand U3054 (N_3054,N_1149,N_243);
nor U3055 (N_3055,N_5,N_555);
or U3056 (N_3056,N_275,N_483);
nor U3057 (N_3057,N_512,N_719);
and U3058 (N_3058,N_1592,N_511);
nand U3059 (N_3059,N_219,N_1705);
and U3060 (N_3060,N_318,N_1613);
xor U3061 (N_3061,N_544,N_529);
or U3062 (N_3062,N_1556,N_245);
xnor U3063 (N_3063,N_1505,N_694);
nor U3064 (N_3064,N_1484,N_98);
nor U3065 (N_3065,N_1911,N_870);
or U3066 (N_3066,N_905,N_1276);
and U3067 (N_3067,N_886,N_1677);
or U3068 (N_3068,N_1364,N_1367);
nand U3069 (N_3069,N_1290,N_492);
nand U3070 (N_3070,N_478,N_386);
nor U3071 (N_3071,N_1491,N_54);
and U3072 (N_3072,N_484,N_1207);
or U3073 (N_3073,N_866,N_469);
nand U3074 (N_3074,N_1865,N_535);
and U3075 (N_3075,N_766,N_693);
nor U3076 (N_3076,N_230,N_994);
nor U3077 (N_3077,N_185,N_468);
and U3078 (N_3078,N_97,N_63);
nand U3079 (N_3079,N_776,N_762);
or U3080 (N_3080,N_1111,N_223);
and U3081 (N_3081,N_1454,N_478);
xnor U3082 (N_3082,N_1733,N_721);
or U3083 (N_3083,N_1517,N_1666);
nand U3084 (N_3084,N_783,N_1252);
nor U3085 (N_3085,N_139,N_1140);
or U3086 (N_3086,N_1339,N_939);
nand U3087 (N_3087,N_803,N_1299);
nand U3088 (N_3088,N_1473,N_286);
nor U3089 (N_3089,N_370,N_1893);
and U3090 (N_3090,N_448,N_88);
nor U3091 (N_3091,N_589,N_683);
or U3092 (N_3092,N_1798,N_852);
nand U3093 (N_3093,N_189,N_1696);
nand U3094 (N_3094,N_1288,N_179);
nand U3095 (N_3095,N_1871,N_480);
nand U3096 (N_3096,N_432,N_1128);
or U3097 (N_3097,N_619,N_28);
nand U3098 (N_3098,N_648,N_1469);
xnor U3099 (N_3099,N_1408,N_34);
nand U3100 (N_3100,N_1065,N_1729);
or U3101 (N_3101,N_746,N_1968);
nand U3102 (N_3102,N_1424,N_1564);
or U3103 (N_3103,N_47,N_1867);
nand U3104 (N_3104,N_72,N_535);
nand U3105 (N_3105,N_180,N_789);
or U3106 (N_3106,N_552,N_132);
nand U3107 (N_3107,N_1678,N_170);
nor U3108 (N_3108,N_112,N_1962);
or U3109 (N_3109,N_655,N_1999);
and U3110 (N_3110,N_363,N_398);
nand U3111 (N_3111,N_525,N_757);
nand U3112 (N_3112,N_1843,N_350);
nor U3113 (N_3113,N_1887,N_1044);
xor U3114 (N_3114,N_437,N_492);
or U3115 (N_3115,N_1004,N_1111);
nand U3116 (N_3116,N_1004,N_520);
nand U3117 (N_3117,N_1886,N_1963);
nand U3118 (N_3118,N_1638,N_347);
and U3119 (N_3119,N_258,N_1817);
xor U3120 (N_3120,N_1240,N_838);
or U3121 (N_3121,N_1541,N_1063);
nand U3122 (N_3122,N_1862,N_671);
nor U3123 (N_3123,N_741,N_877);
or U3124 (N_3124,N_1415,N_1811);
xor U3125 (N_3125,N_1436,N_1205);
nand U3126 (N_3126,N_1742,N_233);
and U3127 (N_3127,N_94,N_66);
xnor U3128 (N_3128,N_1853,N_466);
or U3129 (N_3129,N_1742,N_148);
or U3130 (N_3130,N_1228,N_1352);
and U3131 (N_3131,N_1337,N_1738);
nor U3132 (N_3132,N_1965,N_1209);
and U3133 (N_3133,N_755,N_877);
xnor U3134 (N_3134,N_1123,N_1977);
nand U3135 (N_3135,N_1071,N_36);
and U3136 (N_3136,N_301,N_1630);
or U3137 (N_3137,N_963,N_343);
nor U3138 (N_3138,N_1728,N_582);
and U3139 (N_3139,N_404,N_1746);
and U3140 (N_3140,N_1091,N_1455);
xor U3141 (N_3141,N_578,N_324);
nand U3142 (N_3142,N_319,N_417);
nand U3143 (N_3143,N_1083,N_1241);
and U3144 (N_3144,N_305,N_804);
and U3145 (N_3145,N_1175,N_1576);
nor U3146 (N_3146,N_773,N_1946);
and U3147 (N_3147,N_1373,N_1372);
nand U3148 (N_3148,N_506,N_468);
nand U3149 (N_3149,N_1598,N_1526);
nor U3150 (N_3150,N_1606,N_1464);
or U3151 (N_3151,N_987,N_1745);
or U3152 (N_3152,N_826,N_146);
xor U3153 (N_3153,N_779,N_1788);
xnor U3154 (N_3154,N_371,N_751);
and U3155 (N_3155,N_998,N_1649);
or U3156 (N_3156,N_1667,N_109);
nand U3157 (N_3157,N_23,N_1727);
or U3158 (N_3158,N_639,N_479);
nand U3159 (N_3159,N_1323,N_1741);
nor U3160 (N_3160,N_287,N_1759);
or U3161 (N_3161,N_181,N_608);
nor U3162 (N_3162,N_1564,N_441);
nor U3163 (N_3163,N_1317,N_1603);
xnor U3164 (N_3164,N_1433,N_612);
nand U3165 (N_3165,N_17,N_441);
nor U3166 (N_3166,N_1515,N_344);
nor U3167 (N_3167,N_1747,N_483);
nand U3168 (N_3168,N_744,N_319);
nand U3169 (N_3169,N_1238,N_551);
xnor U3170 (N_3170,N_162,N_111);
and U3171 (N_3171,N_1873,N_1400);
nor U3172 (N_3172,N_1578,N_1366);
nor U3173 (N_3173,N_663,N_1186);
or U3174 (N_3174,N_293,N_588);
nand U3175 (N_3175,N_351,N_1565);
or U3176 (N_3176,N_1899,N_495);
nand U3177 (N_3177,N_1353,N_1066);
and U3178 (N_3178,N_351,N_1038);
xnor U3179 (N_3179,N_1651,N_1423);
or U3180 (N_3180,N_251,N_1055);
xnor U3181 (N_3181,N_317,N_617);
and U3182 (N_3182,N_575,N_19);
and U3183 (N_3183,N_395,N_1909);
and U3184 (N_3184,N_498,N_584);
nor U3185 (N_3185,N_1970,N_103);
and U3186 (N_3186,N_1618,N_445);
and U3187 (N_3187,N_1600,N_921);
nand U3188 (N_3188,N_181,N_337);
nor U3189 (N_3189,N_1437,N_1078);
or U3190 (N_3190,N_1998,N_1906);
nor U3191 (N_3191,N_121,N_136);
or U3192 (N_3192,N_992,N_390);
xnor U3193 (N_3193,N_1619,N_1719);
nand U3194 (N_3194,N_1672,N_1651);
nand U3195 (N_3195,N_968,N_246);
or U3196 (N_3196,N_372,N_994);
xnor U3197 (N_3197,N_1806,N_1366);
nand U3198 (N_3198,N_284,N_112);
xor U3199 (N_3199,N_580,N_1891);
nand U3200 (N_3200,N_1257,N_142);
nor U3201 (N_3201,N_1840,N_15);
nor U3202 (N_3202,N_1022,N_101);
and U3203 (N_3203,N_1230,N_1793);
nand U3204 (N_3204,N_974,N_134);
and U3205 (N_3205,N_629,N_1039);
and U3206 (N_3206,N_824,N_610);
or U3207 (N_3207,N_1425,N_1101);
nand U3208 (N_3208,N_0,N_1796);
and U3209 (N_3209,N_553,N_1686);
nand U3210 (N_3210,N_1207,N_1934);
and U3211 (N_3211,N_249,N_1001);
or U3212 (N_3212,N_32,N_817);
nand U3213 (N_3213,N_1689,N_1028);
and U3214 (N_3214,N_425,N_1610);
or U3215 (N_3215,N_1550,N_811);
and U3216 (N_3216,N_15,N_982);
nor U3217 (N_3217,N_842,N_1916);
or U3218 (N_3218,N_1440,N_403);
and U3219 (N_3219,N_730,N_69);
or U3220 (N_3220,N_1088,N_1141);
nand U3221 (N_3221,N_544,N_758);
nor U3222 (N_3222,N_1633,N_54);
and U3223 (N_3223,N_1448,N_892);
or U3224 (N_3224,N_826,N_1458);
or U3225 (N_3225,N_575,N_1642);
nor U3226 (N_3226,N_217,N_1547);
or U3227 (N_3227,N_305,N_847);
nand U3228 (N_3228,N_335,N_198);
xnor U3229 (N_3229,N_1514,N_278);
nor U3230 (N_3230,N_1028,N_366);
nand U3231 (N_3231,N_1031,N_518);
nand U3232 (N_3232,N_1353,N_114);
or U3233 (N_3233,N_1845,N_1860);
nand U3234 (N_3234,N_1505,N_1672);
and U3235 (N_3235,N_265,N_900);
and U3236 (N_3236,N_1561,N_1071);
or U3237 (N_3237,N_494,N_507);
or U3238 (N_3238,N_1791,N_623);
or U3239 (N_3239,N_1145,N_1201);
and U3240 (N_3240,N_1485,N_1489);
nand U3241 (N_3241,N_1425,N_5);
nand U3242 (N_3242,N_1181,N_1290);
and U3243 (N_3243,N_1616,N_1363);
nand U3244 (N_3244,N_1229,N_1782);
or U3245 (N_3245,N_2,N_1467);
and U3246 (N_3246,N_1651,N_1932);
nand U3247 (N_3247,N_1166,N_685);
or U3248 (N_3248,N_862,N_392);
or U3249 (N_3249,N_1483,N_817);
xnor U3250 (N_3250,N_1179,N_376);
and U3251 (N_3251,N_488,N_82);
or U3252 (N_3252,N_141,N_1650);
or U3253 (N_3253,N_1472,N_1409);
nand U3254 (N_3254,N_1153,N_1691);
and U3255 (N_3255,N_1425,N_562);
nor U3256 (N_3256,N_1432,N_1880);
nand U3257 (N_3257,N_1487,N_365);
and U3258 (N_3258,N_139,N_1365);
nand U3259 (N_3259,N_1769,N_1094);
and U3260 (N_3260,N_521,N_1935);
and U3261 (N_3261,N_91,N_1583);
or U3262 (N_3262,N_386,N_1697);
or U3263 (N_3263,N_1891,N_269);
or U3264 (N_3264,N_1094,N_1074);
nand U3265 (N_3265,N_1218,N_1776);
or U3266 (N_3266,N_1213,N_1643);
nand U3267 (N_3267,N_1376,N_383);
nor U3268 (N_3268,N_269,N_576);
nor U3269 (N_3269,N_434,N_817);
or U3270 (N_3270,N_457,N_596);
nand U3271 (N_3271,N_1831,N_1748);
or U3272 (N_3272,N_1711,N_1410);
nor U3273 (N_3273,N_464,N_365);
and U3274 (N_3274,N_1016,N_403);
and U3275 (N_3275,N_194,N_430);
or U3276 (N_3276,N_1602,N_1170);
or U3277 (N_3277,N_1510,N_470);
or U3278 (N_3278,N_14,N_696);
nand U3279 (N_3279,N_859,N_211);
nand U3280 (N_3280,N_1231,N_209);
and U3281 (N_3281,N_1317,N_1454);
nor U3282 (N_3282,N_1620,N_1804);
or U3283 (N_3283,N_1345,N_329);
nor U3284 (N_3284,N_7,N_942);
nand U3285 (N_3285,N_650,N_1977);
or U3286 (N_3286,N_1638,N_1615);
or U3287 (N_3287,N_1263,N_727);
or U3288 (N_3288,N_962,N_509);
nand U3289 (N_3289,N_377,N_1320);
and U3290 (N_3290,N_403,N_581);
nand U3291 (N_3291,N_461,N_1614);
nand U3292 (N_3292,N_538,N_1245);
xnor U3293 (N_3293,N_1069,N_139);
and U3294 (N_3294,N_235,N_1724);
xor U3295 (N_3295,N_1896,N_667);
and U3296 (N_3296,N_115,N_141);
xnor U3297 (N_3297,N_60,N_1509);
or U3298 (N_3298,N_1800,N_1173);
and U3299 (N_3299,N_353,N_1871);
nand U3300 (N_3300,N_10,N_1451);
nand U3301 (N_3301,N_1734,N_1177);
and U3302 (N_3302,N_10,N_835);
nand U3303 (N_3303,N_804,N_793);
or U3304 (N_3304,N_118,N_1716);
nor U3305 (N_3305,N_525,N_1912);
and U3306 (N_3306,N_390,N_687);
and U3307 (N_3307,N_902,N_1699);
or U3308 (N_3308,N_438,N_129);
nor U3309 (N_3309,N_1945,N_724);
nand U3310 (N_3310,N_798,N_1956);
or U3311 (N_3311,N_64,N_1958);
or U3312 (N_3312,N_1690,N_1760);
nand U3313 (N_3313,N_16,N_701);
or U3314 (N_3314,N_807,N_301);
nand U3315 (N_3315,N_1599,N_1071);
nand U3316 (N_3316,N_1715,N_1336);
and U3317 (N_3317,N_594,N_1141);
xnor U3318 (N_3318,N_934,N_602);
nor U3319 (N_3319,N_1881,N_1428);
or U3320 (N_3320,N_455,N_402);
nand U3321 (N_3321,N_1324,N_931);
and U3322 (N_3322,N_1637,N_12);
and U3323 (N_3323,N_429,N_173);
or U3324 (N_3324,N_71,N_1804);
or U3325 (N_3325,N_1373,N_1420);
xor U3326 (N_3326,N_1249,N_220);
nand U3327 (N_3327,N_1676,N_61);
nand U3328 (N_3328,N_590,N_342);
nor U3329 (N_3329,N_1051,N_701);
or U3330 (N_3330,N_43,N_1648);
and U3331 (N_3331,N_176,N_222);
nor U3332 (N_3332,N_1655,N_1703);
xor U3333 (N_3333,N_22,N_1482);
nor U3334 (N_3334,N_544,N_1766);
nand U3335 (N_3335,N_857,N_921);
and U3336 (N_3336,N_1038,N_967);
nand U3337 (N_3337,N_186,N_1237);
nand U3338 (N_3338,N_1621,N_220);
xor U3339 (N_3339,N_1959,N_46);
nand U3340 (N_3340,N_1754,N_1522);
xor U3341 (N_3341,N_697,N_236);
nor U3342 (N_3342,N_1638,N_796);
nand U3343 (N_3343,N_1126,N_1910);
and U3344 (N_3344,N_1618,N_139);
nand U3345 (N_3345,N_1504,N_1073);
nand U3346 (N_3346,N_1916,N_784);
nor U3347 (N_3347,N_190,N_1766);
nor U3348 (N_3348,N_181,N_508);
or U3349 (N_3349,N_214,N_185);
nand U3350 (N_3350,N_1670,N_194);
nand U3351 (N_3351,N_337,N_1930);
nor U3352 (N_3352,N_1182,N_1066);
and U3353 (N_3353,N_626,N_664);
or U3354 (N_3354,N_1396,N_504);
and U3355 (N_3355,N_1075,N_1391);
xnor U3356 (N_3356,N_1174,N_588);
nor U3357 (N_3357,N_1946,N_1720);
or U3358 (N_3358,N_52,N_1673);
and U3359 (N_3359,N_1939,N_1222);
nor U3360 (N_3360,N_1528,N_763);
or U3361 (N_3361,N_603,N_1695);
nand U3362 (N_3362,N_1774,N_666);
nor U3363 (N_3363,N_906,N_1242);
nand U3364 (N_3364,N_994,N_1857);
and U3365 (N_3365,N_629,N_1311);
and U3366 (N_3366,N_796,N_1931);
nand U3367 (N_3367,N_1792,N_553);
and U3368 (N_3368,N_1016,N_1906);
or U3369 (N_3369,N_269,N_1781);
nor U3370 (N_3370,N_556,N_539);
and U3371 (N_3371,N_1563,N_513);
or U3372 (N_3372,N_6,N_1164);
nand U3373 (N_3373,N_1279,N_1732);
nor U3374 (N_3374,N_1545,N_427);
and U3375 (N_3375,N_1425,N_1355);
and U3376 (N_3376,N_1857,N_1650);
or U3377 (N_3377,N_1179,N_1077);
and U3378 (N_3378,N_1418,N_372);
xnor U3379 (N_3379,N_95,N_1956);
nor U3380 (N_3380,N_1513,N_993);
xor U3381 (N_3381,N_925,N_1095);
nor U3382 (N_3382,N_414,N_483);
nor U3383 (N_3383,N_733,N_1435);
nor U3384 (N_3384,N_1121,N_998);
nor U3385 (N_3385,N_237,N_1758);
or U3386 (N_3386,N_1233,N_1499);
nor U3387 (N_3387,N_1338,N_161);
nor U3388 (N_3388,N_147,N_1037);
or U3389 (N_3389,N_1047,N_394);
and U3390 (N_3390,N_445,N_1548);
and U3391 (N_3391,N_1307,N_530);
and U3392 (N_3392,N_669,N_1933);
and U3393 (N_3393,N_991,N_1098);
nor U3394 (N_3394,N_257,N_103);
nand U3395 (N_3395,N_710,N_368);
or U3396 (N_3396,N_1390,N_1386);
xor U3397 (N_3397,N_103,N_1062);
and U3398 (N_3398,N_472,N_1269);
nor U3399 (N_3399,N_1013,N_185);
xor U3400 (N_3400,N_1608,N_1112);
nand U3401 (N_3401,N_1681,N_1634);
nand U3402 (N_3402,N_44,N_1563);
nand U3403 (N_3403,N_792,N_803);
and U3404 (N_3404,N_283,N_659);
or U3405 (N_3405,N_1686,N_954);
and U3406 (N_3406,N_1501,N_807);
xnor U3407 (N_3407,N_1199,N_828);
xnor U3408 (N_3408,N_852,N_491);
nor U3409 (N_3409,N_1011,N_545);
and U3410 (N_3410,N_1014,N_1747);
or U3411 (N_3411,N_694,N_189);
nand U3412 (N_3412,N_1824,N_438);
and U3413 (N_3413,N_1094,N_1781);
and U3414 (N_3414,N_294,N_1147);
and U3415 (N_3415,N_289,N_1961);
xor U3416 (N_3416,N_1552,N_229);
nand U3417 (N_3417,N_1935,N_1145);
nor U3418 (N_3418,N_1180,N_864);
or U3419 (N_3419,N_1993,N_1835);
nand U3420 (N_3420,N_1092,N_267);
nand U3421 (N_3421,N_1829,N_1600);
nor U3422 (N_3422,N_503,N_1790);
nand U3423 (N_3423,N_941,N_1015);
or U3424 (N_3424,N_1853,N_886);
and U3425 (N_3425,N_777,N_987);
nand U3426 (N_3426,N_258,N_338);
nor U3427 (N_3427,N_1482,N_1002);
nand U3428 (N_3428,N_1169,N_1624);
nor U3429 (N_3429,N_1920,N_932);
nand U3430 (N_3430,N_247,N_1960);
nor U3431 (N_3431,N_35,N_1095);
and U3432 (N_3432,N_1559,N_576);
nand U3433 (N_3433,N_1920,N_214);
or U3434 (N_3434,N_787,N_242);
or U3435 (N_3435,N_1985,N_458);
nor U3436 (N_3436,N_882,N_424);
or U3437 (N_3437,N_1725,N_691);
nor U3438 (N_3438,N_1420,N_1120);
and U3439 (N_3439,N_1304,N_1385);
and U3440 (N_3440,N_1412,N_1580);
or U3441 (N_3441,N_1976,N_870);
and U3442 (N_3442,N_772,N_1150);
or U3443 (N_3443,N_1635,N_1906);
nor U3444 (N_3444,N_1336,N_1730);
nand U3445 (N_3445,N_1193,N_863);
or U3446 (N_3446,N_1505,N_644);
nor U3447 (N_3447,N_1464,N_1078);
nand U3448 (N_3448,N_720,N_331);
nand U3449 (N_3449,N_493,N_1235);
nor U3450 (N_3450,N_1125,N_204);
nand U3451 (N_3451,N_804,N_359);
nand U3452 (N_3452,N_1125,N_1606);
or U3453 (N_3453,N_1988,N_1689);
nor U3454 (N_3454,N_1831,N_655);
nand U3455 (N_3455,N_181,N_738);
or U3456 (N_3456,N_1953,N_547);
nand U3457 (N_3457,N_1987,N_1315);
nor U3458 (N_3458,N_300,N_1603);
nand U3459 (N_3459,N_1742,N_251);
nand U3460 (N_3460,N_1979,N_240);
nand U3461 (N_3461,N_1888,N_1402);
nand U3462 (N_3462,N_1583,N_1611);
or U3463 (N_3463,N_411,N_906);
nor U3464 (N_3464,N_1775,N_986);
xnor U3465 (N_3465,N_9,N_1526);
nand U3466 (N_3466,N_839,N_1832);
nor U3467 (N_3467,N_597,N_1467);
or U3468 (N_3468,N_788,N_794);
or U3469 (N_3469,N_1337,N_1472);
nand U3470 (N_3470,N_1885,N_846);
nand U3471 (N_3471,N_1649,N_590);
or U3472 (N_3472,N_1504,N_600);
nand U3473 (N_3473,N_719,N_1547);
nand U3474 (N_3474,N_1579,N_1117);
and U3475 (N_3475,N_352,N_529);
nand U3476 (N_3476,N_1819,N_1810);
nand U3477 (N_3477,N_1951,N_1244);
and U3478 (N_3478,N_446,N_1177);
and U3479 (N_3479,N_492,N_1041);
or U3480 (N_3480,N_134,N_1931);
xor U3481 (N_3481,N_584,N_1738);
and U3482 (N_3482,N_1794,N_348);
or U3483 (N_3483,N_55,N_727);
xor U3484 (N_3484,N_1527,N_551);
nor U3485 (N_3485,N_1987,N_1114);
nor U3486 (N_3486,N_276,N_1632);
nand U3487 (N_3487,N_1523,N_724);
xnor U3488 (N_3488,N_643,N_1754);
xor U3489 (N_3489,N_275,N_1696);
or U3490 (N_3490,N_540,N_17);
or U3491 (N_3491,N_1474,N_1329);
nand U3492 (N_3492,N_1216,N_1823);
and U3493 (N_3493,N_787,N_229);
nand U3494 (N_3494,N_756,N_1324);
xnor U3495 (N_3495,N_1467,N_621);
or U3496 (N_3496,N_804,N_968);
or U3497 (N_3497,N_1790,N_1099);
xnor U3498 (N_3498,N_94,N_341);
and U3499 (N_3499,N_1730,N_1137);
or U3500 (N_3500,N_1264,N_1440);
nand U3501 (N_3501,N_1290,N_436);
nand U3502 (N_3502,N_758,N_1627);
or U3503 (N_3503,N_723,N_583);
or U3504 (N_3504,N_714,N_100);
nand U3505 (N_3505,N_225,N_1265);
or U3506 (N_3506,N_509,N_266);
nor U3507 (N_3507,N_1018,N_1565);
nor U3508 (N_3508,N_361,N_343);
nor U3509 (N_3509,N_1768,N_300);
nor U3510 (N_3510,N_1148,N_302);
and U3511 (N_3511,N_1752,N_1354);
nand U3512 (N_3512,N_1933,N_354);
nor U3513 (N_3513,N_782,N_1171);
nand U3514 (N_3514,N_782,N_1787);
nand U3515 (N_3515,N_755,N_1078);
or U3516 (N_3516,N_1917,N_315);
and U3517 (N_3517,N_852,N_674);
and U3518 (N_3518,N_305,N_1171);
nand U3519 (N_3519,N_1783,N_1508);
nor U3520 (N_3520,N_1491,N_1269);
nor U3521 (N_3521,N_352,N_1309);
or U3522 (N_3522,N_692,N_1471);
nand U3523 (N_3523,N_1534,N_659);
or U3524 (N_3524,N_125,N_1763);
and U3525 (N_3525,N_1911,N_1386);
and U3526 (N_3526,N_1542,N_1489);
and U3527 (N_3527,N_705,N_1989);
or U3528 (N_3528,N_206,N_970);
or U3529 (N_3529,N_1078,N_954);
nor U3530 (N_3530,N_1508,N_1276);
nand U3531 (N_3531,N_1394,N_1120);
and U3532 (N_3532,N_317,N_1081);
and U3533 (N_3533,N_1671,N_1620);
xnor U3534 (N_3534,N_105,N_1714);
and U3535 (N_3535,N_1459,N_619);
nand U3536 (N_3536,N_472,N_1354);
and U3537 (N_3537,N_1400,N_1884);
nand U3538 (N_3538,N_580,N_1169);
or U3539 (N_3539,N_1724,N_307);
nor U3540 (N_3540,N_409,N_769);
and U3541 (N_3541,N_650,N_31);
nor U3542 (N_3542,N_970,N_1535);
or U3543 (N_3543,N_1837,N_1995);
nor U3544 (N_3544,N_1634,N_1178);
nand U3545 (N_3545,N_1967,N_545);
nor U3546 (N_3546,N_1046,N_1638);
xor U3547 (N_3547,N_643,N_830);
and U3548 (N_3548,N_1201,N_1567);
or U3549 (N_3549,N_856,N_91);
nor U3550 (N_3550,N_581,N_1555);
nand U3551 (N_3551,N_1028,N_1932);
or U3552 (N_3552,N_843,N_1498);
nand U3553 (N_3553,N_809,N_115);
and U3554 (N_3554,N_132,N_834);
or U3555 (N_3555,N_1695,N_1795);
nand U3556 (N_3556,N_738,N_163);
and U3557 (N_3557,N_1176,N_1057);
and U3558 (N_3558,N_769,N_293);
and U3559 (N_3559,N_1886,N_219);
nand U3560 (N_3560,N_367,N_1441);
nand U3561 (N_3561,N_43,N_758);
nand U3562 (N_3562,N_1301,N_358);
nand U3563 (N_3563,N_1065,N_1175);
and U3564 (N_3564,N_160,N_875);
nand U3565 (N_3565,N_1321,N_74);
and U3566 (N_3566,N_30,N_357);
nand U3567 (N_3567,N_1592,N_1517);
nand U3568 (N_3568,N_821,N_1495);
nor U3569 (N_3569,N_750,N_758);
and U3570 (N_3570,N_228,N_1153);
or U3571 (N_3571,N_1922,N_1066);
nand U3572 (N_3572,N_380,N_176);
nor U3573 (N_3573,N_50,N_650);
nand U3574 (N_3574,N_1433,N_137);
and U3575 (N_3575,N_63,N_29);
or U3576 (N_3576,N_1863,N_1307);
nand U3577 (N_3577,N_1064,N_182);
nand U3578 (N_3578,N_453,N_1580);
and U3579 (N_3579,N_992,N_146);
or U3580 (N_3580,N_412,N_639);
or U3581 (N_3581,N_1592,N_51);
nor U3582 (N_3582,N_1851,N_131);
nand U3583 (N_3583,N_483,N_168);
or U3584 (N_3584,N_1485,N_258);
and U3585 (N_3585,N_203,N_709);
or U3586 (N_3586,N_1900,N_1989);
nor U3587 (N_3587,N_1882,N_698);
and U3588 (N_3588,N_555,N_1443);
or U3589 (N_3589,N_1916,N_1922);
nand U3590 (N_3590,N_1553,N_657);
xor U3591 (N_3591,N_388,N_310);
nor U3592 (N_3592,N_1913,N_1045);
and U3593 (N_3593,N_1316,N_972);
nand U3594 (N_3594,N_1102,N_923);
xnor U3595 (N_3595,N_77,N_251);
and U3596 (N_3596,N_321,N_1497);
nor U3597 (N_3597,N_1399,N_660);
or U3598 (N_3598,N_1261,N_686);
nand U3599 (N_3599,N_1178,N_297);
nand U3600 (N_3600,N_1263,N_842);
nand U3601 (N_3601,N_1946,N_944);
nor U3602 (N_3602,N_476,N_57);
or U3603 (N_3603,N_848,N_963);
nor U3604 (N_3604,N_346,N_1051);
and U3605 (N_3605,N_1109,N_702);
and U3606 (N_3606,N_755,N_1137);
nand U3607 (N_3607,N_1746,N_55);
and U3608 (N_3608,N_217,N_1629);
nand U3609 (N_3609,N_1503,N_1288);
nand U3610 (N_3610,N_1851,N_250);
and U3611 (N_3611,N_766,N_628);
or U3612 (N_3612,N_1358,N_1969);
nand U3613 (N_3613,N_559,N_269);
or U3614 (N_3614,N_1693,N_1209);
and U3615 (N_3615,N_1745,N_1396);
xor U3616 (N_3616,N_738,N_91);
nor U3617 (N_3617,N_1877,N_1715);
nand U3618 (N_3618,N_755,N_530);
and U3619 (N_3619,N_1759,N_248);
nor U3620 (N_3620,N_693,N_553);
and U3621 (N_3621,N_609,N_1939);
or U3622 (N_3622,N_912,N_1106);
nor U3623 (N_3623,N_1902,N_593);
nand U3624 (N_3624,N_1390,N_958);
nand U3625 (N_3625,N_1892,N_662);
nand U3626 (N_3626,N_184,N_872);
nand U3627 (N_3627,N_775,N_977);
nand U3628 (N_3628,N_1950,N_229);
nor U3629 (N_3629,N_238,N_1263);
nor U3630 (N_3630,N_293,N_1978);
or U3631 (N_3631,N_1382,N_223);
and U3632 (N_3632,N_1380,N_617);
and U3633 (N_3633,N_893,N_1293);
nand U3634 (N_3634,N_1921,N_1318);
nand U3635 (N_3635,N_990,N_1471);
and U3636 (N_3636,N_1632,N_1013);
xnor U3637 (N_3637,N_619,N_414);
nand U3638 (N_3638,N_1434,N_951);
or U3639 (N_3639,N_529,N_1236);
nor U3640 (N_3640,N_589,N_876);
or U3641 (N_3641,N_1662,N_1596);
xnor U3642 (N_3642,N_724,N_1401);
and U3643 (N_3643,N_1029,N_1346);
nor U3644 (N_3644,N_1410,N_832);
nor U3645 (N_3645,N_1966,N_1410);
nor U3646 (N_3646,N_76,N_275);
nor U3647 (N_3647,N_1836,N_586);
nand U3648 (N_3648,N_243,N_599);
nor U3649 (N_3649,N_1040,N_183);
nand U3650 (N_3650,N_631,N_1336);
and U3651 (N_3651,N_732,N_1314);
and U3652 (N_3652,N_511,N_129);
nand U3653 (N_3653,N_139,N_345);
nand U3654 (N_3654,N_1955,N_682);
xnor U3655 (N_3655,N_466,N_1495);
xor U3656 (N_3656,N_1629,N_121);
nand U3657 (N_3657,N_1159,N_190);
xor U3658 (N_3658,N_582,N_367);
nor U3659 (N_3659,N_31,N_1838);
nor U3660 (N_3660,N_1618,N_1422);
xnor U3661 (N_3661,N_718,N_1705);
nand U3662 (N_3662,N_9,N_246);
or U3663 (N_3663,N_344,N_182);
nor U3664 (N_3664,N_1646,N_400);
xor U3665 (N_3665,N_1872,N_920);
and U3666 (N_3666,N_565,N_746);
nor U3667 (N_3667,N_1197,N_685);
nand U3668 (N_3668,N_1542,N_248);
xnor U3669 (N_3669,N_753,N_1684);
nand U3670 (N_3670,N_1406,N_14);
xnor U3671 (N_3671,N_1009,N_44);
nand U3672 (N_3672,N_1959,N_1522);
nor U3673 (N_3673,N_5,N_767);
or U3674 (N_3674,N_1171,N_831);
xor U3675 (N_3675,N_790,N_624);
or U3676 (N_3676,N_1813,N_946);
nor U3677 (N_3677,N_1208,N_22);
or U3678 (N_3678,N_153,N_398);
xor U3679 (N_3679,N_1993,N_748);
nor U3680 (N_3680,N_317,N_278);
and U3681 (N_3681,N_1010,N_749);
and U3682 (N_3682,N_1351,N_1211);
nor U3683 (N_3683,N_851,N_904);
and U3684 (N_3684,N_1098,N_610);
nand U3685 (N_3685,N_880,N_1698);
xnor U3686 (N_3686,N_945,N_1652);
xor U3687 (N_3687,N_1553,N_1281);
nand U3688 (N_3688,N_587,N_1885);
nor U3689 (N_3689,N_410,N_803);
and U3690 (N_3690,N_201,N_460);
or U3691 (N_3691,N_1542,N_1831);
and U3692 (N_3692,N_178,N_80);
xor U3693 (N_3693,N_255,N_1998);
or U3694 (N_3694,N_1146,N_1626);
xor U3695 (N_3695,N_166,N_865);
nand U3696 (N_3696,N_1483,N_170);
and U3697 (N_3697,N_645,N_552);
and U3698 (N_3698,N_11,N_701);
nand U3699 (N_3699,N_1136,N_1459);
xnor U3700 (N_3700,N_514,N_644);
nor U3701 (N_3701,N_751,N_646);
or U3702 (N_3702,N_1192,N_1166);
xnor U3703 (N_3703,N_1578,N_281);
or U3704 (N_3704,N_645,N_306);
or U3705 (N_3705,N_1314,N_1476);
and U3706 (N_3706,N_984,N_845);
and U3707 (N_3707,N_1713,N_1819);
or U3708 (N_3708,N_167,N_421);
nor U3709 (N_3709,N_324,N_1858);
or U3710 (N_3710,N_1083,N_1563);
nor U3711 (N_3711,N_1998,N_377);
or U3712 (N_3712,N_1688,N_705);
nand U3713 (N_3713,N_393,N_1856);
and U3714 (N_3714,N_1657,N_1905);
and U3715 (N_3715,N_993,N_1214);
nor U3716 (N_3716,N_1269,N_713);
and U3717 (N_3717,N_1865,N_578);
or U3718 (N_3718,N_1931,N_1514);
nor U3719 (N_3719,N_1807,N_639);
nor U3720 (N_3720,N_1374,N_1074);
or U3721 (N_3721,N_792,N_199);
and U3722 (N_3722,N_535,N_538);
xnor U3723 (N_3723,N_1886,N_1839);
nand U3724 (N_3724,N_1150,N_1050);
and U3725 (N_3725,N_913,N_1532);
and U3726 (N_3726,N_1375,N_811);
xnor U3727 (N_3727,N_323,N_1756);
nand U3728 (N_3728,N_106,N_712);
nand U3729 (N_3729,N_1364,N_1217);
and U3730 (N_3730,N_334,N_1449);
or U3731 (N_3731,N_97,N_798);
or U3732 (N_3732,N_1779,N_271);
or U3733 (N_3733,N_519,N_1714);
and U3734 (N_3734,N_789,N_1689);
nand U3735 (N_3735,N_1956,N_736);
nor U3736 (N_3736,N_349,N_457);
and U3737 (N_3737,N_1524,N_87);
and U3738 (N_3738,N_1685,N_1434);
nor U3739 (N_3739,N_1409,N_1732);
and U3740 (N_3740,N_1648,N_1049);
xnor U3741 (N_3741,N_1162,N_1563);
nor U3742 (N_3742,N_606,N_232);
or U3743 (N_3743,N_1082,N_1327);
nand U3744 (N_3744,N_1825,N_262);
or U3745 (N_3745,N_1038,N_113);
xor U3746 (N_3746,N_368,N_851);
and U3747 (N_3747,N_1864,N_722);
and U3748 (N_3748,N_90,N_508);
nand U3749 (N_3749,N_1554,N_423);
or U3750 (N_3750,N_1124,N_1345);
or U3751 (N_3751,N_1704,N_188);
or U3752 (N_3752,N_145,N_590);
and U3753 (N_3753,N_1594,N_1050);
or U3754 (N_3754,N_1321,N_389);
xnor U3755 (N_3755,N_18,N_1464);
xor U3756 (N_3756,N_1381,N_1674);
nor U3757 (N_3757,N_1066,N_1743);
and U3758 (N_3758,N_627,N_842);
nand U3759 (N_3759,N_617,N_447);
and U3760 (N_3760,N_1841,N_1700);
nor U3761 (N_3761,N_326,N_573);
nand U3762 (N_3762,N_284,N_883);
nor U3763 (N_3763,N_1419,N_1507);
nand U3764 (N_3764,N_1686,N_518);
xor U3765 (N_3765,N_4,N_945);
or U3766 (N_3766,N_1406,N_516);
nand U3767 (N_3767,N_1442,N_809);
and U3768 (N_3768,N_1196,N_878);
and U3769 (N_3769,N_1789,N_1705);
or U3770 (N_3770,N_1370,N_1103);
nand U3771 (N_3771,N_1111,N_1134);
or U3772 (N_3772,N_566,N_292);
nand U3773 (N_3773,N_680,N_278);
or U3774 (N_3774,N_871,N_965);
nand U3775 (N_3775,N_1827,N_835);
nor U3776 (N_3776,N_935,N_398);
or U3777 (N_3777,N_1252,N_315);
and U3778 (N_3778,N_631,N_1582);
or U3779 (N_3779,N_312,N_1278);
nand U3780 (N_3780,N_84,N_1753);
and U3781 (N_3781,N_1169,N_1433);
and U3782 (N_3782,N_1844,N_689);
nand U3783 (N_3783,N_1421,N_501);
nor U3784 (N_3784,N_304,N_1160);
and U3785 (N_3785,N_1329,N_1216);
xnor U3786 (N_3786,N_438,N_677);
nand U3787 (N_3787,N_257,N_957);
xnor U3788 (N_3788,N_1160,N_134);
xnor U3789 (N_3789,N_1828,N_1385);
nand U3790 (N_3790,N_954,N_850);
nand U3791 (N_3791,N_478,N_1345);
and U3792 (N_3792,N_422,N_1242);
nand U3793 (N_3793,N_879,N_182);
and U3794 (N_3794,N_952,N_1881);
and U3795 (N_3795,N_381,N_0);
and U3796 (N_3796,N_1914,N_129);
nand U3797 (N_3797,N_1255,N_1412);
nor U3798 (N_3798,N_1114,N_687);
and U3799 (N_3799,N_1826,N_934);
or U3800 (N_3800,N_1634,N_1738);
nand U3801 (N_3801,N_1251,N_1);
and U3802 (N_3802,N_475,N_143);
nor U3803 (N_3803,N_1041,N_643);
and U3804 (N_3804,N_619,N_1708);
and U3805 (N_3805,N_222,N_1381);
or U3806 (N_3806,N_1081,N_502);
nand U3807 (N_3807,N_815,N_1405);
xor U3808 (N_3808,N_350,N_845);
or U3809 (N_3809,N_1319,N_1600);
nor U3810 (N_3810,N_816,N_1939);
nor U3811 (N_3811,N_1626,N_1177);
nand U3812 (N_3812,N_687,N_330);
nor U3813 (N_3813,N_1817,N_638);
nor U3814 (N_3814,N_984,N_1180);
nor U3815 (N_3815,N_412,N_1151);
or U3816 (N_3816,N_604,N_1145);
nor U3817 (N_3817,N_1917,N_466);
and U3818 (N_3818,N_740,N_310);
nor U3819 (N_3819,N_146,N_565);
and U3820 (N_3820,N_1248,N_809);
nor U3821 (N_3821,N_1238,N_1316);
xor U3822 (N_3822,N_1789,N_1584);
nand U3823 (N_3823,N_1780,N_1192);
or U3824 (N_3824,N_938,N_1044);
nand U3825 (N_3825,N_1615,N_656);
and U3826 (N_3826,N_1936,N_1978);
xor U3827 (N_3827,N_743,N_1519);
nor U3828 (N_3828,N_1077,N_443);
xor U3829 (N_3829,N_903,N_1350);
nor U3830 (N_3830,N_913,N_1087);
nand U3831 (N_3831,N_1257,N_1875);
or U3832 (N_3832,N_529,N_777);
and U3833 (N_3833,N_1527,N_1683);
or U3834 (N_3834,N_512,N_1965);
nand U3835 (N_3835,N_1340,N_953);
nor U3836 (N_3836,N_1329,N_784);
nor U3837 (N_3837,N_939,N_1909);
nor U3838 (N_3838,N_1866,N_1801);
xnor U3839 (N_3839,N_419,N_1408);
and U3840 (N_3840,N_1826,N_545);
or U3841 (N_3841,N_29,N_1143);
and U3842 (N_3842,N_861,N_905);
and U3843 (N_3843,N_1397,N_1930);
and U3844 (N_3844,N_1349,N_1225);
nand U3845 (N_3845,N_1195,N_845);
and U3846 (N_3846,N_606,N_1653);
nand U3847 (N_3847,N_685,N_1976);
or U3848 (N_3848,N_201,N_1775);
nor U3849 (N_3849,N_1535,N_693);
nor U3850 (N_3850,N_764,N_1209);
or U3851 (N_3851,N_1659,N_121);
nand U3852 (N_3852,N_1806,N_1638);
nor U3853 (N_3853,N_1374,N_1354);
and U3854 (N_3854,N_1402,N_403);
nand U3855 (N_3855,N_1690,N_126);
or U3856 (N_3856,N_1251,N_1280);
nor U3857 (N_3857,N_1957,N_1647);
nand U3858 (N_3858,N_476,N_1691);
or U3859 (N_3859,N_255,N_75);
and U3860 (N_3860,N_1815,N_31);
and U3861 (N_3861,N_1037,N_248);
xor U3862 (N_3862,N_702,N_1760);
or U3863 (N_3863,N_1929,N_1008);
nor U3864 (N_3864,N_1715,N_400);
nor U3865 (N_3865,N_633,N_1431);
xnor U3866 (N_3866,N_279,N_27);
nand U3867 (N_3867,N_291,N_1105);
nand U3868 (N_3868,N_134,N_1263);
nor U3869 (N_3869,N_1025,N_1333);
xor U3870 (N_3870,N_344,N_1884);
and U3871 (N_3871,N_67,N_1711);
or U3872 (N_3872,N_1031,N_172);
and U3873 (N_3873,N_376,N_664);
or U3874 (N_3874,N_547,N_1532);
nand U3875 (N_3875,N_1579,N_780);
and U3876 (N_3876,N_880,N_1284);
and U3877 (N_3877,N_709,N_107);
nand U3878 (N_3878,N_1849,N_1203);
and U3879 (N_3879,N_1947,N_846);
and U3880 (N_3880,N_581,N_1238);
or U3881 (N_3881,N_965,N_818);
xnor U3882 (N_3882,N_26,N_1228);
and U3883 (N_3883,N_929,N_318);
or U3884 (N_3884,N_1397,N_315);
or U3885 (N_3885,N_1276,N_1495);
nor U3886 (N_3886,N_934,N_1389);
or U3887 (N_3887,N_347,N_318);
and U3888 (N_3888,N_1552,N_1475);
or U3889 (N_3889,N_707,N_1458);
and U3890 (N_3890,N_886,N_1549);
and U3891 (N_3891,N_1860,N_1067);
and U3892 (N_3892,N_822,N_1174);
xnor U3893 (N_3893,N_535,N_1878);
nand U3894 (N_3894,N_1687,N_634);
and U3895 (N_3895,N_1349,N_1297);
nor U3896 (N_3896,N_879,N_1801);
and U3897 (N_3897,N_18,N_1076);
xor U3898 (N_3898,N_1283,N_964);
nand U3899 (N_3899,N_804,N_14);
or U3900 (N_3900,N_447,N_565);
xor U3901 (N_3901,N_1253,N_1010);
or U3902 (N_3902,N_857,N_1982);
nor U3903 (N_3903,N_385,N_371);
and U3904 (N_3904,N_1611,N_654);
and U3905 (N_3905,N_344,N_580);
xnor U3906 (N_3906,N_586,N_1483);
nor U3907 (N_3907,N_859,N_1958);
or U3908 (N_3908,N_804,N_806);
nand U3909 (N_3909,N_1734,N_372);
nand U3910 (N_3910,N_1656,N_1436);
and U3911 (N_3911,N_368,N_71);
nand U3912 (N_3912,N_632,N_796);
and U3913 (N_3913,N_1311,N_1495);
nand U3914 (N_3914,N_1576,N_1594);
nor U3915 (N_3915,N_1586,N_1000);
or U3916 (N_3916,N_902,N_949);
nor U3917 (N_3917,N_1907,N_932);
or U3918 (N_3918,N_874,N_1877);
or U3919 (N_3919,N_1954,N_1912);
nand U3920 (N_3920,N_1925,N_1120);
or U3921 (N_3921,N_875,N_1052);
nor U3922 (N_3922,N_1925,N_626);
nand U3923 (N_3923,N_639,N_1397);
or U3924 (N_3924,N_188,N_584);
xor U3925 (N_3925,N_1640,N_1669);
nor U3926 (N_3926,N_168,N_414);
nor U3927 (N_3927,N_1412,N_557);
and U3928 (N_3928,N_574,N_902);
nor U3929 (N_3929,N_1974,N_457);
or U3930 (N_3930,N_1546,N_1831);
nor U3931 (N_3931,N_882,N_1079);
nand U3932 (N_3932,N_1878,N_505);
and U3933 (N_3933,N_1350,N_1617);
and U3934 (N_3934,N_481,N_1308);
or U3935 (N_3935,N_1410,N_409);
xor U3936 (N_3936,N_712,N_1760);
or U3937 (N_3937,N_1690,N_1905);
or U3938 (N_3938,N_542,N_1777);
xor U3939 (N_3939,N_1918,N_1283);
and U3940 (N_3940,N_1294,N_1586);
or U3941 (N_3941,N_1063,N_539);
and U3942 (N_3942,N_1271,N_137);
and U3943 (N_3943,N_1037,N_1243);
nand U3944 (N_3944,N_503,N_746);
and U3945 (N_3945,N_189,N_1188);
and U3946 (N_3946,N_688,N_1783);
nor U3947 (N_3947,N_935,N_1381);
and U3948 (N_3948,N_1969,N_564);
xor U3949 (N_3949,N_1687,N_421);
nor U3950 (N_3950,N_1454,N_34);
and U3951 (N_3951,N_344,N_471);
nand U3952 (N_3952,N_897,N_732);
nand U3953 (N_3953,N_207,N_1302);
xnor U3954 (N_3954,N_1393,N_1992);
nor U3955 (N_3955,N_1145,N_550);
and U3956 (N_3956,N_1954,N_134);
or U3957 (N_3957,N_1241,N_1691);
or U3958 (N_3958,N_534,N_1647);
or U3959 (N_3959,N_1578,N_1182);
and U3960 (N_3960,N_908,N_1195);
nor U3961 (N_3961,N_123,N_1042);
or U3962 (N_3962,N_622,N_621);
xor U3963 (N_3963,N_1960,N_437);
nand U3964 (N_3964,N_1472,N_731);
xor U3965 (N_3965,N_1044,N_1328);
and U3966 (N_3966,N_563,N_217);
or U3967 (N_3967,N_72,N_1886);
and U3968 (N_3968,N_1531,N_1645);
and U3969 (N_3969,N_1532,N_1521);
xor U3970 (N_3970,N_1673,N_1136);
and U3971 (N_3971,N_1319,N_867);
nor U3972 (N_3972,N_1762,N_824);
nor U3973 (N_3973,N_1143,N_1494);
nor U3974 (N_3974,N_1509,N_1022);
or U3975 (N_3975,N_1766,N_702);
xor U3976 (N_3976,N_1584,N_1136);
nand U3977 (N_3977,N_1354,N_916);
nor U3978 (N_3978,N_252,N_197);
nor U3979 (N_3979,N_967,N_558);
and U3980 (N_3980,N_950,N_1230);
xnor U3981 (N_3981,N_556,N_1289);
nand U3982 (N_3982,N_1347,N_1619);
nor U3983 (N_3983,N_1886,N_445);
or U3984 (N_3984,N_460,N_892);
xnor U3985 (N_3985,N_1643,N_1068);
or U3986 (N_3986,N_241,N_1677);
nand U3987 (N_3987,N_407,N_609);
or U3988 (N_3988,N_499,N_679);
nand U3989 (N_3989,N_984,N_541);
or U3990 (N_3990,N_565,N_1782);
and U3991 (N_3991,N_924,N_1561);
and U3992 (N_3992,N_1641,N_1502);
nand U3993 (N_3993,N_1523,N_500);
nand U3994 (N_3994,N_15,N_147);
xor U3995 (N_3995,N_189,N_150);
or U3996 (N_3996,N_1437,N_896);
or U3997 (N_3997,N_627,N_1612);
nor U3998 (N_3998,N_1597,N_598);
nor U3999 (N_3999,N_846,N_844);
and U4000 (N_4000,N_2233,N_3042);
nand U4001 (N_4001,N_3555,N_3581);
nor U4002 (N_4002,N_2697,N_2553);
or U4003 (N_4003,N_2991,N_2170);
nand U4004 (N_4004,N_2773,N_2192);
nand U4005 (N_4005,N_3604,N_2625);
and U4006 (N_4006,N_3586,N_3423);
xor U4007 (N_4007,N_2535,N_2031);
or U4008 (N_4008,N_2498,N_2672);
xnor U4009 (N_4009,N_3336,N_2075);
xnor U4010 (N_4010,N_2750,N_3598);
and U4011 (N_4011,N_3808,N_2585);
or U4012 (N_4012,N_3457,N_2935);
or U4013 (N_4013,N_2774,N_3637);
or U4014 (N_4014,N_3727,N_3825);
and U4015 (N_4015,N_3146,N_2199);
or U4016 (N_4016,N_3843,N_3588);
or U4017 (N_4017,N_3814,N_2456);
nand U4018 (N_4018,N_3323,N_3160);
nand U4019 (N_4019,N_2307,N_3383);
xnor U4020 (N_4020,N_3246,N_2156);
nand U4021 (N_4021,N_3815,N_3389);
nand U4022 (N_4022,N_3216,N_2927);
and U4023 (N_4023,N_2510,N_3713);
nor U4024 (N_4024,N_3027,N_2355);
nor U4025 (N_4025,N_2589,N_3969);
and U4026 (N_4026,N_3528,N_3517);
and U4027 (N_4027,N_2926,N_2058);
xor U4028 (N_4028,N_3872,N_2978);
nand U4029 (N_4029,N_3023,N_3724);
or U4030 (N_4030,N_2993,N_2753);
xor U4031 (N_4031,N_2896,N_3072);
nand U4032 (N_4032,N_3626,N_2719);
and U4033 (N_4033,N_2410,N_3290);
nor U4034 (N_4034,N_3335,N_3572);
and U4035 (N_4035,N_2570,N_3445);
nor U4036 (N_4036,N_2173,N_3823);
and U4037 (N_4037,N_3178,N_3696);
nand U4038 (N_4038,N_3175,N_2558);
xnor U4039 (N_4039,N_3341,N_2998);
or U4040 (N_4040,N_3931,N_2447);
xor U4041 (N_4041,N_2465,N_3968);
or U4042 (N_4042,N_3653,N_2344);
nand U4043 (N_4043,N_2047,N_2886);
or U4044 (N_4044,N_2113,N_2827);
and U4045 (N_4045,N_3213,N_2651);
nand U4046 (N_4046,N_3743,N_3046);
nand U4047 (N_4047,N_3575,N_3422);
and U4048 (N_4048,N_3390,N_3397);
or U4049 (N_4049,N_2963,N_2612);
nand U4050 (N_4050,N_3613,N_3244);
or U4051 (N_4051,N_3418,N_2483);
nor U4052 (N_4052,N_3742,N_3537);
xnor U4053 (N_4053,N_2791,N_2360);
and U4054 (N_4054,N_2038,N_2150);
nand U4055 (N_4055,N_2761,N_2540);
and U4056 (N_4056,N_2775,N_2841);
or U4057 (N_4057,N_3894,N_2862);
nand U4058 (N_4058,N_3812,N_3120);
or U4059 (N_4059,N_2563,N_2627);
and U4060 (N_4060,N_3097,N_2283);
or U4061 (N_4061,N_3601,N_2736);
or U4062 (N_4062,N_3911,N_3276);
and U4063 (N_4063,N_3171,N_2337);
nand U4064 (N_4064,N_2892,N_2953);
nor U4065 (N_4065,N_3811,N_3631);
and U4066 (N_4066,N_2033,N_2083);
xor U4067 (N_4067,N_3589,N_3786);
nand U4068 (N_4068,N_2036,N_3067);
or U4069 (N_4069,N_3753,N_3229);
or U4070 (N_4070,N_2019,N_3452);
xor U4071 (N_4071,N_2421,N_2347);
or U4072 (N_4072,N_3086,N_3669);
nand U4073 (N_4073,N_3334,N_3510);
nor U4074 (N_4074,N_2388,N_2390);
nand U4075 (N_4075,N_2029,N_2583);
and U4076 (N_4076,N_3520,N_3647);
or U4077 (N_4077,N_3313,N_2037);
or U4078 (N_4078,N_3848,N_3711);
and U4079 (N_4079,N_2802,N_3775);
xnor U4080 (N_4080,N_2165,N_3278);
xnor U4081 (N_4081,N_2155,N_3132);
or U4082 (N_4082,N_3627,N_2505);
or U4083 (N_4083,N_3788,N_2757);
nor U4084 (N_4084,N_2710,N_3990);
xor U4085 (N_4085,N_2392,N_3664);
nor U4086 (N_4086,N_3258,N_2845);
nor U4087 (N_4087,N_3773,N_3438);
and U4088 (N_4088,N_2454,N_2275);
or U4089 (N_4089,N_2222,N_2232);
nor U4090 (N_4090,N_2228,N_2414);
nor U4091 (N_4091,N_3933,N_3944);
or U4092 (N_4092,N_2093,N_2383);
or U4093 (N_4093,N_3054,N_3487);
and U4094 (N_4094,N_3230,N_2471);
nand U4095 (N_4095,N_3243,N_2277);
nor U4096 (N_4096,N_3283,N_3154);
or U4097 (N_4097,N_3509,N_3137);
nand U4098 (N_4098,N_3964,N_3237);
xor U4099 (N_4099,N_3500,N_2145);
and U4100 (N_4100,N_3180,N_2833);
nor U4101 (N_4101,N_3385,N_2618);
nand U4102 (N_4102,N_3095,N_2151);
nand U4103 (N_4103,N_2399,N_3900);
and U4104 (N_4104,N_3411,N_3011);
nor U4105 (N_4105,N_2106,N_2603);
nand U4106 (N_4106,N_3570,N_2330);
nand U4107 (N_4107,N_2634,N_2091);
xnor U4108 (N_4108,N_3923,N_3311);
nand U4109 (N_4109,N_3856,N_3725);
and U4110 (N_4110,N_3198,N_3710);
nor U4111 (N_4111,N_2180,N_2605);
nor U4112 (N_4112,N_2039,N_3646);
nand U4113 (N_4113,N_3462,N_3017);
xor U4114 (N_4114,N_2329,N_3899);
and U4115 (N_4115,N_3443,N_3057);
and U4116 (N_4116,N_3936,N_2321);
nor U4117 (N_4117,N_2726,N_3407);
nor U4118 (N_4118,N_3236,N_2667);
xnor U4119 (N_4119,N_3060,N_2954);
or U4120 (N_4120,N_3794,N_3369);
and U4121 (N_4121,N_2082,N_3671);
xor U4122 (N_4122,N_2599,N_3878);
nand U4123 (N_4123,N_2663,N_3408);
nand U4124 (N_4124,N_3922,N_3015);
nor U4125 (N_4125,N_2482,N_2185);
or U4126 (N_4126,N_3153,N_3701);
and U4127 (N_4127,N_2767,N_3202);
and U4128 (N_4128,N_3567,N_3116);
or U4129 (N_4129,N_2137,N_2308);
and U4130 (N_4130,N_3376,N_2121);
and U4131 (N_4131,N_2818,N_2322);
nor U4132 (N_4132,N_2533,N_3263);
nor U4133 (N_4133,N_2512,N_3281);
nor U4134 (N_4134,N_3368,N_2765);
or U4135 (N_4135,N_3639,N_3974);
or U4136 (N_4136,N_3692,N_3486);
and U4137 (N_4137,N_3558,N_2947);
and U4138 (N_4138,N_2287,N_3616);
nor U4139 (N_4139,N_3867,N_3988);
nand U4140 (N_4140,N_2919,N_3442);
or U4141 (N_4141,N_2879,N_3542);
nand U4142 (N_4142,N_2100,N_2218);
nand U4143 (N_4143,N_3096,N_3420);
nand U4144 (N_4144,N_3667,N_2629);
and U4145 (N_4145,N_2450,N_2851);
or U4146 (N_4146,N_3354,N_2934);
or U4147 (N_4147,N_3952,N_3652);
nand U4148 (N_4148,N_3758,N_3644);
nor U4149 (N_4149,N_2890,N_2402);
nor U4150 (N_4150,N_2056,N_2653);
nor U4151 (N_4151,N_3591,N_3429);
and U4152 (N_4152,N_3037,N_2366);
or U4153 (N_4153,N_2692,N_2472);
nor U4154 (N_4154,N_2468,N_3987);
nor U4155 (N_4155,N_2965,N_2861);
or U4156 (N_4156,N_2486,N_2844);
or U4157 (N_4157,N_3849,N_2497);
nand U4158 (N_4158,N_2986,N_2217);
and U4159 (N_4159,N_3630,N_3184);
nand U4160 (N_4160,N_2898,N_2276);
and U4161 (N_4161,N_2616,N_3951);
nand U4162 (N_4162,N_3884,N_2839);
or U4163 (N_4163,N_3564,N_3228);
xnor U4164 (N_4164,N_2361,N_2557);
or U4165 (N_4165,N_2593,N_2243);
nand U4166 (N_4166,N_2123,N_2567);
xor U4167 (N_4167,N_3139,N_3499);
xor U4168 (N_4168,N_3063,N_3114);
xnor U4169 (N_4169,N_2708,N_3308);
nand U4170 (N_4170,N_3195,N_2258);
nor U4171 (N_4171,N_2054,N_3085);
and U4172 (N_4172,N_3506,N_3032);
and U4173 (N_4173,N_3553,N_3401);
nand U4174 (N_4174,N_3359,N_3001);
xor U4175 (N_4175,N_2732,N_3847);
nand U4176 (N_4176,N_2746,N_3870);
nand U4177 (N_4177,N_2958,N_3650);
or U4178 (N_4178,N_3388,N_3491);
nand U4179 (N_4179,N_2664,N_3746);
nor U4180 (N_4180,N_3417,N_3677);
or U4181 (N_4181,N_2020,N_3285);
nor U4182 (N_4182,N_2216,N_3972);
nand U4183 (N_4183,N_2398,N_3208);
nor U4184 (N_4184,N_3051,N_2528);
nand U4185 (N_4185,N_3778,N_2256);
or U4186 (N_4186,N_2395,N_3143);
xnor U4187 (N_4187,N_2574,N_3993);
or U4188 (N_4188,N_3822,N_2577);
and U4189 (N_4189,N_2000,N_2050);
nand U4190 (N_4190,N_3535,N_3709);
and U4191 (N_4191,N_2828,N_3522);
nor U4192 (N_4192,N_3059,N_2354);
or U4193 (N_4193,N_3594,N_2067);
nor U4194 (N_4194,N_2242,N_3482);
and U4195 (N_4195,N_3934,N_2795);
or U4196 (N_4196,N_2555,N_3241);
nand U4197 (N_4197,N_3862,N_2200);
nor U4198 (N_4198,N_3844,N_3938);
or U4199 (N_4199,N_2077,N_3190);
nand U4200 (N_4200,N_3309,N_3102);
and U4201 (N_4201,N_3127,N_2901);
or U4202 (N_4202,N_3157,N_2566);
xor U4203 (N_4203,N_3955,N_3306);
or U4204 (N_4204,N_2336,N_2872);
and U4205 (N_4205,N_2670,N_3013);
nand U4206 (N_4206,N_3685,N_2545);
or U4207 (N_4207,N_2431,N_3947);
xor U4208 (N_4208,N_2842,N_3882);
or U4209 (N_4209,N_2720,N_2460);
nand U4210 (N_4210,N_3248,N_3905);
xor U4211 (N_4211,N_3170,N_2702);
or U4212 (N_4212,N_2473,N_3764);
and U4213 (N_4213,N_3571,N_2184);
nor U4214 (N_4214,N_2314,N_3574);
nand U4215 (N_4215,N_2956,N_2476);
and U4216 (N_4216,N_2952,N_2126);
or U4217 (N_4217,N_2849,N_3371);
nor U4218 (N_4218,N_3859,N_3643);
nand U4219 (N_4219,N_2789,N_3966);
or U4220 (N_4220,N_2023,N_3118);
and U4221 (N_4221,N_3694,N_3769);
nand U4222 (N_4222,N_3437,N_3210);
nor U4223 (N_4223,N_2974,N_3525);
and U4224 (N_4224,N_3141,N_2193);
xnor U4225 (N_4225,N_3480,N_3759);
and U4226 (N_4226,N_2318,N_2229);
or U4227 (N_4227,N_2763,N_2244);
nand U4228 (N_4228,N_3728,N_3681);
xor U4229 (N_4229,N_3793,N_3386);
or U4230 (N_4230,N_2724,N_3400);
nand U4231 (N_4231,N_2022,N_2440);
nor U4232 (N_4232,N_3559,N_2111);
nand U4233 (N_4233,N_2970,N_3286);
and U4234 (N_4234,N_3274,N_3332);
nand U4235 (N_4235,N_2040,N_2300);
nor U4236 (N_4236,N_3994,N_3062);
xnor U4237 (N_4237,N_2906,N_2120);
nor U4238 (N_4238,N_3860,N_2230);
nand U4239 (N_4239,N_2401,N_3857);
and U4240 (N_4240,N_2536,N_3469);
xor U4241 (N_4241,N_2679,N_2542);
nor U4242 (N_4242,N_2976,N_2334);
or U4243 (N_4243,N_3165,N_2012);
and U4244 (N_4244,N_2573,N_3618);
or U4245 (N_4245,N_2643,N_2508);
or U4246 (N_4246,N_3045,N_3456);
or U4247 (N_4247,N_2061,N_2899);
or U4248 (N_4248,N_3151,N_2264);
and U4249 (N_4249,N_2289,N_2135);
and U4250 (N_4250,N_3777,N_3804);
or U4251 (N_4251,N_2266,N_2358);
and U4252 (N_4252,N_2490,N_3686);
nand U4253 (N_4253,N_2615,N_2018);
nor U4254 (N_4254,N_3737,N_2208);
or U4255 (N_4255,N_3942,N_3748);
and U4256 (N_4256,N_3126,N_2403);
or U4257 (N_4257,N_2857,N_3043);
nor U4258 (N_4258,N_3414,N_3784);
nand U4259 (N_4259,N_3239,N_2118);
nand U4260 (N_4260,N_3318,N_2335);
nor U4261 (N_4261,N_3958,N_3049);
nand U4262 (N_4262,N_3349,N_2798);
nand U4263 (N_4263,N_2804,N_3055);
nor U4264 (N_4264,N_3465,N_3698);
and U4265 (N_4265,N_2560,N_2794);
nand U4266 (N_4266,N_2130,N_3463);
and U4267 (N_4267,N_2831,N_3744);
and U4268 (N_4268,N_2698,N_2214);
nand U4269 (N_4269,N_2522,N_3619);
nor U4270 (N_4270,N_2734,N_2983);
nor U4271 (N_4271,N_2412,N_3582);
or U4272 (N_4272,N_2235,N_2187);
nand U4273 (N_4273,N_3625,N_3679);
nor U4274 (N_4274,N_3003,N_3221);
or U4275 (N_4275,N_2425,N_2371);
nand U4276 (N_4276,N_2640,N_2092);
and U4277 (N_4277,N_2723,N_2838);
and U4278 (N_4278,N_2600,N_3762);
xnor U4279 (N_4279,N_3367,N_2253);
and U4280 (N_4280,N_2587,N_3756);
or U4281 (N_4281,N_2396,N_3666);
nand U4282 (N_4282,N_3519,N_2149);
nand U4283 (N_4283,N_3834,N_3430);
nand U4284 (N_4284,N_2325,N_2727);
and U4285 (N_4285,N_3384,N_2715);
or U4286 (N_4286,N_2808,N_3563);
or U4287 (N_4287,N_2850,N_2772);
nand U4288 (N_4288,N_3215,N_3076);
and U4289 (N_4289,N_2144,N_3755);
nand U4290 (N_4290,N_2094,N_2237);
nor U4291 (N_4291,N_2680,N_2086);
xor U4292 (N_4292,N_2999,N_2864);
nand U4293 (N_4293,N_3416,N_3092);
nand U4294 (N_4294,N_3629,N_3088);
or U4295 (N_4295,N_3640,N_3344);
xnor U4296 (N_4296,N_2282,N_3837);
nor U4297 (N_4297,N_2929,N_3110);
nand U4298 (N_4298,N_2768,N_3431);
or U4299 (N_4299,N_2532,N_3148);
and U4300 (N_4300,N_3730,N_3739);
xor U4301 (N_4301,N_2960,N_2738);
or U4302 (N_4302,N_3454,N_3568);
or U4303 (N_4303,N_2099,N_3339);
and U4304 (N_4304,N_3250,N_3780);
xnor U4305 (N_4305,N_3655,N_3026);
and U4306 (N_4306,N_3223,N_3317);
nor U4307 (N_4307,N_3828,N_3378);
nand U4308 (N_4308,N_3635,N_3470);
and U4309 (N_4309,N_3172,N_2779);
xor U4310 (N_4310,N_3122,N_3119);
nor U4311 (N_4311,N_2493,N_2231);
nor U4312 (N_4312,N_3982,N_3918);
nand U4313 (N_4313,N_2327,N_3464);
and U4314 (N_4314,N_2357,N_3950);
or U4315 (N_4315,N_2805,N_2424);
nand U4316 (N_4316,N_2098,N_2010);
nand U4317 (N_4317,N_2662,N_2552);
xnor U4318 (N_4318,N_2026,N_3134);
or U4319 (N_4319,N_3879,N_2451);
and U4320 (N_4320,N_2815,N_3660);
and U4321 (N_4321,N_3357,N_2417);
or U4322 (N_4322,N_3104,N_2195);
or U4323 (N_4323,N_2996,N_3338);
and U4324 (N_4324,N_2586,N_3426);
nand U4325 (N_4325,N_2320,N_2432);
and U4326 (N_4326,N_3196,N_2968);
or U4327 (N_4327,N_3802,N_2176);
or U4328 (N_4328,N_2140,N_2239);
nand U4329 (N_4329,N_2561,N_3270);
nor U4330 (N_4330,N_3301,N_2796);
nor U4331 (N_4331,N_3851,N_2270);
or U4332 (N_4332,N_2422,N_3676);
nand U4333 (N_4333,N_2513,N_2074);
and U4334 (N_4334,N_2379,N_3580);
or U4335 (N_4335,N_3658,N_2635);
xor U4336 (N_4336,N_3142,N_3289);
nand U4337 (N_4337,N_3047,N_2967);
or U4338 (N_4338,N_2030,N_2220);
nor U4339 (N_4339,N_2368,N_2478);
nor U4340 (N_4340,N_2699,N_2880);
nor U4341 (N_4341,N_2548,N_3018);
and U4342 (N_4342,N_2446,N_2606);
nand U4343 (N_4343,N_3826,N_3916);
and U4344 (N_4344,N_3163,N_3135);
and U4345 (N_4345,N_3226,N_3935);
nor U4346 (N_4346,N_2855,N_3661);
nand U4347 (N_4347,N_3440,N_2584);
xnor U4348 (N_4348,N_2777,N_3704);
and U4349 (N_4349,N_3373,N_2182);
nor U4350 (N_4350,N_3161,N_2286);
nand U4351 (N_4351,N_2261,N_3077);
nand U4352 (N_4352,N_2854,N_3413);
or U4353 (N_4353,N_3747,N_2836);
or U4354 (N_4354,N_2597,N_3893);
or U4355 (N_4355,N_3795,N_3065);
nor U4356 (N_4356,N_3707,N_2939);
nand U4357 (N_4357,N_2613,N_3033);
nand U4358 (N_4358,N_2547,N_2647);
or U4359 (N_4359,N_3881,N_3008);
nand U4360 (N_4360,N_3315,N_2740);
nand U4361 (N_4361,N_2177,N_3261);
xnor U4362 (N_4362,N_2196,N_3566);
and U4363 (N_4363,N_3419,N_2349);
and U4364 (N_4364,N_3654,N_3700);
nand U4365 (N_4365,N_3529,N_2240);
or U4366 (N_4366,N_2526,N_3551);
or U4367 (N_4367,N_2089,N_3502);
nor U4368 (N_4368,N_3673,N_2632);
and U4369 (N_4369,N_2515,N_3949);
xor U4370 (N_4370,N_2620,N_2369);
and U4371 (N_4371,N_3820,N_3355);
nor U4372 (N_4372,N_2021,N_2363);
nand U4373 (N_4373,N_3455,N_2564);
and U4374 (N_4374,N_2311,N_2262);
and U4375 (N_4375,N_2628,N_3929);
and U4376 (N_4376,N_3300,N_2183);
or U4377 (N_4377,N_2810,N_2984);
nor U4378 (N_4378,N_3998,N_3004);
nor U4379 (N_4379,N_3940,N_2549);
nand U4380 (N_4380,N_2933,N_2511);
xnor U4381 (N_4381,N_3501,N_2756);
nor U4382 (N_4382,N_3895,N_3657);
nor U4383 (N_4383,N_2006,N_2829);
or U4384 (N_4384,N_3975,N_3546);
nand U4385 (N_4385,N_2590,N_2197);
nor U4386 (N_4386,N_3565,N_2186);
nand U4387 (N_4387,N_2408,N_2633);
and U4388 (N_4388,N_3410,N_2464);
xor U4389 (N_4389,N_3374,N_2373);
or U4390 (N_4390,N_2032,N_3291);
and U4391 (N_4391,N_2252,N_2718);
and U4392 (N_4392,N_3145,N_2133);
and U4393 (N_4393,N_2387,N_2236);
or U4394 (N_4394,N_2671,N_2066);
and U4395 (N_4395,N_2550,N_2345);
or U4396 (N_4396,N_3056,N_2268);
or U4397 (N_4397,N_2621,N_2821);
and U4398 (N_4398,N_3242,N_2041);
nand U4399 (N_4399,N_2251,N_3296);
nand U4400 (N_4400,N_2400,N_2957);
nand U4401 (N_4401,N_2932,N_3295);
nor U4402 (N_4402,N_2792,N_3797);
or U4403 (N_4403,N_3377,N_2095);
nor U4404 (N_4404,N_2524,N_2797);
and U4405 (N_4405,N_3479,N_3597);
and U4406 (N_4406,N_3268,N_3028);
and U4407 (N_4407,N_3434,N_2104);
and U4408 (N_4408,N_3477,N_3138);
or U4409 (N_4409,N_3642,N_3084);
or U4410 (N_4410,N_2178,N_3035);
nor U4411 (N_4411,N_3304,N_2162);
nor U4412 (N_4412,N_3858,N_2212);
and U4413 (N_4413,N_3706,N_3645);
and U4414 (N_4414,N_3156,N_2376);
nand U4415 (N_4415,N_2920,N_3252);
and U4416 (N_4416,N_2882,N_2843);
or U4417 (N_4417,N_3897,N_2078);
nor U4418 (N_4418,N_2568,N_2985);
nor U4419 (N_4419,N_3053,N_2441);
and U4420 (N_4420,N_3531,N_3699);
nand U4421 (N_4421,N_3101,N_2278);
or U4422 (N_4422,N_3379,N_3830);
nor U4423 (N_4423,N_3817,N_3257);
nand U4424 (N_4424,N_3471,N_2609);
nand U4425 (N_4425,N_3358,N_3016);
or U4426 (N_4426,N_2690,N_2915);
and U4427 (N_4427,N_2364,N_3663);
nor U4428 (N_4428,N_3006,N_2825);
nand U4429 (N_4429,N_3194,N_3850);
xnor U4430 (N_4430,N_2869,N_3372);
nand U4431 (N_4431,N_3314,N_3364);
xnor U4432 (N_4432,N_2631,N_2905);
and U4433 (N_4433,N_2865,N_3863);
nand U4434 (N_4434,N_2940,N_3288);
nor U4435 (N_4435,N_2315,N_3638);
and U4436 (N_4436,N_3515,N_2576);
nor U4437 (N_4437,N_3816,N_2888);
and U4438 (N_4438,N_3350,N_2695);
nand U4439 (N_4439,N_2045,N_2119);
nand U4440 (N_4440,N_3892,N_2474);
nand U4441 (N_4441,N_3209,N_3920);
nor U4442 (N_4442,N_3363,N_3584);
nor U4443 (N_4443,N_2225,N_3220);
nand U4444 (N_4444,N_3312,N_3498);
nand U4445 (N_4445,N_3129,N_3678);
and U4446 (N_4446,N_2648,N_3560);
or U4447 (N_4447,N_2391,N_3492);
nor U4448 (N_4448,N_3917,N_3365);
nand U4449 (N_4449,N_3731,N_2529);
and U4450 (N_4450,N_3996,N_3342);
xnor U4451 (N_4451,N_3474,N_3512);
xor U4452 (N_4452,N_2579,N_3720);
xnor U4453 (N_4453,N_2885,N_3012);
nor U4454 (N_4454,N_3189,N_3821);
and U4455 (N_4455,N_3292,N_2516);
xnor U4456 (N_4456,N_3328,N_3207);
nor U4457 (N_4457,N_3277,N_2614);
and U4458 (N_4458,N_3538,N_2011);
xor U4459 (N_4459,N_3254,N_3287);
nand U4460 (N_4460,N_3712,N_2418);
or U4461 (N_4461,N_3577,N_2108);
nand U4462 (N_4462,N_2346,N_3741);
or U4463 (N_4463,N_3583,N_3977);
nor U4464 (N_4464,N_3595,N_3105);
or U4465 (N_4465,N_2009,N_3675);
and U4466 (N_4466,N_3912,N_3548);
or U4467 (N_4467,N_2445,N_2457);
nor U4468 (N_4468,N_2372,N_2437);
nor U4469 (N_4469,N_2319,N_2972);
and U4470 (N_4470,N_2436,N_2352);
nor U4471 (N_4471,N_3561,N_2607);
or U4472 (N_4472,N_2716,N_2201);
nand U4473 (N_4473,N_3428,N_2877);
or U4474 (N_4474,N_3908,N_3079);
nor U4475 (N_4475,N_2048,N_2580);
nor U4476 (N_4476,N_2669,N_3602);
and U4477 (N_4477,N_2883,N_3351);
nand U4478 (N_4478,N_3532,N_2873);
or U4479 (N_4479,N_3569,N_3549);
or U4480 (N_4480,N_3824,N_3925);
or U4481 (N_4481,N_2226,N_2887);
xnor U4482 (N_4482,N_2989,N_3441);
nand U4483 (N_4483,N_2813,N_2678);
nand U4484 (N_4484,N_3599,N_2987);
or U4485 (N_4485,N_2684,N_3656);
and U4486 (N_4486,N_3521,N_3227);
nor U4487 (N_4487,N_3222,N_2382);
or U4488 (N_4488,N_3050,N_2565);
nand U4489 (N_4489,N_3155,N_3792);
or U4490 (N_4490,N_2453,N_3985);
nor U4491 (N_4491,N_3214,N_3298);
or U4492 (N_4492,N_3370,N_3668);
nor U4493 (N_4493,N_3503,N_3745);
nor U4494 (N_4494,N_3562,N_2623);
or U4495 (N_4495,N_2205,N_3040);
or U4496 (N_4496,N_3984,N_3956);
and U4497 (N_4497,N_3829,N_3391);
xor U4498 (N_4498,N_3796,N_3665);
and U4499 (N_4499,N_3326,N_2323);
and U4500 (N_4500,N_2016,N_3766);
and U4501 (N_4501,N_3159,N_2626);
nor U4502 (N_4502,N_2248,N_2834);
nor U4503 (N_4503,N_2675,N_2630);
nand U4504 (N_4504,N_2809,N_3612);
xor U4505 (N_4505,N_2543,N_3688);
nor U4506 (N_4506,N_2793,N_3107);
xor U4507 (N_4507,N_2189,N_3907);
nand U4508 (N_4508,N_2754,N_2404);
or U4509 (N_4509,N_2116,N_2668);
and U4510 (N_4510,N_3903,N_2814);
nor U4511 (N_4511,N_2338,N_3789);
xor U4512 (N_4512,N_3962,N_2342);
xor U4513 (N_4513,N_3751,N_2333);
nand U4514 (N_4514,N_3224,N_3620);
nor U4515 (N_4515,N_2279,N_2469);
nor U4516 (N_4516,N_3485,N_3986);
nor U4517 (N_4517,N_3064,N_2918);
and U4518 (N_4518,N_2769,N_3472);
or U4519 (N_4519,N_2367,N_3540);
or U4520 (N_4520,N_3147,N_3991);
nand U4521 (N_4521,N_3204,N_3953);
nand U4522 (N_4522,N_2415,N_3361);
nand U4523 (N_4523,N_3305,N_2517);
xor U4524 (N_4524,N_3271,N_2895);
xor U4525 (N_4525,N_3930,N_3760);
nor U4526 (N_4526,N_2990,N_2309);
and U4527 (N_4527,N_2494,N_2739);
nand U4528 (N_4528,N_2015,N_2008);
nand U4529 (N_4529,N_3174,N_3451);
xnor U4530 (N_4530,N_2407,N_3014);
nand U4531 (N_4531,N_3809,N_2824);
nor U4532 (N_4532,N_3275,N_2502);
and U4533 (N_4533,N_2005,N_3507);
and U4534 (N_4534,N_2370,N_2470);
nor U4535 (N_4535,N_2411,N_3946);
nand U4536 (N_4536,N_2081,N_3614);
nand U4537 (N_4537,N_3262,N_2080);
and U4538 (N_4538,N_2575,N_2682);
or U4539 (N_4539,N_3716,N_2676);
nand U4540 (N_4540,N_3831,N_3767);
nand U4541 (N_4541,N_2696,N_3636);
and U4542 (N_4542,N_2745,N_2087);
and U4543 (N_4543,N_3768,N_2705);
nor U4544 (N_4544,N_2112,N_3818);
and U4545 (N_4545,N_3799,N_2743);
or U4546 (N_4546,N_2339,N_2608);
and U4547 (N_4547,N_3203,N_3081);
nor U4548 (N_4548,N_3406,N_2131);
xor U4549 (N_4549,N_3253,N_3721);
nand U4550 (N_4550,N_3150,N_3188);
and U4551 (N_4551,N_3763,N_2127);
or U4552 (N_4552,N_3345,N_3106);
and U4553 (N_4553,N_3125,N_3948);
and U4554 (N_4554,N_2247,N_3468);
nand U4555 (N_4555,N_2304,N_2781);
nand U4556 (N_4556,N_2733,N_2503);
or U4557 (N_4557,N_2689,N_2105);
and U4558 (N_4558,N_3489,N_2578);
nor U4559 (N_4559,N_2541,N_2523);
or U4560 (N_4560,N_2434,N_3191);
nor U4561 (N_4561,N_3130,N_2504);
nand U4562 (N_4562,N_2788,N_3992);
nand U4563 (N_4563,N_2480,N_3539);
and U4564 (N_4564,N_2348,N_3608);
nand U4565 (N_4565,N_2406,N_2782);
nand U4566 (N_4566,N_2556,N_3875);
or U4567 (N_4567,N_2290,N_3115);
nand U4568 (N_4568,N_3587,N_3360);
nor U4569 (N_4569,N_2728,N_2024);
xor U4570 (N_4570,N_2569,N_2365);
nor U4571 (N_4571,N_3623,N_3466);
nor U4572 (N_4572,N_2168,N_3449);
and U4573 (N_4573,N_2717,N_3199);
or U4574 (N_4574,N_3819,N_3117);
or U4575 (N_4575,N_3864,N_2649);
or U4576 (N_4576,N_2259,N_3833);
or U4577 (N_4577,N_2198,N_2784);
and U4578 (N_4578,N_2830,N_3504);
and U4579 (N_4579,N_2452,N_2938);
nor U4580 (N_4580,N_2154,N_2190);
and U4581 (N_4581,N_2819,N_3073);
and U4582 (N_4582,N_2977,N_3622);
xnor U4583 (N_4583,N_3890,N_3779);
nand U4584 (N_4584,N_2495,N_2455);
or U4585 (N_4585,N_2169,N_2281);
nand U4586 (N_4586,N_3340,N_3846);
nand U4587 (N_4587,N_3541,N_3404);
nand U4588 (N_4588,N_3961,N_2982);
nand U4589 (N_4589,N_2046,N_2707);
nor U4590 (N_4590,N_2652,N_3787);
nor U4591 (N_4591,N_2462,N_2950);
or U4592 (N_4592,N_3511,N_2175);
and U4593 (N_4593,N_3375,N_2461);
nor U4594 (N_4594,N_2683,N_2913);
or U4595 (N_4595,N_2713,N_2313);
or U4596 (N_4596,N_2202,N_2530);
nor U4597 (N_4597,N_3919,N_3219);
nor U4598 (N_4598,N_2962,N_2172);
and U4599 (N_4599,N_2302,N_2858);
or U4600 (N_4600,N_2312,N_2866);
nor U4601 (N_4601,N_3481,N_3705);
and U4602 (N_4602,N_3842,N_2088);
nand U4603 (N_4603,N_3596,N_3624);
nand U4604 (N_4604,N_2234,N_2467);
nor U4605 (N_4605,N_3861,N_3366);
nand U4606 (N_4606,N_3891,N_2025);
nand U4607 (N_4607,N_2034,N_2475);
or U4608 (N_4608,N_3898,N_2747);
and U4609 (N_4609,N_2981,N_3393);
and U4610 (N_4610,N_2294,N_3723);
or U4611 (N_4611,N_2181,N_3182);
or U4612 (N_4612,N_3089,N_3526);
or U4613 (N_4613,N_2125,N_3717);
and U4614 (N_4614,N_3910,N_2174);
and U4615 (N_4615,N_2514,N_3593);
and U4616 (N_4616,N_2292,N_2044);
nand U4617 (N_4617,N_3573,N_3080);
and U4618 (N_4618,N_2381,N_2295);
xor U4619 (N_4619,N_3325,N_2458);
and U4620 (N_4620,N_3889,N_2153);
and U4621 (N_4621,N_2594,N_3007);
nand U4622 (N_4622,N_3068,N_2271);
nand U4623 (N_4623,N_2875,N_2288);
nor U4624 (N_4624,N_3495,N_3321);
or U4625 (N_4625,N_2519,N_3691);
nor U4626 (N_4626,N_2114,N_2260);
or U4627 (N_4627,N_2941,N_2752);
nand U4628 (N_4628,N_2637,N_2847);
nor U4629 (N_4629,N_3453,N_2521);
xor U4630 (N_4630,N_2158,N_3885);
nand U4631 (N_4631,N_2007,N_3649);
nand U4632 (N_4632,N_2003,N_3269);
or U4633 (N_4633,N_3600,N_3765);
or U4634 (N_4634,N_3505,N_3031);
nand U4635 (N_4635,N_3460,N_2742);
or U4636 (N_4636,N_2800,N_2876);
nand U4637 (N_4637,N_2762,N_3738);
and U4638 (N_4638,N_3264,N_2912);
xor U4639 (N_4639,N_3483,N_2052);
nor U4640 (N_4640,N_2582,N_3024);
and U4641 (N_4641,N_3954,N_2488);
nor U4642 (N_4642,N_3734,N_2491);
and U4643 (N_4643,N_3781,N_2979);
nand U4644 (N_4644,N_2907,N_2863);
and U4645 (N_4645,N_3835,N_3606);
nand U4646 (N_4646,N_2520,N_3123);
nand U4647 (N_4647,N_3256,N_2062);
and U4648 (N_4648,N_3044,N_3461);
nor U4649 (N_4649,N_3450,N_3527);
and U4650 (N_4650,N_2393,N_2889);
or U4651 (N_4651,N_2601,N_3770);
or U4652 (N_4652,N_2975,N_3557);
nand U4653 (N_4653,N_2152,N_3939);
nand U4654 (N_4654,N_2832,N_3963);
nor U4655 (N_4655,N_2658,N_2722);
xnor U4656 (N_4656,N_3682,N_3536);
or U4657 (N_4657,N_2806,N_2537);
and U4658 (N_4658,N_3238,N_2110);
nand U4659 (N_4659,N_2604,N_3915);
nor U4660 (N_4660,N_3726,N_3981);
or U4661 (N_4661,N_3402,N_2826);
nor U4662 (N_4662,N_3914,N_2096);
and U4663 (N_4663,N_2142,N_2946);
nand U4664 (N_4664,N_3497,N_3534);
or U4665 (N_4665,N_2435,N_2706);
or U4666 (N_4666,N_3836,N_3176);
xor U4667 (N_4667,N_2485,N_2691);
and U4668 (N_4668,N_3544,N_3316);
or U4669 (N_4669,N_2673,N_2188);
nand U4670 (N_4670,N_2785,N_3412);
nor U4671 (N_4671,N_3029,N_3965);
and U4672 (N_4672,N_2909,N_2496);
nand U4673 (N_4673,N_2837,N_2846);
nand U4674 (N_4674,N_3398,N_3757);
nand U4675 (N_4675,N_3000,N_2534);
nand U4676 (N_4676,N_3091,N_3621);
nor U4677 (N_4677,N_2255,N_3552);
and U4678 (N_4678,N_3771,N_3124);
xor U4679 (N_4679,N_3839,N_2980);
or U4680 (N_4680,N_2914,N_2735);
nor U4681 (N_4681,N_2592,N_2922);
nand U4682 (N_4682,N_3144,N_2539);
nor U4683 (N_4683,N_2166,N_3855);
and U4684 (N_4684,N_3754,N_2942);
and U4685 (N_4685,N_2267,N_2477);
nor U4686 (N_4686,N_3075,N_2042);
nor U4687 (N_4687,N_2501,N_3852);
nand U4688 (N_4688,N_2328,N_2729);
nor U4689 (N_4689,N_3260,N_2924);
nor U4690 (N_4690,N_2955,N_2273);
nand U4691 (N_4691,N_3162,N_2655);
nor U4692 (N_4692,N_2598,N_3732);
or U4693 (N_4693,N_2820,N_2164);
nor U4694 (N_4694,N_3783,N_2681);
nand U4695 (N_4695,N_2249,N_2744);
and U4696 (N_4696,N_2870,N_2801);
or U4697 (N_4697,N_3448,N_2492);
and U4698 (N_4698,N_3039,N_3058);
and U4699 (N_4699,N_2053,N_2995);
and U4700 (N_4700,N_3513,N_3048);
and U4701 (N_4701,N_2712,N_3446);
nand U4702 (N_4702,N_3247,N_2254);
nor U4703 (N_4703,N_3853,N_3467);
or U4704 (N_4704,N_2758,N_2102);
or U4705 (N_4705,N_3493,N_3232);
or U4706 (N_4706,N_3547,N_2385);
nor U4707 (N_4707,N_2891,N_3735);
nor U4708 (N_4708,N_3217,N_2969);
nand U4709 (N_4709,N_2572,N_3427);
nand U4710 (N_4710,N_2356,N_3659);
nand U4711 (N_4711,N_3197,N_2701);
and U4712 (N_4712,N_2992,N_3926);
or U4713 (N_4713,N_2951,N_2900);
nand U4714 (N_4714,N_3201,N_2161);
and U4715 (N_4715,N_2076,N_3273);
or U4716 (N_4716,N_2481,N_2171);
xor U4717 (N_4717,N_2741,N_3866);
xor U4718 (N_4718,N_3617,N_3395);
or U4719 (N_4719,N_2448,N_2298);
and U4720 (N_4720,N_3578,N_3052);
nand U4721 (N_4721,N_3684,N_3307);
nor U4722 (N_4722,N_3719,N_2484);
and U4723 (N_4723,N_2822,N_2636);
and U4724 (N_4724,N_2902,N_3874);
and U4725 (N_4725,N_2326,N_3475);
nand U4726 (N_4726,N_2611,N_3302);
nand U4727 (N_4727,N_3133,N_2703);
or U4728 (N_4728,N_3807,N_3609);
and U4729 (N_4729,N_2139,N_2057);
and U4730 (N_4730,N_2317,N_3098);
nand U4731 (N_4731,N_3680,N_3967);
and U4732 (N_4732,N_2079,N_2704);
nand U4733 (N_4733,N_3005,N_3478);
nand U4734 (N_4734,N_2783,N_2811);
and U4735 (N_4735,N_3888,N_3038);
or U4736 (N_4736,N_3173,N_2430);
nand U4737 (N_4737,N_3672,N_3579);
xnor U4738 (N_4738,N_2903,N_3433);
nand U4739 (N_4739,N_3211,N_2219);
nor U4740 (N_4740,N_3069,N_3327);
and U4741 (N_4741,N_3800,N_3205);
or U4742 (N_4742,N_3099,N_2700);
nor U4743 (N_4743,N_3803,N_3231);
or U4744 (N_4744,N_3111,N_2641);
and U4745 (N_4745,N_3832,N_3943);
nor U4746 (N_4746,N_3329,N_2207);
nand U4747 (N_4747,N_3352,N_3319);
xnor U4748 (N_4748,N_2128,N_2544);
xnor U4749 (N_4749,N_3333,N_3083);
xnor U4750 (N_4750,N_3112,N_3484);
nand U4751 (N_4751,N_3473,N_3234);
or U4752 (N_4752,N_3827,N_3206);
nor U4753 (N_4753,N_2945,N_2852);
or U4754 (N_4754,N_3641,N_2645);
nand U4755 (N_4755,N_2163,N_2084);
or U4756 (N_4756,N_3648,N_3019);
nand U4757 (N_4757,N_2359,N_3610);
nor U4758 (N_4758,N_3865,N_2546);
nor U4759 (N_4759,N_2659,N_2638);
and U4760 (N_4760,N_3131,N_2324);
xor U4761 (N_4761,N_2581,N_2916);
nand U4762 (N_4762,N_3380,N_2223);
xnor U4763 (N_4763,N_2617,N_3736);
nor U4764 (N_4764,N_2500,N_3140);
nand U4765 (N_4765,N_2405,N_3508);
or U4766 (N_4766,N_2988,N_3240);
xor U4767 (N_4767,N_2001,N_3394);
or U4768 (N_4768,N_2893,N_3094);
and U4769 (N_4769,N_2035,N_2646);
or U4770 (N_4770,N_3310,N_2443);
nand U4771 (N_4771,N_2378,N_2303);
and U4772 (N_4772,N_2246,N_2043);
and U4773 (N_4773,N_2416,N_3689);
nor U4774 (N_4774,N_3494,N_2103);
nand U4775 (N_4775,N_2426,N_2790);
nor U4776 (N_4776,N_3880,N_2069);
xor U4777 (N_4777,N_3249,N_3200);
or U4778 (N_4778,N_2595,N_3979);
and U4779 (N_4779,N_3074,N_2101);
xnor U4780 (N_4780,N_2911,N_2194);
or U4781 (N_4781,N_2910,N_3324);
and U4782 (N_4782,N_2331,N_2002);
xnor U4783 (N_4783,N_3523,N_2677);
or U4784 (N_4784,N_2284,N_2554);
nand U4785 (N_4785,N_2129,N_3280);
nand U4786 (N_4786,N_2299,N_2375);
nand U4787 (N_4787,N_3776,N_2296);
and U4788 (N_4788,N_3683,N_3322);
and U4789 (N_4789,N_3496,N_2463);
nand U4790 (N_4790,N_3166,N_2274);
or U4791 (N_4791,N_3928,N_2027);
and U4792 (N_4792,N_3886,N_2428);
or U4793 (N_4793,N_3218,N_3871);
and U4794 (N_4794,N_2073,N_2654);
or U4795 (N_4795,N_3337,N_3592);
nand U4796 (N_4796,N_2881,N_2943);
and U4797 (N_4797,N_2971,N_3490);
nor U4798 (N_4798,N_3556,N_3576);
xnor U4799 (N_4799,N_2787,N_2459);
nor U4800 (N_4800,N_3259,N_2596);
nand U4801 (N_4801,N_3703,N_3524);
and U4802 (N_4802,N_3957,N_2353);
xnor U4803 (N_4803,N_3983,N_3436);
and U4804 (N_4804,N_3476,N_2807);
and U4805 (N_4805,N_2211,N_3841);
nor U4806 (N_4806,N_2148,N_2661);
nand U4807 (N_4807,N_2731,N_2559);
nand U4808 (N_4808,N_2499,N_3687);
nand U4809 (N_4809,N_3869,N_2997);
xnor U4810 (N_4810,N_2122,N_3514);
xor U4811 (N_4811,N_3225,N_2310);
and U4812 (N_4812,N_2221,N_2921);
nor U4813 (N_4813,N_2065,N_2380);
nand U4814 (N_4814,N_2419,N_3299);
or U4815 (N_4815,N_2072,N_3932);
xor U4816 (N_4816,N_2571,N_2014);
xnor U4817 (N_4817,N_3387,N_3022);
and U4818 (N_4818,N_3168,N_2134);
nand U4819 (N_4819,N_3235,N_3697);
and U4820 (N_4820,N_2994,N_2224);
nand U4821 (N_4821,N_2444,N_2948);
nand U4822 (N_4822,N_2859,N_3294);
nor U4823 (N_4823,N_3070,N_3708);
nor U4824 (N_4824,N_3034,N_3036);
and U4825 (N_4825,N_3702,N_2622);
or U4826 (N_4826,N_3078,N_3722);
nand U4827 (N_4827,N_3690,N_2936);
nand U4828 (N_4828,N_3733,N_3164);
nor U4829 (N_4829,N_3183,N_2904);
or U4830 (N_4830,N_2937,N_3785);
nand U4831 (N_4831,N_2272,N_2409);
or U4832 (N_4832,N_3179,N_3265);
or U4833 (N_4833,N_3973,N_2803);
or U4834 (N_4834,N_2487,N_2860);
nor U4835 (N_4835,N_2351,N_3989);
or U4836 (N_4836,N_2527,N_3392);
nand U4837 (N_4837,N_2786,N_2749);
nand U4838 (N_4838,N_3980,N_3633);
or U4839 (N_4839,N_3873,N_2004);
and U4840 (N_4840,N_2928,N_2780);
nand U4841 (N_4841,N_2878,N_3108);
and U4842 (N_4842,N_2413,N_2856);
nand U4843 (N_4843,N_3801,N_3293);
nand U4844 (N_4844,N_2853,N_3021);
and U4845 (N_4845,N_2884,N_2709);
nor U4846 (N_4846,N_3999,N_2269);
or U4847 (N_4847,N_3121,N_3010);
and U4848 (N_4848,N_3425,N_3603);
nand U4849 (N_4849,N_2263,N_2209);
nor U4850 (N_4850,N_3187,N_2115);
nand U4851 (N_4851,N_2714,N_3330);
xnor U4852 (N_4852,N_3009,N_2748);
xor U4853 (N_4853,N_3995,N_2923);
nor U4854 (N_4854,N_2213,N_2250);
or U4855 (N_4855,N_2343,N_2759);
or U4856 (N_4856,N_3805,N_3750);
nor U4857 (N_4857,N_3868,N_2362);
nand U4858 (N_4858,N_3020,N_3362);
nor U4859 (N_4859,N_3087,N_2132);
or U4860 (N_4860,N_2874,N_3806);
or U4861 (N_4861,N_3435,N_2687);
and U4862 (N_4862,N_3405,N_3030);
nor U4863 (N_4863,N_2241,N_2894);
and U4864 (N_4864,N_3158,N_3399);
nor U4865 (N_4865,N_3585,N_2433);
and U4866 (N_4866,N_3970,N_3978);
xnor U4867 (N_4867,N_2639,N_3976);
or U4868 (N_4868,N_2931,N_2711);
xnor U4869 (N_4869,N_2764,N_3066);
or U4870 (N_4870,N_2799,N_2297);
and U4871 (N_4871,N_3607,N_3632);
nand U4872 (N_4872,N_2917,N_2386);
and U4873 (N_4873,N_2107,N_2721);
and U4874 (N_4874,N_2291,N_2835);
xor U4875 (N_4875,N_2060,N_2017);
and U4876 (N_4876,N_2397,N_2265);
nand U4877 (N_4877,N_2908,N_3415);
nand U4878 (N_4878,N_3267,N_3605);
xnor U4879 (N_4879,N_3458,N_3152);
or U4880 (N_4880,N_3447,N_2055);
and U4881 (N_4881,N_2525,N_2285);
and U4882 (N_4882,N_3233,N_2028);
nand U4883 (N_4883,N_3941,N_2642);
or U4884 (N_4884,N_2925,N_3444);
and U4885 (N_4885,N_2191,N_2531);
or U4886 (N_4886,N_3674,N_3615);
nand U4887 (N_4887,N_3320,N_3090);
and U4888 (N_4888,N_2610,N_2591);
or U4889 (N_4889,N_3782,N_3348);
and U4890 (N_4890,N_2538,N_3282);
nor U4891 (N_4891,N_3906,N_2871);
nor U4892 (N_4892,N_3774,N_3185);
nor U4893 (N_4893,N_2848,N_3193);
xnor U4894 (N_4894,N_2449,N_2085);
nand U4895 (N_4895,N_3251,N_2227);
xor U4896 (N_4896,N_2602,N_3840);
nand U4897 (N_4897,N_3424,N_3550);
or U4898 (N_4898,N_2117,N_3192);
and U4899 (N_4899,N_3876,N_3002);
nor U4900 (N_4900,N_3662,N_2518);
and U4901 (N_4901,N_2867,N_2961);
nand U4902 (N_4902,N_2688,N_3634);
and U4903 (N_4903,N_2438,N_3740);
or U4904 (N_4904,N_3845,N_2665);
xor U4905 (N_4905,N_2949,N_3245);
nor U4906 (N_4906,N_2215,N_3714);
and U4907 (N_4907,N_3459,N_2694);
and U4908 (N_4908,N_3590,N_2141);
and U4909 (N_4909,N_3297,N_2059);
and U4910 (N_4910,N_2507,N_3149);
nor U4911 (N_4911,N_3272,N_3945);
nor U4912 (N_4912,N_2051,N_3960);
nand U4913 (N_4913,N_2305,N_3854);
and U4914 (N_4914,N_3025,N_3902);
and U4915 (N_4915,N_3904,N_3403);
and U4916 (N_4916,N_3927,N_2340);
nor U4917 (N_4917,N_3439,N_3212);
nor U4918 (N_4918,N_2588,N_2897);
nand U4919 (N_4919,N_2063,N_2068);
nor U4920 (N_4920,N_2377,N_3382);
or U4921 (N_4921,N_3693,N_3347);
xnor U4922 (N_4922,N_2203,N_3061);
nor U4923 (N_4923,N_3303,N_3651);
and U4924 (N_4924,N_2778,N_2760);
or U4925 (N_4925,N_2439,N_3924);
or U4926 (N_4926,N_2685,N_2332);
or U4927 (N_4927,N_3877,N_2816);
and U4928 (N_4928,N_3670,N_2064);
and U4929 (N_4929,N_3971,N_2823);
or U4930 (N_4930,N_3752,N_2257);
or U4931 (N_4931,N_2812,N_2751);
nor U4932 (N_4932,N_3071,N_2506);
nor U4933 (N_4933,N_3518,N_3432);
xnor U4934 (N_4934,N_3921,N_3761);
nor U4935 (N_4935,N_2167,N_2509);
nor U4936 (N_4936,N_2350,N_3103);
xor U4937 (N_4937,N_3266,N_3113);
and U4938 (N_4938,N_3100,N_3353);
and U4939 (N_4939,N_2657,N_2070);
and U4940 (N_4940,N_3093,N_3167);
nand U4941 (N_4941,N_2619,N_2071);
or U4942 (N_4942,N_3396,N_2394);
nand U4943 (N_4943,N_2245,N_3356);
and U4944 (N_4944,N_3181,N_2146);
or U4945 (N_4945,N_2293,N_3611);
nor U4946 (N_4946,N_2389,N_2973);
and U4947 (N_4947,N_2143,N_3887);
or U4948 (N_4948,N_2666,N_3997);
and U4949 (N_4949,N_3530,N_2644);
or U4950 (N_4950,N_3554,N_3695);
xnor U4951 (N_4951,N_3883,N_3937);
nor U4952 (N_4952,N_2316,N_3136);
nand U4953 (N_4953,N_3838,N_2730);
and U4954 (N_4954,N_3628,N_2624);
nand U4955 (N_4955,N_2964,N_3791);
nor U4956 (N_4956,N_2766,N_2944);
nor U4957 (N_4957,N_3543,N_2136);
nand U4958 (N_4958,N_3381,N_2160);
xnor U4959 (N_4959,N_2090,N_3913);
nor U4960 (N_4960,N_2147,N_2466);
nor U4961 (N_4961,N_2429,N_3790);
nand U4962 (N_4962,N_2097,N_2204);
nand U4963 (N_4963,N_3810,N_2109);
nand U4964 (N_4964,N_3896,N_2420);
or U4965 (N_4965,N_2280,N_2159);
nand U4966 (N_4966,N_3715,N_2840);
nor U4967 (N_4967,N_2755,N_2442);
nor U4968 (N_4968,N_2776,N_3718);
and U4969 (N_4969,N_2817,N_2179);
and U4970 (N_4970,N_2138,N_3813);
nand U4971 (N_4971,N_3109,N_2562);
nor U4972 (N_4972,N_2013,N_2656);
or U4973 (N_4973,N_2210,N_3729);
nor U4974 (N_4974,N_3901,N_3409);
or U4975 (N_4975,N_2341,N_3186);
xor U4976 (N_4976,N_3909,N_3343);
xor U4977 (N_4977,N_2686,N_2427);
nand U4978 (N_4978,N_2959,N_3255);
or U4979 (N_4979,N_2725,N_2423);
or U4980 (N_4980,N_3177,N_2551);
or U4981 (N_4981,N_2489,N_3346);
and U4982 (N_4982,N_2238,N_3749);
and U4983 (N_4983,N_2479,N_3331);
and U4984 (N_4984,N_3082,N_2737);
and U4985 (N_4985,N_2049,N_3516);
or U4986 (N_4986,N_3169,N_3041);
nand U4987 (N_4987,N_3545,N_2124);
and U4988 (N_4988,N_2374,N_3533);
nor U4989 (N_4989,N_3488,N_2206);
nor U4990 (N_4990,N_2771,N_2157);
or U4991 (N_4991,N_2930,N_2770);
and U4992 (N_4992,N_3284,N_2384);
and U4993 (N_4993,N_2674,N_2301);
nand U4994 (N_4994,N_2966,N_2693);
nand U4995 (N_4995,N_3421,N_3772);
or U4996 (N_4996,N_2650,N_3959);
nand U4997 (N_4997,N_3798,N_2868);
nand U4998 (N_4998,N_2306,N_3128);
and U4999 (N_4999,N_3279,N_2660);
nor U5000 (N_5000,N_3001,N_2260);
and U5001 (N_5001,N_2478,N_3517);
nor U5002 (N_5002,N_2859,N_3334);
and U5003 (N_5003,N_2169,N_2477);
xor U5004 (N_5004,N_2006,N_2804);
xnor U5005 (N_5005,N_2806,N_2295);
nor U5006 (N_5006,N_2141,N_3117);
nor U5007 (N_5007,N_2760,N_3601);
nand U5008 (N_5008,N_3331,N_3880);
and U5009 (N_5009,N_2899,N_2913);
or U5010 (N_5010,N_2906,N_3550);
and U5011 (N_5011,N_2193,N_3022);
nor U5012 (N_5012,N_3746,N_2721);
nor U5013 (N_5013,N_3463,N_3255);
and U5014 (N_5014,N_3881,N_2136);
nor U5015 (N_5015,N_2248,N_2720);
and U5016 (N_5016,N_2664,N_2732);
and U5017 (N_5017,N_3393,N_3704);
xnor U5018 (N_5018,N_2382,N_2360);
and U5019 (N_5019,N_2123,N_3986);
or U5020 (N_5020,N_3777,N_2388);
or U5021 (N_5021,N_3011,N_2532);
nor U5022 (N_5022,N_3398,N_2676);
or U5023 (N_5023,N_3951,N_2051);
or U5024 (N_5024,N_3520,N_3142);
or U5025 (N_5025,N_3208,N_3045);
nor U5026 (N_5026,N_3975,N_3014);
and U5027 (N_5027,N_2429,N_3245);
and U5028 (N_5028,N_2749,N_3907);
or U5029 (N_5029,N_2567,N_3144);
nand U5030 (N_5030,N_3024,N_3851);
and U5031 (N_5031,N_2544,N_2159);
and U5032 (N_5032,N_2639,N_3750);
nand U5033 (N_5033,N_2640,N_3768);
xnor U5034 (N_5034,N_3420,N_2263);
or U5035 (N_5035,N_2220,N_3789);
nand U5036 (N_5036,N_2109,N_3485);
and U5037 (N_5037,N_2395,N_3631);
and U5038 (N_5038,N_2212,N_3211);
and U5039 (N_5039,N_2575,N_3587);
and U5040 (N_5040,N_3034,N_3892);
nand U5041 (N_5041,N_2144,N_3101);
and U5042 (N_5042,N_3830,N_2182);
nor U5043 (N_5043,N_2883,N_2335);
and U5044 (N_5044,N_3132,N_2536);
nand U5045 (N_5045,N_3291,N_3730);
nand U5046 (N_5046,N_2621,N_3078);
nand U5047 (N_5047,N_3655,N_2203);
nor U5048 (N_5048,N_3912,N_2911);
and U5049 (N_5049,N_3012,N_2644);
or U5050 (N_5050,N_2913,N_3322);
and U5051 (N_5051,N_3419,N_3797);
or U5052 (N_5052,N_3248,N_3796);
nand U5053 (N_5053,N_3430,N_2265);
xnor U5054 (N_5054,N_2510,N_3031);
nand U5055 (N_5055,N_2537,N_3064);
nor U5056 (N_5056,N_2978,N_3841);
nand U5057 (N_5057,N_2548,N_3582);
and U5058 (N_5058,N_3301,N_3194);
nor U5059 (N_5059,N_3411,N_2609);
or U5060 (N_5060,N_3199,N_3063);
or U5061 (N_5061,N_2637,N_3399);
or U5062 (N_5062,N_3641,N_3875);
nand U5063 (N_5063,N_2839,N_2286);
and U5064 (N_5064,N_2346,N_3677);
and U5065 (N_5065,N_2743,N_2193);
or U5066 (N_5066,N_3803,N_2038);
nor U5067 (N_5067,N_3657,N_2769);
nor U5068 (N_5068,N_2143,N_3745);
nand U5069 (N_5069,N_3967,N_2726);
nor U5070 (N_5070,N_3837,N_2315);
nand U5071 (N_5071,N_2901,N_3819);
and U5072 (N_5072,N_2990,N_3597);
nand U5073 (N_5073,N_2460,N_2465);
and U5074 (N_5074,N_3309,N_3576);
or U5075 (N_5075,N_2089,N_3711);
or U5076 (N_5076,N_2925,N_2069);
or U5077 (N_5077,N_2023,N_3451);
nor U5078 (N_5078,N_3639,N_3762);
nand U5079 (N_5079,N_2569,N_2613);
or U5080 (N_5080,N_2834,N_2546);
xnor U5081 (N_5081,N_3668,N_2034);
xnor U5082 (N_5082,N_2409,N_2615);
xor U5083 (N_5083,N_3740,N_3820);
xnor U5084 (N_5084,N_2757,N_2294);
nand U5085 (N_5085,N_3456,N_3403);
or U5086 (N_5086,N_3413,N_2845);
or U5087 (N_5087,N_2146,N_3884);
nor U5088 (N_5088,N_3996,N_2404);
nand U5089 (N_5089,N_2386,N_2761);
nor U5090 (N_5090,N_3386,N_2784);
nand U5091 (N_5091,N_2689,N_3583);
nor U5092 (N_5092,N_2622,N_3187);
nand U5093 (N_5093,N_2545,N_2323);
nor U5094 (N_5094,N_3501,N_2961);
or U5095 (N_5095,N_3820,N_3188);
nand U5096 (N_5096,N_3601,N_2696);
nor U5097 (N_5097,N_2312,N_2831);
nor U5098 (N_5098,N_2462,N_3091);
and U5099 (N_5099,N_3026,N_2565);
and U5100 (N_5100,N_3465,N_2701);
nor U5101 (N_5101,N_3833,N_2379);
nand U5102 (N_5102,N_2700,N_2513);
nand U5103 (N_5103,N_2370,N_3091);
and U5104 (N_5104,N_3505,N_3158);
or U5105 (N_5105,N_2929,N_2362);
or U5106 (N_5106,N_2452,N_3415);
and U5107 (N_5107,N_3453,N_3687);
nand U5108 (N_5108,N_3799,N_3143);
nand U5109 (N_5109,N_2647,N_3463);
nor U5110 (N_5110,N_2063,N_3714);
nor U5111 (N_5111,N_3134,N_2029);
or U5112 (N_5112,N_2458,N_3546);
nand U5113 (N_5113,N_2323,N_3745);
nor U5114 (N_5114,N_2818,N_2905);
nor U5115 (N_5115,N_2911,N_2779);
and U5116 (N_5116,N_3004,N_3037);
nand U5117 (N_5117,N_2801,N_2262);
xor U5118 (N_5118,N_2457,N_2540);
nor U5119 (N_5119,N_2377,N_3331);
nand U5120 (N_5120,N_2598,N_2942);
nand U5121 (N_5121,N_3858,N_3528);
nand U5122 (N_5122,N_2094,N_2987);
nor U5123 (N_5123,N_2621,N_2754);
nor U5124 (N_5124,N_3780,N_3195);
xnor U5125 (N_5125,N_3684,N_2596);
or U5126 (N_5126,N_3249,N_2306);
or U5127 (N_5127,N_2651,N_3274);
nand U5128 (N_5128,N_3406,N_3633);
nand U5129 (N_5129,N_3573,N_2729);
nand U5130 (N_5130,N_3466,N_3151);
and U5131 (N_5131,N_2317,N_3678);
or U5132 (N_5132,N_3846,N_3636);
nand U5133 (N_5133,N_2167,N_2976);
nor U5134 (N_5134,N_3646,N_2307);
xor U5135 (N_5135,N_3928,N_2572);
xor U5136 (N_5136,N_3515,N_3152);
and U5137 (N_5137,N_3912,N_2079);
nand U5138 (N_5138,N_3824,N_3657);
nand U5139 (N_5139,N_2128,N_2507);
nand U5140 (N_5140,N_3435,N_2470);
nand U5141 (N_5141,N_2891,N_2832);
nand U5142 (N_5142,N_3181,N_2224);
nor U5143 (N_5143,N_2698,N_3628);
or U5144 (N_5144,N_2886,N_3975);
nor U5145 (N_5145,N_3065,N_2250);
nor U5146 (N_5146,N_2976,N_3165);
xor U5147 (N_5147,N_3827,N_2812);
nand U5148 (N_5148,N_3175,N_2310);
nor U5149 (N_5149,N_3648,N_2945);
nand U5150 (N_5150,N_2261,N_3030);
and U5151 (N_5151,N_3344,N_3708);
or U5152 (N_5152,N_3934,N_3951);
or U5153 (N_5153,N_3532,N_2397);
nand U5154 (N_5154,N_3481,N_2967);
or U5155 (N_5155,N_2598,N_3630);
or U5156 (N_5156,N_3423,N_2962);
nor U5157 (N_5157,N_3330,N_2970);
and U5158 (N_5158,N_3883,N_2302);
nor U5159 (N_5159,N_3084,N_2376);
nor U5160 (N_5160,N_3295,N_3945);
nand U5161 (N_5161,N_2053,N_2335);
nor U5162 (N_5162,N_2656,N_3364);
nor U5163 (N_5163,N_2203,N_2778);
and U5164 (N_5164,N_3289,N_3550);
nand U5165 (N_5165,N_2737,N_3435);
and U5166 (N_5166,N_3115,N_2343);
xor U5167 (N_5167,N_3918,N_2729);
nand U5168 (N_5168,N_3106,N_3999);
and U5169 (N_5169,N_2074,N_3938);
and U5170 (N_5170,N_2899,N_3870);
and U5171 (N_5171,N_3045,N_3249);
nor U5172 (N_5172,N_2125,N_3169);
xnor U5173 (N_5173,N_3393,N_3729);
xnor U5174 (N_5174,N_2110,N_2855);
nand U5175 (N_5175,N_3324,N_3812);
or U5176 (N_5176,N_2883,N_2652);
nand U5177 (N_5177,N_3030,N_2726);
or U5178 (N_5178,N_3864,N_2556);
and U5179 (N_5179,N_3858,N_3255);
and U5180 (N_5180,N_3592,N_3144);
nor U5181 (N_5181,N_2316,N_3025);
nor U5182 (N_5182,N_2476,N_3044);
and U5183 (N_5183,N_2701,N_2166);
nand U5184 (N_5184,N_3871,N_3819);
nor U5185 (N_5185,N_2929,N_3523);
nor U5186 (N_5186,N_3175,N_3019);
nor U5187 (N_5187,N_3403,N_3011);
and U5188 (N_5188,N_2849,N_3252);
nand U5189 (N_5189,N_2343,N_3477);
nand U5190 (N_5190,N_2273,N_2193);
nand U5191 (N_5191,N_3190,N_3313);
nand U5192 (N_5192,N_3812,N_3597);
nor U5193 (N_5193,N_3510,N_2649);
nand U5194 (N_5194,N_2349,N_2410);
nor U5195 (N_5195,N_3605,N_2660);
nand U5196 (N_5196,N_3642,N_2413);
nand U5197 (N_5197,N_3562,N_2461);
and U5198 (N_5198,N_3497,N_2859);
nor U5199 (N_5199,N_2928,N_2455);
or U5200 (N_5200,N_2541,N_3360);
nor U5201 (N_5201,N_3244,N_2360);
nor U5202 (N_5202,N_2948,N_2071);
nand U5203 (N_5203,N_2630,N_2043);
or U5204 (N_5204,N_3277,N_3889);
or U5205 (N_5205,N_2664,N_2600);
xor U5206 (N_5206,N_3197,N_2898);
nor U5207 (N_5207,N_3847,N_2544);
nor U5208 (N_5208,N_2550,N_3855);
nand U5209 (N_5209,N_2434,N_2208);
and U5210 (N_5210,N_2007,N_3658);
nand U5211 (N_5211,N_2260,N_3939);
and U5212 (N_5212,N_3770,N_2226);
or U5213 (N_5213,N_3961,N_3874);
or U5214 (N_5214,N_2545,N_2501);
xnor U5215 (N_5215,N_2476,N_2982);
or U5216 (N_5216,N_3571,N_3515);
nor U5217 (N_5217,N_3613,N_3697);
or U5218 (N_5218,N_3251,N_2155);
nand U5219 (N_5219,N_2376,N_3042);
or U5220 (N_5220,N_2138,N_3255);
xor U5221 (N_5221,N_3228,N_3191);
nor U5222 (N_5222,N_3204,N_2512);
nor U5223 (N_5223,N_2641,N_3601);
xnor U5224 (N_5224,N_3446,N_3989);
or U5225 (N_5225,N_2229,N_2178);
or U5226 (N_5226,N_3978,N_2296);
nand U5227 (N_5227,N_3150,N_3969);
and U5228 (N_5228,N_3741,N_2140);
nor U5229 (N_5229,N_3686,N_3631);
nand U5230 (N_5230,N_2584,N_3667);
and U5231 (N_5231,N_2134,N_3576);
and U5232 (N_5232,N_2363,N_3384);
and U5233 (N_5233,N_2990,N_2436);
nor U5234 (N_5234,N_2269,N_3882);
and U5235 (N_5235,N_3237,N_2324);
or U5236 (N_5236,N_2690,N_3015);
nand U5237 (N_5237,N_2901,N_2622);
or U5238 (N_5238,N_2656,N_3828);
nor U5239 (N_5239,N_3907,N_3102);
nand U5240 (N_5240,N_3794,N_3611);
nand U5241 (N_5241,N_2781,N_2694);
or U5242 (N_5242,N_3602,N_2032);
xnor U5243 (N_5243,N_3887,N_2986);
or U5244 (N_5244,N_3679,N_2695);
and U5245 (N_5245,N_2649,N_2594);
xnor U5246 (N_5246,N_2016,N_2294);
or U5247 (N_5247,N_2896,N_2285);
or U5248 (N_5248,N_2417,N_2283);
or U5249 (N_5249,N_3575,N_3055);
nand U5250 (N_5250,N_3808,N_2624);
nand U5251 (N_5251,N_3245,N_2421);
nor U5252 (N_5252,N_2373,N_2542);
nand U5253 (N_5253,N_2068,N_2161);
and U5254 (N_5254,N_2882,N_2542);
and U5255 (N_5255,N_3273,N_2078);
nor U5256 (N_5256,N_2565,N_2704);
and U5257 (N_5257,N_3888,N_3184);
nor U5258 (N_5258,N_3353,N_2043);
and U5259 (N_5259,N_2075,N_2041);
xnor U5260 (N_5260,N_2606,N_2191);
nor U5261 (N_5261,N_2036,N_3369);
nand U5262 (N_5262,N_3902,N_3952);
nand U5263 (N_5263,N_3378,N_2016);
nor U5264 (N_5264,N_2627,N_2808);
or U5265 (N_5265,N_3805,N_3181);
nand U5266 (N_5266,N_2356,N_2637);
nor U5267 (N_5267,N_3022,N_3917);
and U5268 (N_5268,N_3964,N_2830);
and U5269 (N_5269,N_3468,N_2654);
or U5270 (N_5270,N_2771,N_2500);
nand U5271 (N_5271,N_3769,N_2788);
or U5272 (N_5272,N_2888,N_3271);
xnor U5273 (N_5273,N_3185,N_2088);
and U5274 (N_5274,N_2813,N_2681);
nor U5275 (N_5275,N_3315,N_3439);
nor U5276 (N_5276,N_3853,N_2751);
nor U5277 (N_5277,N_2793,N_2655);
and U5278 (N_5278,N_3470,N_3052);
and U5279 (N_5279,N_2595,N_2246);
nand U5280 (N_5280,N_2465,N_3251);
or U5281 (N_5281,N_3716,N_2464);
and U5282 (N_5282,N_3051,N_2503);
nand U5283 (N_5283,N_2642,N_2676);
and U5284 (N_5284,N_2983,N_2015);
or U5285 (N_5285,N_3234,N_3127);
or U5286 (N_5286,N_3293,N_3881);
and U5287 (N_5287,N_2119,N_3770);
xor U5288 (N_5288,N_2148,N_3563);
nor U5289 (N_5289,N_3259,N_3415);
nand U5290 (N_5290,N_2573,N_3502);
xor U5291 (N_5291,N_3752,N_2239);
xnor U5292 (N_5292,N_3114,N_2554);
nand U5293 (N_5293,N_2298,N_2840);
and U5294 (N_5294,N_3868,N_3744);
nand U5295 (N_5295,N_2718,N_3956);
nor U5296 (N_5296,N_3425,N_2570);
nand U5297 (N_5297,N_2175,N_2768);
nor U5298 (N_5298,N_3923,N_3340);
nor U5299 (N_5299,N_3735,N_3391);
nand U5300 (N_5300,N_3560,N_3802);
and U5301 (N_5301,N_2727,N_3769);
nor U5302 (N_5302,N_2184,N_2692);
nand U5303 (N_5303,N_3466,N_3929);
or U5304 (N_5304,N_3881,N_2296);
nor U5305 (N_5305,N_2169,N_2018);
nor U5306 (N_5306,N_2572,N_2728);
or U5307 (N_5307,N_3276,N_3324);
and U5308 (N_5308,N_3385,N_2392);
nor U5309 (N_5309,N_2161,N_3015);
or U5310 (N_5310,N_2949,N_3172);
xor U5311 (N_5311,N_2102,N_3714);
nand U5312 (N_5312,N_3247,N_2152);
and U5313 (N_5313,N_2442,N_3818);
or U5314 (N_5314,N_2292,N_3079);
and U5315 (N_5315,N_2503,N_2343);
nor U5316 (N_5316,N_2525,N_2291);
xnor U5317 (N_5317,N_3983,N_3927);
or U5318 (N_5318,N_3042,N_3287);
nand U5319 (N_5319,N_2909,N_2830);
xnor U5320 (N_5320,N_2669,N_2253);
or U5321 (N_5321,N_2593,N_2534);
or U5322 (N_5322,N_2793,N_2684);
nand U5323 (N_5323,N_2669,N_3348);
xnor U5324 (N_5324,N_3869,N_3924);
nand U5325 (N_5325,N_3773,N_3040);
or U5326 (N_5326,N_3279,N_2659);
and U5327 (N_5327,N_3057,N_2606);
or U5328 (N_5328,N_3506,N_3271);
nand U5329 (N_5329,N_2005,N_3197);
nand U5330 (N_5330,N_2591,N_2409);
nand U5331 (N_5331,N_3408,N_2307);
or U5332 (N_5332,N_2594,N_2974);
and U5333 (N_5333,N_3699,N_3834);
or U5334 (N_5334,N_3717,N_2279);
or U5335 (N_5335,N_3745,N_2902);
and U5336 (N_5336,N_2355,N_2079);
or U5337 (N_5337,N_3543,N_3037);
nand U5338 (N_5338,N_3727,N_3399);
xor U5339 (N_5339,N_3550,N_2098);
nor U5340 (N_5340,N_3501,N_2109);
nand U5341 (N_5341,N_3918,N_3574);
nand U5342 (N_5342,N_2949,N_3578);
xor U5343 (N_5343,N_3387,N_2752);
or U5344 (N_5344,N_3064,N_2482);
nor U5345 (N_5345,N_3786,N_2791);
and U5346 (N_5346,N_3937,N_2697);
and U5347 (N_5347,N_2245,N_2647);
nor U5348 (N_5348,N_3992,N_3977);
or U5349 (N_5349,N_3875,N_3607);
nand U5350 (N_5350,N_2530,N_3587);
and U5351 (N_5351,N_2234,N_2392);
xor U5352 (N_5352,N_3802,N_3767);
nand U5353 (N_5353,N_2264,N_2960);
or U5354 (N_5354,N_2853,N_2574);
nor U5355 (N_5355,N_2020,N_2726);
or U5356 (N_5356,N_3303,N_3468);
nand U5357 (N_5357,N_2769,N_3253);
nor U5358 (N_5358,N_2980,N_3237);
or U5359 (N_5359,N_2233,N_3990);
xor U5360 (N_5360,N_2916,N_3799);
and U5361 (N_5361,N_3872,N_2935);
or U5362 (N_5362,N_3162,N_2866);
nand U5363 (N_5363,N_3237,N_3899);
and U5364 (N_5364,N_2709,N_3669);
and U5365 (N_5365,N_3197,N_2380);
nand U5366 (N_5366,N_2020,N_3408);
or U5367 (N_5367,N_2006,N_2639);
nand U5368 (N_5368,N_2056,N_2586);
nand U5369 (N_5369,N_3831,N_2375);
nor U5370 (N_5370,N_3800,N_3969);
and U5371 (N_5371,N_2509,N_2961);
or U5372 (N_5372,N_2598,N_3228);
or U5373 (N_5373,N_3421,N_2199);
and U5374 (N_5374,N_2526,N_3853);
and U5375 (N_5375,N_3800,N_2248);
nor U5376 (N_5376,N_3179,N_2089);
or U5377 (N_5377,N_2200,N_2208);
and U5378 (N_5378,N_2435,N_2974);
nor U5379 (N_5379,N_2054,N_3783);
nand U5380 (N_5380,N_3817,N_3883);
nor U5381 (N_5381,N_3181,N_2227);
or U5382 (N_5382,N_2554,N_2240);
nand U5383 (N_5383,N_3685,N_2344);
nand U5384 (N_5384,N_2960,N_3099);
nand U5385 (N_5385,N_3236,N_3963);
nor U5386 (N_5386,N_3691,N_2976);
nand U5387 (N_5387,N_3142,N_2898);
and U5388 (N_5388,N_3344,N_2204);
nor U5389 (N_5389,N_2328,N_3354);
nor U5390 (N_5390,N_2536,N_3171);
nor U5391 (N_5391,N_3375,N_2612);
nand U5392 (N_5392,N_3558,N_3933);
nand U5393 (N_5393,N_3223,N_3413);
nor U5394 (N_5394,N_3713,N_2910);
or U5395 (N_5395,N_2116,N_2557);
nor U5396 (N_5396,N_3379,N_2983);
and U5397 (N_5397,N_3455,N_3170);
nor U5398 (N_5398,N_3391,N_3321);
or U5399 (N_5399,N_2143,N_2003);
and U5400 (N_5400,N_2437,N_3940);
nand U5401 (N_5401,N_2579,N_2879);
and U5402 (N_5402,N_3300,N_3685);
and U5403 (N_5403,N_2382,N_2401);
or U5404 (N_5404,N_3906,N_3937);
nand U5405 (N_5405,N_2899,N_2281);
nand U5406 (N_5406,N_3989,N_3210);
nor U5407 (N_5407,N_3797,N_2892);
nor U5408 (N_5408,N_2649,N_3757);
xor U5409 (N_5409,N_3967,N_2540);
nor U5410 (N_5410,N_2598,N_2534);
nor U5411 (N_5411,N_2288,N_3897);
and U5412 (N_5412,N_2323,N_3884);
xnor U5413 (N_5413,N_3095,N_3330);
xnor U5414 (N_5414,N_3650,N_3893);
or U5415 (N_5415,N_3701,N_3336);
nor U5416 (N_5416,N_2004,N_2069);
or U5417 (N_5417,N_3140,N_2730);
nand U5418 (N_5418,N_2518,N_2888);
nand U5419 (N_5419,N_3010,N_3888);
or U5420 (N_5420,N_3244,N_2579);
nor U5421 (N_5421,N_3811,N_2064);
or U5422 (N_5422,N_2071,N_2803);
and U5423 (N_5423,N_2223,N_3201);
nor U5424 (N_5424,N_3384,N_3568);
nor U5425 (N_5425,N_3460,N_3015);
xnor U5426 (N_5426,N_3221,N_2478);
nor U5427 (N_5427,N_3314,N_3050);
nand U5428 (N_5428,N_3892,N_2232);
and U5429 (N_5429,N_2860,N_2025);
nand U5430 (N_5430,N_2632,N_3288);
nand U5431 (N_5431,N_3735,N_3745);
or U5432 (N_5432,N_3941,N_3267);
or U5433 (N_5433,N_3097,N_2203);
or U5434 (N_5434,N_2147,N_3385);
and U5435 (N_5435,N_3880,N_3865);
or U5436 (N_5436,N_2033,N_3762);
or U5437 (N_5437,N_3985,N_3540);
nor U5438 (N_5438,N_3643,N_2315);
xnor U5439 (N_5439,N_2694,N_2267);
and U5440 (N_5440,N_3099,N_3428);
xor U5441 (N_5441,N_3061,N_2966);
and U5442 (N_5442,N_2211,N_2613);
nor U5443 (N_5443,N_2624,N_2085);
and U5444 (N_5444,N_2998,N_2571);
and U5445 (N_5445,N_2301,N_3798);
nand U5446 (N_5446,N_3081,N_2563);
xor U5447 (N_5447,N_3633,N_2785);
or U5448 (N_5448,N_3268,N_3194);
or U5449 (N_5449,N_2063,N_3024);
nand U5450 (N_5450,N_3334,N_3297);
or U5451 (N_5451,N_3517,N_2533);
nand U5452 (N_5452,N_3916,N_2472);
or U5453 (N_5453,N_2443,N_3990);
and U5454 (N_5454,N_3182,N_3853);
or U5455 (N_5455,N_3226,N_3642);
nor U5456 (N_5456,N_2559,N_3450);
nand U5457 (N_5457,N_3137,N_2791);
nand U5458 (N_5458,N_2077,N_3942);
and U5459 (N_5459,N_3567,N_2389);
and U5460 (N_5460,N_2586,N_2685);
or U5461 (N_5461,N_2352,N_3191);
nor U5462 (N_5462,N_2728,N_2226);
nand U5463 (N_5463,N_2589,N_3307);
or U5464 (N_5464,N_3687,N_2895);
nor U5465 (N_5465,N_2230,N_2702);
nand U5466 (N_5466,N_2110,N_2269);
or U5467 (N_5467,N_2643,N_3369);
nand U5468 (N_5468,N_3833,N_3234);
or U5469 (N_5469,N_2189,N_3593);
xor U5470 (N_5470,N_3819,N_3220);
nor U5471 (N_5471,N_2989,N_3543);
nor U5472 (N_5472,N_2930,N_3897);
and U5473 (N_5473,N_3136,N_2551);
nand U5474 (N_5474,N_2583,N_2869);
nor U5475 (N_5475,N_2808,N_2935);
or U5476 (N_5476,N_3065,N_3801);
and U5477 (N_5477,N_3935,N_3115);
and U5478 (N_5478,N_2937,N_2788);
nor U5479 (N_5479,N_2313,N_2728);
and U5480 (N_5480,N_2424,N_3846);
nand U5481 (N_5481,N_3829,N_2239);
nor U5482 (N_5482,N_2940,N_3584);
or U5483 (N_5483,N_2934,N_2941);
nor U5484 (N_5484,N_3535,N_2196);
and U5485 (N_5485,N_3328,N_3254);
or U5486 (N_5486,N_2579,N_3602);
or U5487 (N_5487,N_2883,N_3670);
nand U5488 (N_5488,N_2240,N_2664);
nand U5489 (N_5489,N_3494,N_2852);
nand U5490 (N_5490,N_3631,N_2556);
xor U5491 (N_5491,N_2949,N_3043);
or U5492 (N_5492,N_3433,N_3591);
nand U5493 (N_5493,N_2985,N_3055);
xor U5494 (N_5494,N_2593,N_3887);
nor U5495 (N_5495,N_3040,N_2357);
nor U5496 (N_5496,N_2802,N_3683);
nor U5497 (N_5497,N_2982,N_3405);
or U5498 (N_5498,N_2197,N_3553);
or U5499 (N_5499,N_2354,N_3962);
or U5500 (N_5500,N_2491,N_2252);
nor U5501 (N_5501,N_2866,N_2388);
and U5502 (N_5502,N_2269,N_3726);
nor U5503 (N_5503,N_3886,N_2358);
xnor U5504 (N_5504,N_3313,N_3706);
nor U5505 (N_5505,N_3100,N_3498);
nor U5506 (N_5506,N_2442,N_3297);
nand U5507 (N_5507,N_2874,N_2452);
nor U5508 (N_5508,N_2640,N_3925);
or U5509 (N_5509,N_2444,N_3882);
nand U5510 (N_5510,N_3801,N_2503);
nor U5511 (N_5511,N_2960,N_3115);
or U5512 (N_5512,N_3903,N_2218);
nor U5513 (N_5513,N_2530,N_3079);
or U5514 (N_5514,N_2571,N_2324);
or U5515 (N_5515,N_3145,N_2473);
nor U5516 (N_5516,N_3719,N_2637);
and U5517 (N_5517,N_2469,N_2991);
and U5518 (N_5518,N_2846,N_3612);
xor U5519 (N_5519,N_2407,N_3192);
nand U5520 (N_5520,N_3307,N_3517);
nor U5521 (N_5521,N_2218,N_2254);
and U5522 (N_5522,N_3380,N_2050);
xnor U5523 (N_5523,N_3728,N_2681);
nor U5524 (N_5524,N_3227,N_2347);
nor U5525 (N_5525,N_2705,N_3318);
and U5526 (N_5526,N_3407,N_2969);
and U5527 (N_5527,N_3056,N_3682);
or U5528 (N_5528,N_2043,N_3756);
xor U5529 (N_5529,N_3732,N_2801);
or U5530 (N_5530,N_3009,N_3908);
or U5531 (N_5531,N_2991,N_2075);
and U5532 (N_5532,N_3040,N_3447);
nor U5533 (N_5533,N_2730,N_2390);
and U5534 (N_5534,N_2625,N_3468);
or U5535 (N_5535,N_2347,N_2018);
nand U5536 (N_5536,N_2005,N_2322);
or U5537 (N_5537,N_2660,N_2369);
or U5538 (N_5538,N_3398,N_2408);
and U5539 (N_5539,N_2260,N_2663);
or U5540 (N_5540,N_3576,N_3233);
nand U5541 (N_5541,N_3356,N_3824);
nor U5542 (N_5542,N_2150,N_3734);
nand U5543 (N_5543,N_2877,N_2664);
nor U5544 (N_5544,N_3494,N_2767);
nand U5545 (N_5545,N_3421,N_2610);
nor U5546 (N_5546,N_3612,N_2188);
and U5547 (N_5547,N_3818,N_2990);
or U5548 (N_5548,N_3384,N_3066);
and U5549 (N_5549,N_3484,N_2830);
and U5550 (N_5550,N_3242,N_2527);
nand U5551 (N_5551,N_2391,N_3877);
or U5552 (N_5552,N_3606,N_3290);
or U5553 (N_5553,N_3057,N_3083);
or U5554 (N_5554,N_3764,N_3964);
or U5555 (N_5555,N_2526,N_2381);
nand U5556 (N_5556,N_2578,N_3675);
nand U5557 (N_5557,N_2695,N_2550);
and U5558 (N_5558,N_2730,N_3104);
nor U5559 (N_5559,N_3089,N_3733);
and U5560 (N_5560,N_3346,N_3896);
xnor U5561 (N_5561,N_3628,N_3048);
and U5562 (N_5562,N_3592,N_2851);
xnor U5563 (N_5563,N_3121,N_3658);
or U5564 (N_5564,N_3609,N_3790);
nand U5565 (N_5565,N_3551,N_2277);
or U5566 (N_5566,N_2768,N_2966);
nor U5567 (N_5567,N_3372,N_2389);
and U5568 (N_5568,N_2731,N_3124);
nand U5569 (N_5569,N_2806,N_2379);
and U5570 (N_5570,N_2160,N_3652);
nor U5571 (N_5571,N_3366,N_3684);
or U5572 (N_5572,N_3149,N_2141);
nor U5573 (N_5573,N_2038,N_3640);
nand U5574 (N_5574,N_2861,N_2249);
nor U5575 (N_5575,N_2231,N_2166);
and U5576 (N_5576,N_2130,N_3077);
nand U5577 (N_5577,N_3459,N_3207);
nor U5578 (N_5578,N_2410,N_3047);
and U5579 (N_5579,N_2918,N_3945);
nor U5580 (N_5580,N_2392,N_3435);
nand U5581 (N_5581,N_2707,N_3864);
nor U5582 (N_5582,N_3896,N_3398);
or U5583 (N_5583,N_2657,N_3868);
nor U5584 (N_5584,N_3718,N_2899);
nand U5585 (N_5585,N_2187,N_3577);
or U5586 (N_5586,N_3277,N_2927);
nand U5587 (N_5587,N_3722,N_3898);
and U5588 (N_5588,N_3011,N_2293);
and U5589 (N_5589,N_2023,N_3383);
xnor U5590 (N_5590,N_3219,N_2926);
nand U5591 (N_5591,N_2513,N_3280);
nor U5592 (N_5592,N_2944,N_3034);
nand U5593 (N_5593,N_2371,N_3754);
or U5594 (N_5594,N_2556,N_3654);
or U5595 (N_5595,N_2890,N_3208);
nor U5596 (N_5596,N_2761,N_3446);
nand U5597 (N_5597,N_2107,N_2369);
and U5598 (N_5598,N_2343,N_2401);
nor U5599 (N_5599,N_2840,N_2845);
or U5600 (N_5600,N_2125,N_3250);
xnor U5601 (N_5601,N_2246,N_3719);
nand U5602 (N_5602,N_3299,N_2854);
nand U5603 (N_5603,N_2458,N_2467);
nor U5604 (N_5604,N_3213,N_2043);
and U5605 (N_5605,N_3045,N_3620);
nor U5606 (N_5606,N_3771,N_2353);
nand U5607 (N_5607,N_2600,N_3911);
nand U5608 (N_5608,N_2230,N_3034);
nor U5609 (N_5609,N_2500,N_3184);
and U5610 (N_5610,N_2440,N_3691);
and U5611 (N_5611,N_2244,N_3019);
or U5612 (N_5612,N_2980,N_2507);
nand U5613 (N_5613,N_2982,N_2622);
nand U5614 (N_5614,N_3286,N_2553);
nand U5615 (N_5615,N_2670,N_3052);
xor U5616 (N_5616,N_2534,N_2304);
and U5617 (N_5617,N_3595,N_3644);
or U5618 (N_5618,N_2105,N_2494);
xor U5619 (N_5619,N_2581,N_2206);
nor U5620 (N_5620,N_3616,N_3002);
nor U5621 (N_5621,N_2173,N_2760);
and U5622 (N_5622,N_2252,N_2854);
or U5623 (N_5623,N_2740,N_3049);
or U5624 (N_5624,N_2418,N_3812);
nor U5625 (N_5625,N_3083,N_2399);
or U5626 (N_5626,N_2265,N_2981);
or U5627 (N_5627,N_3653,N_3170);
or U5628 (N_5628,N_3148,N_3128);
nand U5629 (N_5629,N_2488,N_3007);
and U5630 (N_5630,N_2082,N_3837);
nand U5631 (N_5631,N_3782,N_3891);
and U5632 (N_5632,N_3272,N_2668);
and U5633 (N_5633,N_3568,N_3473);
or U5634 (N_5634,N_2171,N_2553);
and U5635 (N_5635,N_2169,N_2176);
nand U5636 (N_5636,N_3307,N_3392);
or U5637 (N_5637,N_2559,N_2957);
nor U5638 (N_5638,N_3570,N_2540);
and U5639 (N_5639,N_2999,N_3458);
and U5640 (N_5640,N_3881,N_3908);
nand U5641 (N_5641,N_3163,N_2015);
xor U5642 (N_5642,N_3400,N_2339);
nand U5643 (N_5643,N_3953,N_3092);
and U5644 (N_5644,N_3494,N_2076);
nor U5645 (N_5645,N_2265,N_2238);
nand U5646 (N_5646,N_3252,N_3498);
nor U5647 (N_5647,N_3372,N_3922);
or U5648 (N_5648,N_3877,N_3064);
or U5649 (N_5649,N_2079,N_3604);
xnor U5650 (N_5650,N_2651,N_3622);
nor U5651 (N_5651,N_3473,N_2789);
or U5652 (N_5652,N_3268,N_2824);
or U5653 (N_5653,N_3549,N_3618);
nor U5654 (N_5654,N_3228,N_2774);
and U5655 (N_5655,N_2667,N_2910);
and U5656 (N_5656,N_2426,N_2211);
nand U5657 (N_5657,N_3476,N_3908);
and U5658 (N_5658,N_3571,N_2636);
nor U5659 (N_5659,N_3361,N_2755);
or U5660 (N_5660,N_3165,N_3788);
nand U5661 (N_5661,N_2767,N_2839);
nand U5662 (N_5662,N_3304,N_2152);
nor U5663 (N_5663,N_3804,N_2858);
xnor U5664 (N_5664,N_2343,N_3740);
or U5665 (N_5665,N_2638,N_3769);
nand U5666 (N_5666,N_2604,N_3174);
xor U5667 (N_5667,N_2081,N_3628);
and U5668 (N_5668,N_2573,N_2702);
or U5669 (N_5669,N_3884,N_2698);
and U5670 (N_5670,N_2191,N_2539);
nand U5671 (N_5671,N_2734,N_2628);
or U5672 (N_5672,N_2502,N_2023);
nand U5673 (N_5673,N_2281,N_3007);
and U5674 (N_5674,N_3454,N_2643);
nor U5675 (N_5675,N_2737,N_2869);
and U5676 (N_5676,N_2272,N_3251);
nor U5677 (N_5677,N_3320,N_3520);
or U5678 (N_5678,N_2270,N_3042);
or U5679 (N_5679,N_2693,N_3873);
and U5680 (N_5680,N_2154,N_3212);
nand U5681 (N_5681,N_2730,N_2714);
or U5682 (N_5682,N_3896,N_2788);
nand U5683 (N_5683,N_2597,N_2361);
nand U5684 (N_5684,N_2448,N_3890);
and U5685 (N_5685,N_3124,N_2314);
nor U5686 (N_5686,N_3027,N_2182);
and U5687 (N_5687,N_2165,N_3263);
and U5688 (N_5688,N_3998,N_2418);
nor U5689 (N_5689,N_2211,N_2183);
or U5690 (N_5690,N_3062,N_3726);
xnor U5691 (N_5691,N_3043,N_2132);
nor U5692 (N_5692,N_3245,N_2251);
nand U5693 (N_5693,N_2463,N_3680);
nand U5694 (N_5694,N_3929,N_3514);
and U5695 (N_5695,N_2358,N_3595);
or U5696 (N_5696,N_2403,N_3410);
and U5697 (N_5697,N_3734,N_3926);
nor U5698 (N_5698,N_3115,N_2929);
nor U5699 (N_5699,N_2433,N_2738);
nor U5700 (N_5700,N_3490,N_2403);
and U5701 (N_5701,N_2909,N_3658);
and U5702 (N_5702,N_3914,N_2983);
xor U5703 (N_5703,N_2364,N_2686);
or U5704 (N_5704,N_3050,N_3471);
or U5705 (N_5705,N_2810,N_2233);
nand U5706 (N_5706,N_3488,N_2382);
and U5707 (N_5707,N_3249,N_2258);
nor U5708 (N_5708,N_2548,N_3928);
nand U5709 (N_5709,N_3844,N_2002);
nand U5710 (N_5710,N_2975,N_3161);
nand U5711 (N_5711,N_3534,N_2880);
and U5712 (N_5712,N_2116,N_3946);
and U5713 (N_5713,N_2839,N_3665);
and U5714 (N_5714,N_3527,N_3925);
or U5715 (N_5715,N_2772,N_3967);
nand U5716 (N_5716,N_2207,N_2754);
and U5717 (N_5717,N_2291,N_2428);
nand U5718 (N_5718,N_3904,N_3725);
and U5719 (N_5719,N_2319,N_3834);
xnor U5720 (N_5720,N_2982,N_3107);
nand U5721 (N_5721,N_2654,N_3491);
nor U5722 (N_5722,N_3120,N_2560);
nand U5723 (N_5723,N_2046,N_2769);
and U5724 (N_5724,N_2794,N_2330);
xor U5725 (N_5725,N_2135,N_2008);
nor U5726 (N_5726,N_3223,N_3403);
and U5727 (N_5727,N_2808,N_3089);
nand U5728 (N_5728,N_3931,N_3346);
xor U5729 (N_5729,N_2768,N_2433);
nand U5730 (N_5730,N_3648,N_2868);
nand U5731 (N_5731,N_2000,N_2200);
nor U5732 (N_5732,N_2542,N_3057);
or U5733 (N_5733,N_2801,N_3833);
nor U5734 (N_5734,N_3955,N_3200);
nand U5735 (N_5735,N_3555,N_2889);
nor U5736 (N_5736,N_2878,N_3165);
or U5737 (N_5737,N_2570,N_3420);
or U5738 (N_5738,N_2170,N_2185);
or U5739 (N_5739,N_3095,N_2667);
nor U5740 (N_5740,N_3222,N_3658);
xnor U5741 (N_5741,N_3318,N_3030);
nor U5742 (N_5742,N_2500,N_2268);
or U5743 (N_5743,N_3295,N_2791);
and U5744 (N_5744,N_2227,N_2555);
or U5745 (N_5745,N_3445,N_2753);
xor U5746 (N_5746,N_3356,N_3567);
or U5747 (N_5747,N_3203,N_2373);
and U5748 (N_5748,N_2693,N_2939);
nor U5749 (N_5749,N_3666,N_2640);
or U5750 (N_5750,N_3921,N_3845);
nor U5751 (N_5751,N_2887,N_2126);
nor U5752 (N_5752,N_3721,N_2036);
and U5753 (N_5753,N_2959,N_3262);
xnor U5754 (N_5754,N_3248,N_3327);
and U5755 (N_5755,N_3868,N_2522);
nor U5756 (N_5756,N_3821,N_2163);
nand U5757 (N_5757,N_2396,N_2229);
nor U5758 (N_5758,N_2225,N_2390);
nor U5759 (N_5759,N_2312,N_2834);
nand U5760 (N_5760,N_2794,N_3905);
or U5761 (N_5761,N_2769,N_2530);
nand U5762 (N_5762,N_3031,N_2938);
nand U5763 (N_5763,N_3061,N_3275);
nor U5764 (N_5764,N_2592,N_2653);
xnor U5765 (N_5765,N_3337,N_3276);
nand U5766 (N_5766,N_3529,N_2476);
nand U5767 (N_5767,N_3676,N_2701);
and U5768 (N_5768,N_3241,N_2567);
nor U5769 (N_5769,N_3224,N_3605);
or U5770 (N_5770,N_3381,N_3144);
nand U5771 (N_5771,N_2855,N_2664);
or U5772 (N_5772,N_2663,N_3511);
xor U5773 (N_5773,N_3876,N_3745);
and U5774 (N_5774,N_3950,N_3330);
nand U5775 (N_5775,N_2650,N_3154);
nor U5776 (N_5776,N_3035,N_2746);
and U5777 (N_5777,N_3841,N_2511);
and U5778 (N_5778,N_3736,N_2227);
nand U5779 (N_5779,N_2077,N_2234);
or U5780 (N_5780,N_3675,N_2669);
nand U5781 (N_5781,N_2080,N_2205);
xor U5782 (N_5782,N_2765,N_3765);
or U5783 (N_5783,N_2146,N_3160);
nor U5784 (N_5784,N_3597,N_2473);
and U5785 (N_5785,N_2027,N_2623);
xor U5786 (N_5786,N_2416,N_2315);
or U5787 (N_5787,N_3469,N_2847);
xor U5788 (N_5788,N_3304,N_3951);
or U5789 (N_5789,N_3227,N_2835);
nand U5790 (N_5790,N_2121,N_3821);
or U5791 (N_5791,N_3124,N_2605);
nor U5792 (N_5792,N_2348,N_3991);
and U5793 (N_5793,N_3600,N_2670);
nand U5794 (N_5794,N_2501,N_3965);
nand U5795 (N_5795,N_3458,N_3379);
xor U5796 (N_5796,N_2336,N_2596);
xor U5797 (N_5797,N_2985,N_3232);
and U5798 (N_5798,N_2874,N_2191);
nand U5799 (N_5799,N_2659,N_3163);
and U5800 (N_5800,N_2801,N_3201);
nor U5801 (N_5801,N_2421,N_3923);
nand U5802 (N_5802,N_3584,N_3324);
nand U5803 (N_5803,N_2679,N_2544);
nand U5804 (N_5804,N_2094,N_3613);
and U5805 (N_5805,N_2552,N_3056);
or U5806 (N_5806,N_3365,N_2283);
or U5807 (N_5807,N_3506,N_2580);
and U5808 (N_5808,N_2855,N_2530);
nor U5809 (N_5809,N_2723,N_2702);
or U5810 (N_5810,N_3565,N_2552);
and U5811 (N_5811,N_3350,N_3872);
and U5812 (N_5812,N_3994,N_2487);
nor U5813 (N_5813,N_2055,N_2908);
nor U5814 (N_5814,N_2288,N_3674);
xnor U5815 (N_5815,N_3977,N_2770);
nand U5816 (N_5816,N_3186,N_2822);
or U5817 (N_5817,N_2844,N_3359);
nand U5818 (N_5818,N_2500,N_3283);
nand U5819 (N_5819,N_2757,N_3474);
and U5820 (N_5820,N_3358,N_3211);
xor U5821 (N_5821,N_3416,N_2252);
or U5822 (N_5822,N_3149,N_2131);
nor U5823 (N_5823,N_3539,N_2278);
nor U5824 (N_5824,N_3225,N_3246);
and U5825 (N_5825,N_2459,N_2592);
xor U5826 (N_5826,N_3488,N_3694);
or U5827 (N_5827,N_3767,N_3058);
nor U5828 (N_5828,N_3115,N_3426);
or U5829 (N_5829,N_2621,N_3914);
nor U5830 (N_5830,N_2077,N_3847);
or U5831 (N_5831,N_3045,N_2314);
nor U5832 (N_5832,N_3199,N_3286);
nand U5833 (N_5833,N_3107,N_2387);
nand U5834 (N_5834,N_3436,N_3583);
nor U5835 (N_5835,N_3539,N_2538);
or U5836 (N_5836,N_3695,N_2449);
nand U5837 (N_5837,N_2409,N_2334);
xnor U5838 (N_5838,N_2364,N_2541);
nand U5839 (N_5839,N_2977,N_3937);
nor U5840 (N_5840,N_2494,N_2132);
nand U5841 (N_5841,N_2460,N_2101);
or U5842 (N_5842,N_2359,N_2281);
or U5843 (N_5843,N_3565,N_3957);
nand U5844 (N_5844,N_2181,N_2485);
and U5845 (N_5845,N_2608,N_3484);
or U5846 (N_5846,N_3560,N_3833);
nand U5847 (N_5847,N_3492,N_3379);
or U5848 (N_5848,N_3210,N_3377);
nand U5849 (N_5849,N_3087,N_3953);
nand U5850 (N_5850,N_3855,N_2282);
nand U5851 (N_5851,N_2064,N_2767);
nor U5852 (N_5852,N_3191,N_3500);
and U5853 (N_5853,N_3385,N_3940);
nor U5854 (N_5854,N_2459,N_2980);
nor U5855 (N_5855,N_2154,N_3917);
and U5856 (N_5856,N_3816,N_2083);
and U5857 (N_5857,N_2234,N_2208);
nor U5858 (N_5858,N_2271,N_3222);
nor U5859 (N_5859,N_2002,N_3114);
or U5860 (N_5860,N_2985,N_3381);
and U5861 (N_5861,N_3793,N_3905);
nand U5862 (N_5862,N_2087,N_3775);
and U5863 (N_5863,N_3201,N_2595);
nand U5864 (N_5864,N_2456,N_3861);
nand U5865 (N_5865,N_2539,N_3515);
or U5866 (N_5866,N_2949,N_3353);
nor U5867 (N_5867,N_2606,N_2941);
xor U5868 (N_5868,N_3425,N_3606);
nand U5869 (N_5869,N_2271,N_2468);
nand U5870 (N_5870,N_3175,N_3755);
nand U5871 (N_5871,N_3889,N_2397);
nor U5872 (N_5872,N_2514,N_2763);
nand U5873 (N_5873,N_2702,N_2108);
and U5874 (N_5874,N_3869,N_2854);
nor U5875 (N_5875,N_3372,N_3339);
nor U5876 (N_5876,N_3380,N_2477);
nor U5877 (N_5877,N_2527,N_3847);
and U5878 (N_5878,N_2834,N_2130);
xnor U5879 (N_5879,N_3024,N_3097);
or U5880 (N_5880,N_2569,N_3210);
and U5881 (N_5881,N_3018,N_2240);
nand U5882 (N_5882,N_2763,N_3867);
and U5883 (N_5883,N_2388,N_3504);
nor U5884 (N_5884,N_3421,N_3018);
nand U5885 (N_5885,N_3141,N_3516);
or U5886 (N_5886,N_2746,N_3043);
nand U5887 (N_5887,N_2556,N_3680);
nand U5888 (N_5888,N_3934,N_2434);
xnor U5889 (N_5889,N_3256,N_3119);
or U5890 (N_5890,N_3407,N_3784);
or U5891 (N_5891,N_3562,N_3621);
or U5892 (N_5892,N_3763,N_2846);
and U5893 (N_5893,N_3408,N_3208);
or U5894 (N_5894,N_2828,N_3667);
and U5895 (N_5895,N_2617,N_2468);
and U5896 (N_5896,N_2426,N_2503);
nor U5897 (N_5897,N_2256,N_2111);
and U5898 (N_5898,N_3075,N_3796);
and U5899 (N_5899,N_2273,N_2349);
nand U5900 (N_5900,N_3764,N_2125);
and U5901 (N_5901,N_3618,N_2162);
or U5902 (N_5902,N_2257,N_2076);
or U5903 (N_5903,N_3927,N_3933);
and U5904 (N_5904,N_3213,N_2983);
xor U5905 (N_5905,N_2570,N_2913);
xnor U5906 (N_5906,N_2705,N_3626);
or U5907 (N_5907,N_2044,N_2187);
or U5908 (N_5908,N_2674,N_3139);
nor U5909 (N_5909,N_2626,N_3397);
nand U5910 (N_5910,N_2553,N_2600);
and U5911 (N_5911,N_3837,N_3782);
and U5912 (N_5912,N_3314,N_2348);
nand U5913 (N_5913,N_3362,N_2945);
nor U5914 (N_5914,N_2376,N_3838);
nand U5915 (N_5915,N_2350,N_2552);
nor U5916 (N_5916,N_3132,N_2009);
nor U5917 (N_5917,N_3371,N_3483);
xor U5918 (N_5918,N_3321,N_2054);
nand U5919 (N_5919,N_3019,N_3521);
nor U5920 (N_5920,N_2889,N_3961);
xor U5921 (N_5921,N_3867,N_2472);
nor U5922 (N_5922,N_3302,N_3608);
nor U5923 (N_5923,N_3545,N_3560);
xor U5924 (N_5924,N_3093,N_2782);
xor U5925 (N_5925,N_2159,N_3186);
and U5926 (N_5926,N_3527,N_3355);
or U5927 (N_5927,N_3778,N_3114);
nor U5928 (N_5928,N_3232,N_2682);
nor U5929 (N_5929,N_2360,N_2112);
nor U5930 (N_5930,N_2733,N_2788);
nor U5931 (N_5931,N_2656,N_3602);
or U5932 (N_5932,N_2361,N_3428);
xnor U5933 (N_5933,N_3923,N_3094);
nor U5934 (N_5934,N_2914,N_3118);
xnor U5935 (N_5935,N_3272,N_2598);
nand U5936 (N_5936,N_3139,N_2568);
and U5937 (N_5937,N_3551,N_3216);
nand U5938 (N_5938,N_3469,N_3245);
nor U5939 (N_5939,N_3779,N_2422);
or U5940 (N_5940,N_3916,N_3544);
xnor U5941 (N_5941,N_3994,N_3071);
or U5942 (N_5942,N_3893,N_2192);
nand U5943 (N_5943,N_3366,N_3143);
nor U5944 (N_5944,N_2496,N_2749);
and U5945 (N_5945,N_2158,N_2723);
and U5946 (N_5946,N_3155,N_3041);
xor U5947 (N_5947,N_3101,N_2921);
and U5948 (N_5948,N_3301,N_2471);
xnor U5949 (N_5949,N_3235,N_3617);
nor U5950 (N_5950,N_2986,N_2031);
nor U5951 (N_5951,N_3703,N_3910);
or U5952 (N_5952,N_2483,N_2273);
or U5953 (N_5953,N_3109,N_2017);
or U5954 (N_5954,N_2637,N_3417);
or U5955 (N_5955,N_3685,N_3268);
nand U5956 (N_5956,N_3760,N_3066);
xor U5957 (N_5957,N_2111,N_3464);
nand U5958 (N_5958,N_2986,N_3166);
xor U5959 (N_5959,N_2851,N_2223);
xor U5960 (N_5960,N_3839,N_3561);
or U5961 (N_5961,N_3414,N_2669);
nand U5962 (N_5962,N_3097,N_2214);
nor U5963 (N_5963,N_3220,N_2636);
and U5964 (N_5964,N_2957,N_3095);
and U5965 (N_5965,N_2341,N_2924);
xnor U5966 (N_5966,N_3802,N_2411);
nor U5967 (N_5967,N_2083,N_3089);
nor U5968 (N_5968,N_3360,N_3199);
nand U5969 (N_5969,N_2061,N_2534);
nand U5970 (N_5970,N_2817,N_3242);
or U5971 (N_5971,N_2578,N_2793);
or U5972 (N_5972,N_3037,N_2896);
nand U5973 (N_5973,N_3101,N_3092);
nand U5974 (N_5974,N_2806,N_3018);
and U5975 (N_5975,N_3337,N_3310);
xor U5976 (N_5976,N_3862,N_3796);
nor U5977 (N_5977,N_3128,N_2396);
or U5978 (N_5978,N_2942,N_3349);
nor U5979 (N_5979,N_2631,N_3807);
or U5980 (N_5980,N_3917,N_3834);
nor U5981 (N_5981,N_2980,N_3505);
and U5982 (N_5982,N_2746,N_3397);
or U5983 (N_5983,N_2478,N_3472);
nor U5984 (N_5984,N_2360,N_2338);
xor U5985 (N_5985,N_2460,N_3632);
nor U5986 (N_5986,N_3581,N_2211);
nand U5987 (N_5987,N_3810,N_2969);
nor U5988 (N_5988,N_3383,N_2977);
and U5989 (N_5989,N_2096,N_2353);
nor U5990 (N_5990,N_3257,N_2962);
nor U5991 (N_5991,N_3093,N_2320);
or U5992 (N_5992,N_3711,N_2610);
nor U5993 (N_5993,N_2868,N_2502);
and U5994 (N_5994,N_2722,N_3189);
nand U5995 (N_5995,N_3417,N_2393);
and U5996 (N_5996,N_3320,N_2622);
nand U5997 (N_5997,N_2427,N_3352);
nand U5998 (N_5998,N_3357,N_3647);
nand U5999 (N_5999,N_3168,N_2695);
nor U6000 (N_6000,N_5670,N_4102);
or U6001 (N_6001,N_4092,N_5992);
nand U6002 (N_6002,N_4011,N_5952);
and U6003 (N_6003,N_4649,N_5667);
nand U6004 (N_6004,N_4030,N_4930);
and U6005 (N_6005,N_4853,N_4432);
or U6006 (N_6006,N_4358,N_4320);
nor U6007 (N_6007,N_4577,N_4200);
nand U6008 (N_6008,N_5844,N_4059);
nand U6009 (N_6009,N_5440,N_4933);
and U6010 (N_6010,N_5086,N_5102);
and U6011 (N_6011,N_5025,N_4614);
xor U6012 (N_6012,N_4325,N_4311);
and U6013 (N_6013,N_5807,N_5292);
or U6014 (N_6014,N_5480,N_5868);
and U6015 (N_6015,N_5788,N_5057);
xor U6016 (N_6016,N_5545,N_4406);
and U6017 (N_6017,N_4694,N_4162);
nand U6018 (N_6018,N_4967,N_5023);
nand U6019 (N_6019,N_4673,N_4426);
xnor U6020 (N_6020,N_5448,N_4374);
and U6021 (N_6021,N_4107,N_4377);
xor U6022 (N_6022,N_5339,N_4443);
or U6023 (N_6023,N_4921,N_4245);
nor U6024 (N_6024,N_5192,N_5510);
nor U6025 (N_6025,N_5481,N_4344);
nor U6026 (N_6026,N_5065,N_5866);
nand U6027 (N_6027,N_4366,N_5600);
nor U6028 (N_6028,N_4462,N_5648);
nand U6029 (N_6029,N_4345,N_5218);
or U6030 (N_6030,N_5508,N_4945);
and U6031 (N_6031,N_4562,N_5161);
or U6032 (N_6032,N_5073,N_4598);
nor U6033 (N_6033,N_5454,N_4466);
nand U6034 (N_6034,N_4719,N_4353);
or U6035 (N_6035,N_4746,N_4331);
and U6036 (N_6036,N_5721,N_4919);
nor U6037 (N_6037,N_4439,N_4826);
or U6038 (N_6038,N_5553,N_5886);
and U6039 (N_6039,N_5512,N_4809);
and U6040 (N_6040,N_4517,N_4398);
nor U6041 (N_6041,N_5053,N_5944);
and U6042 (N_6042,N_4052,N_4916);
and U6043 (N_6043,N_4729,N_4646);
or U6044 (N_6044,N_5305,N_4487);
nand U6045 (N_6045,N_5706,N_5675);
nand U6046 (N_6046,N_5831,N_4101);
nand U6047 (N_6047,N_5131,N_5628);
nor U6048 (N_6048,N_5079,N_5599);
or U6049 (N_6049,N_4530,N_4913);
nand U6050 (N_6050,N_4996,N_5804);
and U6051 (N_6051,N_4096,N_4400);
nand U6052 (N_6052,N_5109,N_4832);
nand U6053 (N_6053,N_5841,N_4416);
and U6054 (N_6054,N_5496,N_5463);
or U6055 (N_6055,N_4221,N_5573);
and U6056 (N_6056,N_5296,N_5612);
nor U6057 (N_6057,N_5313,N_4015);
nor U6058 (N_6058,N_4678,N_4802);
nor U6059 (N_6059,N_4359,N_4278);
and U6060 (N_6060,N_4784,N_5040);
xor U6061 (N_6061,N_4485,N_5130);
xor U6062 (N_6062,N_5554,N_4910);
nand U6063 (N_6063,N_4733,N_4013);
and U6064 (N_6064,N_4552,N_5244);
nand U6065 (N_6065,N_5862,N_5453);
nor U6066 (N_6066,N_4493,N_4483);
nand U6067 (N_6067,N_5096,N_5605);
and U6068 (N_6068,N_5071,N_5253);
nand U6069 (N_6069,N_5124,N_4566);
xor U6070 (N_6070,N_4243,N_5252);
nor U6071 (N_6071,N_4237,N_4866);
or U6072 (N_6072,N_4363,N_4925);
or U6073 (N_6073,N_5084,N_5276);
and U6074 (N_6074,N_4189,N_5728);
or U6075 (N_6075,N_5098,N_5829);
and U6076 (N_6076,N_5591,N_5441);
nand U6077 (N_6077,N_4644,N_4988);
nand U6078 (N_6078,N_4506,N_5673);
and U6079 (N_6079,N_4137,N_4563);
nor U6080 (N_6080,N_5691,N_5877);
nor U6081 (N_6081,N_4034,N_4509);
and U6082 (N_6082,N_4260,N_5078);
and U6083 (N_6083,N_5217,N_4687);
or U6084 (N_6084,N_4434,N_5796);
nand U6085 (N_6085,N_4965,N_4968);
nor U6086 (N_6086,N_5513,N_5462);
nor U6087 (N_6087,N_5662,N_4801);
and U6088 (N_6088,N_5774,N_5215);
xor U6089 (N_6089,N_5989,N_5826);
or U6090 (N_6090,N_4078,N_5257);
nand U6091 (N_6091,N_4632,N_4149);
and U6092 (N_6092,N_5901,N_4427);
or U6093 (N_6093,N_5751,N_5621);
nor U6094 (N_6094,N_5248,N_4507);
and U6095 (N_6095,N_4732,N_4839);
and U6096 (N_6096,N_5821,N_4706);
nand U6097 (N_6097,N_5528,N_4717);
and U6098 (N_6098,N_4846,N_4159);
nand U6099 (N_6099,N_5926,N_5091);
nand U6100 (N_6100,N_4182,N_4823);
and U6101 (N_6101,N_5753,N_4389);
or U6102 (N_6102,N_4835,N_5645);
or U6103 (N_6103,N_5024,N_5747);
and U6104 (N_6104,N_4749,N_5754);
or U6105 (N_6105,N_4455,N_4753);
and U6106 (N_6106,N_4126,N_5061);
nor U6107 (N_6107,N_5939,N_4428);
and U6108 (N_6108,N_4738,N_4728);
and U6109 (N_6109,N_4272,N_5447);
or U6110 (N_6110,N_4279,N_4587);
nor U6111 (N_6111,N_4589,N_4219);
and U6112 (N_6112,N_4539,N_4519);
and U6113 (N_6113,N_5082,N_5785);
and U6114 (N_6114,N_4373,N_5711);
and U6115 (N_6115,N_5769,N_4225);
nor U6116 (N_6116,N_4583,N_4384);
nand U6117 (N_6117,N_4018,N_4019);
or U6118 (N_6118,N_5189,N_4613);
or U6119 (N_6119,N_5506,N_5050);
or U6120 (N_6120,N_5460,N_4236);
xnor U6121 (N_6121,N_5861,N_4893);
nor U6122 (N_6122,N_5163,N_4634);
nor U6123 (N_6123,N_4656,N_4847);
nor U6124 (N_6124,N_4783,N_5013);
nand U6125 (N_6125,N_4346,N_5104);
and U6126 (N_6126,N_5772,N_4870);
and U6127 (N_6127,N_4280,N_4553);
nor U6128 (N_6128,N_5731,N_5762);
nand U6129 (N_6129,N_4457,N_4037);
nand U6130 (N_6130,N_5879,N_5402);
nor U6131 (N_6131,N_5390,N_5306);
or U6132 (N_6132,N_4618,N_4548);
or U6133 (N_6133,N_4477,N_5113);
or U6134 (N_6134,N_4603,N_5727);
and U6135 (N_6135,N_5611,N_4249);
xnor U6136 (N_6136,N_5855,N_4222);
and U6137 (N_6137,N_4660,N_4799);
and U6138 (N_6138,N_4318,N_4668);
and U6139 (N_6139,N_5786,N_4025);
and U6140 (N_6140,N_5603,N_4216);
and U6141 (N_6141,N_4431,N_5887);
and U6142 (N_6142,N_4610,N_5555);
nand U6143 (N_6143,N_4172,N_5043);
and U6144 (N_6144,N_5570,N_4051);
nand U6145 (N_6145,N_4291,N_5535);
or U6146 (N_6146,N_4302,N_4565);
or U6147 (N_6147,N_4999,N_5719);
or U6148 (N_6148,N_5498,N_5968);
and U6149 (N_6149,N_5661,N_5911);
nor U6150 (N_6150,N_4240,N_4662);
xor U6151 (N_6151,N_5548,N_4873);
xnor U6152 (N_6152,N_4621,N_4557);
nor U6153 (N_6153,N_4735,N_4830);
nor U6154 (N_6154,N_4607,N_4368);
nand U6155 (N_6155,N_4737,N_4689);
and U6156 (N_6156,N_5272,N_5202);
xor U6157 (N_6157,N_4062,N_5196);
nor U6158 (N_6158,N_4760,N_5229);
nand U6159 (N_6159,N_4138,N_5461);
and U6160 (N_6160,N_5677,N_4057);
nor U6161 (N_6161,N_4622,N_5515);
or U6162 (N_6162,N_5699,N_5596);
nand U6163 (N_6163,N_5622,N_4141);
nand U6164 (N_6164,N_4765,N_5914);
and U6165 (N_6165,N_4984,N_5490);
nor U6166 (N_6166,N_5994,N_5046);
and U6167 (N_6167,N_4683,N_4265);
or U6168 (N_6168,N_4989,N_4702);
and U6169 (N_6169,N_4761,N_4212);
and U6170 (N_6170,N_5995,N_4947);
nand U6171 (N_6171,N_5795,N_4350);
and U6172 (N_6172,N_5290,N_4804);
xnor U6173 (N_6173,N_4616,N_4536);
and U6174 (N_6174,N_4827,N_4108);
or U6175 (N_6175,N_5630,N_5950);
xor U6176 (N_6176,N_4578,N_5300);
nor U6177 (N_6177,N_5544,N_5059);
nor U6178 (N_6178,N_4444,N_4424);
nand U6179 (N_6179,N_5503,N_5070);
or U6180 (N_6180,N_4874,N_4150);
xnor U6181 (N_6181,N_4667,N_5589);
and U6182 (N_6182,N_5889,N_4652);
or U6183 (N_6183,N_5108,N_4648);
and U6184 (N_6184,N_4892,N_5003);
nand U6185 (N_6185,N_5588,N_5616);
nor U6186 (N_6186,N_4542,N_5443);
nand U6187 (N_6187,N_5654,N_5167);
nor U6188 (N_6188,N_4045,N_4147);
nand U6189 (N_6189,N_5755,N_4779);
or U6190 (N_6190,N_4329,N_5316);
or U6191 (N_6191,N_5803,N_4602);
xnor U6192 (N_6192,N_5689,N_4215);
or U6193 (N_6193,N_5170,N_4355);
and U6194 (N_6194,N_4731,N_4757);
nor U6195 (N_6195,N_5761,N_4911);
nand U6196 (N_6196,N_5575,N_4135);
nor U6197 (N_6197,N_5814,N_5625);
or U6198 (N_6198,N_5107,N_4971);
or U6199 (N_6199,N_5551,N_4679);
nor U6200 (N_6200,N_4590,N_4361);
nand U6201 (N_6201,N_5429,N_4089);
nand U6202 (N_6202,N_4861,N_4768);
nor U6203 (N_6203,N_4480,N_4695);
nand U6204 (N_6204,N_4049,N_4104);
and U6205 (N_6205,N_5019,N_5343);
nand U6206 (N_6206,N_4198,N_4484);
xnor U6207 (N_6207,N_5606,N_4501);
and U6208 (N_6208,N_5372,N_5008);
xnor U6209 (N_6209,N_4187,N_5993);
nand U6210 (N_6210,N_4213,N_4588);
nor U6211 (N_6211,N_4651,N_5226);
nor U6212 (N_6212,N_5851,N_4937);
or U6213 (N_6213,N_4513,N_4633);
xnor U6214 (N_6214,N_5864,N_4824);
nor U6215 (N_6215,N_5045,N_5210);
xnor U6216 (N_6216,N_5798,N_4254);
nand U6217 (N_6217,N_4448,N_5634);
or U6218 (N_6218,N_5959,N_5004);
nand U6219 (N_6219,N_4914,N_5933);
nor U6220 (N_6220,N_5095,N_5935);
nor U6221 (N_6221,N_5367,N_5188);
xor U6222 (N_6222,N_5720,N_5847);
nand U6223 (N_6223,N_5485,N_5391);
nand U6224 (N_6224,N_4164,N_4401);
nor U6225 (N_6225,N_5876,N_5707);
nor U6226 (N_6226,N_4975,N_4849);
nor U6227 (N_6227,N_5705,N_4568);
and U6228 (N_6228,N_4540,N_4171);
nor U6229 (N_6229,N_4489,N_4756);
or U6230 (N_6230,N_5771,N_4816);
or U6231 (N_6231,N_4028,N_4008);
nand U6232 (N_6232,N_5668,N_4641);
xnor U6233 (N_6233,N_5119,N_5690);
and U6234 (N_6234,N_4617,N_5543);
nand U6235 (N_6235,N_5259,N_4039);
nor U6236 (N_6236,N_5903,N_4923);
xor U6237 (N_6237,N_4604,N_5309);
nand U6238 (N_6238,N_4379,N_4985);
and U6239 (N_6239,N_5235,N_5917);
nand U6240 (N_6240,N_5379,N_5007);
nor U6241 (N_6241,N_4258,N_5484);
xor U6242 (N_6242,N_4136,N_4357);
nor U6243 (N_6243,N_5863,N_5694);
nor U6244 (N_6244,N_4388,N_4145);
nor U6245 (N_6245,N_5414,N_4759);
xnor U6246 (N_6246,N_4956,N_5464);
xor U6247 (N_6247,N_4907,N_4356);
nand U6248 (N_6248,N_5348,N_5209);
and U6249 (N_6249,N_5934,N_4592);
nor U6250 (N_6250,N_4076,N_5805);
nand U6251 (N_6251,N_4467,N_5326);
nand U6252 (N_6252,N_5979,N_4844);
or U6253 (N_6253,N_4313,N_4825);
nand U6254 (N_6254,N_4920,N_4251);
nor U6255 (N_6255,N_4369,N_5439);
nor U6256 (N_6256,N_4814,N_4625);
and U6257 (N_6257,N_5501,N_5427);
nor U6258 (N_6258,N_4896,N_5121);
or U6259 (N_6259,N_5384,N_4098);
nor U6260 (N_6260,N_5650,N_4859);
nand U6261 (N_6261,N_4990,N_5353);
xor U6262 (N_6262,N_4567,N_5445);
nor U6263 (N_6263,N_4751,N_4954);
and U6264 (N_6264,N_5729,N_5524);
or U6265 (N_6265,N_5009,N_4421);
nor U6266 (N_6266,N_5041,N_5878);
or U6267 (N_6267,N_4772,N_5604);
nand U6268 (N_6268,N_5936,N_5155);
or U6269 (N_6269,N_4936,N_5870);
or U6270 (N_6270,N_4130,N_5001);
nand U6271 (N_6271,N_4471,N_5764);
nor U6272 (N_6272,N_4951,N_5139);
and U6273 (N_6273,N_4263,N_4569);
nand U6274 (N_6274,N_4837,N_4067);
or U6275 (N_6275,N_5976,N_4160);
nor U6276 (N_6276,N_4611,N_5468);
nand U6277 (N_6277,N_5514,N_4433);
or U6278 (N_6278,N_5981,N_5406);
and U6279 (N_6279,N_4776,N_5087);
or U6280 (N_6280,N_4273,N_5327);
nor U6281 (N_6281,N_5373,N_5444);
and U6282 (N_6282,N_5802,N_5618);
or U6283 (N_6283,N_4410,N_4606);
and U6284 (N_6284,N_4383,N_5451);
nor U6285 (N_6285,N_4054,N_4877);
and U6286 (N_6286,N_4858,N_5334);
or U6287 (N_6287,N_4447,N_5853);
nand U6288 (N_6288,N_4630,N_4420);
nor U6289 (N_6289,N_4704,N_5808);
and U6290 (N_6290,N_5476,N_5291);
nand U6291 (N_6291,N_4883,N_4643);
nor U6292 (N_6292,N_4006,N_4066);
or U6293 (N_6293,N_5197,N_5956);
nor U6294 (N_6294,N_5817,N_5710);
nor U6295 (N_6295,N_4500,N_4661);
and U6296 (N_6296,N_4571,N_4390);
nand U6297 (N_6297,N_5269,N_5146);
nor U6298 (N_6298,N_5638,N_4880);
nand U6299 (N_6299,N_5479,N_4119);
nand U6300 (N_6300,N_5255,N_4675);
nand U6301 (N_6301,N_4293,N_4033);
and U6302 (N_6302,N_5585,N_4157);
nor U6303 (N_6303,N_4942,N_5303);
nor U6304 (N_6304,N_5449,N_4232);
and U6305 (N_6305,N_4980,N_5657);
nand U6306 (N_6306,N_5093,N_4855);
nor U6307 (N_6307,N_4820,N_5062);
nand U6308 (N_6308,N_5288,N_4440);
nor U6309 (N_6309,N_4790,N_4591);
nor U6310 (N_6310,N_5322,N_4949);
and U6311 (N_6311,N_5321,N_5643);
nand U6312 (N_6312,N_5518,N_4741);
nand U6313 (N_6313,N_5295,N_4686);
nand U6314 (N_6314,N_4262,N_4798);
and U6315 (N_6315,N_4560,N_4475);
xnor U6316 (N_6316,N_4977,N_4065);
nand U6317 (N_6317,N_5308,N_4179);
nor U6318 (N_6318,N_4904,N_4669);
nand U6319 (N_6319,N_4983,N_5610);
nor U6320 (N_6320,N_5159,N_4758);
nand U6321 (N_6321,N_4304,N_5266);
nand U6322 (N_6322,N_4723,N_4183);
or U6323 (N_6323,N_4762,N_5874);
nand U6324 (N_6324,N_4796,N_4378);
xor U6325 (N_6325,N_5568,N_4438);
and U6326 (N_6326,N_4367,N_5112);
nor U6327 (N_6327,N_5247,N_5374);
nor U6328 (N_6328,N_5756,N_4123);
nand U6329 (N_6329,N_5401,N_5265);
or U6330 (N_6330,N_5712,N_5679);
or U6331 (N_6331,N_5219,N_4868);
xor U6332 (N_6332,N_5270,N_4446);
xnor U6333 (N_6333,N_5627,N_4288);
nor U6334 (N_6334,N_5442,N_5824);
or U6335 (N_6335,N_5538,N_5652);
nor U6336 (N_6336,N_5663,N_4364);
or U6337 (N_6337,N_4319,N_5651);
xnor U6338 (N_6338,N_5642,N_5016);
nor U6339 (N_6339,N_4554,N_4408);
nor U6340 (N_6340,N_4525,N_4654);
and U6341 (N_6341,N_5665,N_4450);
and U6342 (N_6342,N_4995,N_5150);
nor U6343 (N_6343,N_5176,N_4156);
or U6344 (N_6344,N_5048,N_5974);
and U6345 (N_6345,N_4125,N_4711);
nor U6346 (N_6346,N_5416,N_4218);
or U6347 (N_6347,N_4312,N_5422);
nor U6348 (N_6348,N_5845,N_4642);
xnor U6349 (N_6349,N_5032,N_5595);
or U6350 (N_6350,N_5483,N_5355);
nand U6351 (N_6351,N_4586,N_5533);
nand U6352 (N_6352,N_5058,N_5368);
nor U6353 (N_6353,N_5369,N_4274);
nand U6354 (N_6354,N_4161,N_4952);
and U6355 (N_6355,N_5649,N_5701);
nor U6356 (N_6356,N_5977,N_4908);
or U6357 (N_6357,N_5763,N_5105);
nand U6358 (N_6358,N_5629,N_5681);
or U6359 (N_6359,N_4698,N_5280);
xnor U6360 (N_6360,N_5521,N_5632);
nand U6361 (N_6361,N_4939,N_4195);
or U6362 (N_6362,N_5998,N_5283);
nor U6363 (N_6363,N_5225,N_5403);
and U6364 (N_6364,N_5659,N_5686);
nand U6365 (N_6365,N_4547,N_4998);
nor U6366 (N_6366,N_4193,N_4834);
and U6367 (N_6367,N_5475,N_5896);
or U6368 (N_6368,N_4685,N_5624);
and U6369 (N_6369,N_5325,N_4931);
nand U6370 (N_6370,N_4202,N_5819);
nor U6371 (N_6371,N_5885,N_4511);
xnor U6372 (N_6372,N_5888,N_5094);
nor U6373 (N_6373,N_4812,N_4502);
or U6374 (N_6374,N_4808,N_5825);
nand U6375 (N_6375,N_5173,N_5378);
nor U6376 (N_6376,N_4640,N_4255);
nor U6377 (N_6377,N_4710,N_5672);
and U6378 (N_6378,N_5574,N_5471);
nand U6379 (N_6379,N_5399,N_4865);
or U6380 (N_6380,N_5973,N_4918);
nor U6381 (N_6381,N_5848,N_4142);
nand U6382 (N_6382,N_4397,N_5738);
xnor U6383 (N_6383,N_5818,N_4214);
and U6384 (N_6384,N_4958,N_5787);
nor U6385 (N_6385,N_5386,N_4974);
nor U6386 (N_6386,N_4680,N_4112);
or U6387 (N_6387,N_4653,N_4626);
nand U6388 (N_6388,N_4692,N_5012);
and U6389 (N_6389,N_5740,N_5777);
and U6390 (N_6390,N_5773,N_4442);
nand U6391 (N_6391,N_4664,N_5636);
or U6392 (N_6392,N_5647,N_5069);
and U6393 (N_6393,N_5609,N_5482);
and U6394 (N_6394,N_5988,N_5264);
xor U6395 (N_6395,N_4774,N_4414);
nand U6396 (N_6396,N_4290,N_4572);
nand U6397 (N_6397,N_4370,N_4516);
nor U6398 (N_6398,N_4780,N_5274);
xnor U6399 (N_6399,N_4600,N_5838);
and U6400 (N_6400,N_5990,N_4556);
nor U6401 (N_6401,N_4890,N_4575);
nand U6402 (N_6402,N_4842,N_4863);
nand U6403 (N_6403,N_5493,N_4479);
and U6404 (N_6404,N_4038,N_4724);
nand U6405 (N_6405,N_4789,N_4806);
nor U6406 (N_6406,N_4982,N_4003);
nand U6407 (N_6407,N_4481,N_4340);
xor U6408 (N_6408,N_4310,N_4470);
and U6409 (N_6409,N_5592,N_5597);
xnor U6410 (N_6410,N_5465,N_5117);
xor U6411 (N_6411,N_5867,N_5983);
nor U6412 (N_6412,N_4259,N_4884);
or U6413 (N_6413,N_4095,N_4869);
nor U6414 (N_6414,N_5986,N_4701);
nand U6415 (N_6415,N_5669,N_4385);
xor U6416 (N_6416,N_4058,N_5431);
nor U6417 (N_6417,N_5921,N_5033);
nor U6418 (N_6418,N_5230,N_5972);
or U6419 (N_6419,N_5232,N_4528);
nor U6420 (N_6420,N_5797,N_5458);
nor U6421 (N_6421,N_4336,N_4453);
nand U6422 (N_6422,N_5947,N_4518);
nand U6423 (N_6423,N_5810,N_4194);
or U6424 (N_6424,N_4026,N_4029);
or U6425 (N_6425,N_5608,N_4301);
xnor U6426 (N_6426,N_5347,N_5351);
nor U6427 (N_6427,N_5893,N_4393);
nor U6428 (N_6428,N_4793,N_4561);
nand U6429 (N_6429,N_4449,N_4227);
or U6430 (N_6430,N_4253,N_4636);
nor U6431 (N_6431,N_4878,N_4520);
or U6432 (N_6432,N_4168,N_5338);
nor U6433 (N_6433,N_5122,N_5822);
and U6434 (N_6434,N_4508,N_5766);
nor U6435 (N_6435,N_4430,N_4209);
nor U6436 (N_6436,N_5038,N_4286);
xor U6437 (N_6437,N_4697,N_5915);
and U6438 (N_6438,N_4053,N_4360);
and U6439 (N_6439,N_4707,N_4871);
nand U6440 (N_6440,N_4551,N_4122);
nand U6441 (N_6441,N_4088,N_5026);
xnor U6442 (N_6442,N_5948,N_4852);
xnor U6443 (N_6443,N_4371,N_5450);
nand U6444 (N_6444,N_4787,N_5341);
and U6445 (N_6445,N_5587,N_4682);
nor U6446 (N_6446,N_5897,N_4307);
and U6447 (N_6447,N_5030,N_4792);
nor U6448 (N_6448,N_5671,N_5298);
or U6449 (N_6449,N_5172,N_5421);
and U6450 (N_6450,N_4332,N_5164);
and U6451 (N_6451,N_4581,N_5700);
nand U6452 (N_6452,N_4022,N_4843);
xor U6453 (N_6453,N_5268,N_4409);
and U6454 (N_6454,N_5066,N_4817);
nand U6455 (N_6455,N_4811,N_5310);
nand U6456 (N_6456,N_5835,N_5037);
nand U6457 (N_6457,N_4238,N_4014);
xnor U6458 (N_6458,N_4217,N_5660);
nor U6459 (N_6459,N_5913,N_5836);
or U6460 (N_6460,N_4545,N_4337);
and U6461 (N_6461,N_5278,N_5405);
nand U6462 (N_6462,N_4615,N_5800);
nand U6463 (N_6463,N_4620,N_5615);
and U6464 (N_6464,N_4382,N_4867);
or U6465 (N_6465,N_5491,N_5285);
xor U6466 (N_6466,N_5881,N_5426);
or U6467 (N_6467,N_5181,N_5626);
and U6468 (N_6468,N_5584,N_5183);
nor U6469 (N_6469,N_4016,N_5722);
and U6470 (N_6470,N_4645,N_4308);
nor U6471 (N_6471,N_5531,N_4693);
or U6472 (N_6472,N_5745,N_4754);
or U6473 (N_6473,N_5466,N_5193);
nor U6474 (N_6474,N_4978,N_4206);
nand U6475 (N_6475,N_4419,N_4314);
xnor U6476 (N_6476,N_4010,N_4836);
nand U6477 (N_6477,N_4392,N_4208);
xnor U6478 (N_6478,N_4742,N_4534);
xnor U6479 (N_6479,N_5143,N_4103);
nand U6480 (N_6480,N_4872,N_5891);
nor U6481 (N_6481,N_4856,N_5567);
nand U6482 (N_6482,N_5653,N_4056);
or U6483 (N_6483,N_4231,N_5221);
or U6484 (N_6484,N_4663,N_5175);
nor U6485 (N_6485,N_5145,N_4167);
nor U6486 (N_6486,N_5582,N_4838);
and U6487 (N_6487,N_4321,N_5415);
nand U6488 (N_6488,N_5237,N_5101);
nand U6489 (N_6489,N_5100,N_5340);
or U6490 (N_6490,N_5171,N_5558);
xor U6491 (N_6491,N_5502,N_5577);
or U6492 (N_6492,N_4128,N_4417);
or U6493 (N_6493,N_4326,N_5495);
and U6494 (N_6494,N_5141,N_5909);
nand U6495 (N_6495,N_5277,N_5907);
or U6496 (N_6496,N_5494,N_4987);
nor U6497 (N_6497,N_4372,N_5942);
xnor U6498 (N_6498,N_5397,N_4478);
and U6499 (N_6499,N_4476,N_5412);
xor U6500 (N_6500,N_5961,N_5579);
or U6501 (N_6501,N_5200,N_4177);
or U6502 (N_6502,N_5035,N_5564);
nand U6503 (N_6503,N_4073,N_5837);
or U6504 (N_6504,N_4570,N_5191);
nand U6505 (N_6505,N_5980,N_5828);
nor U6506 (N_6506,N_4953,N_4124);
or U6507 (N_6507,N_4743,N_4229);
and U6508 (N_6508,N_5790,N_4897);
and U6509 (N_6509,N_4396,N_4418);
nor U6510 (N_6510,N_5331,N_5261);
nand U6511 (N_6511,N_5433,N_5083);
xor U6512 (N_6512,N_4496,N_5457);
and U6513 (N_6513,N_4468,N_4786);
nor U6514 (N_6514,N_5299,N_4647);
xor U6515 (N_6515,N_5906,N_5438);
nand U6516 (N_6516,N_5613,N_4474);
or U6517 (N_6517,N_4185,N_4174);
or U6518 (N_6518,N_4031,N_4807);
nor U6519 (N_6519,N_5750,N_5931);
nor U6520 (N_6520,N_5080,N_4559);
and U6521 (N_6521,N_4233,N_5975);
nor U6522 (N_6522,N_5254,N_5256);
and U6523 (N_6523,N_5865,N_4699);
xor U6524 (N_6524,N_4887,N_4458);
and U6525 (N_6525,N_4579,N_4411);
nand U6526 (N_6526,N_5063,N_4635);
or U6527 (N_6527,N_4097,N_4081);
and U6528 (N_6528,N_4129,N_4009);
and U6529 (N_6529,N_5811,N_5898);
nor U6530 (N_6530,N_5525,N_5206);
nand U6531 (N_6531,N_5704,N_5946);
nor U6532 (N_6532,N_4000,N_5644);
or U6533 (N_6533,N_4079,N_5938);
nor U6534 (N_6534,N_5923,N_4241);
nor U6535 (N_6535,N_4690,N_5364);
nor U6536 (N_6536,N_5530,N_5034);
nor U6537 (N_6537,N_5216,N_5850);
nor U6538 (N_6538,N_4805,N_4086);
nand U6539 (N_6539,N_4387,N_5598);
and U6540 (N_6540,N_5469,N_4558);
or U6541 (N_6541,N_4001,N_5735);
or U6542 (N_6542,N_5039,N_5149);
or U6543 (N_6543,N_4188,N_4317);
nand U6544 (N_6544,N_5852,N_4504);
nand U6545 (N_6545,N_5162,N_4785);
or U6546 (N_6546,N_4955,N_5869);
or U6547 (N_6547,N_4061,N_4845);
nor U6548 (N_6548,N_5128,N_5581);
nand U6549 (N_6549,N_4170,N_5736);
or U6550 (N_6550,N_5580,N_5954);
nor U6551 (N_6551,N_4048,N_5920);
nor U6552 (N_6552,N_5781,N_4526);
or U6553 (N_6553,N_5151,N_5383);
nor U6554 (N_6554,N_5474,N_4599);
and U6555 (N_6555,N_5859,N_4461);
or U6556 (N_6556,N_4800,N_4854);
xor U6557 (N_6557,N_5178,N_5715);
nor U6558 (N_6558,N_4349,N_5919);
or U6559 (N_6559,N_5044,N_4175);
nand U6560 (N_6560,N_5180,N_4275);
nor U6561 (N_6561,N_4531,N_4778);
nand U6562 (N_6562,N_5488,N_5420);
and U6563 (N_6563,N_5546,N_5077);
and U6564 (N_6564,N_5791,N_4303);
and U6565 (N_6565,N_4864,N_4541);
xnor U6566 (N_6566,N_5036,N_4163);
or U6567 (N_6567,N_4109,N_4072);
nor U6568 (N_6568,N_5714,N_5963);
xnor U6569 (N_6569,N_4684,N_5526);
nor U6570 (N_6570,N_5054,N_5741);
nor U6571 (N_6571,N_4334,N_4220);
nor U6572 (N_6572,N_4084,N_4060);
xor U6573 (N_6573,N_4234,N_4099);
or U6574 (N_6574,N_5987,N_5446);
nand U6575 (N_6575,N_5144,N_5177);
and U6576 (N_6576,N_5425,N_5072);
nor U6577 (N_6577,N_5435,N_4494);
and U6578 (N_6578,N_4451,N_4752);
nand U6579 (N_6579,N_5231,N_5060);
and U6580 (N_6580,N_5246,N_4903);
nor U6581 (N_6581,N_4862,N_5860);
or U6582 (N_6582,N_4691,N_5168);
nor U6583 (N_6583,N_5970,N_4464);
and U6584 (N_6584,N_4268,N_5569);
or U6585 (N_6585,N_4422,N_5815);
xor U6586 (N_6586,N_5111,N_4726);
nand U6587 (N_6587,N_5536,N_4248);
nor U6588 (N_6588,N_4505,N_4205);
or U6589 (N_6589,N_5724,N_4585);
nor U6590 (N_6590,N_5014,N_4573);
nand U6591 (N_6591,N_4722,N_5011);
nand U6592 (N_6592,N_5294,N_5408);
or U6593 (N_6593,N_5284,N_5090);
and U6594 (N_6594,N_4395,N_5213);
or U6595 (N_6595,N_4950,N_4328);
nand U6596 (N_6596,N_5693,N_5241);
nor U6597 (N_6597,N_5487,N_4899);
or U6598 (N_6598,N_5359,N_4375);
nor U6599 (N_6599,N_4744,N_4252);
nand U6600 (N_6600,N_5842,N_5335);
or U6601 (N_6601,N_4323,N_4981);
or U6602 (N_6602,N_5388,N_5153);
or U6603 (N_6603,N_5097,N_5583);
nor U6604 (N_6604,N_4239,N_5262);
xor U6605 (N_6605,N_5413,N_5801);
nand U6606 (N_6606,N_5392,N_4169);
nor U6607 (N_6607,N_4224,N_4180);
or U6608 (N_6608,N_5744,N_4782);
nor U6609 (N_6609,N_4889,N_4544);
xnor U6610 (N_6610,N_4376,N_5547);
nand U6611 (N_6611,N_4718,N_4339);
and U6612 (N_6612,N_4829,N_4549);
and U6613 (N_6613,N_4972,N_5717);
and U6614 (N_6614,N_4927,N_5398);
nand U6615 (N_6615,N_5138,N_5430);
nand U6616 (N_6616,N_4075,N_5436);
or U6617 (N_6617,N_5002,N_5937);
or U6618 (N_6618,N_5725,N_4004);
xor U6619 (N_6619,N_5382,N_4495);
nor U6620 (N_6620,N_4007,N_5778);
nand U6621 (N_6621,N_5830,N_5472);
or U6622 (N_6622,N_5932,N_4244);
and U6623 (N_6623,N_4550,N_4860);
nand U6624 (N_6624,N_4196,N_4810);
nor U6625 (N_6625,N_4210,N_4445);
and U6626 (N_6626,N_5233,N_4623);
nand U6627 (N_6627,N_5214,N_5456);
xnor U6628 (N_6628,N_5195,N_5984);
and U6629 (N_6629,N_4204,N_5813);
nor U6630 (N_6630,N_5027,N_4902);
and U6631 (N_6631,N_4247,N_5238);
or U6632 (N_6632,N_5301,N_4524);
nand U6633 (N_6633,N_5511,N_4962);
nor U6634 (N_6634,N_5319,N_4909);
or U6635 (N_6635,N_5563,N_5623);
nand U6636 (N_6636,N_4270,N_4771);
nor U6637 (N_6637,N_4386,N_4938);
or U6638 (N_6638,N_4659,N_4969);
nor U6639 (N_6639,N_5251,N_5275);
nor U6640 (N_6640,N_5519,N_4333);
nand U6641 (N_6641,N_4881,N_4935);
or U6642 (N_6642,N_5832,N_4399);
and U6643 (N_6643,N_5419,N_5198);
xnor U6644 (N_6644,N_4402,N_5165);
or U6645 (N_6645,N_5884,N_5875);
nor U6646 (N_6646,N_4134,N_4619);
nand U6647 (N_6647,N_4677,N_4658);
or U6648 (N_6648,N_5344,N_4117);
nand U6649 (N_6649,N_4412,N_4282);
nor U6650 (N_6650,N_5930,N_4605);
nor U6651 (N_6651,N_4341,N_4192);
nand U6652 (N_6652,N_4223,N_4584);
or U6653 (N_6653,N_5185,N_5208);
and U6654 (N_6654,N_5212,N_4672);
nor U6655 (N_6655,N_4730,N_4482);
xnor U6656 (N_6656,N_5540,N_4973);
nand U6657 (N_6657,N_5949,N_4297);
and U6658 (N_6658,N_4083,N_4354);
nand U6659 (N_6659,N_5417,N_5918);
xnor U6660 (N_6660,N_4797,N_5330);
nand U6661 (N_6661,N_5356,N_4638);
nand U6662 (N_6662,N_5106,N_5179);
and U6663 (N_6663,N_5542,N_5697);
nand U6664 (N_6664,N_5021,N_4281);
and U6665 (N_6665,N_5201,N_4875);
nor U6666 (N_6666,N_5539,N_4404);
or U6667 (N_6667,N_5953,N_5590);
nand U6668 (N_6668,N_5571,N_4242);
or U6669 (N_6669,N_5962,N_5158);
and U6670 (N_6670,N_5666,N_4121);
nand U6671 (N_6671,N_5680,N_4041);
nand U6672 (N_6672,N_4437,N_4093);
xnor U6673 (N_6673,N_5263,N_5115);
nand U6674 (N_6674,N_4514,N_5357);
nor U6675 (N_6675,N_5137,N_5267);
and U6676 (N_6676,N_5955,N_5646);
or U6677 (N_6677,N_4503,N_5380);
nand U6678 (N_6678,N_4963,N_4696);
nor U6679 (N_6679,N_5236,N_4555);
xor U6680 (N_6680,N_4077,N_4486);
or U6681 (N_6681,N_5220,N_5748);
nand U6682 (N_6682,N_4322,N_5056);
or U6683 (N_6683,N_5696,N_5997);
nor U6684 (N_6684,N_5234,N_4069);
nor U6685 (N_6685,N_5127,N_4499);
nor U6686 (N_6686,N_5509,N_5240);
or U6687 (N_6687,N_5996,N_4090);
nand U6688 (N_6688,N_4199,N_4891);
nand U6689 (N_6689,N_4957,N_4144);
nor U6690 (N_6690,N_5929,N_4885);
and U6691 (N_6691,N_5370,N_5194);
or U6692 (N_6692,N_4739,N_5051);
nand U6693 (N_6693,N_5849,N_5812);
nor U6694 (N_6694,N_5396,N_4250);
nor U6695 (N_6695,N_5132,N_5110);
nor U6696 (N_6696,N_4498,N_5418);
nand U6697 (N_6697,N_4324,N_4068);
or U6698 (N_6698,N_4721,N_4715);
or U6699 (N_6699,N_4803,N_4943);
nand U6700 (N_6700,N_4023,N_5187);
nand U6701 (N_6701,N_5752,N_4639);
and U6702 (N_6702,N_5840,N_5562);
and U6703 (N_6703,N_5809,N_5991);
and U6704 (N_6704,N_4627,N_5892);
or U6705 (N_6705,N_5927,N_5074);
or U6706 (N_6706,N_5739,N_5537);
nand U6707 (N_6707,N_4991,N_5204);
nand U6708 (N_6708,N_4795,N_5352);
or U6709 (N_6709,N_4841,N_5000);
nor U6710 (N_6710,N_4287,N_4986);
nor U6711 (N_6711,N_5010,N_4094);
nand U6712 (N_6712,N_5730,N_4298);
nand U6713 (N_6713,N_4284,N_5969);
or U6714 (N_6714,N_5366,N_4655);
nand U6715 (N_6715,N_5088,N_4289);
nand U6716 (N_6716,N_4681,N_4497);
xnor U6717 (N_6717,N_4813,N_5223);
nor U6718 (N_6718,N_5779,N_4405);
and U6719 (N_6719,N_5806,N_4533);
and U6720 (N_6720,N_4012,N_4966);
and U6721 (N_6721,N_4351,N_4926);
nand U6722 (N_6722,N_5905,N_4044);
or U6723 (N_6723,N_4436,N_4888);
nand U6724 (N_6724,N_5478,N_4674);
or U6725 (N_6725,N_5081,N_5504);
or U6726 (N_6726,N_4197,N_4113);
or U6727 (N_6727,N_5982,N_4593);
xnor U6728 (N_6728,N_4612,N_5678);
nand U6729 (N_6729,N_5978,N_4465);
nand U6730 (N_6730,N_5311,N_4292);
and U6731 (N_6731,N_5297,N_5064);
nand U6732 (N_6732,N_5857,N_5375);
and U6733 (N_6733,N_5925,N_5228);
nand U6734 (N_6734,N_5363,N_5839);
and U6735 (N_6735,N_4050,N_5092);
nor U6736 (N_6736,N_5685,N_5260);
nor U6737 (N_6737,N_4922,N_5674);
nor U6738 (N_6738,N_5523,N_4201);
nor U6739 (N_6739,N_5602,N_4211);
and U6740 (N_6740,N_4002,N_4934);
and U6741 (N_6741,N_5068,N_4111);
nand U6742 (N_6742,N_4929,N_4788);
nor U6743 (N_6743,N_5637,N_4960);
nor U6744 (N_6744,N_4700,N_5307);
nand U6745 (N_6745,N_5395,N_5134);
or U6746 (N_6746,N_5902,N_5273);
and U6747 (N_6747,N_5186,N_5890);
xor U6748 (N_6748,N_5042,N_5965);
or U6749 (N_6749,N_4940,N_5641);
and U6750 (N_6750,N_5732,N_5529);
nand U6751 (N_6751,N_5682,N_4348);
and U6752 (N_6752,N_5656,N_4173);
and U6753 (N_6753,N_4105,N_4415);
and U6754 (N_6754,N_4347,N_5639);
or U6755 (N_6755,N_4527,N_4488);
nand U6756 (N_6756,N_5578,N_4979);
or U6757 (N_6757,N_4708,N_5489);
nand U6758 (N_6758,N_5709,N_5028);
nor U6759 (N_6759,N_4133,N_4491);
and U6760 (N_6760,N_5289,N_5614);
nor U6761 (N_6761,N_5174,N_5318);
or U6762 (N_6762,N_4764,N_5620);
or U6763 (N_6763,N_4665,N_5549);
and U6764 (N_6764,N_5089,N_4454);
and U6765 (N_6765,N_5015,N_5916);
nor U6766 (N_6766,N_5393,N_4155);
nor U6767 (N_6767,N_5967,N_5792);
nor U6768 (N_6768,N_5345,N_4035);
nor U6769 (N_6769,N_5723,N_5854);
or U6770 (N_6770,N_5757,N_4763);
nor U6771 (N_6771,N_5133,N_5286);
nand U6772 (N_6772,N_5816,N_5452);
or U6773 (N_6773,N_4261,N_5103);
and U6774 (N_6774,N_4970,N_5958);
or U6775 (N_6775,N_5635,N_4781);
xor U6776 (N_6776,N_4459,N_5361);
or U6777 (N_6777,N_4898,N_4176);
and U6778 (N_6778,N_4535,N_5320);
nand U6779 (N_6779,N_5249,N_5827);
nor U6780 (N_6780,N_5142,N_4748);
xnor U6781 (N_6781,N_5895,N_4676);
or U6782 (N_6782,N_4257,N_4352);
nor U6783 (N_6783,N_4184,N_4720);
and U6784 (N_6784,N_5565,N_5302);
and U6785 (N_6785,N_5767,N_5550);
nand U6786 (N_6786,N_4305,N_5776);
and U6787 (N_6787,N_5619,N_4522);
and U6788 (N_6788,N_4315,N_5843);
nor U6789 (N_6789,N_5031,N_4879);
nor U6790 (N_6790,N_5780,N_4948);
nand U6791 (N_6791,N_4595,N_5943);
or U6792 (N_6792,N_5640,N_5499);
nand U6793 (N_6793,N_5410,N_5467);
xnor U6794 (N_6794,N_4851,N_4127);
or U6795 (N_6795,N_5698,N_5293);
nor U6796 (N_6796,N_5607,N_5354);
or U6797 (N_6797,N_5349,N_4857);
nand U6798 (N_6798,N_4609,N_4624);
or U6799 (N_6799,N_5067,N_5250);
nor U6800 (N_6800,N_5434,N_5928);
or U6801 (N_6801,N_5336,N_5957);
nor U6802 (N_6802,N_4166,N_5075);
and U6803 (N_6803,N_5742,N_5085);
or U6804 (N_6804,N_4564,N_5017);
nand U6805 (N_6805,N_4190,N_4734);
and U6806 (N_6806,N_4523,N_5703);
or U6807 (N_6807,N_4828,N_4532);
and U6808 (N_6808,N_5020,N_4766);
and U6809 (N_6809,N_5099,N_5586);
nor U6810 (N_6810,N_4670,N_5424);
or U6811 (N_6811,N_4992,N_5055);
and U6812 (N_6812,N_4203,N_4146);
nor U6813 (N_6813,N_5522,N_4071);
nor U6814 (N_6814,N_5423,N_4153);
nor U6815 (N_6815,N_4713,N_5005);
or U6816 (N_6816,N_5116,N_4688);
nand U6817 (N_6817,N_5737,N_4131);
or U6818 (N_6818,N_4120,N_4714);
and U6819 (N_6819,N_4021,N_5473);
nor U6820 (N_6820,N_5157,N_5702);
or U6821 (N_6821,N_5317,N_4906);
nand U6822 (N_6822,N_5601,N_5125);
and U6823 (N_6823,N_4596,N_4380);
nor U6824 (N_6824,N_5169,N_4608);
xnor U6825 (N_6825,N_5683,N_4894);
or U6826 (N_6826,N_5971,N_4178);
xor U6827 (N_6827,N_5794,N_5135);
nand U6828 (N_6828,N_5633,N_4895);
nand U6829 (N_6829,N_5820,N_5594);
xnor U6830 (N_6830,N_5360,N_4574);
xor U6831 (N_6831,N_4330,N_5455);
nor U6832 (N_6832,N_4327,N_5470);
nor U6833 (N_6833,N_4594,N_5716);
and U6834 (N_6834,N_5784,N_4005);
nand U6835 (N_6835,N_4158,N_5904);
nand U6836 (N_6836,N_4946,N_5566);
and U6837 (N_6837,N_4546,N_5328);
nor U6838 (N_6838,N_5880,N_4912);
or U6839 (N_6839,N_4961,N_5910);
or U6840 (N_6840,N_5541,N_5557);
nand U6841 (N_6841,N_4151,N_5520);
nand U6842 (N_6842,N_5258,N_5224);
or U6843 (N_6843,N_4460,N_4381);
and U6844 (N_6844,N_5492,N_4228);
and U6845 (N_6845,N_4650,N_5765);
nor U6846 (N_6846,N_4047,N_5951);
nand U6847 (N_6847,N_5695,N_5516);
and U6848 (N_6848,N_5966,N_4063);
nand U6849 (N_6849,N_4152,N_5243);
nand U6850 (N_6850,N_5687,N_4819);
and U6851 (N_6851,N_5329,N_4472);
nor U6852 (N_6852,N_5655,N_5676);
nand U6853 (N_6853,N_4343,N_4391);
or U6854 (N_6854,N_4024,N_5734);
nor U6855 (N_6855,N_5156,N_4087);
nor U6856 (N_6856,N_4628,N_5411);
nor U6857 (N_6857,N_5324,N_5126);
and U6858 (N_6858,N_5823,N_5658);
or U6859 (N_6859,N_5076,N_5517);
or U6860 (N_6860,N_5140,N_5534);
nand U6861 (N_6861,N_4959,N_4976);
nand U6862 (N_6862,N_4207,N_4055);
nand U6863 (N_6863,N_5783,N_5350);
or U6864 (N_6864,N_5199,N_4267);
nor U6865 (N_6865,N_5505,N_5486);
nand U6866 (N_6866,N_4091,N_4080);
or U6867 (N_6867,N_5407,N_5572);
nor U6868 (N_6868,N_4256,N_4705);
nor U6869 (N_6869,N_4473,N_5304);
or U6870 (N_6870,N_4070,N_4521);
nand U6871 (N_6871,N_5497,N_5775);
nor U6872 (N_6872,N_5985,N_5560);
nor U6873 (N_6873,N_5782,N_5377);
nand U6874 (N_6874,N_4043,N_5271);
and U6875 (N_6875,N_4815,N_4543);
and U6876 (N_6876,N_5912,N_4423);
or U6877 (N_6877,N_4818,N_5708);
and U6878 (N_6878,N_5692,N_5856);
nor U6879 (N_6879,N_4601,N_5337);
and U6880 (N_6880,N_4736,N_5314);
xnor U6881 (N_6881,N_4703,N_5371);
and U6882 (N_6882,N_4582,N_5207);
and U6883 (N_6883,N_4299,N_4492);
nor U6884 (N_6884,N_4271,N_4725);
or U6885 (N_6885,N_5561,N_4032);
nand U6886 (N_6886,N_4106,N_5160);
or U6887 (N_6887,N_4394,N_5222);
nor U6888 (N_6888,N_5123,N_4115);
nor U6889 (N_6889,N_4512,N_4266);
xor U6890 (N_6890,N_4490,N_4901);
xnor U6891 (N_6891,N_5279,N_5631);
nor U6892 (N_6892,N_5894,N_4510);
and U6893 (N_6893,N_5924,N_5726);
xor U6894 (N_6894,N_4747,N_4040);
nand U6895 (N_6895,N_5190,N_5385);
or U6896 (N_6896,N_5459,N_5428);
nor U6897 (N_6897,N_5733,N_4017);
and U6898 (N_6898,N_5148,N_5908);
nand U6899 (N_6899,N_5400,N_5559);
or U6900 (N_6900,N_5047,N_4148);
or U6901 (N_6901,N_4456,N_5018);
or U6902 (N_6902,N_4657,N_5203);
nor U6903 (N_6903,N_4666,N_4139);
nor U6904 (N_6904,N_5960,N_4769);
xor U6905 (N_6905,N_4082,N_5684);
or U6906 (N_6906,N_4629,N_5999);
xor U6907 (N_6907,N_5552,N_4100);
xnor U6908 (N_6908,N_4709,N_4316);
nor U6909 (N_6909,N_5789,N_4745);
and U6910 (N_6910,N_5768,N_5507);
nand U6911 (N_6911,N_4283,N_4306);
nand U6912 (N_6912,N_4294,N_4309);
and U6913 (N_6913,N_4132,N_5758);
xor U6914 (N_6914,N_4775,N_4074);
or U6915 (N_6915,N_4529,N_5900);
nand U6916 (N_6916,N_5746,N_4773);
nor U6917 (N_6917,N_4295,N_4848);
or U6918 (N_6918,N_5749,N_5282);
nand U6919 (N_6919,N_5688,N_4822);
and U6920 (N_6920,N_4143,N_4924);
and U6921 (N_6921,N_5940,N_5287);
and U6922 (N_6922,N_4085,N_4191);
or U6923 (N_6923,N_5394,N_5205);
nand U6924 (N_6924,N_5846,N_5152);
or U6925 (N_6925,N_4932,N_4755);
nor U6926 (N_6926,N_4767,N_4230);
nand U6927 (N_6927,N_4064,N_4821);
or U6928 (N_6928,N_5281,N_4915);
and U6929 (N_6929,N_4365,N_5333);
nor U6930 (N_6930,N_4850,N_4338);
xor U6931 (N_6931,N_4046,N_4269);
nor U6932 (N_6932,N_5129,N_5899);
or U6933 (N_6933,N_4186,N_5049);
and U6934 (N_6934,N_4840,N_5713);
nand U6935 (N_6935,N_4463,N_5362);
nor U6936 (N_6936,N_4917,N_5147);
nor U6937 (N_6937,N_5437,N_4403);
nand U6938 (N_6938,N_4435,N_4425);
nand U6939 (N_6939,N_4777,N_5404);
or U6940 (N_6940,N_4335,N_5312);
and U6941 (N_6941,N_5022,N_5387);
nor U6942 (N_6942,N_4671,N_5964);
xor U6943 (N_6943,N_4712,N_5593);
or U6944 (N_6944,N_4276,N_5365);
xor U6945 (N_6945,N_4165,N_4794);
nand U6946 (N_6946,N_4637,N_5532);
nand U6947 (N_6947,N_4576,N_5184);
or U6948 (N_6948,N_5432,N_5743);
nand U6949 (N_6949,N_5664,N_5052);
nor U6950 (N_6950,N_5006,N_4441);
or U6951 (N_6951,N_5477,N_4235);
or U6952 (N_6952,N_4413,N_5136);
and U6953 (N_6953,N_4452,N_5760);
nor U6954 (N_6954,N_4886,N_4140);
nand U6955 (N_6955,N_5834,N_5858);
or U6956 (N_6956,N_4833,N_5381);
and U6957 (N_6957,N_5793,N_5770);
nand U6958 (N_6958,N_4110,N_5245);
or U6959 (N_6959,N_4118,N_5376);
or U6960 (N_6960,N_4300,N_5120);
or U6961 (N_6961,N_4407,N_5166);
and U6962 (N_6962,N_4362,N_5617);
and U6963 (N_6963,N_5118,N_5211);
nand U6964 (N_6964,N_4538,N_4941);
nand U6965 (N_6965,N_4226,N_4580);
nor U6966 (N_6966,N_4631,N_5883);
nand U6967 (N_6967,N_4770,N_5941);
nand U6968 (N_6968,N_4246,N_4285);
nor U6969 (N_6969,N_4469,N_4036);
nand U6970 (N_6970,N_4964,N_5556);
nand U6971 (N_6971,N_4928,N_4727);
or U6972 (N_6972,N_4882,N_4537);
and U6973 (N_6973,N_4597,N_5346);
nor U6974 (N_6974,N_4831,N_5799);
and U6975 (N_6975,N_4900,N_5527);
or U6976 (N_6976,N_5242,N_5323);
nor U6977 (N_6977,N_5718,N_5154);
and U6978 (N_6978,N_4027,N_4042);
or U6979 (N_6979,N_5239,N_4716);
and U6980 (N_6980,N_5872,N_5358);
xnor U6981 (N_6981,N_4116,N_4993);
nor U6982 (N_6982,N_5029,N_4876);
nor U6983 (N_6983,N_4181,N_5227);
nand U6984 (N_6984,N_4905,N_5182);
or U6985 (N_6985,N_4740,N_5873);
xor U6986 (N_6986,N_4429,N_5500);
or U6987 (N_6987,N_4994,N_4750);
or U6988 (N_6988,N_4997,N_4277);
nor U6989 (N_6989,N_5922,N_4515);
nand U6990 (N_6990,N_4154,N_5945);
nand U6991 (N_6991,N_5342,N_4114);
and U6992 (N_6992,N_5833,N_5409);
and U6993 (N_6993,N_5332,N_5882);
nor U6994 (N_6994,N_5576,N_4296);
nand U6995 (N_6995,N_4264,N_5389);
nor U6996 (N_6996,N_4342,N_4020);
nor U6997 (N_6997,N_4791,N_5315);
nor U6998 (N_6998,N_4944,N_5871);
nor U6999 (N_6999,N_5114,N_5759);
or U7000 (N_7000,N_5752,N_5391);
and U7001 (N_7001,N_5220,N_5649);
or U7002 (N_7002,N_4561,N_4590);
nand U7003 (N_7003,N_4808,N_5978);
nand U7004 (N_7004,N_4799,N_4858);
xor U7005 (N_7005,N_4698,N_5281);
or U7006 (N_7006,N_4421,N_5224);
or U7007 (N_7007,N_5809,N_4355);
xnor U7008 (N_7008,N_5793,N_5556);
and U7009 (N_7009,N_5626,N_4667);
or U7010 (N_7010,N_4178,N_4436);
and U7011 (N_7011,N_4890,N_5849);
nor U7012 (N_7012,N_5846,N_5140);
or U7013 (N_7013,N_5101,N_5971);
nor U7014 (N_7014,N_5451,N_4096);
nor U7015 (N_7015,N_5113,N_4189);
nand U7016 (N_7016,N_5846,N_5340);
nor U7017 (N_7017,N_5582,N_4356);
or U7018 (N_7018,N_5790,N_4882);
or U7019 (N_7019,N_5204,N_4802);
nand U7020 (N_7020,N_4393,N_4299);
nand U7021 (N_7021,N_5746,N_5521);
or U7022 (N_7022,N_5940,N_5319);
or U7023 (N_7023,N_5032,N_5261);
xnor U7024 (N_7024,N_5519,N_5604);
and U7025 (N_7025,N_4028,N_4503);
nor U7026 (N_7026,N_4574,N_5105);
nor U7027 (N_7027,N_5546,N_5455);
nor U7028 (N_7028,N_5920,N_4312);
xnor U7029 (N_7029,N_4009,N_4446);
nor U7030 (N_7030,N_4799,N_4978);
nor U7031 (N_7031,N_4412,N_4705);
nor U7032 (N_7032,N_5304,N_4575);
or U7033 (N_7033,N_4837,N_4582);
xor U7034 (N_7034,N_5993,N_4365);
and U7035 (N_7035,N_4397,N_4181);
and U7036 (N_7036,N_4604,N_5758);
nand U7037 (N_7037,N_4625,N_4219);
nand U7038 (N_7038,N_5685,N_4275);
or U7039 (N_7039,N_4479,N_5290);
or U7040 (N_7040,N_4776,N_4148);
and U7041 (N_7041,N_5875,N_4973);
or U7042 (N_7042,N_5261,N_5966);
and U7043 (N_7043,N_4261,N_5878);
and U7044 (N_7044,N_5742,N_4675);
and U7045 (N_7045,N_5560,N_4208);
or U7046 (N_7046,N_4533,N_4627);
nor U7047 (N_7047,N_4715,N_5108);
and U7048 (N_7048,N_4778,N_4602);
nor U7049 (N_7049,N_5053,N_5197);
and U7050 (N_7050,N_4821,N_5232);
nor U7051 (N_7051,N_4944,N_4357);
and U7052 (N_7052,N_5108,N_4985);
and U7053 (N_7053,N_5942,N_4262);
nand U7054 (N_7054,N_4338,N_4400);
and U7055 (N_7055,N_5619,N_4639);
or U7056 (N_7056,N_5185,N_5491);
nor U7057 (N_7057,N_4907,N_4760);
nand U7058 (N_7058,N_5630,N_4155);
nand U7059 (N_7059,N_4803,N_5254);
or U7060 (N_7060,N_4909,N_4564);
nor U7061 (N_7061,N_4186,N_5402);
nor U7062 (N_7062,N_5780,N_5224);
and U7063 (N_7063,N_4810,N_4293);
nand U7064 (N_7064,N_4995,N_4094);
nand U7065 (N_7065,N_5591,N_5293);
xor U7066 (N_7066,N_5032,N_5123);
nor U7067 (N_7067,N_4130,N_5047);
or U7068 (N_7068,N_4914,N_4664);
xnor U7069 (N_7069,N_5769,N_4315);
xor U7070 (N_7070,N_4734,N_5248);
or U7071 (N_7071,N_5456,N_5547);
nand U7072 (N_7072,N_5553,N_4274);
xor U7073 (N_7073,N_5563,N_5778);
nor U7074 (N_7074,N_4648,N_4529);
nor U7075 (N_7075,N_4677,N_4762);
xnor U7076 (N_7076,N_5460,N_4701);
xnor U7077 (N_7077,N_5768,N_5869);
or U7078 (N_7078,N_5628,N_5943);
nor U7079 (N_7079,N_4472,N_5357);
and U7080 (N_7080,N_4669,N_5799);
or U7081 (N_7081,N_4655,N_4324);
xor U7082 (N_7082,N_5049,N_5933);
nand U7083 (N_7083,N_4796,N_5709);
or U7084 (N_7084,N_5482,N_4785);
or U7085 (N_7085,N_5097,N_4839);
or U7086 (N_7086,N_5308,N_5387);
nand U7087 (N_7087,N_4629,N_4627);
nand U7088 (N_7088,N_4647,N_4746);
and U7089 (N_7089,N_4752,N_4255);
nand U7090 (N_7090,N_4626,N_4334);
or U7091 (N_7091,N_4341,N_4679);
nand U7092 (N_7092,N_4547,N_4623);
or U7093 (N_7093,N_4281,N_4495);
or U7094 (N_7094,N_4967,N_5788);
and U7095 (N_7095,N_4152,N_5721);
nor U7096 (N_7096,N_4023,N_5817);
nand U7097 (N_7097,N_5977,N_4246);
and U7098 (N_7098,N_5115,N_5653);
nand U7099 (N_7099,N_4233,N_4704);
and U7100 (N_7100,N_5882,N_4808);
nor U7101 (N_7101,N_5435,N_4910);
and U7102 (N_7102,N_4243,N_5132);
nand U7103 (N_7103,N_5390,N_4300);
nand U7104 (N_7104,N_5069,N_4790);
nor U7105 (N_7105,N_5708,N_5292);
and U7106 (N_7106,N_5150,N_5885);
nor U7107 (N_7107,N_4031,N_4778);
xnor U7108 (N_7108,N_5541,N_5331);
and U7109 (N_7109,N_4562,N_5974);
nand U7110 (N_7110,N_4908,N_5345);
or U7111 (N_7111,N_4731,N_4134);
or U7112 (N_7112,N_4066,N_5363);
nor U7113 (N_7113,N_4059,N_4448);
nand U7114 (N_7114,N_4310,N_4196);
and U7115 (N_7115,N_5331,N_5544);
or U7116 (N_7116,N_5352,N_5825);
or U7117 (N_7117,N_5460,N_4995);
and U7118 (N_7118,N_5808,N_4521);
and U7119 (N_7119,N_4649,N_5763);
and U7120 (N_7120,N_5356,N_4296);
and U7121 (N_7121,N_4139,N_4885);
nand U7122 (N_7122,N_5881,N_5091);
nand U7123 (N_7123,N_4557,N_4173);
nor U7124 (N_7124,N_4369,N_5702);
or U7125 (N_7125,N_4469,N_5609);
nor U7126 (N_7126,N_4092,N_5976);
or U7127 (N_7127,N_4098,N_5924);
nand U7128 (N_7128,N_4304,N_4108);
or U7129 (N_7129,N_5653,N_4335);
or U7130 (N_7130,N_4746,N_5814);
nand U7131 (N_7131,N_5549,N_5515);
nand U7132 (N_7132,N_5712,N_5051);
xnor U7133 (N_7133,N_4141,N_5883);
nand U7134 (N_7134,N_5908,N_5333);
nor U7135 (N_7135,N_5689,N_4856);
nor U7136 (N_7136,N_5071,N_4082);
nand U7137 (N_7137,N_5857,N_4667);
nand U7138 (N_7138,N_4723,N_5028);
nand U7139 (N_7139,N_4167,N_5594);
and U7140 (N_7140,N_5712,N_5026);
and U7141 (N_7141,N_5798,N_4147);
xnor U7142 (N_7142,N_5274,N_5781);
nor U7143 (N_7143,N_4196,N_5696);
and U7144 (N_7144,N_5887,N_5675);
nand U7145 (N_7145,N_5942,N_5207);
nand U7146 (N_7146,N_5104,N_5830);
and U7147 (N_7147,N_4113,N_4462);
nand U7148 (N_7148,N_5614,N_5556);
nor U7149 (N_7149,N_5279,N_4465);
or U7150 (N_7150,N_4845,N_4036);
and U7151 (N_7151,N_4000,N_4249);
nor U7152 (N_7152,N_4000,N_4444);
xor U7153 (N_7153,N_5487,N_5235);
and U7154 (N_7154,N_5708,N_5281);
or U7155 (N_7155,N_4677,N_4079);
or U7156 (N_7156,N_5598,N_4476);
xnor U7157 (N_7157,N_4115,N_4200);
nand U7158 (N_7158,N_4123,N_5343);
xnor U7159 (N_7159,N_5684,N_5955);
nor U7160 (N_7160,N_5424,N_4918);
and U7161 (N_7161,N_4710,N_5771);
or U7162 (N_7162,N_4043,N_5171);
or U7163 (N_7163,N_4580,N_5464);
nor U7164 (N_7164,N_5659,N_4507);
nor U7165 (N_7165,N_4626,N_4760);
nor U7166 (N_7166,N_5761,N_4052);
nor U7167 (N_7167,N_5072,N_4316);
nor U7168 (N_7168,N_5305,N_4542);
and U7169 (N_7169,N_4669,N_4895);
or U7170 (N_7170,N_4412,N_5091);
nand U7171 (N_7171,N_5087,N_5106);
xor U7172 (N_7172,N_5518,N_5850);
xnor U7173 (N_7173,N_4202,N_4133);
or U7174 (N_7174,N_5513,N_5245);
nand U7175 (N_7175,N_4179,N_4155);
or U7176 (N_7176,N_5740,N_5308);
nand U7177 (N_7177,N_5260,N_4870);
nand U7178 (N_7178,N_5206,N_4729);
nor U7179 (N_7179,N_5750,N_4041);
nand U7180 (N_7180,N_4992,N_5466);
and U7181 (N_7181,N_4608,N_4849);
or U7182 (N_7182,N_5880,N_5837);
or U7183 (N_7183,N_4771,N_4256);
or U7184 (N_7184,N_5149,N_5193);
and U7185 (N_7185,N_4717,N_5271);
or U7186 (N_7186,N_4832,N_4308);
and U7187 (N_7187,N_4803,N_4931);
nor U7188 (N_7188,N_5931,N_4753);
and U7189 (N_7189,N_4021,N_5427);
or U7190 (N_7190,N_4107,N_5276);
nor U7191 (N_7191,N_5000,N_5684);
nor U7192 (N_7192,N_4813,N_4705);
or U7193 (N_7193,N_4802,N_4086);
nor U7194 (N_7194,N_5074,N_5160);
or U7195 (N_7195,N_4165,N_4628);
and U7196 (N_7196,N_5332,N_5377);
or U7197 (N_7197,N_5866,N_4236);
nor U7198 (N_7198,N_4653,N_4264);
xnor U7199 (N_7199,N_4619,N_4648);
and U7200 (N_7200,N_4032,N_5157);
or U7201 (N_7201,N_4614,N_5763);
nand U7202 (N_7202,N_4953,N_4264);
nor U7203 (N_7203,N_5659,N_5746);
nand U7204 (N_7204,N_4507,N_5335);
nor U7205 (N_7205,N_5200,N_5206);
xnor U7206 (N_7206,N_4850,N_4493);
nor U7207 (N_7207,N_5529,N_4179);
or U7208 (N_7208,N_4129,N_5348);
or U7209 (N_7209,N_4822,N_4957);
nor U7210 (N_7210,N_4576,N_4267);
or U7211 (N_7211,N_5394,N_4361);
or U7212 (N_7212,N_5537,N_5357);
nor U7213 (N_7213,N_5912,N_4732);
or U7214 (N_7214,N_5976,N_4877);
nand U7215 (N_7215,N_5861,N_5202);
nand U7216 (N_7216,N_5844,N_4436);
xnor U7217 (N_7217,N_4965,N_5299);
and U7218 (N_7218,N_5394,N_4937);
nor U7219 (N_7219,N_5930,N_5359);
xor U7220 (N_7220,N_4319,N_4985);
or U7221 (N_7221,N_4762,N_4591);
nor U7222 (N_7222,N_5039,N_5009);
nand U7223 (N_7223,N_4984,N_4083);
and U7224 (N_7224,N_4701,N_4888);
nor U7225 (N_7225,N_5707,N_5480);
and U7226 (N_7226,N_5957,N_4576);
or U7227 (N_7227,N_5137,N_4062);
or U7228 (N_7228,N_5667,N_5450);
and U7229 (N_7229,N_4770,N_5795);
or U7230 (N_7230,N_4924,N_4065);
and U7231 (N_7231,N_5912,N_5723);
xor U7232 (N_7232,N_5483,N_5328);
nor U7233 (N_7233,N_5603,N_4033);
nand U7234 (N_7234,N_5823,N_4189);
nand U7235 (N_7235,N_4867,N_5997);
and U7236 (N_7236,N_5621,N_5994);
nand U7237 (N_7237,N_5055,N_4385);
nand U7238 (N_7238,N_5931,N_5275);
and U7239 (N_7239,N_4704,N_5955);
and U7240 (N_7240,N_5112,N_5883);
and U7241 (N_7241,N_5585,N_5764);
nand U7242 (N_7242,N_4451,N_4637);
nor U7243 (N_7243,N_5916,N_4111);
and U7244 (N_7244,N_4515,N_4967);
or U7245 (N_7245,N_4639,N_4046);
nor U7246 (N_7246,N_4366,N_5077);
or U7247 (N_7247,N_4368,N_4761);
and U7248 (N_7248,N_4242,N_5324);
and U7249 (N_7249,N_5961,N_4200);
or U7250 (N_7250,N_5812,N_4454);
and U7251 (N_7251,N_5822,N_4508);
and U7252 (N_7252,N_5555,N_4806);
nor U7253 (N_7253,N_5888,N_5790);
and U7254 (N_7254,N_4943,N_5985);
and U7255 (N_7255,N_4102,N_4042);
nor U7256 (N_7256,N_5005,N_5217);
nand U7257 (N_7257,N_4291,N_4220);
nor U7258 (N_7258,N_4916,N_5995);
and U7259 (N_7259,N_5076,N_5943);
xnor U7260 (N_7260,N_4589,N_4146);
nand U7261 (N_7261,N_4123,N_4516);
and U7262 (N_7262,N_4079,N_4905);
xor U7263 (N_7263,N_4656,N_4207);
nor U7264 (N_7264,N_5387,N_5285);
or U7265 (N_7265,N_4169,N_4090);
nor U7266 (N_7266,N_4839,N_5240);
nor U7267 (N_7267,N_5231,N_5456);
or U7268 (N_7268,N_4920,N_5186);
nor U7269 (N_7269,N_4113,N_4258);
xor U7270 (N_7270,N_4734,N_5553);
or U7271 (N_7271,N_5127,N_5797);
and U7272 (N_7272,N_4640,N_5200);
nand U7273 (N_7273,N_5807,N_4331);
xnor U7274 (N_7274,N_4122,N_5297);
and U7275 (N_7275,N_4785,N_5826);
xnor U7276 (N_7276,N_4840,N_5779);
nor U7277 (N_7277,N_5932,N_4703);
nand U7278 (N_7278,N_5209,N_5970);
or U7279 (N_7279,N_5947,N_4467);
or U7280 (N_7280,N_4204,N_5920);
or U7281 (N_7281,N_4799,N_4520);
and U7282 (N_7282,N_4442,N_5665);
and U7283 (N_7283,N_5184,N_5591);
nor U7284 (N_7284,N_5611,N_5463);
nand U7285 (N_7285,N_4777,N_5555);
nand U7286 (N_7286,N_4769,N_5070);
and U7287 (N_7287,N_4990,N_4022);
and U7288 (N_7288,N_5100,N_5143);
and U7289 (N_7289,N_4136,N_4837);
nand U7290 (N_7290,N_4704,N_4460);
nand U7291 (N_7291,N_5103,N_4507);
or U7292 (N_7292,N_4844,N_4041);
or U7293 (N_7293,N_4236,N_4473);
or U7294 (N_7294,N_5584,N_4952);
nand U7295 (N_7295,N_4187,N_4067);
xnor U7296 (N_7296,N_5285,N_5051);
nand U7297 (N_7297,N_5589,N_4756);
xor U7298 (N_7298,N_4245,N_4132);
or U7299 (N_7299,N_4854,N_5451);
nand U7300 (N_7300,N_4140,N_4085);
and U7301 (N_7301,N_5984,N_5465);
and U7302 (N_7302,N_5128,N_5205);
nor U7303 (N_7303,N_4837,N_5927);
nor U7304 (N_7304,N_4714,N_5020);
or U7305 (N_7305,N_4469,N_4815);
or U7306 (N_7306,N_4461,N_4593);
or U7307 (N_7307,N_4143,N_5909);
or U7308 (N_7308,N_5808,N_4273);
and U7309 (N_7309,N_4077,N_5455);
nand U7310 (N_7310,N_5427,N_4720);
nor U7311 (N_7311,N_4332,N_4539);
or U7312 (N_7312,N_4153,N_5019);
nor U7313 (N_7313,N_4560,N_4400);
or U7314 (N_7314,N_5608,N_4512);
or U7315 (N_7315,N_5971,N_4714);
xor U7316 (N_7316,N_4342,N_4415);
nand U7317 (N_7317,N_5582,N_4143);
nor U7318 (N_7318,N_5885,N_4253);
nand U7319 (N_7319,N_4083,N_4686);
and U7320 (N_7320,N_4336,N_4179);
or U7321 (N_7321,N_5172,N_5455);
nand U7322 (N_7322,N_5664,N_5149);
xor U7323 (N_7323,N_4138,N_4162);
and U7324 (N_7324,N_4767,N_5246);
nand U7325 (N_7325,N_5797,N_5724);
xnor U7326 (N_7326,N_4637,N_4433);
nand U7327 (N_7327,N_5755,N_4785);
nor U7328 (N_7328,N_5435,N_4480);
nand U7329 (N_7329,N_5423,N_4462);
nor U7330 (N_7330,N_5731,N_4102);
or U7331 (N_7331,N_5926,N_4552);
nand U7332 (N_7332,N_5326,N_4890);
or U7333 (N_7333,N_4618,N_4573);
nand U7334 (N_7334,N_5661,N_4629);
xor U7335 (N_7335,N_5903,N_5985);
nand U7336 (N_7336,N_5357,N_5567);
and U7337 (N_7337,N_5742,N_5198);
nor U7338 (N_7338,N_5094,N_5280);
nor U7339 (N_7339,N_4631,N_5908);
nor U7340 (N_7340,N_4422,N_5770);
nor U7341 (N_7341,N_4399,N_4924);
nor U7342 (N_7342,N_4651,N_4821);
nand U7343 (N_7343,N_5829,N_5891);
nor U7344 (N_7344,N_4116,N_5277);
nand U7345 (N_7345,N_4981,N_4575);
nor U7346 (N_7346,N_5264,N_4575);
and U7347 (N_7347,N_5016,N_5080);
nand U7348 (N_7348,N_4075,N_5578);
nand U7349 (N_7349,N_5818,N_4191);
and U7350 (N_7350,N_5020,N_5062);
or U7351 (N_7351,N_4759,N_5691);
and U7352 (N_7352,N_5589,N_5306);
and U7353 (N_7353,N_4920,N_4043);
and U7354 (N_7354,N_5540,N_4809);
and U7355 (N_7355,N_5541,N_5041);
xnor U7356 (N_7356,N_4044,N_5732);
nor U7357 (N_7357,N_5868,N_5805);
nor U7358 (N_7358,N_4592,N_4565);
or U7359 (N_7359,N_5256,N_4448);
nor U7360 (N_7360,N_5742,N_5338);
nand U7361 (N_7361,N_4273,N_5656);
and U7362 (N_7362,N_4248,N_4347);
nand U7363 (N_7363,N_5554,N_5690);
xor U7364 (N_7364,N_5012,N_4591);
and U7365 (N_7365,N_5540,N_4100);
nor U7366 (N_7366,N_4508,N_5397);
and U7367 (N_7367,N_4768,N_4251);
nand U7368 (N_7368,N_4723,N_4715);
nand U7369 (N_7369,N_5968,N_5654);
nor U7370 (N_7370,N_4858,N_4344);
or U7371 (N_7371,N_5837,N_5489);
and U7372 (N_7372,N_4157,N_5913);
or U7373 (N_7373,N_5761,N_5638);
xor U7374 (N_7374,N_5372,N_4671);
nor U7375 (N_7375,N_4343,N_4686);
nand U7376 (N_7376,N_5432,N_5569);
or U7377 (N_7377,N_4793,N_5495);
xnor U7378 (N_7378,N_5798,N_5187);
or U7379 (N_7379,N_4642,N_4946);
or U7380 (N_7380,N_5227,N_4657);
nand U7381 (N_7381,N_5333,N_5073);
nor U7382 (N_7382,N_5944,N_5636);
or U7383 (N_7383,N_5521,N_4567);
xnor U7384 (N_7384,N_5777,N_4491);
and U7385 (N_7385,N_5169,N_4400);
nand U7386 (N_7386,N_5386,N_4734);
or U7387 (N_7387,N_4725,N_5934);
and U7388 (N_7388,N_5021,N_4004);
and U7389 (N_7389,N_5811,N_4208);
nand U7390 (N_7390,N_4197,N_5629);
or U7391 (N_7391,N_5152,N_5816);
nand U7392 (N_7392,N_4678,N_4212);
nand U7393 (N_7393,N_4110,N_5403);
nor U7394 (N_7394,N_4698,N_4157);
nand U7395 (N_7395,N_4686,N_5669);
nand U7396 (N_7396,N_5624,N_4788);
nand U7397 (N_7397,N_4116,N_4099);
nor U7398 (N_7398,N_4751,N_4249);
and U7399 (N_7399,N_5445,N_4535);
or U7400 (N_7400,N_5969,N_4694);
xnor U7401 (N_7401,N_4727,N_4474);
and U7402 (N_7402,N_4305,N_5480);
nor U7403 (N_7403,N_5055,N_4587);
and U7404 (N_7404,N_5730,N_5207);
nand U7405 (N_7405,N_5765,N_5188);
and U7406 (N_7406,N_5512,N_4838);
nor U7407 (N_7407,N_5926,N_5681);
and U7408 (N_7408,N_4481,N_4265);
or U7409 (N_7409,N_5084,N_5584);
nor U7410 (N_7410,N_5911,N_5527);
xnor U7411 (N_7411,N_5271,N_4707);
and U7412 (N_7412,N_5489,N_4747);
xnor U7413 (N_7413,N_5709,N_4236);
xor U7414 (N_7414,N_4262,N_4035);
or U7415 (N_7415,N_5231,N_5108);
or U7416 (N_7416,N_4739,N_5233);
and U7417 (N_7417,N_4246,N_4260);
xnor U7418 (N_7418,N_4074,N_5390);
nand U7419 (N_7419,N_4869,N_4099);
nor U7420 (N_7420,N_4744,N_4603);
and U7421 (N_7421,N_5025,N_5870);
or U7422 (N_7422,N_5021,N_5487);
nand U7423 (N_7423,N_5100,N_4860);
nand U7424 (N_7424,N_5160,N_4482);
nor U7425 (N_7425,N_5239,N_4945);
and U7426 (N_7426,N_4550,N_5059);
or U7427 (N_7427,N_5820,N_5042);
nor U7428 (N_7428,N_4185,N_5597);
and U7429 (N_7429,N_4641,N_4738);
xor U7430 (N_7430,N_5992,N_5841);
nand U7431 (N_7431,N_4545,N_5730);
nand U7432 (N_7432,N_5435,N_4018);
and U7433 (N_7433,N_5416,N_5840);
and U7434 (N_7434,N_4752,N_5375);
nor U7435 (N_7435,N_4847,N_5105);
nand U7436 (N_7436,N_5536,N_4801);
or U7437 (N_7437,N_4870,N_4631);
or U7438 (N_7438,N_5106,N_5684);
xor U7439 (N_7439,N_5246,N_4772);
and U7440 (N_7440,N_5528,N_5780);
and U7441 (N_7441,N_4828,N_5183);
nand U7442 (N_7442,N_5035,N_5595);
and U7443 (N_7443,N_4202,N_4436);
nor U7444 (N_7444,N_5742,N_5139);
or U7445 (N_7445,N_4107,N_4554);
and U7446 (N_7446,N_4994,N_5851);
or U7447 (N_7447,N_5381,N_4880);
or U7448 (N_7448,N_5615,N_5052);
nor U7449 (N_7449,N_5599,N_4761);
nor U7450 (N_7450,N_4019,N_4893);
nor U7451 (N_7451,N_4292,N_4290);
or U7452 (N_7452,N_5645,N_4074);
nor U7453 (N_7453,N_5006,N_5706);
or U7454 (N_7454,N_4771,N_5983);
nor U7455 (N_7455,N_5191,N_5343);
or U7456 (N_7456,N_4720,N_5688);
and U7457 (N_7457,N_4316,N_5873);
nor U7458 (N_7458,N_5406,N_5626);
nor U7459 (N_7459,N_5324,N_5398);
nand U7460 (N_7460,N_5404,N_4262);
nand U7461 (N_7461,N_5837,N_5652);
xnor U7462 (N_7462,N_5138,N_5616);
and U7463 (N_7463,N_5113,N_4535);
nor U7464 (N_7464,N_5080,N_4018);
nor U7465 (N_7465,N_5633,N_5860);
nand U7466 (N_7466,N_5978,N_4035);
nand U7467 (N_7467,N_5866,N_4159);
nand U7468 (N_7468,N_4276,N_4900);
nand U7469 (N_7469,N_5403,N_4318);
or U7470 (N_7470,N_4123,N_4741);
nor U7471 (N_7471,N_4662,N_4198);
and U7472 (N_7472,N_4663,N_5742);
nor U7473 (N_7473,N_4554,N_4781);
or U7474 (N_7474,N_5793,N_5822);
xnor U7475 (N_7475,N_4706,N_5221);
nor U7476 (N_7476,N_5819,N_5607);
or U7477 (N_7477,N_4082,N_4085);
or U7478 (N_7478,N_5341,N_4220);
xnor U7479 (N_7479,N_5661,N_5142);
nor U7480 (N_7480,N_4769,N_4783);
nand U7481 (N_7481,N_5263,N_4114);
or U7482 (N_7482,N_5627,N_5439);
and U7483 (N_7483,N_4240,N_4985);
xnor U7484 (N_7484,N_5513,N_4648);
nand U7485 (N_7485,N_4303,N_5585);
or U7486 (N_7486,N_5891,N_5757);
and U7487 (N_7487,N_4214,N_4450);
or U7488 (N_7488,N_4773,N_4714);
or U7489 (N_7489,N_4498,N_4529);
or U7490 (N_7490,N_4260,N_4924);
nand U7491 (N_7491,N_4639,N_5991);
and U7492 (N_7492,N_4507,N_4192);
xnor U7493 (N_7493,N_4608,N_4553);
nand U7494 (N_7494,N_4760,N_5711);
nor U7495 (N_7495,N_5413,N_5312);
nand U7496 (N_7496,N_4819,N_5452);
xor U7497 (N_7497,N_5717,N_5943);
nor U7498 (N_7498,N_5660,N_5504);
or U7499 (N_7499,N_5078,N_5262);
and U7500 (N_7500,N_4799,N_4842);
nor U7501 (N_7501,N_4206,N_5238);
and U7502 (N_7502,N_5715,N_4023);
nor U7503 (N_7503,N_5254,N_5621);
nor U7504 (N_7504,N_4032,N_4301);
and U7505 (N_7505,N_5982,N_4692);
xor U7506 (N_7506,N_5333,N_4375);
or U7507 (N_7507,N_4895,N_4392);
and U7508 (N_7508,N_5773,N_4098);
and U7509 (N_7509,N_5801,N_5761);
nor U7510 (N_7510,N_4814,N_5188);
xnor U7511 (N_7511,N_5366,N_5930);
nand U7512 (N_7512,N_5525,N_5338);
nor U7513 (N_7513,N_4094,N_5200);
xor U7514 (N_7514,N_5446,N_4499);
xnor U7515 (N_7515,N_5457,N_4129);
xor U7516 (N_7516,N_5866,N_5226);
xnor U7517 (N_7517,N_5025,N_4051);
nand U7518 (N_7518,N_4981,N_5373);
nand U7519 (N_7519,N_4348,N_5610);
nor U7520 (N_7520,N_5875,N_5567);
nand U7521 (N_7521,N_4521,N_5402);
nor U7522 (N_7522,N_4105,N_5350);
or U7523 (N_7523,N_4604,N_4228);
or U7524 (N_7524,N_5602,N_5779);
nand U7525 (N_7525,N_4559,N_5881);
and U7526 (N_7526,N_5224,N_5534);
and U7527 (N_7527,N_5610,N_5655);
nor U7528 (N_7528,N_4236,N_4128);
nand U7529 (N_7529,N_5570,N_4625);
nand U7530 (N_7530,N_4956,N_5379);
nor U7531 (N_7531,N_5547,N_4588);
xor U7532 (N_7532,N_5011,N_5147);
nor U7533 (N_7533,N_5244,N_5148);
nand U7534 (N_7534,N_4914,N_4967);
nand U7535 (N_7535,N_4456,N_5874);
xor U7536 (N_7536,N_4358,N_5155);
xnor U7537 (N_7537,N_5073,N_5438);
and U7538 (N_7538,N_5271,N_5466);
nor U7539 (N_7539,N_5808,N_5492);
nor U7540 (N_7540,N_4172,N_5681);
xnor U7541 (N_7541,N_4611,N_5813);
xor U7542 (N_7542,N_4309,N_4712);
nor U7543 (N_7543,N_5922,N_5314);
and U7544 (N_7544,N_4445,N_5614);
nor U7545 (N_7545,N_5196,N_4306);
nand U7546 (N_7546,N_4625,N_4726);
or U7547 (N_7547,N_5260,N_4680);
nor U7548 (N_7548,N_4575,N_4209);
and U7549 (N_7549,N_5171,N_5466);
nand U7550 (N_7550,N_4397,N_4468);
or U7551 (N_7551,N_5508,N_4943);
or U7552 (N_7552,N_5506,N_5710);
or U7553 (N_7553,N_5054,N_4027);
nor U7554 (N_7554,N_5827,N_4608);
nor U7555 (N_7555,N_5680,N_4828);
and U7556 (N_7556,N_4477,N_4910);
or U7557 (N_7557,N_5371,N_4002);
nand U7558 (N_7558,N_4906,N_4413);
nand U7559 (N_7559,N_4905,N_4519);
and U7560 (N_7560,N_4293,N_4459);
and U7561 (N_7561,N_4658,N_4678);
nand U7562 (N_7562,N_4262,N_5480);
and U7563 (N_7563,N_5252,N_5525);
nor U7564 (N_7564,N_4781,N_5042);
or U7565 (N_7565,N_5205,N_5640);
and U7566 (N_7566,N_4928,N_5244);
nand U7567 (N_7567,N_4376,N_5758);
or U7568 (N_7568,N_5765,N_4613);
nor U7569 (N_7569,N_5975,N_5115);
nor U7570 (N_7570,N_4077,N_5472);
nand U7571 (N_7571,N_5650,N_5003);
nand U7572 (N_7572,N_4691,N_5749);
or U7573 (N_7573,N_5459,N_4273);
nor U7574 (N_7574,N_4744,N_4962);
or U7575 (N_7575,N_4398,N_5561);
nand U7576 (N_7576,N_4394,N_4021);
nor U7577 (N_7577,N_5750,N_4212);
and U7578 (N_7578,N_4523,N_5266);
and U7579 (N_7579,N_4446,N_4597);
or U7580 (N_7580,N_4859,N_4332);
nor U7581 (N_7581,N_5220,N_4325);
nand U7582 (N_7582,N_4006,N_4414);
nor U7583 (N_7583,N_5610,N_5906);
or U7584 (N_7584,N_4096,N_4171);
nor U7585 (N_7585,N_5308,N_4047);
nand U7586 (N_7586,N_4103,N_4390);
or U7587 (N_7587,N_5609,N_4888);
nand U7588 (N_7588,N_4145,N_5901);
or U7589 (N_7589,N_4769,N_5541);
nand U7590 (N_7590,N_5655,N_4664);
nand U7591 (N_7591,N_4136,N_5653);
and U7592 (N_7592,N_5808,N_5295);
or U7593 (N_7593,N_5118,N_4410);
nor U7594 (N_7594,N_5872,N_4487);
nor U7595 (N_7595,N_4235,N_4536);
or U7596 (N_7596,N_5606,N_4220);
nand U7597 (N_7597,N_5137,N_5633);
nand U7598 (N_7598,N_4759,N_5070);
and U7599 (N_7599,N_4661,N_5991);
nand U7600 (N_7600,N_4770,N_5059);
or U7601 (N_7601,N_5337,N_4348);
or U7602 (N_7602,N_5771,N_4068);
xnor U7603 (N_7603,N_4519,N_4631);
nand U7604 (N_7604,N_5219,N_4547);
and U7605 (N_7605,N_4039,N_4864);
nand U7606 (N_7606,N_4157,N_4652);
xnor U7607 (N_7607,N_5903,N_4327);
nor U7608 (N_7608,N_4650,N_4450);
and U7609 (N_7609,N_5256,N_4976);
nand U7610 (N_7610,N_5308,N_5528);
and U7611 (N_7611,N_5861,N_5473);
nand U7612 (N_7612,N_4382,N_4752);
nor U7613 (N_7613,N_4058,N_5309);
nand U7614 (N_7614,N_5941,N_5566);
or U7615 (N_7615,N_5592,N_5119);
or U7616 (N_7616,N_5669,N_5677);
or U7617 (N_7617,N_5882,N_5554);
nor U7618 (N_7618,N_4755,N_5115);
and U7619 (N_7619,N_5165,N_5825);
nand U7620 (N_7620,N_5349,N_5085);
nand U7621 (N_7621,N_5942,N_5423);
xnor U7622 (N_7622,N_4444,N_4222);
and U7623 (N_7623,N_5470,N_4686);
nor U7624 (N_7624,N_4495,N_4564);
nand U7625 (N_7625,N_4676,N_4009);
and U7626 (N_7626,N_4197,N_4828);
nand U7627 (N_7627,N_4038,N_4255);
nor U7628 (N_7628,N_4421,N_5188);
or U7629 (N_7629,N_5557,N_4557);
and U7630 (N_7630,N_5723,N_5803);
and U7631 (N_7631,N_5029,N_5372);
nand U7632 (N_7632,N_4057,N_5177);
or U7633 (N_7633,N_4692,N_5094);
nor U7634 (N_7634,N_5481,N_4600);
and U7635 (N_7635,N_5891,N_4844);
nand U7636 (N_7636,N_4520,N_5103);
or U7637 (N_7637,N_5210,N_5918);
and U7638 (N_7638,N_4183,N_5484);
and U7639 (N_7639,N_4888,N_5940);
and U7640 (N_7640,N_5715,N_5519);
or U7641 (N_7641,N_5798,N_5416);
or U7642 (N_7642,N_5743,N_4548);
and U7643 (N_7643,N_4753,N_5258);
or U7644 (N_7644,N_5775,N_4576);
nand U7645 (N_7645,N_4658,N_4456);
nand U7646 (N_7646,N_4138,N_5927);
xnor U7647 (N_7647,N_5145,N_5000);
or U7648 (N_7648,N_5968,N_4053);
nor U7649 (N_7649,N_5124,N_5858);
nor U7650 (N_7650,N_4875,N_4468);
and U7651 (N_7651,N_4295,N_5828);
and U7652 (N_7652,N_5678,N_5262);
xor U7653 (N_7653,N_5835,N_5340);
nand U7654 (N_7654,N_4758,N_4679);
or U7655 (N_7655,N_5603,N_4454);
and U7656 (N_7656,N_4449,N_5847);
nand U7657 (N_7657,N_4658,N_5621);
nand U7658 (N_7658,N_5099,N_4761);
nand U7659 (N_7659,N_5142,N_5224);
and U7660 (N_7660,N_5602,N_4763);
and U7661 (N_7661,N_4626,N_4047);
or U7662 (N_7662,N_4531,N_5885);
and U7663 (N_7663,N_5777,N_5723);
nand U7664 (N_7664,N_5369,N_4176);
xnor U7665 (N_7665,N_5288,N_5151);
and U7666 (N_7666,N_5772,N_5755);
and U7667 (N_7667,N_4938,N_4710);
nor U7668 (N_7668,N_5641,N_4006);
and U7669 (N_7669,N_5549,N_4304);
nand U7670 (N_7670,N_5456,N_4384);
nand U7671 (N_7671,N_5838,N_4976);
xor U7672 (N_7672,N_5892,N_5333);
nand U7673 (N_7673,N_5312,N_4431);
xor U7674 (N_7674,N_4601,N_4540);
and U7675 (N_7675,N_5443,N_5904);
nand U7676 (N_7676,N_4174,N_5946);
or U7677 (N_7677,N_4073,N_5289);
and U7678 (N_7678,N_4347,N_5400);
nor U7679 (N_7679,N_4950,N_5985);
and U7680 (N_7680,N_4094,N_5209);
nor U7681 (N_7681,N_5163,N_5555);
nand U7682 (N_7682,N_4115,N_5512);
and U7683 (N_7683,N_4708,N_4365);
nor U7684 (N_7684,N_4555,N_4107);
nand U7685 (N_7685,N_4802,N_5826);
nand U7686 (N_7686,N_5729,N_5571);
or U7687 (N_7687,N_4900,N_5725);
xor U7688 (N_7688,N_5701,N_4477);
or U7689 (N_7689,N_5143,N_5371);
and U7690 (N_7690,N_4767,N_4768);
or U7691 (N_7691,N_4774,N_5052);
xnor U7692 (N_7692,N_5959,N_4614);
xnor U7693 (N_7693,N_5858,N_5214);
or U7694 (N_7694,N_5576,N_5137);
and U7695 (N_7695,N_5057,N_4380);
nor U7696 (N_7696,N_4449,N_5194);
nand U7697 (N_7697,N_5555,N_4386);
nand U7698 (N_7698,N_5508,N_4059);
or U7699 (N_7699,N_5352,N_4106);
nand U7700 (N_7700,N_5897,N_4962);
and U7701 (N_7701,N_5557,N_5613);
nand U7702 (N_7702,N_5541,N_5156);
nand U7703 (N_7703,N_5479,N_5710);
xnor U7704 (N_7704,N_5818,N_4463);
xor U7705 (N_7705,N_5821,N_4794);
nor U7706 (N_7706,N_4942,N_4860);
or U7707 (N_7707,N_5836,N_4408);
nand U7708 (N_7708,N_4008,N_4445);
and U7709 (N_7709,N_4106,N_4301);
and U7710 (N_7710,N_5205,N_4387);
or U7711 (N_7711,N_5189,N_4675);
xnor U7712 (N_7712,N_4255,N_4843);
or U7713 (N_7713,N_4436,N_5485);
or U7714 (N_7714,N_5774,N_5637);
nor U7715 (N_7715,N_4440,N_4897);
xor U7716 (N_7716,N_4173,N_5729);
and U7717 (N_7717,N_5707,N_5322);
or U7718 (N_7718,N_5720,N_5208);
and U7719 (N_7719,N_4496,N_5667);
nor U7720 (N_7720,N_4687,N_5864);
or U7721 (N_7721,N_4641,N_4463);
nand U7722 (N_7722,N_5252,N_4971);
or U7723 (N_7723,N_4345,N_5796);
xor U7724 (N_7724,N_4634,N_4812);
nand U7725 (N_7725,N_5495,N_5118);
nand U7726 (N_7726,N_4753,N_4135);
or U7727 (N_7727,N_5217,N_5289);
nand U7728 (N_7728,N_5918,N_5867);
or U7729 (N_7729,N_4099,N_4982);
and U7730 (N_7730,N_4664,N_4009);
and U7731 (N_7731,N_4350,N_5671);
and U7732 (N_7732,N_5504,N_4844);
or U7733 (N_7733,N_5991,N_5715);
nand U7734 (N_7734,N_5866,N_4184);
and U7735 (N_7735,N_5993,N_5557);
and U7736 (N_7736,N_4842,N_5801);
nand U7737 (N_7737,N_4007,N_4141);
or U7738 (N_7738,N_4683,N_5212);
xnor U7739 (N_7739,N_5551,N_5573);
or U7740 (N_7740,N_5854,N_5316);
and U7741 (N_7741,N_5845,N_4231);
xnor U7742 (N_7742,N_5580,N_5355);
and U7743 (N_7743,N_4293,N_4353);
and U7744 (N_7744,N_5135,N_4762);
and U7745 (N_7745,N_4724,N_5429);
xor U7746 (N_7746,N_5375,N_4460);
or U7747 (N_7747,N_5851,N_5433);
or U7748 (N_7748,N_4641,N_5978);
nor U7749 (N_7749,N_4709,N_5054);
or U7750 (N_7750,N_5587,N_5736);
or U7751 (N_7751,N_4366,N_4806);
xor U7752 (N_7752,N_5912,N_5951);
nand U7753 (N_7753,N_5165,N_5293);
and U7754 (N_7754,N_4275,N_4101);
or U7755 (N_7755,N_4155,N_4631);
xor U7756 (N_7756,N_5838,N_5153);
and U7757 (N_7757,N_4170,N_4209);
or U7758 (N_7758,N_5590,N_5858);
xnor U7759 (N_7759,N_5314,N_5270);
xor U7760 (N_7760,N_5954,N_5703);
nor U7761 (N_7761,N_4479,N_4626);
nand U7762 (N_7762,N_4034,N_5834);
and U7763 (N_7763,N_4392,N_5520);
nor U7764 (N_7764,N_4121,N_4823);
xnor U7765 (N_7765,N_5209,N_4022);
or U7766 (N_7766,N_4115,N_4962);
nor U7767 (N_7767,N_5376,N_4544);
or U7768 (N_7768,N_4760,N_5541);
nand U7769 (N_7769,N_4964,N_5050);
nand U7770 (N_7770,N_5506,N_5354);
nand U7771 (N_7771,N_4018,N_4793);
nand U7772 (N_7772,N_5584,N_4091);
nor U7773 (N_7773,N_4210,N_4086);
and U7774 (N_7774,N_4454,N_4167);
or U7775 (N_7775,N_5679,N_4345);
or U7776 (N_7776,N_5660,N_4022);
nand U7777 (N_7777,N_5203,N_4176);
nor U7778 (N_7778,N_5951,N_5578);
nor U7779 (N_7779,N_4846,N_4633);
nand U7780 (N_7780,N_5741,N_5785);
nand U7781 (N_7781,N_5550,N_4624);
nand U7782 (N_7782,N_4701,N_4547);
and U7783 (N_7783,N_4005,N_4661);
and U7784 (N_7784,N_4756,N_4780);
xnor U7785 (N_7785,N_4530,N_5218);
nand U7786 (N_7786,N_4014,N_5833);
or U7787 (N_7787,N_5693,N_5734);
xor U7788 (N_7788,N_5042,N_4643);
nand U7789 (N_7789,N_4518,N_5591);
nand U7790 (N_7790,N_4824,N_4513);
nor U7791 (N_7791,N_4321,N_4102);
or U7792 (N_7792,N_5952,N_5406);
and U7793 (N_7793,N_5342,N_4373);
and U7794 (N_7794,N_4876,N_4160);
or U7795 (N_7795,N_5808,N_5857);
nand U7796 (N_7796,N_4704,N_5107);
or U7797 (N_7797,N_5281,N_4688);
nor U7798 (N_7798,N_5359,N_5574);
xor U7799 (N_7799,N_5743,N_4098);
and U7800 (N_7800,N_4115,N_5299);
or U7801 (N_7801,N_5460,N_5761);
or U7802 (N_7802,N_4884,N_4648);
nor U7803 (N_7803,N_5376,N_5266);
nand U7804 (N_7804,N_4453,N_5268);
xnor U7805 (N_7805,N_4532,N_4098);
and U7806 (N_7806,N_4891,N_4950);
xor U7807 (N_7807,N_5974,N_4468);
nor U7808 (N_7808,N_5212,N_5271);
xor U7809 (N_7809,N_4790,N_5551);
nor U7810 (N_7810,N_5670,N_5231);
and U7811 (N_7811,N_5094,N_5429);
and U7812 (N_7812,N_5447,N_4045);
nor U7813 (N_7813,N_5516,N_5606);
or U7814 (N_7814,N_4758,N_4650);
or U7815 (N_7815,N_5039,N_4991);
nand U7816 (N_7816,N_5288,N_5921);
and U7817 (N_7817,N_4986,N_5224);
nand U7818 (N_7818,N_4124,N_5303);
and U7819 (N_7819,N_5455,N_4146);
or U7820 (N_7820,N_4046,N_4459);
nor U7821 (N_7821,N_4501,N_4611);
and U7822 (N_7822,N_5982,N_4888);
nand U7823 (N_7823,N_5463,N_5808);
and U7824 (N_7824,N_4148,N_5426);
nor U7825 (N_7825,N_4004,N_4308);
nor U7826 (N_7826,N_4466,N_4574);
nor U7827 (N_7827,N_4729,N_4014);
xnor U7828 (N_7828,N_4827,N_4840);
and U7829 (N_7829,N_5018,N_5122);
nand U7830 (N_7830,N_5767,N_4126);
and U7831 (N_7831,N_4835,N_5490);
nand U7832 (N_7832,N_4858,N_4326);
nand U7833 (N_7833,N_4982,N_4085);
nand U7834 (N_7834,N_4355,N_5704);
nand U7835 (N_7835,N_4924,N_4402);
nand U7836 (N_7836,N_4886,N_5549);
nor U7837 (N_7837,N_4150,N_4429);
or U7838 (N_7838,N_4751,N_5864);
nand U7839 (N_7839,N_5164,N_5291);
xor U7840 (N_7840,N_4472,N_5819);
or U7841 (N_7841,N_5211,N_4362);
and U7842 (N_7842,N_4156,N_4952);
nand U7843 (N_7843,N_4557,N_5184);
and U7844 (N_7844,N_4879,N_4556);
xor U7845 (N_7845,N_5108,N_5475);
and U7846 (N_7846,N_4645,N_5631);
nor U7847 (N_7847,N_4997,N_5154);
nor U7848 (N_7848,N_4930,N_4112);
nor U7849 (N_7849,N_4124,N_5327);
and U7850 (N_7850,N_4046,N_5386);
or U7851 (N_7851,N_5768,N_5838);
nand U7852 (N_7852,N_4570,N_4613);
nor U7853 (N_7853,N_5133,N_4776);
and U7854 (N_7854,N_4828,N_5755);
and U7855 (N_7855,N_5196,N_4075);
or U7856 (N_7856,N_4389,N_4762);
xnor U7857 (N_7857,N_4809,N_4193);
and U7858 (N_7858,N_5048,N_5773);
nand U7859 (N_7859,N_4387,N_5494);
nor U7860 (N_7860,N_5259,N_4883);
nand U7861 (N_7861,N_5152,N_5658);
nor U7862 (N_7862,N_4476,N_5978);
and U7863 (N_7863,N_4418,N_5926);
or U7864 (N_7864,N_5113,N_5108);
and U7865 (N_7865,N_4560,N_5066);
or U7866 (N_7866,N_4914,N_5051);
or U7867 (N_7867,N_4665,N_5300);
nand U7868 (N_7868,N_5624,N_4089);
and U7869 (N_7869,N_4930,N_4882);
and U7870 (N_7870,N_4286,N_5937);
xnor U7871 (N_7871,N_5727,N_5563);
and U7872 (N_7872,N_5656,N_5125);
and U7873 (N_7873,N_4038,N_5058);
xnor U7874 (N_7874,N_4378,N_5846);
or U7875 (N_7875,N_4264,N_5227);
nand U7876 (N_7876,N_4295,N_5717);
nand U7877 (N_7877,N_4607,N_5301);
xor U7878 (N_7878,N_4117,N_5669);
nand U7879 (N_7879,N_5976,N_4949);
or U7880 (N_7880,N_4621,N_4309);
nor U7881 (N_7881,N_5924,N_4298);
nand U7882 (N_7882,N_5586,N_4435);
nor U7883 (N_7883,N_4175,N_4473);
nand U7884 (N_7884,N_4270,N_4279);
xnor U7885 (N_7885,N_4547,N_4679);
nand U7886 (N_7886,N_5275,N_5840);
and U7887 (N_7887,N_5931,N_4472);
and U7888 (N_7888,N_4445,N_5681);
and U7889 (N_7889,N_5085,N_4954);
xnor U7890 (N_7890,N_5834,N_4945);
and U7891 (N_7891,N_4178,N_5305);
nand U7892 (N_7892,N_5927,N_4151);
and U7893 (N_7893,N_4353,N_4128);
and U7894 (N_7894,N_5766,N_5168);
and U7895 (N_7895,N_5487,N_4333);
and U7896 (N_7896,N_4183,N_5136);
nor U7897 (N_7897,N_5588,N_4901);
or U7898 (N_7898,N_4351,N_5733);
xor U7899 (N_7899,N_5504,N_4597);
nand U7900 (N_7900,N_5984,N_5457);
nand U7901 (N_7901,N_5713,N_4780);
and U7902 (N_7902,N_4484,N_4028);
and U7903 (N_7903,N_5378,N_5750);
nand U7904 (N_7904,N_4534,N_4364);
xnor U7905 (N_7905,N_5118,N_5452);
xor U7906 (N_7906,N_5330,N_5743);
and U7907 (N_7907,N_4094,N_5538);
xnor U7908 (N_7908,N_5985,N_4460);
and U7909 (N_7909,N_4248,N_4980);
and U7910 (N_7910,N_5033,N_4893);
xnor U7911 (N_7911,N_5287,N_5870);
nor U7912 (N_7912,N_4912,N_4088);
nand U7913 (N_7913,N_4442,N_5548);
xor U7914 (N_7914,N_4177,N_5095);
nand U7915 (N_7915,N_4517,N_5749);
or U7916 (N_7916,N_4005,N_4610);
and U7917 (N_7917,N_5084,N_4643);
and U7918 (N_7918,N_5427,N_5075);
xor U7919 (N_7919,N_5678,N_4089);
or U7920 (N_7920,N_5873,N_4180);
and U7921 (N_7921,N_4943,N_4742);
nor U7922 (N_7922,N_4454,N_5161);
nand U7923 (N_7923,N_5707,N_5768);
and U7924 (N_7924,N_4454,N_5702);
and U7925 (N_7925,N_4534,N_5517);
nand U7926 (N_7926,N_4391,N_5649);
nand U7927 (N_7927,N_4357,N_4269);
nor U7928 (N_7928,N_5306,N_4013);
nor U7929 (N_7929,N_5205,N_4293);
nor U7930 (N_7930,N_5389,N_5234);
or U7931 (N_7931,N_4036,N_5304);
and U7932 (N_7932,N_5719,N_4954);
xor U7933 (N_7933,N_5189,N_4518);
or U7934 (N_7934,N_4446,N_4367);
and U7935 (N_7935,N_4772,N_4070);
and U7936 (N_7936,N_5602,N_5761);
nand U7937 (N_7937,N_4546,N_4657);
xnor U7938 (N_7938,N_4517,N_4302);
nand U7939 (N_7939,N_5468,N_5615);
and U7940 (N_7940,N_5314,N_5056);
or U7941 (N_7941,N_5698,N_4267);
or U7942 (N_7942,N_5066,N_5555);
xor U7943 (N_7943,N_4532,N_5780);
nor U7944 (N_7944,N_5054,N_5824);
nor U7945 (N_7945,N_5158,N_4490);
nor U7946 (N_7946,N_4488,N_4760);
or U7947 (N_7947,N_5705,N_5312);
and U7948 (N_7948,N_4411,N_5338);
nor U7949 (N_7949,N_5680,N_5621);
nor U7950 (N_7950,N_4232,N_5673);
and U7951 (N_7951,N_5165,N_4744);
or U7952 (N_7952,N_5218,N_4011);
or U7953 (N_7953,N_4324,N_5949);
or U7954 (N_7954,N_5819,N_5943);
or U7955 (N_7955,N_5566,N_4504);
and U7956 (N_7956,N_4603,N_5308);
and U7957 (N_7957,N_5355,N_4686);
or U7958 (N_7958,N_4873,N_5962);
nor U7959 (N_7959,N_4479,N_4539);
or U7960 (N_7960,N_4877,N_5458);
and U7961 (N_7961,N_5248,N_4121);
and U7962 (N_7962,N_4158,N_4985);
and U7963 (N_7963,N_4400,N_4465);
nor U7964 (N_7964,N_5394,N_5867);
nor U7965 (N_7965,N_4627,N_4785);
and U7966 (N_7966,N_4866,N_4596);
nand U7967 (N_7967,N_4720,N_4979);
or U7968 (N_7968,N_4484,N_5546);
xnor U7969 (N_7969,N_5748,N_4227);
and U7970 (N_7970,N_5119,N_5128);
nand U7971 (N_7971,N_5214,N_5916);
and U7972 (N_7972,N_4109,N_5774);
or U7973 (N_7973,N_4323,N_5193);
or U7974 (N_7974,N_5278,N_4389);
or U7975 (N_7975,N_4888,N_5557);
nor U7976 (N_7976,N_5924,N_4201);
and U7977 (N_7977,N_5353,N_5151);
or U7978 (N_7978,N_5938,N_4933);
xnor U7979 (N_7979,N_4180,N_4900);
or U7980 (N_7980,N_4631,N_4857);
xnor U7981 (N_7981,N_4729,N_5353);
and U7982 (N_7982,N_4139,N_5873);
and U7983 (N_7983,N_5544,N_4534);
nor U7984 (N_7984,N_4919,N_5688);
xor U7985 (N_7985,N_5728,N_4933);
or U7986 (N_7986,N_4249,N_5089);
nor U7987 (N_7987,N_5370,N_4274);
or U7988 (N_7988,N_5802,N_5484);
or U7989 (N_7989,N_4582,N_5874);
and U7990 (N_7990,N_5559,N_5005);
nand U7991 (N_7991,N_5626,N_4440);
nand U7992 (N_7992,N_4079,N_4467);
nor U7993 (N_7993,N_5895,N_4282);
xnor U7994 (N_7994,N_5635,N_5690);
or U7995 (N_7995,N_5376,N_4111);
nor U7996 (N_7996,N_4816,N_4452);
nor U7997 (N_7997,N_5399,N_5443);
nor U7998 (N_7998,N_5284,N_4323);
nand U7999 (N_7999,N_5275,N_5107);
nor U8000 (N_8000,N_6076,N_6704);
xnor U8001 (N_8001,N_6953,N_6813);
or U8002 (N_8002,N_6656,N_7410);
or U8003 (N_8003,N_6051,N_6184);
or U8004 (N_8004,N_7068,N_6015);
or U8005 (N_8005,N_7241,N_7009);
nand U8006 (N_8006,N_6189,N_7132);
or U8007 (N_8007,N_6312,N_7151);
nand U8008 (N_8008,N_7976,N_6479);
nor U8009 (N_8009,N_7780,N_6745);
nor U8010 (N_8010,N_7094,N_6415);
nand U8011 (N_8011,N_7271,N_7943);
nor U8012 (N_8012,N_6730,N_7682);
nor U8013 (N_8013,N_6451,N_7750);
xnor U8014 (N_8014,N_7303,N_6787);
nor U8015 (N_8015,N_6885,N_7001);
or U8016 (N_8016,N_7678,N_7979);
nand U8017 (N_8017,N_7801,N_7518);
nor U8018 (N_8018,N_6582,N_7730);
xnor U8019 (N_8019,N_6464,N_6134);
nand U8020 (N_8020,N_6249,N_7244);
nor U8021 (N_8021,N_6401,N_7665);
or U8022 (N_8022,N_7030,N_7528);
nor U8023 (N_8023,N_7337,N_6904);
or U8024 (N_8024,N_6431,N_7738);
or U8025 (N_8025,N_6417,N_7647);
or U8026 (N_8026,N_7951,N_6499);
and U8027 (N_8027,N_7343,N_7186);
and U8028 (N_8028,N_6388,N_6253);
or U8029 (N_8029,N_7114,N_6889);
or U8030 (N_8030,N_7486,N_7855);
nor U8031 (N_8031,N_7416,N_7973);
or U8032 (N_8032,N_7853,N_7421);
nand U8033 (N_8033,N_7459,N_7002);
nor U8034 (N_8034,N_6827,N_7636);
or U8035 (N_8035,N_7150,N_6516);
nor U8036 (N_8036,N_6177,N_6303);
and U8037 (N_8037,N_6360,N_7883);
xnor U8038 (N_8038,N_7296,N_6569);
nor U8039 (N_8039,N_7452,N_7352);
nor U8040 (N_8040,N_6794,N_6489);
nor U8041 (N_8041,N_6172,N_6914);
and U8042 (N_8042,N_7185,N_7417);
xor U8043 (N_8043,N_6040,N_6135);
nand U8044 (N_8044,N_7274,N_7909);
or U8045 (N_8045,N_6206,N_7335);
nor U8046 (N_8046,N_7003,N_6300);
nor U8047 (N_8047,N_7993,N_6701);
or U8048 (N_8048,N_7530,N_6363);
nor U8049 (N_8049,N_7564,N_7884);
xor U8050 (N_8050,N_6507,N_7413);
nor U8051 (N_8051,N_7802,N_6061);
nor U8052 (N_8052,N_6221,N_6096);
and U8053 (N_8053,N_6728,N_6549);
and U8054 (N_8054,N_7793,N_6553);
or U8055 (N_8055,N_7015,N_6307);
nor U8056 (N_8056,N_7775,N_6833);
or U8057 (N_8057,N_7549,N_6630);
nand U8058 (N_8058,N_7907,N_6317);
nand U8059 (N_8059,N_6325,N_6374);
nand U8060 (N_8060,N_7349,N_7773);
and U8061 (N_8061,N_7426,N_7872);
or U8062 (N_8062,N_7378,N_7714);
nand U8063 (N_8063,N_6054,N_6931);
nand U8064 (N_8064,N_6808,N_6824);
and U8065 (N_8065,N_6205,N_6441);
or U8066 (N_8066,N_6683,N_7927);
nand U8067 (N_8067,N_7514,N_7763);
or U8068 (N_8068,N_6998,N_6757);
and U8069 (N_8069,N_7240,N_6367);
or U8070 (N_8070,N_6688,N_6844);
nand U8071 (N_8071,N_7341,N_7161);
or U8072 (N_8072,N_6547,N_6445);
nor U8073 (N_8073,N_7886,N_7948);
and U8074 (N_8074,N_6793,N_6493);
or U8075 (N_8075,N_6088,N_7147);
nor U8076 (N_8076,N_6660,N_7854);
nand U8077 (N_8077,N_6602,N_7539);
and U8078 (N_8078,N_7955,N_7061);
nor U8079 (N_8079,N_6125,N_6494);
and U8080 (N_8080,N_7901,N_6562);
and U8081 (N_8081,N_6501,N_7338);
nor U8082 (N_8082,N_7867,N_6101);
nand U8083 (N_8083,N_6724,N_6532);
or U8084 (N_8084,N_6257,N_7461);
and U8085 (N_8085,N_6284,N_7965);
and U8086 (N_8086,N_7744,N_7175);
nor U8087 (N_8087,N_7471,N_6544);
nor U8088 (N_8088,N_6848,N_7829);
or U8089 (N_8089,N_7612,N_6925);
nor U8090 (N_8090,N_6213,N_7038);
xor U8091 (N_8091,N_6606,N_7447);
and U8092 (N_8092,N_6839,N_6503);
nand U8093 (N_8093,N_7593,N_7861);
xnor U8094 (N_8094,N_7467,N_6954);
or U8095 (N_8095,N_6675,N_6027);
nand U8096 (N_8096,N_7039,N_7155);
or U8097 (N_8097,N_7138,N_6796);
or U8098 (N_8098,N_6255,N_6756);
nand U8099 (N_8099,N_7637,N_7814);
nor U8100 (N_8100,N_6302,N_6639);
nand U8101 (N_8101,N_6613,N_7042);
or U8102 (N_8102,N_6879,N_6905);
and U8103 (N_8103,N_6845,N_7990);
nand U8104 (N_8104,N_7328,N_6603);
nand U8105 (N_8105,N_7056,N_6585);
nand U8106 (N_8106,N_6222,N_6747);
xnor U8107 (N_8107,N_7975,N_6416);
nand U8108 (N_8108,N_7293,N_6368);
or U8109 (N_8109,N_6165,N_7810);
nand U8110 (N_8110,N_6800,N_6315);
nor U8111 (N_8111,N_6310,N_6472);
nand U8112 (N_8112,N_7429,N_7210);
and U8113 (N_8113,N_7894,N_7893);
nor U8114 (N_8114,N_6557,N_6163);
or U8115 (N_8115,N_7627,N_7401);
and U8116 (N_8116,N_6060,N_6968);
nor U8117 (N_8117,N_7857,N_6413);
nand U8118 (N_8118,N_6427,N_6668);
nand U8119 (N_8119,N_6939,N_6778);
nand U8120 (N_8120,N_6950,N_7017);
and U8121 (N_8121,N_6220,N_6862);
and U8122 (N_8122,N_7294,N_6311);
xor U8123 (N_8123,N_6575,N_7928);
xor U8124 (N_8124,N_7562,N_7610);
nand U8125 (N_8125,N_7758,N_7960);
xor U8126 (N_8126,N_7237,N_6999);
or U8127 (N_8127,N_7195,N_6232);
xor U8128 (N_8128,N_7897,N_7712);
nor U8129 (N_8129,N_7676,N_7922);
nand U8130 (N_8130,N_6560,N_7183);
and U8131 (N_8131,N_6790,N_7501);
and U8132 (N_8132,N_6622,N_6801);
nand U8133 (N_8133,N_6275,N_7279);
and U8134 (N_8134,N_6289,N_7914);
nor U8135 (N_8135,N_6011,N_6971);
nor U8136 (N_8136,N_7313,N_7760);
nor U8137 (N_8137,N_6565,N_6330);
nor U8138 (N_8138,N_6842,N_6989);
nor U8139 (N_8139,N_7092,N_7356);
nand U8140 (N_8140,N_7011,N_6434);
or U8141 (N_8141,N_7949,N_6267);
and U8142 (N_8142,N_6880,N_6488);
and U8143 (N_8143,N_6577,N_7298);
xnor U8144 (N_8144,N_6429,N_6835);
nand U8145 (N_8145,N_6916,N_6157);
and U8146 (N_8146,N_6952,N_7776);
nor U8147 (N_8147,N_6053,N_7756);
and U8148 (N_8148,N_6710,N_6063);
nor U8149 (N_8149,N_7531,N_7603);
or U8150 (N_8150,N_6026,N_6002);
nor U8151 (N_8151,N_6293,N_7715);
or U8152 (N_8152,N_7439,N_7351);
or U8153 (N_8153,N_7433,N_7815);
or U8154 (N_8154,N_7534,N_6722);
or U8155 (N_8155,N_7281,N_6779);
and U8156 (N_8156,N_7905,N_7100);
nand U8157 (N_8157,N_7060,N_7028);
and U8158 (N_8158,N_6143,N_7283);
and U8159 (N_8159,N_6509,N_7632);
or U8160 (N_8160,N_6226,N_6521);
nand U8161 (N_8161,N_6929,N_7947);
or U8162 (N_8162,N_7107,N_6452);
nor U8163 (N_8163,N_6881,N_6346);
nand U8164 (N_8164,N_6713,N_7704);
nor U8165 (N_8165,N_7212,N_6500);
or U8166 (N_8166,N_6637,N_6139);
and U8167 (N_8167,N_6438,N_7910);
xor U8168 (N_8168,N_6681,N_7059);
nor U8169 (N_8169,N_7157,N_6198);
and U8170 (N_8170,N_7639,N_7348);
xnor U8171 (N_8171,N_6913,N_7222);
nand U8172 (N_8172,N_6748,N_7661);
nor U8173 (N_8173,N_7784,N_7101);
and U8174 (N_8174,N_7253,N_7911);
nor U8175 (N_8175,N_7048,N_6963);
and U8176 (N_8176,N_6631,N_7657);
nand U8177 (N_8177,N_7889,N_6277);
xnor U8178 (N_8178,N_7996,N_7950);
and U8179 (N_8179,N_6930,N_6477);
or U8180 (N_8180,N_6283,N_7076);
nand U8181 (N_8181,N_7305,N_6446);
nor U8182 (N_8182,N_7405,N_6349);
nand U8183 (N_8183,N_6102,N_6715);
xor U8184 (N_8184,N_7934,N_6404);
xnor U8185 (N_8185,N_7765,N_7248);
and U8186 (N_8186,N_7063,N_6254);
nor U8187 (N_8187,N_7192,N_6647);
nand U8188 (N_8188,N_7747,N_6679);
and U8189 (N_8189,N_7862,N_6943);
and U8190 (N_8190,N_6000,N_7967);
and U8191 (N_8191,N_6884,N_7314);
nor U8192 (N_8192,N_7696,N_7211);
and U8193 (N_8193,N_7770,N_6240);
nor U8194 (N_8194,N_7504,N_7956);
and U8195 (N_8195,N_7983,N_6822);
or U8196 (N_8196,N_6362,N_7187);
nand U8197 (N_8197,N_6084,N_7790);
and U8198 (N_8198,N_7488,N_6552);
and U8199 (N_8199,N_7172,N_6290);
xor U8200 (N_8200,N_7573,N_7450);
nor U8201 (N_8201,N_7353,N_7615);
or U8202 (N_8202,N_7444,N_7440);
nor U8203 (N_8203,N_6181,N_7340);
and U8204 (N_8204,N_7617,N_6457);
nand U8205 (N_8205,N_6854,N_7134);
nand U8206 (N_8206,N_7600,N_6122);
nor U8207 (N_8207,N_7200,N_7394);
and U8208 (N_8208,N_6397,N_7848);
or U8209 (N_8209,N_7685,N_6294);
nand U8210 (N_8210,N_7912,N_6448);
nand U8211 (N_8211,N_6495,N_7268);
and U8212 (N_8212,N_7840,N_7247);
or U8213 (N_8213,N_7601,N_7299);
and U8214 (N_8214,N_7767,N_6234);
or U8215 (N_8215,N_6230,N_7843);
or U8216 (N_8216,N_7710,N_6995);
nor U8217 (N_8217,N_6481,N_7135);
or U8218 (N_8218,N_7424,N_7936);
xor U8219 (N_8219,N_6531,N_6536);
xor U8220 (N_8220,N_7532,N_6354);
and U8221 (N_8221,N_6804,N_7988);
nand U8222 (N_8222,N_7691,N_6528);
or U8223 (N_8223,N_6737,N_7871);
or U8224 (N_8224,N_7850,N_7629);
nor U8225 (N_8225,N_7336,N_6832);
or U8226 (N_8226,N_6204,N_6539);
nand U8227 (N_8227,N_6803,N_6512);
nor U8228 (N_8228,N_6849,N_6454);
or U8229 (N_8229,N_6771,N_6347);
nand U8230 (N_8230,N_7519,N_6020);
or U8231 (N_8231,N_7548,N_6773);
nor U8232 (N_8232,N_6807,N_6447);
nor U8233 (N_8233,N_6893,N_6323);
and U8234 (N_8234,N_7156,N_7230);
or U8235 (N_8235,N_6915,N_6717);
or U8236 (N_8236,N_6716,N_6145);
nor U8237 (N_8237,N_6308,N_7998);
nor U8238 (N_8238,N_7705,N_7473);
nor U8239 (N_8239,N_6497,N_7823);
xnor U8240 (N_8240,N_6373,N_6402);
or U8241 (N_8241,N_7014,N_6077);
or U8242 (N_8242,N_6933,N_6295);
and U8243 (N_8243,N_7596,N_6540);
nor U8244 (N_8244,N_7529,N_6705);
nand U8245 (N_8245,N_7201,N_6065);
nand U8246 (N_8246,N_6338,N_6333);
xor U8247 (N_8247,N_7372,N_7903);
nor U8248 (N_8248,N_6714,N_7194);
xor U8249 (N_8249,N_6612,N_6772);
nor U8250 (N_8250,N_7819,N_7844);
or U8251 (N_8251,N_7097,N_6523);
xor U8252 (N_8252,N_7751,N_7231);
nand U8253 (N_8253,N_7668,N_7485);
and U8254 (N_8254,N_6093,N_6467);
or U8255 (N_8255,N_6594,N_7484);
and U8256 (N_8256,N_7992,N_7800);
nand U8257 (N_8257,N_7083,N_6085);
xnor U8258 (N_8258,N_7160,N_7512);
and U8259 (N_8259,N_7130,N_7737);
nor U8260 (N_8260,N_6389,N_7755);
and U8261 (N_8261,N_6957,N_6406);
and U8262 (N_8262,N_7383,N_6187);
nand U8263 (N_8263,N_7969,N_6623);
xor U8264 (N_8264,N_6109,N_6689);
or U8265 (N_8265,N_7785,N_6899);
or U8266 (N_8266,N_6997,N_7970);
nand U8267 (N_8267,N_7584,N_6644);
nor U8268 (N_8268,N_7839,N_7812);
and U8269 (N_8269,N_7154,N_7189);
nor U8270 (N_8270,N_6242,N_7168);
nand U8271 (N_8271,N_6774,N_7689);
nand U8272 (N_8272,N_7641,N_6788);
nand U8273 (N_8273,N_7376,N_6058);
and U8274 (N_8274,N_7834,N_6551);
nor U8275 (N_8275,N_6066,N_6471);
nor U8276 (N_8276,N_7285,N_6048);
nand U8277 (N_8277,N_6906,N_6150);
nand U8278 (N_8278,N_7888,N_6579);
nor U8279 (N_8279,N_6241,N_7193);
or U8280 (N_8280,N_6130,N_7560);
nand U8281 (N_8281,N_6318,N_6046);
nor U8282 (N_8282,N_7749,N_7733);
nor U8283 (N_8283,N_6657,N_7631);
or U8284 (N_8284,N_7635,N_7255);
and U8285 (N_8285,N_7547,N_6956);
and U8286 (N_8286,N_7624,N_7618);
and U8287 (N_8287,N_7620,N_6455);
and U8288 (N_8288,N_6331,N_7355);
or U8289 (N_8289,N_6381,N_6856);
and U8290 (N_8290,N_7490,N_7781);
and U8291 (N_8291,N_6940,N_7430);
nor U8292 (N_8292,N_7436,N_7267);
nor U8293 (N_8293,N_7406,N_7939);
nand U8294 (N_8294,N_6475,N_7004);
nor U8295 (N_8295,N_7671,N_6991);
xnor U8296 (N_8296,N_7646,N_6740);
nor U8297 (N_8297,N_6269,N_7523);
nand U8298 (N_8298,N_7441,N_6760);
and U8299 (N_8299,N_7718,N_6684);
and U8300 (N_8300,N_7713,N_6836);
nor U8301 (N_8301,N_6083,N_6282);
or U8302 (N_8302,N_7968,N_6239);
and U8303 (N_8303,N_6245,N_6062);
xor U8304 (N_8304,N_7178,N_6256);
or U8305 (N_8305,N_6821,N_7721);
nor U8306 (N_8306,N_7581,N_7541);
nand U8307 (N_8307,N_6922,N_6511);
and U8308 (N_8308,N_6013,N_6600);
nor U8309 (N_8309,N_6233,N_6932);
nor U8310 (N_8310,N_6351,N_7380);
nand U8311 (N_8311,N_7792,N_7724);
or U8312 (N_8312,N_6113,N_6677);
xor U8313 (N_8313,N_7110,N_6628);
and U8314 (N_8314,N_6319,N_6520);
nand U8315 (N_8315,N_6754,N_7246);
nor U8316 (N_8316,N_7622,N_7043);
and U8317 (N_8317,N_7044,N_7027);
xor U8318 (N_8318,N_6098,N_7062);
or U8319 (N_8319,N_7373,N_6203);
or U8320 (N_8320,N_7206,N_7437);
and U8321 (N_8321,N_7209,N_7041);
nor U8322 (N_8322,N_6791,N_6414);
or U8323 (N_8323,N_7202,N_6951);
nor U8324 (N_8324,N_7125,N_7025);
or U8325 (N_8325,N_7128,N_6023);
nand U8326 (N_8326,N_7895,N_6871);
nand U8327 (N_8327,N_7270,N_6108);
and U8328 (N_8328,N_7408,N_6545);
or U8329 (N_8329,N_7732,N_7933);
nand U8330 (N_8330,N_6876,N_6610);
xor U8331 (N_8331,N_6410,N_7981);
nand U8332 (N_8332,N_7196,N_6418);
and U8333 (N_8333,N_7418,N_6453);
or U8334 (N_8334,N_6902,N_6120);
nor U8335 (N_8335,N_6605,N_6168);
nand U8336 (N_8336,N_6525,N_7264);
nand U8337 (N_8337,N_6529,N_6372);
nor U8338 (N_8338,N_6841,N_7904);
nor U8339 (N_8339,N_6753,N_7929);
nand U8340 (N_8340,N_7753,N_7215);
nand U8341 (N_8341,N_6498,N_7788);
or U8342 (N_8342,N_6296,N_7489);
or U8343 (N_8343,N_6342,N_7051);
or U8344 (N_8344,N_7120,N_6875);
nor U8345 (N_8345,N_6900,N_6025);
nor U8346 (N_8346,N_7687,N_7010);
nand U8347 (N_8347,N_7860,N_7799);
and U8348 (N_8348,N_7681,N_7482);
or U8349 (N_8349,N_6141,N_6752);
nand U8350 (N_8350,N_6285,N_7858);
or U8351 (N_8351,N_7502,N_7422);
nand U8352 (N_8352,N_6422,N_7284);
or U8353 (N_8353,N_6201,N_7851);
nand U8354 (N_8354,N_6124,N_6478);
nor U8355 (N_8355,N_7164,N_7694);
or U8356 (N_8356,N_7731,N_7602);
nand U8357 (N_8357,N_7390,N_6288);
xor U8358 (N_8358,N_6625,N_7728);
nand U8359 (N_8359,N_6056,N_6082);
or U8360 (N_8360,N_6041,N_6016);
nor U8361 (N_8361,N_6857,N_6712);
and U8362 (N_8362,N_6567,N_6969);
or U8363 (N_8363,N_7554,N_7937);
and U8364 (N_8364,N_7371,N_6185);
nand U8365 (N_8365,N_7845,N_7654);
and U8366 (N_8366,N_6167,N_6783);
and U8367 (N_8367,N_7260,N_7908);
nor U8368 (N_8368,N_7289,N_6659);
or U8369 (N_8369,N_7446,N_7675);
nor U8370 (N_8370,N_7594,N_7058);
nand U8371 (N_8371,N_6199,N_7959);
or U8372 (N_8372,N_7925,N_7497);
or U8373 (N_8373,N_7772,N_6112);
nor U8374 (N_8374,N_7590,N_6948);
nor U8375 (N_8375,N_7265,N_7509);
nor U8376 (N_8376,N_7677,N_7403);
or U8377 (N_8377,N_7327,N_7366);
nand U8378 (N_8378,N_6209,N_7761);
nor U8379 (N_8379,N_7725,N_7966);
nor U8380 (N_8380,N_6433,N_7404);
nor U8381 (N_8381,N_7842,N_6571);
or U8382 (N_8382,N_6151,N_7055);
nor U8383 (N_8383,N_7377,N_7346);
nor U8384 (N_8384,N_7849,N_6298);
or U8385 (N_8385,N_6069,N_6105);
nor U8386 (N_8386,N_6247,N_7859);
or U8387 (N_8387,N_6767,N_6248);
nor U8388 (N_8388,N_6459,N_6891);
and U8389 (N_8389,N_7766,N_7953);
xnor U8390 (N_8390,N_7614,N_7940);
and U8391 (N_8391,N_6812,N_7503);
nand U8392 (N_8392,N_6042,N_6476);
nor U8393 (N_8393,N_7229,N_7708);
or U8394 (N_8394,N_7971,N_6817);
nand U8395 (N_8395,N_7263,N_6286);
nor U8396 (N_8396,N_6361,N_7419);
nand U8397 (N_8397,N_6805,N_7278);
nor U8398 (N_8398,N_7451,N_7638);
and U8399 (N_8399,N_7238,N_7239);
nor U8400 (N_8400,N_6648,N_6994);
nand U8401 (N_8401,N_6001,N_6262);
nor U8402 (N_8402,N_6019,N_7827);
and U8403 (N_8403,N_7464,N_7479);
nand U8404 (N_8404,N_7930,N_6661);
or U8405 (N_8405,N_6744,N_6736);
nor U8406 (N_8406,N_7599,N_6215);
or U8407 (N_8407,N_6735,N_6483);
nand U8408 (N_8408,N_6797,N_6179);
nor U8409 (N_8409,N_7536,N_6502);
nand U8410 (N_8410,N_6806,N_7660);
and U8411 (N_8411,N_7566,N_7249);
nor U8412 (N_8412,N_6538,N_6961);
nand U8413 (N_8413,N_6510,N_7300);
or U8414 (N_8414,N_6522,N_7588);
or U8415 (N_8415,N_7958,N_6126);
or U8416 (N_8416,N_6263,N_7923);
or U8417 (N_8417,N_6384,N_6364);
nor U8418 (N_8418,N_7986,N_6894);
nor U8419 (N_8419,N_7047,N_6009);
xor U8420 (N_8420,N_6877,N_7207);
or U8421 (N_8421,N_6670,N_6169);
and U8422 (N_8422,N_7029,N_7124);
xor U8423 (N_8423,N_7115,N_6383);
and U8424 (N_8424,N_7386,N_6359);
xnor U8425 (N_8425,N_7666,N_6586);
and U8426 (N_8426,N_6775,N_7317);
or U8427 (N_8427,N_6170,N_6784);
and U8428 (N_8428,N_7324,N_6550);
nand U8429 (N_8429,N_7099,N_6707);
nand U8430 (N_8430,N_7621,N_7865);
and U8431 (N_8431,N_6261,N_6635);
xor U8432 (N_8432,N_6443,N_6449);
and U8433 (N_8433,N_7081,N_7686);
or U8434 (N_8434,N_6225,N_7640);
or U8435 (N_8435,N_7980,N_6385);
nor U8436 (N_8436,N_7989,N_6238);
and U8437 (N_8437,N_6986,N_7697);
nand U8438 (N_8438,N_6674,N_6799);
or U8439 (N_8439,N_6087,N_6814);
or U8440 (N_8440,N_6634,N_7159);
xor U8441 (N_8441,N_7468,N_6345);
and U8442 (N_8442,N_7820,N_6343);
or U8443 (N_8443,N_7499,N_6685);
and U8444 (N_8444,N_6336,N_6075);
and U8445 (N_8445,N_6726,N_6175);
nor U8446 (N_8446,N_7117,N_6104);
nand U8447 (N_8447,N_6686,N_7902);
and U8448 (N_8448,N_6561,N_7310);
or U8449 (N_8449,N_6942,N_6297);
and U8450 (N_8450,N_7589,N_6955);
nor U8451 (N_8451,N_6918,N_6160);
nand U8452 (N_8452,N_6371,N_6162);
and U8453 (N_8453,N_6469,N_6356);
nor U8454 (N_8454,N_6131,N_6067);
and U8455 (N_8455,N_6078,N_6543);
nand U8456 (N_8456,N_7236,N_7064);
and U8457 (N_8457,N_6838,N_6265);
or U8458 (N_8458,N_6641,N_7587);
nand U8459 (N_8459,N_6466,N_6589);
and U8460 (N_8460,N_7716,N_6669);
and U8461 (N_8461,N_6616,N_6959);
nand U8462 (N_8462,N_7301,N_6541);
or U8463 (N_8463,N_6627,N_6021);
nand U8464 (N_8464,N_7495,N_6161);
xnor U8465 (N_8465,N_7762,N_7304);
nand U8466 (N_8466,N_6387,N_6461);
and U8467 (N_8467,N_7650,N_6344);
and U8468 (N_8468,N_6340,N_7875);
nor U8469 (N_8469,N_7277,N_7516);
or U8470 (N_8470,N_7515,N_6287);
nor U8471 (N_8471,N_7932,N_6985);
nor U8472 (N_8472,N_7828,N_6530);
or U8473 (N_8473,N_7651,N_7522);
nand U8474 (N_8474,N_6268,N_6910);
nor U8475 (N_8475,N_7498,N_6036);
and U8476 (N_8476,N_6430,N_7742);
and U8477 (N_8477,N_6566,N_6264);
nor U8478 (N_8478,N_6320,N_6858);
and U8479 (N_8479,N_6508,N_6878);
xor U8480 (N_8480,N_6620,N_6166);
nand U8481 (N_8481,N_6873,N_7942);
nor U8482 (N_8482,N_7803,N_7090);
nor U8483 (N_8483,N_7754,N_7242);
nand U8484 (N_8484,N_7556,N_6158);
nand U8485 (N_8485,N_7050,N_6355);
or U8486 (N_8486,N_7659,N_6299);
nor U8487 (N_8487,N_6785,N_7302);
or U8488 (N_8488,N_7619,N_7095);
nand U8489 (N_8489,N_6171,N_6780);
xnor U8490 (N_8490,N_6618,N_7846);
nor U8491 (N_8491,N_7112,N_7891);
nand U8492 (N_8492,N_6895,N_6458);
nand U8493 (N_8493,N_7088,N_6535);
nor U8494 (N_8494,N_6119,N_7272);
nor U8495 (N_8495,N_7521,N_7357);
xnor U8496 (N_8496,N_7818,N_6123);
nor U8497 (N_8497,N_6743,N_6305);
or U8498 (N_8498,N_6682,N_7570);
or U8499 (N_8499,N_6259,N_7679);
nand U8500 (N_8500,N_6080,N_6014);
or U8501 (N_8501,N_6766,N_7778);
or U8502 (N_8502,N_7276,N_6941);
nor U8503 (N_8503,N_6115,N_7688);
or U8504 (N_8504,N_7162,N_7524);
or U8505 (N_8505,N_7188,N_7796);
nand U8506 (N_8506,N_7362,N_6004);
xnor U8507 (N_8507,N_6764,N_6938);
nand U8508 (N_8508,N_6935,N_7852);
and U8509 (N_8509,N_7007,N_7642);
or U8510 (N_8510,N_6534,N_7535);
or U8511 (N_8511,N_6974,N_6867);
and U8512 (N_8512,N_6008,N_7994);
or U8513 (N_8513,N_7174,N_7311);
nor U8514 (N_8514,N_7887,N_6850);
nor U8515 (N_8515,N_6546,N_7291);
nand U8516 (N_8516,N_7466,N_7127);
or U8517 (N_8517,N_6224,N_6038);
nor U8518 (N_8518,N_7626,N_6564);
or U8519 (N_8519,N_7184,N_7129);
nand U8520 (N_8520,N_7706,N_7572);
or U8521 (N_8521,N_6407,N_7312);
nor U8522 (N_8522,N_7077,N_6465);
nand U8523 (N_8523,N_7709,N_6568);
nand U8524 (N_8524,N_6409,N_6770);
nor U8525 (N_8525,N_6629,N_6155);
or U8526 (N_8526,N_6353,N_7768);
xor U8527 (N_8527,N_6010,N_7435);
and U8528 (N_8528,N_6419,N_6907);
or U8529 (N_8529,N_6029,N_7214);
nand U8530 (N_8530,N_7397,N_7809);
nor U8531 (N_8531,N_7935,N_6127);
and U8532 (N_8532,N_6202,N_7363);
and U8533 (N_8533,N_7034,N_7711);
or U8534 (N_8534,N_7567,N_7074);
nand U8535 (N_8535,N_6815,N_7333);
or U8536 (N_8536,N_6272,N_7173);
nor U8537 (N_8537,N_7552,N_7525);
and U8538 (N_8538,N_7952,N_6655);
nand U8539 (N_8539,N_7385,N_7580);
or U8540 (N_8540,N_6651,N_6217);
nor U8541 (N_8541,N_7663,N_7121);
or U8542 (N_8542,N_6164,N_6049);
and U8543 (N_8543,N_6834,N_7727);
nor U8544 (N_8544,N_7257,N_6376);
or U8545 (N_8545,N_6246,N_6052);
xor U8546 (N_8546,N_6855,N_7743);
and U8547 (N_8547,N_7111,N_7542);
nand U8548 (N_8548,N_6005,N_7656);
or U8549 (N_8549,N_7838,N_6828);
or U8550 (N_8550,N_7306,N_7119);
and U8551 (N_8551,N_6671,N_6375);
and U8552 (N_8552,N_6983,N_6742);
and U8553 (N_8553,N_7961,N_6378);
or U8554 (N_8554,N_7469,N_7374);
nor U8555 (N_8555,N_7455,N_6426);
nand U8556 (N_8556,N_6456,N_7103);
and U8557 (N_8557,N_6136,N_6099);
and U8558 (N_8558,N_6090,N_6033);
nor U8559 (N_8559,N_6395,N_7067);
and U8560 (N_8560,N_7093,N_7224);
nand U8561 (N_8561,N_6485,N_6695);
xnor U8562 (N_8562,N_7227,N_7251);
or U8563 (N_8563,N_6444,N_7391);
nand U8564 (N_8564,N_7347,N_7821);
nor U8565 (N_8565,N_7364,N_6927);
or U8566 (N_8566,N_7393,N_6114);
or U8567 (N_8567,N_6826,N_6652);
nand U8568 (N_8568,N_7442,N_6964);
or U8569 (N_8569,N_7275,N_6776);
xnor U8570 (N_8570,N_7329,N_7576);
or U8571 (N_8571,N_6223,N_6709);
nor U8572 (N_8572,N_6846,N_7483);
and U8573 (N_8573,N_7645,N_7662);
and U8574 (N_8574,N_6598,N_7680);
and U8575 (N_8575,N_6673,N_6182);
xor U8576 (N_8576,N_6727,N_7608);
nand U8577 (N_8577,N_6604,N_6632);
and U8578 (N_8578,N_6352,N_6738);
nor U8579 (N_8579,N_6967,N_6975);
nand U8580 (N_8580,N_6798,N_7527);
nand U8581 (N_8581,N_7794,N_6092);
nor U8582 (N_8582,N_6391,N_7334);
nand U8583 (N_8583,N_6193,N_6412);
nand U8584 (N_8584,N_7644,N_7182);
nand U8585 (N_8585,N_6183,N_7804);
or U8586 (N_8586,N_7049,N_6823);
or U8587 (N_8587,N_7037,N_7997);
and U8588 (N_8588,N_7825,N_6400);
or U8589 (N_8589,N_6420,N_7574);
nand U8590 (N_8590,N_7673,N_7457);
nor U8591 (N_8591,N_6990,N_7633);
or U8592 (N_8592,N_6006,N_7791);
and U8593 (N_8593,N_6909,N_7745);
or U8594 (N_8594,N_6200,N_7358);
xor U8595 (N_8595,N_7280,N_7102);
and U8596 (N_8596,N_7693,N_7609);
nand U8597 (N_8597,N_6408,N_6116);
or U8598 (N_8598,N_7170,N_7919);
and U8599 (N_8599,N_7764,N_6188);
nor U8600 (N_8600,N_6617,N_6482);
xor U8601 (N_8601,N_7089,N_6527);
or U8602 (N_8602,N_7604,N_7605);
nand U8603 (N_8603,N_6663,N_6094);
or U8604 (N_8604,N_6337,N_6936);
nand U8605 (N_8605,N_7667,N_7434);
and U8606 (N_8606,N_7517,N_6646);
nand U8607 (N_8607,N_6022,N_6313);
nand U8608 (N_8608,N_6339,N_7035);
or U8609 (N_8609,N_7384,N_6140);
or U8610 (N_8610,N_7414,N_6984);
nand U8611 (N_8611,N_6570,N_7944);
nand U8612 (N_8612,N_7075,N_6146);
or U8613 (N_8613,N_6491,N_6110);
nor U8614 (N_8614,N_7777,N_7079);
nand U8615 (N_8615,N_6474,N_6227);
and U8616 (N_8616,N_6070,N_6073);
nand U8617 (N_8617,N_7769,N_7389);
or U8618 (N_8618,N_6281,N_7142);
or U8619 (N_8619,N_7208,N_6291);
nor U8620 (N_8620,N_7165,N_7545);
nor U8621 (N_8621,N_6057,N_6252);
and U8622 (N_8622,N_6435,N_7892);
and U8623 (N_8623,N_7606,N_7287);
xor U8624 (N_8624,N_7292,N_7831);
and U8625 (N_8625,N_6152,N_7890);
nor U8626 (N_8626,N_7866,N_6229);
and U8627 (N_8627,N_7456,N_7899);
or U8628 (N_8628,N_7964,N_6820);
nand U8629 (N_8629,N_6919,N_6869);
or U8630 (N_8630,N_7991,N_6690);
and U8631 (N_8631,N_7084,N_7719);
nor U8632 (N_8632,N_6920,N_7729);
or U8633 (N_8633,N_6274,N_6729);
and U8634 (N_8634,N_7233,N_7438);
nand U8635 (N_8635,N_6421,N_6072);
nor U8636 (N_8636,N_6672,N_7649);
or U8637 (N_8637,N_7533,N_7683);
or U8638 (N_8638,N_7835,N_6390);
or U8639 (N_8639,N_7630,N_7826);
and U8640 (N_8640,N_7837,N_6746);
or U8641 (N_8641,N_6792,N_7546);
and U8642 (N_8642,N_6874,N_6432);
or U8643 (N_8643,N_6786,N_6156);
and U8644 (N_8644,N_6696,N_6097);
nand U8645 (N_8645,N_7140,N_6519);
xnor U8646 (N_8646,N_7022,N_7962);
nand U8647 (N_8647,N_6513,N_6591);
and U8648 (N_8648,N_6324,N_6089);
nor U8649 (N_8649,N_6208,N_7783);
nand U8650 (N_8650,N_6601,N_6450);
nor U8651 (N_8651,N_7722,N_6843);
nor U8652 (N_8652,N_6496,N_7322);
nor U8653 (N_8653,N_7013,N_7918);
or U8654 (N_8654,N_6037,N_6638);
xor U8655 (N_8655,N_7428,N_7342);
nand U8656 (N_8656,N_7774,N_7611);
nand U8657 (N_8657,N_6864,N_7513);
nand U8658 (N_8658,N_7046,N_7863);
xor U8659 (N_8659,N_7868,N_7219);
nor U8660 (N_8660,N_6463,N_7585);
nand U8661 (N_8661,N_7204,N_6818);
nor U8662 (N_8662,N_7592,N_7613);
xnor U8663 (N_8663,N_7152,N_7472);
and U8664 (N_8664,N_7878,N_6555);
nand U8665 (N_8665,N_7454,N_7558);
nor U8666 (N_8666,N_6619,N_6332);
nand U8667 (N_8667,N_6860,N_6244);
and U8668 (N_8668,N_6816,N_6852);
and U8669 (N_8669,N_7757,N_6437);
nor U8670 (N_8670,N_7344,N_6825);
and U8671 (N_8671,N_7308,N_7012);
nand U8672 (N_8672,N_7474,N_6190);
and U8673 (N_8673,N_7000,N_6768);
or U8674 (N_8674,N_7261,N_6278);
nor U8675 (N_8675,N_6423,N_6693);
or U8676 (N_8676,N_7396,N_6694);
nand U8677 (N_8677,N_6440,N_7786);
and U8678 (N_8678,N_6210,N_6106);
or U8679 (N_8679,N_6720,N_6865);
nand U8680 (N_8680,N_6958,N_6732);
or U8681 (N_8681,N_7203,N_7586);
and U8682 (N_8682,N_6645,N_7748);
and U8683 (N_8683,N_6059,N_7559);
or U8684 (N_8684,N_6678,N_6718);
nor U8685 (N_8685,N_6607,N_7431);
nor U8686 (N_8686,N_6007,N_7258);
xor U8687 (N_8687,N_7571,N_7551);
or U8688 (N_8688,N_6934,N_6982);
and U8689 (N_8689,N_7033,N_6191);
nor U8690 (N_8690,N_7096,N_7146);
and U8691 (N_8691,N_6365,N_7917);
and U8692 (N_8692,N_6819,N_7579);
nor U8693 (N_8693,N_6548,N_6937);
nor U8694 (N_8694,N_6650,N_6595);
or U8695 (N_8695,N_6993,N_6396);
and U8696 (N_8696,N_7669,N_7021);
xor U8697 (N_8697,N_6271,N_7698);
and U8698 (N_8698,N_7078,N_6692);
xor U8699 (N_8699,N_6149,N_7018);
and U8700 (N_8700,N_7295,N_6988);
and U8701 (N_8701,N_7974,N_7597);
nor U8702 (N_8702,N_7286,N_6572);
or U8703 (N_8703,N_7520,N_6978);
nor U8704 (N_8704,N_7053,N_7443);
and U8705 (N_8705,N_7795,N_7583);
nor U8706 (N_8706,N_6830,N_6996);
or U8707 (N_8707,N_6012,N_6580);
and U8708 (N_8708,N_7080,N_6194);
or U8709 (N_8709,N_6556,N_6851);
or U8710 (N_8710,N_7475,N_7369);
nor U8711 (N_8711,N_7256,N_7381);
and U8712 (N_8712,N_7205,N_6327);
nor U8713 (N_8713,N_6615,N_6329);
nor U8714 (N_8714,N_6235,N_6691);
xor U8715 (N_8715,N_7217,N_7118);
and U8716 (N_8716,N_6107,N_7166);
or U8717 (N_8717,N_7811,N_6301);
nand U8718 (N_8718,N_7190,N_6370);
nand U8719 (N_8719,N_7087,N_7739);
and U8720 (N_8720,N_7141,N_7882);
xor U8721 (N_8721,N_6809,N_7316);
nor U8722 (N_8722,N_7412,N_6861);
nor U8723 (N_8723,N_7507,N_7752);
nor U8724 (N_8724,N_7652,N_7420);
nand U8725 (N_8725,N_6912,N_6148);
xnor U8726 (N_8726,N_7982,N_7643);
and U8727 (N_8727,N_6866,N_6981);
and U8728 (N_8728,N_6128,N_6810);
and U8729 (N_8729,N_7847,N_6765);
or U8730 (N_8730,N_7379,N_7822);
nand U8731 (N_8731,N_7139,N_6436);
and U8732 (N_8732,N_7807,N_7538);
and U8733 (N_8733,N_6394,N_6515);
xor U8734 (N_8734,N_6972,N_7395);
or U8735 (N_8735,N_6176,N_6608);
nand U8736 (N_8736,N_7898,N_6237);
nor U8737 (N_8737,N_6017,N_7149);
nor U8738 (N_8738,N_6335,N_6924);
or U8739 (N_8739,N_7321,N_7575);
and U8740 (N_8740,N_7361,N_6590);
and U8741 (N_8741,N_6129,N_7144);
nor U8742 (N_8742,N_6917,N_6218);
nand U8743 (N_8743,N_6517,N_7553);
nand U8744 (N_8744,N_6047,N_6926);
or U8745 (N_8745,N_6626,N_6697);
and U8746 (N_8746,N_7832,N_7510);
nor U8747 (N_8747,N_6795,N_7198);
nor U8748 (N_8748,N_6399,N_7307);
nor U8749 (N_8749,N_7670,N_6762);
or U8750 (N_8750,N_6699,N_6366);
or U8751 (N_8751,N_6970,N_6593);
or U8752 (N_8752,N_7537,N_7463);
and U8753 (N_8753,N_7506,N_6174);
and U8754 (N_8754,N_7915,N_7108);
nor U8755 (N_8755,N_6486,N_6928);
and U8756 (N_8756,N_6279,N_6611);
and U8757 (N_8757,N_6649,N_7568);
and U8758 (N_8758,N_6563,N_7113);
nor U8759 (N_8759,N_6840,N_7478);
and U8760 (N_8760,N_7319,N_7137);
nand U8761 (N_8761,N_6700,N_6091);
nand U8762 (N_8762,N_7069,N_6470);
or U8763 (N_8763,N_6386,N_6032);
xor U8764 (N_8764,N_6460,N_7808);
nor U8765 (N_8765,N_6403,N_6811);
nand U8766 (N_8766,N_6309,N_7625);
nor U8767 (N_8767,N_7879,N_7323);
nor U8768 (N_8768,N_6533,N_7180);
xor U8769 (N_8769,N_6292,N_7577);
or U8770 (N_8770,N_6411,N_6837);
or U8771 (N_8771,N_7005,N_6147);
nand U8772 (N_8772,N_7221,N_6640);
nor U8773 (N_8773,N_7496,N_6962);
or U8774 (N_8774,N_6658,N_6979);
and U8775 (N_8775,N_6236,N_6276);
or U8776 (N_8776,N_6118,N_6250);
nor U8777 (N_8777,N_7492,N_6947);
and U8778 (N_8778,N_6358,N_6596);
nor U8779 (N_8779,N_6280,N_7318);
nand U8780 (N_8780,N_6853,N_6750);
xor U8781 (N_8781,N_6518,N_7557);
and U8782 (N_8782,N_7741,N_6064);
xnor U8783 (N_8783,N_7073,N_6676);
nor U8784 (N_8784,N_6196,N_6424);
xnor U8785 (N_8785,N_7787,N_7540);
nand U8786 (N_8786,N_7169,N_6369);
or U8787 (N_8787,N_6890,N_7703);
nand U8788 (N_8788,N_7282,N_7086);
nand U8789 (N_8789,N_7565,N_7266);
and U8790 (N_8790,N_6666,N_7817);
or U8791 (N_8791,N_6973,N_6380);
nand U8792 (N_8792,N_7331,N_6079);
nor U8793 (N_8793,N_6473,N_7026);
nor U8794 (N_8794,N_6018,N_6306);
and U8795 (N_8795,N_7511,N_7269);
or U8796 (N_8796,N_7288,N_7398);
nand U8797 (N_8797,N_7040,N_6480);
nand U8798 (N_8798,N_6758,N_6621);
and U8799 (N_8799,N_7824,N_7065);
nand U8800 (N_8800,N_6966,N_6030);
or U8801 (N_8801,N_6180,N_6653);
nor U8802 (N_8802,N_7008,N_6043);
and U8803 (N_8803,N_6142,N_7813);
xnor U8804 (N_8804,N_7325,N_7595);
and U8805 (N_8805,N_6524,N_7582);
and U8806 (N_8806,N_6428,N_6863);
and U8807 (N_8807,N_7921,N_7126);
nor U8808 (N_8808,N_7945,N_6304);
and U8809 (N_8809,N_7984,N_7655);
nand U8810 (N_8810,N_7692,N_7700);
xor U8811 (N_8811,N_6055,N_7019);
and U8812 (N_8812,N_6086,N_7684);
nor U8813 (N_8813,N_7977,N_6687);
nor U8814 (N_8814,N_6643,N_6680);
or U8815 (N_8815,N_7735,N_6228);
or U8816 (N_8816,N_6044,N_6599);
or U8817 (N_8817,N_7148,N_6578);
nor U8818 (N_8818,N_7924,N_7158);
and U8819 (N_8819,N_7896,N_6992);
nand U8820 (N_8820,N_6945,N_6506);
or U8821 (N_8821,N_7916,N_7493);
or U8822 (N_8822,N_7104,N_7409);
or U8823 (N_8823,N_6719,N_6462);
xor U8824 (N_8824,N_7880,N_6781);
nand U8825 (N_8825,N_7082,N_7798);
nor U8826 (N_8826,N_6392,N_7098);
and U8827 (N_8827,N_6769,N_6074);
xor U8828 (N_8828,N_7105,N_6903);
nor U8829 (N_8829,N_6633,N_7999);
nand U8830 (N_8830,N_7458,N_7816);
or U8831 (N_8831,N_6071,N_7740);
nor U8832 (N_8832,N_6870,N_7674);
nor U8833 (N_8833,N_7177,N_7734);
xnor U8834 (N_8834,N_7106,N_7411);
nand U8835 (N_8835,N_7225,N_7402);
xnor U8836 (N_8836,N_6897,N_7031);
or U8837 (N_8837,N_7453,N_7400);
and U8838 (N_8838,N_6081,N_6212);
nor U8839 (N_8839,N_6377,N_7234);
or U8840 (N_8840,N_7163,N_6144);
nor U8841 (N_8841,N_6490,N_7382);
and U8842 (N_8842,N_6960,N_7957);
nand U8843 (N_8843,N_7873,N_6706);
or U8844 (N_8844,N_6642,N_6946);
nand U8845 (N_8845,N_7563,N_6944);
or U8846 (N_8846,N_6662,N_6883);
or U8847 (N_8847,N_7181,N_7555);
or U8848 (N_8848,N_7223,N_6211);
nor U8849 (N_8849,N_7836,N_6698);
and U8850 (N_8850,N_7145,N_7197);
nand U8851 (N_8851,N_7273,N_7423);
nor U8852 (N_8852,N_7491,N_7954);
nor U8853 (N_8853,N_6192,N_7856);
and U8854 (N_8854,N_7320,N_7427);
xor U8855 (N_8855,N_7167,N_7578);
nor U8856 (N_8856,N_6505,N_7941);
and U8857 (N_8857,N_7505,N_6741);
nor U8858 (N_8858,N_7020,N_7448);
or U8859 (N_8859,N_7250,N_6003);
nand U8860 (N_8860,N_7771,N_7449);
and U8861 (N_8861,N_7544,N_7425);
nor U8862 (N_8862,N_6892,N_7699);
nor U8863 (N_8863,N_7806,N_6439);
and U8864 (N_8864,N_6702,N_6654);
nor U8865 (N_8865,N_6755,N_6405);
or U8866 (N_8866,N_6911,N_6782);
and U8867 (N_8867,N_6251,N_7481);
nand U8868 (N_8868,N_7070,N_7972);
nor U8869 (N_8869,N_7116,N_7717);
and U8870 (N_8870,N_7634,N_6111);
and U8871 (N_8871,N_7877,N_7978);
nand U8872 (N_8872,N_7066,N_6314);
or U8873 (N_8873,N_7938,N_6328);
nor U8874 (N_8874,N_7339,N_7876);
or U8875 (N_8875,N_6197,N_6537);
and U8876 (N_8876,N_7779,N_7243);
or U8877 (N_8877,N_7628,N_7462);
or U8878 (N_8878,N_7032,N_6487);
or U8879 (N_8879,N_6260,N_6103);
nand U8880 (N_8880,N_6761,N_6526);
nand U8881 (N_8881,N_7543,N_7736);
or U8882 (N_8882,N_6258,N_7226);
nor U8883 (N_8883,N_6734,N_6583);
nor U8884 (N_8884,N_7695,N_6214);
and U8885 (N_8885,N_7782,N_6117);
and U8886 (N_8886,N_6316,N_6725);
or U8887 (N_8887,N_6554,N_7350);
or U8888 (N_8888,N_6665,N_7365);
nor U8889 (N_8889,N_7131,N_6492);
nand U8890 (N_8890,N_6965,N_7913);
and U8891 (N_8891,N_6886,N_6896);
and U8892 (N_8892,N_6348,N_7616);
or U8893 (N_8893,N_6636,N_7354);
and U8894 (N_8894,N_7259,N_7830);
nand U8895 (N_8895,N_7985,N_7375);
xor U8896 (N_8896,N_7841,N_6273);
nor U8897 (N_8897,N_6504,N_7931);
or U8898 (N_8898,N_6379,N_7387);
nand U8899 (N_8899,N_7926,N_7176);
xor U8900 (N_8900,N_7476,N_6266);
and U8901 (N_8901,N_7388,N_7024);
xnor U8902 (N_8902,N_6068,N_6901);
and U8903 (N_8903,N_6739,N_6219);
xnor U8904 (N_8904,N_7797,N_6977);
nand U8905 (N_8905,N_7432,N_7006);
and U8906 (N_8906,N_6341,N_7359);
nor U8907 (N_8907,N_6923,N_6243);
xnor U8908 (N_8908,N_6132,N_6882);
nand U8909 (N_8909,N_7054,N_6576);
nor U8910 (N_8910,N_7946,N_6035);
or U8911 (N_8911,N_7407,N_7561);
and U8912 (N_8912,N_7235,N_7881);
or U8913 (N_8913,N_7071,N_6723);
nand U8914 (N_8914,N_7415,N_7664);
nor U8915 (N_8915,N_7171,N_7213);
nor U8916 (N_8916,N_6542,N_6887);
nand U8917 (N_8917,N_7920,N_6153);
nand U8918 (N_8918,N_6588,N_6024);
nand U8919 (N_8919,N_7133,N_7672);
xor U8920 (N_8920,N_7569,N_7701);
xnor U8921 (N_8921,N_7658,N_6334);
nor U8922 (N_8922,N_7290,N_7508);
xnor U8923 (N_8923,N_6231,N_7399);
or U8924 (N_8924,N_6831,N_7085);
nor U8925 (N_8925,N_6095,N_6980);
nand U8926 (N_8926,N_6350,N_7445);
xnor U8927 (N_8927,N_6558,N_7392);
nor U8928 (N_8928,N_6322,N_7216);
and U8929 (N_8929,N_7091,N_7368);
nand U8930 (N_8930,N_7218,N_6777);
and U8931 (N_8931,N_7057,N_7345);
xnor U8932 (N_8932,N_6624,N_6442);
nor U8933 (N_8933,N_6703,N_6195);
nand U8934 (N_8934,N_7864,N_7315);
nor U8935 (N_8935,N_6028,N_6045);
nor U8936 (N_8936,N_6326,N_6609);
nor U8937 (N_8937,N_7370,N_7252);
nor U8938 (N_8938,N_7623,N_7746);
nand U8939 (N_8939,N_7045,N_6789);
xnor U8940 (N_8940,N_7016,N_7720);
nor U8941 (N_8941,N_6216,N_6949);
or U8942 (N_8942,N_6159,N_6270);
nand U8943 (N_8943,N_7805,N_7900);
or U8944 (N_8944,N_7199,N_7245);
or U8945 (N_8945,N_6829,N_6039);
or U8946 (N_8946,N_7367,N_6868);
xor U8947 (N_8947,N_7153,N_6398);
and U8948 (N_8948,N_7123,N_6733);
or U8949 (N_8949,N_7494,N_6847);
and U8950 (N_8950,N_7870,N_6908);
and U8951 (N_8951,N_6711,N_7648);
and U8952 (N_8952,N_7707,N_7477);
or U8953 (N_8953,N_6138,N_7228);
or U8954 (N_8954,N_6137,N_6100);
and U8955 (N_8955,N_6898,N_6173);
nor U8956 (N_8956,N_7254,N_6708);
nor U8957 (N_8957,N_7500,N_7143);
and U8958 (N_8958,N_6031,N_7326);
nor U8959 (N_8959,N_6559,N_6207);
nor U8960 (N_8960,N_6976,N_6802);
nor U8961 (N_8961,N_7723,N_6357);
nor U8962 (N_8962,N_7465,N_7550);
or U8963 (N_8963,N_7309,N_6133);
nand U8964 (N_8964,N_7995,N_6763);
nand U8965 (N_8965,N_6514,N_7789);
and U8966 (N_8966,N_6749,N_7653);
nor U8967 (N_8967,N_7833,N_7470);
or U8968 (N_8968,N_7607,N_6667);
nand U8969 (N_8969,N_7036,N_6872);
nand U8970 (N_8970,N_6178,N_6721);
and U8971 (N_8971,N_7480,N_7591);
nor U8972 (N_8972,N_6484,N_6731);
nor U8973 (N_8973,N_7330,N_7297);
xnor U8974 (N_8974,N_7262,N_7052);
and U8975 (N_8975,N_6574,N_6664);
or U8976 (N_8976,N_6759,N_7598);
nor U8977 (N_8977,N_6587,N_6751);
nand U8978 (N_8978,N_7179,N_6425);
xnor U8979 (N_8979,N_7232,N_7690);
nor U8980 (N_8980,N_6121,N_6382);
or U8981 (N_8981,N_6468,N_7109);
nand U8982 (N_8982,N_6393,N_6888);
nor U8983 (N_8983,N_6597,N_7360);
and U8984 (N_8984,N_7122,N_7702);
or U8985 (N_8985,N_6573,N_7759);
nor U8986 (N_8986,N_7487,N_7191);
xor U8987 (N_8987,N_6921,N_6592);
xnor U8988 (N_8988,N_6581,N_7963);
nand U8989 (N_8989,N_7220,N_6034);
nand U8990 (N_8990,N_6154,N_7023);
nor U8991 (N_8991,N_7072,N_6614);
nor U8992 (N_8992,N_7987,N_7136);
nor U8993 (N_8993,N_7460,N_6321);
nor U8994 (N_8994,N_6859,N_7906);
nand U8995 (N_8995,N_7726,N_7885);
and U8996 (N_8996,N_7526,N_7869);
nor U8997 (N_8997,N_6186,N_7874);
nor U8998 (N_8998,N_7332,N_6584);
or U8999 (N_8999,N_6050,N_6987);
xor U9000 (N_9000,N_6304,N_7384);
nor U9001 (N_9001,N_6087,N_7144);
and U9002 (N_9002,N_7120,N_6256);
and U9003 (N_9003,N_7186,N_7573);
or U9004 (N_9004,N_6399,N_6658);
nand U9005 (N_9005,N_6571,N_7785);
or U9006 (N_9006,N_7181,N_6363);
nor U9007 (N_9007,N_6674,N_6098);
and U9008 (N_9008,N_6757,N_6063);
nand U9009 (N_9009,N_7978,N_6820);
nand U9010 (N_9010,N_7162,N_7709);
nor U9011 (N_9011,N_6586,N_7194);
nand U9012 (N_9012,N_6190,N_7829);
nor U9013 (N_9013,N_7217,N_7122);
and U9014 (N_9014,N_6497,N_7728);
or U9015 (N_9015,N_7849,N_6075);
and U9016 (N_9016,N_7842,N_6707);
xnor U9017 (N_9017,N_6000,N_7052);
and U9018 (N_9018,N_7318,N_7930);
xnor U9019 (N_9019,N_6247,N_7142);
and U9020 (N_9020,N_7281,N_7962);
xnor U9021 (N_9021,N_7426,N_7653);
nand U9022 (N_9022,N_7930,N_6742);
xor U9023 (N_9023,N_7176,N_6946);
nand U9024 (N_9024,N_6027,N_6586);
nor U9025 (N_9025,N_6277,N_7704);
or U9026 (N_9026,N_6930,N_6874);
and U9027 (N_9027,N_6178,N_7694);
or U9028 (N_9028,N_7353,N_6045);
or U9029 (N_9029,N_7999,N_7556);
nand U9030 (N_9030,N_6293,N_7799);
nand U9031 (N_9031,N_6497,N_7398);
xor U9032 (N_9032,N_7455,N_7275);
and U9033 (N_9033,N_7709,N_6866);
and U9034 (N_9034,N_6437,N_6897);
or U9035 (N_9035,N_7285,N_6390);
nor U9036 (N_9036,N_6397,N_6615);
and U9037 (N_9037,N_7370,N_6407);
nand U9038 (N_9038,N_7980,N_6641);
nor U9039 (N_9039,N_6159,N_6487);
nor U9040 (N_9040,N_7100,N_7831);
nor U9041 (N_9041,N_7996,N_7449);
or U9042 (N_9042,N_7692,N_6491);
and U9043 (N_9043,N_7273,N_7497);
or U9044 (N_9044,N_6500,N_7754);
nand U9045 (N_9045,N_6694,N_7147);
nor U9046 (N_9046,N_6537,N_6652);
nor U9047 (N_9047,N_7646,N_6026);
or U9048 (N_9048,N_6081,N_6528);
or U9049 (N_9049,N_7122,N_7360);
nor U9050 (N_9050,N_7072,N_6652);
nand U9051 (N_9051,N_7158,N_6062);
nor U9052 (N_9052,N_6030,N_6088);
nor U9053 (N_9053,N_6147,N_7062);
nor U9054 (N_9054,N_6134,N_6917);
nand U9055 (N_9055,N_7681,N_6565);
nor U9056 (N_9056,N_6116,N_6859);
or U9057 (N_9057,N_7637,N_7471);
or U9058 (N_9058,N_6052,N_7728);
nand U9059 (N_9059,N_6778,N_7240);
nor U9060 (N_9060,N_6048,N_6341);
xnor U9061 (N_9061,N_7058,N_7314);
nor U9062 (N_9062,N_6685,N_6891);
nor U9063 (N_9063,N_7686,N_6535);
and U9064 (N_9064,N_6247,N_6580);
or U9065 (N_9065,N_6177,N_7493);
and U9066 (N_9066,N_6690,N_6388);
nor U9067 (N_9067,N_7786,N_7710);
nor U9068 (N_9068,N_6088,N_6477);
nand U9069 (N_9069,N_7183,N_6394);
nand U9070 (N_9070,N_6562,N_6194);
nand U9071 (N_9071,N_6181,N_7138);
or U9072 (N_9072,N_6317,N_7176);
xnor U9073 (N_9073,N_7436,N_7303);
or U9074 (N_9074,N_6709,N_7816);
nand U9075 (N_9075,N_6017,N_6054);
nand U9076 (N_9076,N_7818,N_7622);
nor U9077 (N_9077,N_6254,N_7503);
or U9078 (N_9078,N_6735,N_7583);
xnor U9079 (N_9079,N_6722,N_7213);
nor U9080 (N_9080,N_6344,N_6276);
or U9081 (N_9081,N_7497,N_6647);
nor U9082 (N_9082,N_6987,N_6017);
xor U9083 (N_9083,N_7429,N_6551);
nand U9084 (N_9084,N_6712,N_7212);
xor U9085 (N_9085,N_7673,N_6228);
nand U9086 (N_9086,N_6268,N_7774);
nor U9087 (N_9087,N_7219,N_6835);
nor U9088 (N_9088,N_7774,N_7924);
nor U9089 (N_9089,N_6098,N_7866);
or U9090 (N_9090,N_7258,N_6757);
and U9091 (N_9091,N_7580,N_6799);
xnor U9092 (N_9092,N_6843,N_7591);
and U9093 (N_9093,N_7868,N_6806);
and U9094 (N_9094,N_7637,N_6256);
and U9095 (N_9095,N_7361,N_6119);
nand U9096 (N_9096,N_6053,N_7942);
xor U9097 (N_9097,N_7928,N_7492);
nand U9098 (N_9098,N_6631,N_7936);
xnor U9099 (N_9099,N_6597,N_6932);
nor U9100 (N_9100,N_7720,N_6734);
nor U9101 (N_9101,N_6110,N_6388);
or U9102 (N_9102,N_7289,N_6970);
or U9103 (N_9103,N_7712,N_7750);
and U9104 (N_9104,N_7291,N_7248);
or U9105 (N_9105,N_7946,N_6961);
or U9106 (N_9106,N_6088,N_6169);
nand U9107 (N_9107,N_6106,N_6824);
or U9108 (N_9108,N_7604,N_6234);
nor U9109 (N_9109,N_7856,N_6924);
nand U9110 (N_9110,N_7057,N_6626);
nor U9111 (N_9111,N_7481,N_6221);
and U9112 (N_9112,N_6588,N_7568);
or U9113 (N_9113,N_7896,N_7962);
or U9114 (N_9114,N_6138,N_6348);
and U9115 (N_9115,N_7120,N_6199);
or U9116 (N_9116,N_7631,N_6445);
and U9117 (N_9117,N_6514,N_7087);
nand U9118 (N_9118,N_6018,N_7313);
or U9119 (N_9119,N_7812,N_6182);
xnor U9120 (N_9120,N_6594,N_7040);
nand U9121 (N_9121,N_7504,N_6979);
xor U9122 (N_9122,N_7499,N_6239);
or U9123 (N_9123,N_6219,N_7063);
nand U9124 (N_9124,N_6643,N_6243);
and U9125 (N_9125,N_7805,N_7810);
nor U9126 (N_9126,N_7677,N_6323);
nor U9127 (N_9127,N_7227,N_7374);
or U9128 (N_9128,N_7037,N_6989);
xnor U9129 (N_9129,N_6038,N_6396);
nor U9130 (N_9130,N_6692,N_7941);
or U9131 (N_9131,N_6024,N_7165);
nand U9132 (N_9132,N_7790,N_7884);
and U9133 (N_9133,N_6075,N_7423);
or U9134 (N_9134,N_6920,N_6416);
and U9135 (N_9135,N_6118,N_6714);
and U9136 (N_9136,N_7149,N_6507);
or U9137 (N_9137,N_6805,N_7501);
or U9138 (N_9138,N_6703,N_7041);
nor U9139 (N_9139,N_7559,N_6541);
nor U9140 (N_9140,N_6491,N_6809);
and U9141 (N_9141,N_6415,N_6114);
nor U9142 (N_9142,N_7110,N_6168);
nand U9143 (N_9143,N_7241,N_7402);
or U9144 (N_9144,N_6916,N_7097);
nand U9145 (N_9145,N_7773,N_6371);
nor U9146 (N_9146,N_7249,N_6568);
nor U9147 (N_9147,N_6613,N_6233);
nand U9148 (N_9148,N_7098,N_6016);
nand U9149 (N_9149,N_7866,N_6164);
nand U9150 (N_9150,N_6245,N_7600);
and U9151 (N_9151,N_7501,N_6742);
nand U9152 (N_9152,N_7622,N_7443);
nor U9153 (N_9153,N_7384,N_7904);
nand U9154 (N_9154,N_7081,N_6955);
nand U9155 (N_9155,N_6010,N_7002);
nor U9156 (N_9156,N_7250,N_6680);
or U9157 (N_9157,N_6261,N_6325);
and U9158 (N_9158,N_6806,N_6910);
or U9159 (N_9159,N_6668,N_7970);
nor U9160 (N_9160,N_7692,N_6305);
and U9161 (N_9161,N_7194,N_6226);
or U9162 (N_9162,N_7086,N_6708);
nand U9163 (N_9163,N_7779,N_6153);
nand U9164 (N_9164,N_7310,N_6628);
nand U9165 (N_9165,N_7342,N_7652);
nand U9166 (N_9166,N_7145,N_7229);
and U9167 (N_9167,N_6512,N_6126);
or U9168 (N_9168,N_7073,N_6899);
or U9169 (N_9169,N_7853,N_6123);
or U9170 (N_9170,N_6784,N_6951);
and U9171 (N_9171,N_7742,N_6387);
and U9172 (N_9172,N_6950,N_7509);
nor U9173 (N_9173,N_6035,N_7078);
or U9174 (N_9174,N_6463,N_7465);
and U9175 (N_9175,N_7244,N_6075);
and U9176 (N_9176,N_7679,N_6835);
and U9177 (N_9177,N_7858,N_7927);
or U9178 (N_9178,N_6217,N_7051);
or U9179 (N_9179,N_7100,N_7315);
nand U9180 (N_9180,N_6477,N_7272);
nor U9181 (N_9181,N_6340,N_6329);
nand U9182 (N_9182,N_7116,N_7132);
and U9183 (N_9183,N_6480,N_6468);
nand U9184 (N_9184,N_6424,N_7594);
nor U9185 (N_9185,N_6695,N_6945);
or U9186 (N_9186,N_7045,N_7559);
or U9187 (N_9187,N_6598,N_6024);
or U9188 (N_9188,N_6854,N_7811);
xor U9189 (N_9189,N_6130,N_6009);
or U9190 (N_9190,N_7562,N_7802);
and U9191 (N_9191,N_6228,N_6779);
nand U9192 (N_9192,N_7178,N_7538);
nand U9193 (N_9193,N_6452,N_7913);
or U9194 (N_9194,N_7728,N_7759);
nor U9195 (N_9195,N_7483,N_6116);
or U9196 (N_9196,N_6984,N_6740);
nor U9197 (N_9197,N_7457,N_7199);
xor U9198 (N_9198,N_7293,N_6272);
and U9199 (N_9199,N_7474,N_7964);
nand U9200 (N_9200,N_6887,N_7770);
xor U9201 (N_9201,N_7081,N_6695);
or U9202 (N_9202,N_7563,N_7714);
nor U9203 (N_9203,N_6833,N_7780);
nand U9204 (N_9204,N_7027,N_6964);
nand U9205 (N_9205,N_6934,N_7322);
nand U9206 (N_9206,N_6485,N_6746);
nand U9207 (N_9207,N_6759,N_7043);
and U9208 (N_9208,N_7412,N_6985);
nand U9209 (N_9209,N_6349,N_7681);
nand U9210 (N_9210,N_7614,N_6102);
or U9211 (N_9211,N_6372,N_7978);
nand U9212 (N_9212,N_6554,N_6009);
and U9213 (N_9213,N_6631,N_7838);
and U9214 (N_9214,N_7178,N_6067);
nand U9215 (N_9215,N_6624,N_7497);
and U9216 (N_9216,N_7944,N_7770);
and U9217 (N_9217,N_6639,N_6751);
and U9218 (N_9218,N_6684,N_7133);
xnor U9219 (N_9219,N_7444,N_7002);
and U9220 (N_9220,N_7075,N_6234);
and U9221 (N_9221,N_7059,N_6554);
or U9222 (N_9222,N_7155,N_6031);
nand U9223 (N_9223,N_6542,N_6724);
or U9224 (N_9224,N_7772,N_6180);
and U9225 (N_9225,N_7560,N_6102);
xnor U9226 (N_9226,N_6300,N_7185);
nand U9227 (N_9227,N_6759,N_6717);
nor U9228 (N_9228,N_6732,N_7660);
xnor U9229 (N_9229,N_7841,N_6078);
nand U9230 (N_9230,N_7440,N_7016);
or U9231 (N_9231,N_6464,N_7707);
nor U9232 (N_9232,N_7124,N_6054);
nor U9233 (N_9233,N_7893,N_6972);
and U9234 (N_9234,N_6537,N_6554);
nand U9235 (N_9235,N_6752,N_6253);
and U9236 (N_9236,N_6852,N_6862);
nand U9237 (N_9237,N_7438,N_7882);
nand U9238 (N_9238,N_6435,N_6546);
and U9239 (N_9239,N_6246,N_6172);
nand U9240 (N_9240,N_7356,N_7921);
nand U9241 (N_9241,N_7818,N_7176);
or U9242 (N_9242,N_6525,N_7829);
nor U9243 (N_9243,N_6971,N_7658);
nor U9244 (N_9244,N_7686,N_7730);
nand U9245 (N_9245,N_6796,N_7654);
nor U9246 (N_9246,N_7937,N_6821);
nand U9247 (N_9247,N_7208,N_6901);
nand U9248 (N_9248,N_7026,N_6113);
and U9249 (N_9249,N_6876,N_6899);
nand U9250 (N_9250,N_6440,N_7153);
and U9251 (N_9251,N_7675,N_6995);
nand U9252 (N_9252,N_6921,N_7385);
and U9253 (N_9253,N_6323,N_6344);
or U9254 (N_9254,N_6907,N_7529);
nand U9255 (N_9255,N_7127,N_6573);
or U9256 (N_9256,N_7039,N_7886);
and U9257 (N_9257,N_6894,N_6170);
and U9258 (N_9258,N_7424,N_6359);
nor U9259 (N_9259,N_7845,N_6017);
xor U9260 (N_9260,N_7267,N_7090);
nor U9261 (N_9261,N_7126,N_7917);
nor U9262 (N_9262,N_6900,N_6087);
xor U9263 (N_9263,N_6963,N_6990);
or U9264 (N_9264,N_7655,N_6087);
or U9265 (N_9265,N_6057,N_6361);
nand U9266 (N_9266,N_6221,N_6447);
nor U9267 (N_9267,N_6449,N_6321);
xor U9268 (N_9268,N_7959,N_7903);
and U9269 (N_9269,N_7054,N_7234);
and U9270 (N_9270,N_6626,N_6232);
and U9271 (N_9271,N_6599,N_6480);
or U9272 (N_9272,N_6264,N_6472);
xor U9273 (N_9273,N_6331,N_6366);
nand U9274 (N_9274,N_7129,N_6506);
nand U9275 (N_9275,N_6087,N_6321);
nand U9276 (N_9276,N_7676,N_6737);
or U9277 (N_9277,N_7490,N_7373);
nand U9278 (N_9278,N_6172,N_7702);
or U9279 (N_9279,N_7502,N_7441);
or U9280 (N_9280,N_7923,N_6806);
nand U9281 (N_9281,N_6856,N_7801);
and U9282 (N_9282,N_6010,N_6278);
or U9283 (N_9283,N_7353,N_6257);
nor U9284 (N_9284,N_7730,N_6830);
nor U9285 (N_9285,N_6079,N_6255);
nand U9286 (N_9286,N_7241,N_6798);
or U9287 (N_9287,N_6927,N_6380);
nand U9288 (N_9288,N_6681,N_7062);
and U9289 (N_9289,N_7508,N_6559);
or U9290 (N_9290,N_7830,N_7633);
or U9291 (N_9291,N_6198,N_7695);
nor U9292 (N_9292,N_7611,N_7025);
nand U9293 (N_9293,N_6977,N_6456);
or U9294 (N_9294,N_7177,N_6581);
nor U9295 (N_9295,N_7867,N_6532);
nand U9296 (N_9296,N_6314,N_7567);
nand U9297 (N_9297,N_6728,N_6700);
or U9298 (N_9298,N_7983,N_7186);
xnor U9299 (N_9299,N_7321,N_7129);
and U9300 (N_9300,N_6566,N_7679);
nor U9301 (N_9301,N_6488,N_7124);
nor U9302 (N_9302,N_6613,N_6927);
xor U9303 (N_9303,N_6304,N_6496);
and U9304 (N_9304,N_6800,N_6942);
nor U9305 (N_9305,N_6107,N_7753);
or U9306 (N_9306,N_6693,N_7094);
nand U9307 (N_9307,N_6278,N_6154);
nor U9308 (N_9308,N_6744,N_7790);
nand U9309 (N_9309,N_6631,N_6295);
or U9310 (N_9310,N_6772,N_7272);
nor U9311 (N_9311,N_6010,N_7949);
and U9312 (N_9312,N_6534,N_7828);
or U9313 (N_9313,N_7705,N_7927);
nand U9314 (N_9314,N_6526,N_6884);
nand U9315 (N_9315,N_7596,N_7878);
nor U9316 (N_9316,N_7472,N_7266);
or U9317 (N_9317,N_7179,N_7735);
or U9318 (N_9318,N_6518,N_7597);
xnor U9319 (N_9319,N_6509,N_6593);
nand U9320 (N_9320,N_6002,N_7410);
nor U9321 (N_9321,N_6289,N_6412);
xnor U9322 (N_9322,N_7114,N_6946);
and U9323 (N_9323,N_7322,N_7447);
or U9324 (N_9324,N_6524,N_7783);
xor U9325 (N_9325,N_7193,N_7432);
nor U9326 (N_9326,N_6858,N_6483);
xnor U9327 (N_9327,N_6463,N_7322);
nor U9328 (N_9328,N_6628,N_7808);
or U9329 (N_9329,N_7655,N_6890);
and U9330 (N_9330,N_6538,N_7786);
nand U9331 (N_9331,N_6776,N_7365);
nand U9332 (N_9332,N_7323,N_6713);
nand U9333 (N_9333,N_6659,N_7155);
nor U9334 (N_9334,N_7181,N_6975);
or U9335 (N_9335,N_7632,N_7523);
or U9336 (N_9336,N_7865,N_7214);
nor U9337 (N_9337,N_7694,N_6224);
and U9338 (N_9338,N_6149,N_6455);
nor U9339 (N_9339,N_6154,N_7767);
nand U9340 (N_9340,N_7650,N_6054);
and U9341 (N_9341,N_7488,N_6740);
and U9342 (N_9342,N_6650,N_7033);
or U9343 (N_9343,N_6382,N_6746);
nor U9344 (N_9344,N_6829,N_7599);
and U9345 (N_9345,N_7800,N_7876);
xor U9346 (N_9346,N_6976,N_6303);
nand U9347 (N_9347,N_7054,N_6427);
nand U9348 (N_9348,N_6583,N_7722);
nor U9349 (N_9349,N_6250,N_7285);
nand U9350 (N_9350,N_7305,N_7523);
nand U9351 (N_9351,N_6142,N_6212);
nor U9352 (N_9352,N_6134,N_7668);
nand U9353 (N_9353,N_6225,N_6539);
or U9354 (N_9354,N_7554,N_6716);
nand U9355 (N_9355,N_6138,N_7721);
nand U9356 (N_9356,N_6091,N_6728);
nor U9357 (N_9357,N_7042,N_6733);
or U9358 (N_9358,N_7171,N_6529);
or U9359 (N_9359,N_6986,N_6612);
nand U9360 (N_9360,N_7410,N_6889);
nand U9361 (N_9361,N_6351,N_7487);
nor U9362 (N_9362,N_7353,N_7264);
or U9363 (N_9363,N_6040,N_6538);
or U9364 (N_9364,N_7581,N_6444);
nor U9365 (N_9365,N_7527,N_7310);
nor U9366 (N_9366,N_6728,N_6922);
nand U9367 (N_9367,N_6941,N_6759);
nor U9368 (N_9368,N_6094,N_7754);
and U9369 (N_9369,N_6560,N_6254);
xor U9370 (N_9370,N_6379,N_7241);
xnor U9371 (N_9371,N_6115,N_6455);
nand U9372 (N_9372,N_7650,N_7257);
and U9373 (N_9373,N_7346,N_6736);
or U9374 (N_9374,N_6098,N_6046);
or U9375 (N_9375,N_7518,N_7103);
or U9376 (N_9376,N_7780,N_6592);
or U9377 (N_9377,N_6670,N_6640);
nor U9378 (N_9378,N_7778,N_6295);
nand U9379 (N_9379,N_6837,N_7336);
nand U9380 (N_9380,N_7319,N_7831);
or U9381 (N_9381,N_6311,N_7142);
nand U9382 (N_9382,N_7164,N_7721);
or U9383 (N_9383,N_7410,N_7917);
and U9384 (N_9384,N_7504,N_7312);
xnor U9385 (N_9385,N_7288,N_6529);
or U9386 (N_9386,N_6157,N_7593);
xor U9387 (N_9387,N_6231,N_7277);
or U9388 (N_9388,N_7857,N_7797);
or U9389 (N_9389,N_6477,N_6508);
and U9390 (N_9390,N_7737,N_7621);
or U9391 (N_9391,N_6561,N_6404);
nand U9392 (N_9392,N_6365,N_6928);
or U9393 (N_9393,N_7383,N_6009);
or U9394 (N_9394,N_7535,N_7715);
nand U9395 (N_9395,N_6085,N_6274);
nand U9396 (N_9396,N_7927,N_7427);
nand U9397 (N_9397,N_6389,N_7100);
nor U9398 (N_9398,N_7172,N_6579);
nand U9399 (N_9399,N_6293,N_7302);
and U9400 (N_9400,N_7950,N_6750);
nand U9401 (N_9401,N_7849,N_6272);
nor U9402 (N_9402,N_6221,N_6923);
and U9403 (N_9403,N_6633,N_7136);
nor U9404 (N_9404,N_7650,N_7526);
or U9405 (N_9405,N_6524,N_6520);
nor U9406 (N_9406,N_6689,N_6676);
nand U9407 (N_9407,N_6779,N_6888);
nor U9408 (N_9408,N_7467,N_7798);
nor U9409 (N_9409,N_7486,N_7976);
xor U9410 (N_9410,N_6250,N_6721);
or U9411 (N_9411,N_7947,N_6567);
and U9412 (N_9412,N_6855,N_7322);
or U9413 (N_9413,N_6790,N_6128);
nor U9414 (N_9414,N_7769,N_6329);
nor U9415 (N_9415,N_6724,N_6533);
nor U9416 (N_9416,N_7622,N_7831);
nor U9417 (N_9417,N_6213,N_7107);
or U9418 (N_9418,N_6731,N_6375);
or U9419 (N_9419,N_6087,N_6741);
nor U9420 (N_9420,N_6556,N_6751);
nor U9421 (N_9421,N_7359,N_7843);
and U9422 (N_9422,N_7430,N_6446);
or U9423 (N_9423,N_7499,N_7805);
and U9424 (N_9424,N_6107,N_6904);
nand U9425 (N_9425,N_7876,N_6582);
or U9426 (N_9426,N_6747,N_7508);
and U9427 (N_9427,N_7320,N_6864);
nand U9428 (N_9428,N_7372,N_6499);
and U9429 (N_9429,N_6826,N_6754);
xor U9430 (N_9430,N_7895,N_7929);
nand U9431 (N_9431,N_6891,N_7832);
nand U9432 (N_9432,N_7924,N_7809);
nand U9433 (N_9433,N_6776,N_7903);
or U9434 (N_9434,N_7413,N_7146);
or U9435 (N_9435,N_7162,N_7440);
nand U9436 (N_9436,N_7312,N_6679);
or U9437 (N_9437,N_7788,N_7187);
or U9438 (N_9438,N_7348,N_6667);
and U9439 (N_9439,N_7265,N_7662);
nand U9440 (N_9440,N_6569,N_6953);
and U9441 (N_9441,N_7607,N_6940);
nor U9442 (N_9442,N_7533,N_7848);
xor U9443 (N_9443,N_7348,N_7277);
nand U9444 (N_9444,N_6594,N_6677);
and U9445 (N_9445,N_7555,N_6740);
nand U9446 (N_9446,N_7880,N_7179);
and U9447 (N_9447,N_6384,N_6035);
nand U9448 (N_9448,N_7049,N_7804);
xnor U9449 (N_9449,N_6108,N_6330);
or U9450 (N_9450,N_6023,N_6281);
or U9451 (N_9451,N_7492,N_6195);
or U9452 (N_9452,N_6076,N_7135);
nand U9453 (N_9453,N_7345,N_7378);
nor U9454 (N_9454,N_6618,N_7886);
xnor U9455 (N_9455,N_7784,N_6653);
or U9456 (N_9456,N_7108,N_7843);
and U9457 (N_9457,N_6037,N_7524);
nor U9458 (N_9458,N_6489,N_7553);
and U9459 (N_9459,N_7413,N_7791);
or U9460 (N_9460,N_7117,N_7030);
nor U9461 (N_9461,N_7880,N_7264);
nand U9462 (N_9462,N_6539,N_7506);
nand U9463 (N_9463,N_6148,N_7751);
and U9464 (N_9464,N_6805,N_6872);
nand U9465 (N_9465,N_7304,N_6881);
nand U9466 (N_9466,N_7335,N_6827);
and U9467 (N_9467,N_7991,N_6909);
and U9468 (N_9468,N_6547,N_7950);
nor U9469 (N_9469,N_6844,N_6657);
and U9470 (N_9470,N_6650,N_6986);
or U9471 (N_9471,N_7049,N_7374);
nand U9472 (N_9472,N_6921,N_6456);
or U9473 (N_9473,N_6825,N_7665);
and U9474 (N_9474,N_7774,N_6958);
nand U9475 (N_9475,N_7873,N_7485);
nor U9476 (N_9476,N_6141,N_6603);
nand U9477 (N_9477,N_6316,N_7133);
or U9478 (N_9478,N_7995,N_6310);
and U9479 (N_9479,N_7661,N_6636);
or U9480 (N_9480,N_6123,N_7432);
nor U9481 (N_9481,N_7223,N_7983);
nor U9482 (N_9482,N_7837,N_6065);
and U9483 (N_9483,N_6463,N_6292);
xnor U9484 (N_9484,N_7107,N_6192);
or U9485 (N_9485,N_7814,N_6229);
and U9486 (N_9486,N_6215,N_6747);
nor U9487 (N_9487,N_6195,N_6936);
nor U9488 (N_9488,N_6558,N_7764);
nor U9489 (N_9489,N_7071,N_7431);
nor U9490 (N_9490,N_6891,N_6325);
and U9491 (N_9491,N_7009,N_7674);
and U9492 (N_9492,N_7364,N_7206);
or U9493 (N_9493,N_6252,N_7572);
nor U9494 (N_9494,N_7530,N_6995);
nor U9495 (N_9495,N_7615,N_6921);
nor U9496 (N_9496,N_7215,N_7195);
or U9497 (N_9497,N_6535,N_6778);
and U9498 (N_9498,N_6291,N_6516);
or U9499 (N_9499,N_6120,N_7956);
or U9500 (N_9500,N_6630,N_7641);
xnor U9501 (N_9501,N_6967,N_7296);
or U9502 (N_9502,N_7382,N_7933);
nor U9503 (N_9503,N_6837,N_7795);
nand U9504 (N_9504,N_7297,N_6565);
or U9505 (N_9505,N_7269,N_6509);
nor U9506 (N_9506,N_6564,N_7547);
or U9507 (N_9507,N_7451,N_6436);
or U9508 (N_9508,N_7879,N_6955);
and U9509 (N_9509,N_6260,N_7145);
nor U9510 (N_9510,N_7323,N_6228);
and U9511 (N_9511,N_6706,N_7702);
or U9512 (N_9512,N_7912,N_7497);
or U9513 (N_9513,N_7392,N_6109);
nor U9514 (N_9514,N_6054,N_6606);
xor U9515 (N_9515,N_6913,N_6045);
xor U9516 (N_9516,N_7355,N_6296);
xnor U9517 (N_9517,N_7180,N_6473);
and U9518 (N_9518,N_7888,N_6022);
nand U9519 (N_9519,N_7045,N_6225);
nor U9520 (N_9520,N_6298,N_6676);
or U9521 (N_9521,N_7560,N_6386);
nand U9522 (N_9522,N_6082,N_6503);
nor U9523 (N_9523,N_7111,N_7910);
and U9524 (N_9524,N_6185,N_6652);
nor U9525 (N_9525,N_6054,N_6505);
and U9526 (N_9526,N_6190,N_7737);
nor U9527 (N_9527,N_7958,N_7244);
and U9528 (N_9528,N_7858,N_7989);
nand U9529 (N_9529,N_7058,N_7400);
nand U9530 (N_9530,N_6676,N_7700);
nor U9531 (N_9531,N_7315,N_6306);
nand U9532 (N_9532,N_6905,N_6144);
nor U9533 (N_9533,N_7872,N_6863);
and U9534 (N_9534,N_7944,N_6738);
nand U9535 (N_9535,N_6819,N_6210);
xnor U9536 (N_9536,N_7064,N_6402);
and U9537 (N_9537,N_6831,N_6141);
xnor U9538 (N_9538,N_7097,N_7045);
nand U9539 (N_9539,N_7568,N_6698);
nand U9540 (N_9540,N_6614,N_7394);
and U9541 (N_9541,N_7358,N_7271);
or U9542 (N_9542,N_6214,N_6209);
or U9543 (N_9543,N_6650,N_6835);
and U9544 (N_9544,N_6936,N_6194);
and U9545 (N_9545,N_6562,N_6162);
or U9546 (N_9546,N_7203,N_6388);
xor U9547 (N_9547,N_7973,N_7397);
nor U9548 (N_9548,N_6185,N_7776);
xor U9549 (N_9549,N_6709,N_6011);
xnor U9550 (N_9550,N_6017,N_6013);
or U9551 (N_9551,N_7435,N_6699);
nand U9552 (N_9552,N_6881,N_6953);
nand U9553 (N_9553,N_6563,N_7116);
and U9554 (N_9554,N_7702,N_6429);
or U9555 (N_9555,N_7089,N_6641);
or U9556 (N_9556,N_7903,N_7179);
or U9557 (N_9557,N_6782,N_7121);
nand U9558 (N_9558,N_7699,N_7857);
and U9559 (N_9559,N_6894,N_6093);
nor U9560 (N_9560,N_7657,N_6539);
nand U9561 (N_9561,N_6856,N_6957);
or U9562 (N_9562,N_7879,N_6140);
nand U9563 (N_9563,N_7190,N_7279);
xnor U9564 (N_9564,N_7642,N_7525);
nor U9565 (N_9565,N_6716,N_6790);
nand U9566 (N_9566,N_7572,N_6173);
or U9567 (N_9567,N_7242,N_7590);
nand U9568 (N_9568,N_6935,N_6561);
and U9569 (N_9569,N_6210,N_6048);
or U9570 (N_9570,N_6265,N_7649);
xnor U9571 (N_9571,N_6381,N_6880);
nand U9572 (N_9572,N_6686,N_6302);
nand U9573 (N_9573,N_7121,N_6118);
nand U9574 (N_9574,N_6991,N_7322);
or U9575 (N_9575,N_6284,N_7969);
nor U9576 (N_9576,N_6621,N_7926);
or U9577 (N_9577,N_6393,N_7417);
nand U9578 (N_9578,N_6507,N_6697);
nor U9579 (N_9579,N_6968,N_6138);
and U9580 (N_9580,N_6544,N_6605);
nand U9581 (N_9581,N_6307,N_7693);
or U9582 (N_9582,N_6901,N_6578);
nand U9583 (N_9583,N_7561,N_6170);
nand U9584 (N_9584,N_6947,N_6493);
nand U9585 (N_9585,N_7159,N_7395);
nand U9586 (N_9586,N_7554,N_7411);
nand U9587 (N_9587,N_7159,N_6533);
nor U9588 (N_9588,N_7058,N_6237);
nor U9589 (N_9589,N_7276,N_6402);
nor U9590 (N_9590,N_7864,N_7016);
or U9591 (N_9591,N_7929,N_7362);
and U9592 (N_9592,N_6860,N_7964);
nand U9593 (N_9593,N_7898,N_7344);
nor U9594 (N_9594,N_6084,N_6584);
and U9595 (N_9595,N_7939,N_6100);
and U9596 (N_9596,N_6768,N_7108);
and U9597 (N_9597,N_7960,N_6997);
or U9598 (N_9598,N_7024,N_7451);
or U9599 (N_9599,N_7718,N_7446);
nand U9600 (N_9600,N_7984,N_6700);
or U9601 (N_9601,N_7318,N_6042);
xor U9602 (N_9602,N_7339,N_7156);
or U9603 (N_9603,N_7844,N_7321);
nor U9604 (N_9604,N_7239,N_6668);
or U9605 (N_9605,N_6233,N_6750);
or U9606 (N_9606,N_7017,N_6719);
and U9607 (N_9607,N_7559,N_6348);
or U9608 (N_9608,N_7390,N_6871);
or U9609 (N_9609,N_6286,N_7490);
and U9610 (N_9610,N_6502,N_6721);
nand U9611 (N_9611,N_7601,N_7274);
or U9612 (N_9612,N_6472,N_7750);
xor U9613 (N_9613,N_6234,N_6008);
and U9614 (N_9614,N_6926,N_7943);
xor U9615 (N_9615,N_7159,N_7300);
or U9616 (N_9616,N_6563,N_6865);
and U9617 (N_9617,N_6868,N_6447);
nand U9618 (N_9618,N_6873,N_7518);
or U9619 (N_9619,N_7434,N_7061);
or U9620 (N_9620,N_6755,N_7242);
nand U9621 (N_9621,N_7036,N_7131);
and U9622 (N_9622,N_6714,N_6096);
nor U9623 (N_9623,N_7104,N_7745);
or U9624 (N_9624,N_6250,N_6495);
or U9625 (N_9625,N_7090,N_6138);
nand U9626 (N_9626,N_7040,N_7381);
nand U9627 (N_9627,N_7337,N_6668);
nor U9628 (N_9628,N_7535,N_6794);
nor U9629 (N_9629,N_6684,N_6380);
and U9630 (N_9630,N_7100,N_6799);
nand U9631 (N_9631,N_7817,N_6254);
nor U9632 (N_9632,N_6861,N_6075);
nor U9633 (N_9633,N_6832,N_7817);
or U9634 (N_9634,N_6825,N_7325);
or U9635 (N_9635,N_6642,N_6470);
and U9636 (N_9636,N_7306,N_6994);
and U9637 (N_9637,N_7728,N_7587);
or U9638 (N_9638,N_7760,N_6105);
and U9639 (N_9639,N_7840,N_7645);
or U9640 (N_9640,N_6381,N_6544);
nand U9641 (N_9641,N_6238,N_7346);
or U9642 (N_9642,N_7960,N_7998);
and U9643 (N_9643,N_6319,N_7060);
or U9644 (N_9644,N_7126,N_7683);
and U9645 (N_9645,N_7143,N_6281);
nand U9646 (N_9646,N_7340,N_7379);
nand U9647 (N_9647,N_7084,N_6037);
xnor U9648 (N_9648,N_7037,N_7873);
nor U9649 (N_9649,N_7902,N_6827);
or U9650 (N_9650,N_7015,N_6893);
or U9651 (N_9651,N_7710,N_7191);
nor U9652 (N_9652,N_6963,N_6354);
or U9653 (N_9653,N_6309,N_7467);
and U9654 (N_9654,N_6972,N_7867);
and U9655 (N_9655,N_6556,N_6606);
nor U9656 (N_9656,N_6635,N_6961);
or U9657 (N_9657,N_7514,N_6531);
nor U9658 (N_9658,N_7189,N_7571);
and U9659 (N_9659,N_7149,N_7618);
nor U9660 (N_9660,N_6520,N_7218);
nor U9661 (N_9661,N_6475,N_7127);
xor U9662 (N_9662,N_7355,N_7748);
or U9663 (N_9663,N_6091,N_6719);
and U9664 (N_9664,N_7782,N_6031);
xor U9665 (N_9665,N_7921,N_6056);
or U9666 (N_9666,N_6190,N_6098);
xor U9667 (N_9667,N_7174,N_7266);
xnor U9668 (N_9668,N_6477,N_7021);
nand U9669 (N_9669,N_7900,N_6829);
nor U9670 (N_9670,N_6735,N_7691);
and U9671 (N_9671,N_6331,N_7146);
nor U9672 (N_9672,N_6069,N_7638);
or U9673 (N_9673,N_7935,N_6530);
and U9674 (N_9674,N_6444,N_6323);
nor U9675 (N_9675,N_7937,N_7193);
and U9676 (N_9676,N_7442,N_6897);
nor U9677 (N_9677,N_6928,N_6318);
or U9678 (N_9678,N_7079,N_6324);
xnor U9679 (N_9679,N_7762,N_7526);
nand U9680 (N_9680,N_6872,N_7915);
nor U9681 (N_9681,N_6090,N_7823);
xnor U9682 (N_9682,N_7562,N_6929);
nand U9683 (N_9683,N_6229,N_6902);
nor U9684 (N_9684,N_7917,N_7232);
and U9685 (N_9685,N_7059,N_7872);
and U9686 (N_9686,N_7505,N_6946);
xor U9687 (N_9687,N_6993,N_6557);
or U9688 (N_9688,N_6758,N_6080);
and U9689 (N_9689,N_6206,N_7639);
xnor U9690 (N_9690,N_7020,N_6936);
or U9691 (N_9691,N_7731,N_6754);
nor U9692 (N_9692,N_6514,N_6728);
nor U9693 (N_9693,N_6639,N_7245);
and U9694 (N_9694,N_7096,N_7242);
nor U9695 (N_9695,N_7867,N_7982);
nor U9696 (N_9696,N_7661,N_6754);
nor U9697 (N_9697,N_6829,N_7960);
and U9698 (N_9698,N_6125,N_6814);
nor U9699 (N_9699,N_7453,N_6518);
or U9700 (N_9700,N_7378,N_6570);
or U9701 (N_9701,N_6877,N_6480);
or U9702 (N_9702,N_6699,N_6289);
nor U9703 (N_9703,N_7097,N_7400);
nor U9704 (N_9704,N_6978,N_6549);
or U9705 (N_9705,N_6286,N_6897);
and U9706 (N_9706,N_7088,N_7561);
nand U9707 (N_9707,N_6035,N_7258);
xnor U9708 (N_9708,N_7671,N_6995);
and U9709 (N_9709,N_7242,N_6837);
nor U9710 (N_9710,N_7449,N_6921);
nor U9711 (N_9711,N_7629,N_6452);
or U9712 (N_9712,N_6245,N_6658);
or U9713 (N_9713,N_7134,N_6281);
and U9714 (N_9714,N_6010,N_7610);
nand U9715 (N_9715,N_6520,N_7129);
and U9716 (N_9716,N_7472,N_6474);
xor U9717 (N_9717,N_7287,N_7279);
nand U9718 (N_9718,N_6610,N_6351);
nand U9719 (N_9719,N_7892,N_6211);
nand U9720 (N_9720,N_7261,N_7865);
or U9721 (N_9721,N_6353,N_6566);
and U9722 (N_9722,N_7258,N_6395);
nand U9723 (N_9723,N_6222,N_7206);
or U9724 (N_9724,N_7092,N_7127);
or U9725 (N_9725,N_7290,N_7571);
or U9726 (N_9726,N_6833,N_6495);
and U9727 (N_9727,N_6814,N_7321);
nand U9728 (N_9728,N_7906,N_6250);
nand U9729 (N_9729,N_6512,N_7342);
nor U9730 (N_9730,N_6319,N_7280);
nor U9731 (N_9731,N_7498,N_6943);
xnor U9732 (N_9732,N_7183,N_6412);
and U9733 (N_9733,N_7099,N_6790);
xnor U9734 (N_9734,N_7364,N_7104);
xor U9735 (N_9735,N_7831,N_6406);
nand U9736 (N_9736,N_6012,N_7007);
or U9737 (N_9737,N_6093,N_7830);
or U9738 (N_9738,N_6945,N_7848);
nor U9739 (N_9739,N_6759,N_6598);
nand U9740 (N_9740,N_6206,N_7770);
nor U9741 (N_9741,N_6744,N_6340);
or U9742 (N_9742,N_6130,N_6855);
or U9743 (N_9743,N_7218,N_6894);
nand U9744 (N_9744,N_7179,N_6833);
or U9745 (N_9745,N_6002,N_7472);
xnor U9746 (N_9746,N_6789,N_7249);
nand U9747 (N_9747,N_7390,N_6887);
nor U9748 (N_9748,N_7986,N_7753);
or U9749 (N_9749,N_6977,N_7002);
nand U9750 (N_9750,N_7258,N_7375);
and U9751 (N_9751,N_7800,N_7188);
or U9752 (N_9752,N_6046,N_7721);
and U9753 (N_9753,N_7672,N_6921);
or U9754 (N_9754,N_6848,N_7511);
nand U9755 (N_9755,N_7857,N_7941);
nor U9756 (N_9756,N_6224,N_6157);
and U9757 (N_9757,N_7043,N_6399);
nor U9758 (N_9758,N_6906,N_6087);
and U9759 (N_9759,N_6795,N_7840);
nand U9760 (N_9760,N_6342,N_7660);
or U9761 (N_9761,N_6423,N_7427);
and U9762 (N_9762,N_7193,N_6927);
or U9763 (N_9763,N_6495,N_7407);
nor U9764 (N_9764,N_7153,N_7386);
nand U9765 (N_9765,N_6001,N_7456);
nand U9766 (N_9766,N_7774,N_6872);
nor U9767 (N_9767,N_7479,N_6726);
xnor U9768 (N_9768,N_7130,N_6696);
nor U9769 (N_9769,N_6136,N_6583);
and U9770 (N_9770,N_6086,N_6297);
nor U9771 (N_9771,N_6726,N_7316);
or U9772 (N_9772,N_7151,N_7830);
xor U9773 (N_9773,N_6952,N_6701);
and U9774 (N_9774,N_6898,N_6541);
and U9775 (N_9775,N_6292,N_7364);
and U9776 (N_9776,N_7339,N_7565);
nand U9777 (N_9777,N_7213,N_7972);
xor U9778 (N_9778,N_6721,N_7633);
or U9779 (N_9779,N_7488,N_7151);
or U9780 (N_9780,N_6990,N_6215);
nand U9781 (N_9781,N_6997,N_7231);
nor U9782 (N_9782,N_6444,N_7634);
or U9783 (N_9783,N_7670,N_7598);
and U9784 (N_9784,N_6172,N_7685);
nor U9785 (N_9785,N_6843,N_7039);
nand U9786 (N_9786,N_6471,N_7970);
and U9787 (N_9787,N_6432,N_7652);
or U9788 (N_9788,N_7884,N_7817);
or U9789 (N_9789,N_6563,N_7305);
nand U9790 (N_9790,N_7165,N_6846);
nand U9791 (N_9791,N_7166,N_7705);
nand U9792 (N_9792,N_6511,N_6961);
nand U9793 (N_9793,N_6126,N_7101);
nor U9794 (N_9794,N_6722,N_7421);
or U9795 (N_9795,N_7422,N_6391);
or U9796 (N_9796,N_6073,N_6619);
xnor U9797 (N_9797,N_6335,N_6323);
nor U9798 (N_9798,N_7886,N_6980);
and U9799 (N_9799,N_6182,N_7081);
and U9800 (N_9800,N_7108,N_7281);
or U9801 (N_9801,N_7441,N_6338);
nand U9802 (N_9802,N_7328,N_7867);
or U9803 (N_9803,N_7328,N_7290);
xnor U9804 (N_9804,N_7135,N_7172);
or U9805 (N_9805,N_6613,N_7201);
nand U9806 (N_9806,N_6372,N_7081);
nand U9807 (N_9807,N_6135,N_6872);
nand U9808 (N_9808,N_6266,N_6312);
and U9809 (N_9809,N_6733,N_6232);
or U9810 (N_9810,N_7283,N_6448);
and U9811 (N_9811,N_7919,N_6347);
or U9812 (N_9812,N_7092,N_6286);
or U9813 (N_9813,N_7496,N_7626);
nand U9814 (N_9814,N_6983,N_6665);
and U9815 (N_9815,N_7170,N_7310);
or U9816 (N_9816,N_6934,N_7079);
nor U9817 (N_9817,N_7534,N_7850);
and U9818 (N_9818,N_6893,N_7505);
or U9819 (N_9819,N_7781,N_6665);
xor U9820 (N_9820,N_6174,N_7246);
and U9821 (N_9821,N_6325,N_6286);
nor U9822 (N_9822,N_7313,N_6482);
nand U9823 (N_9823,N_6319,N_7901);
and U9824 (N_9824,N_6090,N_6887);
and U9825 (N_9825,N_7445,N_7929);
or U9826 (N_9826,N_6593,N_6546);
and U9827 (N_9827,N_6163,N_7752);
or U9828 (N_9828,N_7427,N_7281);
nand U9829 (N_9829,N_6377,N_7960);
nand U9830 (N_9830,N_6255,N_6163);
nor U9831 (N_9831,N_7854,N_6151);
nor U9832 (N_9832,N_7852,N_6752);
and U9833 (N_9833,N_6709,N_7133);
nor U9834 (N_9834,N_6227,N_6599);
nand U9835 (N_9835,N_6618,N_7505);
nand U9836 (N_9836,N_6182,N_7352);
xnor U9837 (N_9837,N_7283,N_6172);
nand U9838 (N_9838,N_7570,N_7420);
and U9839 (N_9839,N_7141,N_6677);
xor U9840 (N_9840,N_6979,N_7803);
or U9841 (N_9841,N_6886,N_6648);
nor U9842 (N_9842,N_7679,N_6153);
or U9843 (N_9843,N_7135,N_6746);
nor U9844 (N_9844,N_7578,N_6994);
nand U9845 (N_9845,N_7297,N_7103);
and U9846 (N_9846,N_6192,N_7211);
and U9847 (N_9847,N_7326,N_7319);
and U9848 (N_9848,N_7057,N_6052);
and U9849 (N_9849,N_6296,N_7048);
and U9850 (N_9850,N_6504,N_6934);
nand U9851 (N_9851,N_7797,N_7408);
nand U9852 (N_9852,N_7269,N_6371);
nand U9853 (N_9853,N_6935,N_7691);
nor U9854 (N_9854,N_6971,N_6977);
nor U9855 (N_9855,N_6151,N_7209);
xnor U9856 (N_9856,N_7694,N_7921);
nor U9857 (N_9857,N_6658,N_6079);
xnor U9858 (N_9858,N_6336,N_7265);
nor U9859 (N_9859,N_7566,N_7255);
nor U9860 (N_9860,N_6998,N_6599);
or U9861 (N_9861,N_7381,N_6920);
nand U9862 (N_9862,N_6319,N_6506);
nor U9863 (N_9863,N_7166,N_7524);
nor U9864 (N_9864,N_6256,N_6986);
and U9865 (N_9865,N_6121,N_7717);
and U9866 (N_9866,N_7267,N_6730);
nor U9867 (N_9867,N_7548,N_6924);
nor U9868 (N_9868,N_7990,N_6054);
and U9869 (N_9869,N_7696,N_6755);
nand U9870 (N_9870,N_7925,N_7475);
or U9871 (N_9871,N_7513,N_7037);
xor U9872 (N_9872,N_6854,N_6090);
nand U9873 (N_9873,N_7344,N_7743);
nand U9874 (N_9874,N_7544,N_6014);
or U9875 (N_9875,N_6897,N_6831);
nand U9876 (N_9876,N_7720,N_7977);
or U9877 (N_9877,N_7910,N_6651);
nor U9878 (N_9878,N_6782,N_6120);
nand U9879 (N_9879,N_6667,N_6956);
and U9880 (N_9880,N_6186,N_6459);
or U9881 (N_9881,N_6078,N_7401);
and U9882 (N_9882,N_6147,N_6494);
and U9883 (N_9883,N_7450,N_6722);
and U9884 (N_9884,N_7650,N_7532);
nor U9885 (N_9885,N_7975,N_7255);
xor U9886 (N_9886,N_6192,N_6328);
or U9887 (N_9887,N_6092,N_7497);
and U9888 (N_9888,N_6115,N_6920);
or U9889 (N_9889,N_6088,N_6101);
or U9890 (N_9890,N_6788,N_7921);
and U9891 (N_9891,N_6503,N_6923);
nand U9892 (N_9892,N_7533,N_7708);
nand U9893 (N_9893,N_7182,N_6314);
nand U9894 (N_9894,N_7138,N_7690);
xnor U9895 (N_9895,N_6609,N_7085);
nand U9896 (N_9896,N_7393,N_7476);
nor U9897 (N_9897,N_7824,N_6415);
xor U9898 (N_9898,N_6938,N_7555);
nand U9899 (N_9899,N_7112,N_6020);
or U9900 (N_9900,N_7783,N_6339);
and U9901 (N_9901,N_7767,N_7662);
nand U9902 (N_9902,N_6142,N_6548);
nor U9903 (N_9903,N_6875,N_7784);
or U9904 (N_9904,N_7828,N_6316);
or U9905 (N_9905,N_6002,N_7919);
or U9906 (N_9906,N_7098,N_6937);
nand U9907 (N_9907,N_6077,N_6487);
nand U9908 (N_9908,N_6708,N_7036);
or U9909 (N_9909,N_7905,N_7998);
nor U9910 (N_9910,N_7813,N_6278);
nand U9911 (N_9911,N_6426,N_6918);
or U9912 (N_9912,N_6489,N_7680);
or U9913 (N_9913,N_6033,N_7764);
and U9914 (N_9914,N_7991,N_7689);
xnor U9915 (N_9915,N_7171,N_6245);
or U9916 (N_9916,N_6795,N_6454);
or U9917 (N_9917,N_6459,N_7468);
nor U9918 (N_9918,N_6714,N_7298);
nand U9919 (N_9919,N_6540,N_6203);
nand U9920 (N_9920,N_7235,N_7911);
nand U9921 (N_9921,N_7201,N_7347);
or U9922 (N_9922,N_6093,N_7868);
or U9923 (N_9923,N_6372,N_7951);
and U9924 (N_9924,N_7612,N_6827);
or U9925 (N_9925,N_6214,N_7902);
xnor U9926 (N_9926,N_6619,N_6435);
nor U9927 (N_9927,N_7967,N_6632);
or U9928 (N_9928,N_7998,N_6069);
nand U9929 (N_9929,N_7844,N_6382);
nand U9930 (N_9930,N_7363,N_6727);
nand U9931 (N_9931,N_7181,N_7339);
or U9932 (N_9932,N_7058,N_7526);
or U9933 (N_9933,N_7561,N_6362);
or U9934 (N_9934,N_7071,N_7119);
or U9935 (N_9935,N_6604,N_6308);
nor U9936 (N_9936,N_6970,N_6185);
nor U9937 (N_9937,N_6899,N_7178);
nand U9938 (N_9938,N_6597,N_7575);
nand U9939 (N_9939,N_6105,N_6303);
or U9940 (N_9940,N_7135,N_6924);
nand U9941 (N_9941,N_7825,N_7283);
and U9942 (N_9942,N_7127,N_6700);
or U9943 (N_9943,N_6664,N_7081);
or U9944 (N_9944,N_6074,N_6231);
nand U9945 (N_9945,N_6391,N_6435);
and U9946 (N_9946,N_7268,N_6607);
nand U9947 (N_9947,N_7528,N_6597);
nand U9948 (N_9948,N_7702,N_6757);
or U9949 (N_9949,N_6745,N_6793);
and U9950 (N_9950,N_7676,N_7895);
nor U9951 (N_9951,N_6413,N_6769);
xnor U9952 (N_9952,N_6977,N_6138);
or U9953 (N_9953,N_6630,N_6282);
nand U9954 (N_9954,N_6607,N_7199);
or U9955 (N_9955,N_6089,N_7139);
nor U9956 (N_9956,N_6146,N_6477);
nand U9957 (N_9957,N_7827,N_6098);
nor U9958 (N_9958,N_6443,N_6842);
nand U9959 (N_9959,N_6038,N_6941);
or U9960 (N_9960,N_6132,N_7170);
and U9961 (N_9961,N_6668,N_6814);
nand U9962 (N_9962,N_7688,N_7061);
or U9963 (N_9963,N_6038,N_7685);
and U9964 (N_9964,N_7150,N_6652);
and U9965 (N_9965,N_6477,N_7197);
and U9966 (N_9966,N_6316,N_7857);
nor U9967 (N_9967,N_7259,N_7210);
xnor U9968 (N_9968,N_6297,N_6133);
nor U9969 (N_9969,N_7291,N_6628);
nand U9970 (N_9970,N_7267,N_7435);
and U9971 (N_9971,N_6220,N_7654);
xor U9972 (N_9972,N_7241,N_6719);
nand U9973 (N_9973,N_7719,N_7806);
or U9974 (N_9974,N_7893,N_7547);
and U9975 (N_9975,N_7773,N_7322);
or U9976 (N_9976,N_7901,N_7807);
xor U9977 (N_9977,N_6607,N_7126);
nor U9978 (N_9978,N_6772,N_7693);
nand U9979 (N_9979,N_6472,N_7809);
xor U9980 (N_9980,N_6377,N_7363);
and U9981 (N_9981,N_7099,N_7865);
nor U9982 (N_9982,N_7904,N_6157);
nand U9983 (N_9983,N_6862,N_6504);
nor U9984 (N_9984,N_7934,N_6537);
nor U9985 (N_9985,N_6611,N_6641);
nand U9986 (N_9986,N_7881,N_6185);
nor U9987 (N_9987,N_6933,N_6174);
and U9988 (N_9988,N_6162,N_6662);
nor U9989 (N_9989,N_7872,N_6143);
xor U9990 (N_9990,N_6066,N_7492);
and U9991 (N_9991,N_6735,N_7377);
and U9992 (N_9992,N_7243,N_7200);
xor U9993 (N_9993,N_7431,N_7717);
and U9994 (N_9994,N_6495,N_6043);
nor U9995 (N_9995,N_7277,N_6914);
nand U9996 (N_9996,N_7901,N_6006);
and U9997 (N_9997,N_6999,N_7086);
nand U9998 (N_9998,N_7453,N_6836);
or U9999 (N_9999,N_7396,N_6236);
nand UO_0 (O_0,N_8914,N_9385);
or UO_1 (O_1,N_8203,N_8920);
and UO_2 (O_2,N_9571,N_9956);
nand UO_3 (O_3,N_8083,N_9941);
and UO_4 (O_4,N_9328,N_8285);
and UO_5 (O_5,N_8307,N_9917);
and UO_6 (O_6,N_9340,N_9862);
xnor UO_7 (O_7,N_9009,N_8032);
xnor UO_8 (O_8,N_8792,N_8516);
or UO_9 (O_9,N_8949,N_9545);
or UO_10 (O_10,N_9275,N_9828);
or UO_11 (O_11,N_8765,N_9909);
or UO_12 (O_12,N_9918,N_8634);
nand UO_13 (O_13,N_9536,N_9310);
and UO_14 (O_14,N_8110,N_8863);
or UO_15 (O_15,N_9826,N_8311);
and UO_16 (O_16,N_9611,N_9282);
or UO_17 (O_17,N_8630,N_8539);
nor UO_18 (O_18,N_9914,N_9790);
or UO_19 (O_19,N_8713,N_9699);
and UO_20 (O_20,N_9147,N_8996);
or UO_21 (O_21,N_8173,N_8979);
or UO_22 (O_22,N_8118,N_8332);
and UO_23 (O_23,N_9840,N_8484);
and UO_24 (O_24,N_8229,N_9540);
or UO_25 (O_25,N_8559,N_9601);
nand UO_26 (O_26,N_9749,N_8432);
xor UO_27 (O_27,N_8702,N_9367);
xnor UO_28 (O_28,N_9621,N_9966);
xor UO_29 (O_29,N_9818,N_9911);
or UO_30 (O_30,N_8799,N_8771);
nand UO_31 (O_31,N_9085,N_9779);
and UO_32 (O_32,N_9153,N_8971);
nor UO_33 (O_33,N_8718,N_9078);
or UO_34 (O_34,N_8859,N_9423);
or UO_35 (O_35,N_8839,N_9746);
xor UO_36 (O_36,N_9199,N_8717);
and UO_37 (O_37,N_9365,N_9025);
or UO_38 (O_38,N_9172,N_8105);
nor UO_39 (O_39,N_9823,N_8942);
xnor UO_40 (O_40,N_8330,N_8073);
xnor UO_41 (O_41,N_8564,N_9894);
nand UO_42 (O_42,N_8127,N_9234);
nand UO_43 (O_43,N_8106,N_9727);
nor UO_44 (O_44,N_9656,N_9572);
xnor UO_45 (O_45,N_9748,N_9564);
xor UO_46 (O_46,N_8829,N_8759);
xnor UO_47 (O_47,N_9520,N_8838);
nor UO_48 (O_48,N_8807,N_9170);
nand UO_49 (O_49,N_8678,N_8235);
nor UO_50 (O_50,N_8514,N_9119);
and UO_51 (O_51,N_8376,N_8109);
and UO_52 (O_52,N_9235,N_9167);
nand UO_53 (O_53,N_8134,N_9675);
nor UO_54 (O_54,N_9408,N_8036);
nor UO_55 (O_55,N_9210,N_9121);
nor UO_56 (O_56,N_8269,N_8247);
nand UO_57 (O_57,N_8748,N_8305);
and UO_58 (O_58,N_9500,N_8511);
or UO_59 (O_59,N_8868,N_8703);
or UO_60 (O_60,N_9975,N_9178);
nor UO_61 (O_61,N_8457,N_8414);
nor UO_62 (O_62,N_8858,N_9904);
or UO_63 (O_63,N_8010,N_8842);
nand UO_64 (O_64,N_8260,N_9453);
xnor UO_65 (O_65,N_9583,N_9627);
nand UO_66 (O_66,N_8673,N_8007);
nand UO_67 (O_67,N_8591,N_8356);
xnor UO_68 (O_68,N_8348,N_8277);
nand UO_69 (O_69,N_9922,N_8796);
nor UO_70 (O_70,N_9796,N_9057);
and UO_71 (O_71,N_8560,N_8142);
and UO_72 (O_72,N_9496,N_8872);
and UO_73 (O_73,N_9303,N_8533);
nor UO_74 (O_74,N_9546,N_9593);
nand UO_75 (O_75,N_8855,N_8308);
nand UO_76 (O_76,N_8454,N_8263);
and UO_77 (O_77,N_8515,N_9512);
nand UO_78 (O_78,N_8629,N_8853);
nand UO_79 (O_79,N_9401,N_9008);
and UO_80 (O_80,N_9849,N_9100);
nand UO_81 (O_81,N_8207,N_9442);
xnor UO_82 (O_82,N_8760,N_9413);
nand UO_83 (O_83,N_8383,N_9197);
xor UO_84 (O_84,N_9420,N_8289);
nor UO_85 (O_85,N_9964,N_8068);
xor UO_86 (O_86,N_8174,N_9873);
nor UO_87 (O_87,N_8985,N_8567);
or UO_88 (O_88,N_9785,N_9291);
nor UO_89 (O_89,N_8278,N_9763);
nand UO_90 (O_90,N_8508,N_9990);
nor UO_91 (O_91,N_8584,N_8562);
or UO_92 (O_92,N_8120,N_8738);
nor UO_93 (O_93,N_8077,N_9380);
or UO_94 (O_94,N_8500,N_9800);
nand UO_95 (O_95,N_8350,N_9148);
and UO_96 (O_96,N_8531,N_8322);
or UO_97 (O_97,N_9359,N_9700);
nor UO_98 (O_98,N_9897,N_8825);
and UO_99 (O_99,N_8343,N_8845);
nor UO_100 (O_100,N_8181,N_9971);
and UO_101 (O_101,N_9266,N_9216);
nor UO_102 (O_102,N_9523,N_8455);
and UO_103 (O_103,N_8947,N_9010);
nand UO_104 (O_104,N_9864,N_8076);
or UO_105 (O_105,N_9932,N_9969);
nor UO_106 (O_106,N_8766,N_9226);
nand UO_107 (O_107,N_9351,N_9726);
or UO_108 (O_108,N_9537,N_9510);
xor UO_109 (O_109,N_9631,N_8873);
and UO_110 (O_110,N_8312,N_8418);
nor UO_111 (O_111,N_9999,N_8100);
nor UO_112 (O_112,N_9610,N_8783);
nand UO_113 (O_113,N_9947,N_9400);
or UO_114 (O_114,N_9690,N_8085);
nor UO_115 (O_115,N_9972,N_9138);
and UO_116 (O_116,N_9033,N_8283);
nor UO_117 (O_117,N_8900,N_8304);
nand UO_118 (O_118,N_9125,N_8927);
xnor UO_119 (O_119,N_9005,N_8980);
xor UO_120 (O_120,N_8395,N_8719);
xnor UO_121 (O_121,N_9946,N_9083);
nor UO_122 (O_122,N_9110,N_8575);
xor UO_123 (O_123,N_8546,N_9084);
nand UO_124 (O_124,N_9669,N_8023);
and UO_125 (O_125,N_9052,N_9437);
and UO_126 (O_126,N_9741,N_9866);
nor UO_127 (O_127,N_8059,N_8574);
nor UO_128 (O_128,N_8427,N_8102);
and UO_129 (O_129,N_9835,N_9115);
xor UO_130 (O_130,N_9075,N_8213);
nand UO_131 (O_131,N_9534,N_9375);
xor UO_132 (O_132,N_8195,N_9880);
nand UO_133 (O_133,N_8468,N_8699);
nor UO_134 (O_134,N_9103,N_9089);
or UO_135 (O_135,N_9740,N_8282);
and UO_136 (O_136,N_9087,N_9668);
and UO_137 (O_137,N_9633,N_9097);
nor UO_138 (O_138,N_9134,N_9939);
nor UO_139 (O_139,N_9223,N_9146);
nor UO_140 (O_140,N_9230,N_8530);
or UO_141 (O_141,N_8870,N_8126);
and UO_142 (O_142,N_9092,N_9637);
and UO_143 (O_143,N_9739,N_9541);
nor UO_144 (O_144,N_9166,N_9012);
or UO_145 (O_145,N_9577,N_9244);
nor UO_146 (O_146,N_8103,N_8415);
nand UO_147 (O_147,N_9182,N_8162);
and UO_148 (O_148,N_8815,N_9935);
nand UO_149 (O_149,N_8180,N_8769);
xnor UO_150 (O_150,N_9908,N_9614);
nand UO_151 (O_151,N_9639,N_9979);
or UO_152 (O_152,N_8513,N_8258);
and UO_153 (O_153,N_9618,N_8431);
and UO_154 (O_154,N_8294,N_8074);
nand UO_155 (O_155,N_8166,N_9588);
nand UO_156 (O_156,N_8501,N_9492);
nor UO_157 (O_157,N_9186,N_9483);
or UO_158 (O_158,N_9308,N_9987);
nand UO_159 (O_159,N_9058,N_9901);
and UO_160 (O_160,N_8000,N_8885);
xnor UO_161 (O_161,N_9837,N_9836);
nand UO_162 (O_162,N_8217,N_9776);
nand UO_163 (O_163,N_9550,N_8117);
nand UO_164 (O_164,N_9416,N_8646);
nand UO_165 (O_165,N_9160,N_9710);
or UO_166 (O_166,N_8071,N_8236);
nand UO_167 (O_167,N_9176,N_9686);
and UO_168 (O_168,N_8152,N_8208);
or UO_169 (O_169,N_8913,N_9558);
xnor UO_170 (O_170,N_9723,N_8688);
or UO_171 (O_171,N_8416,N_8877);
nand UO_172 (O_172,N_9991,N_9355);
and UO_173 (O_173,N_9219,N_8136);
or UO_174 (O_174,N_8806,N_8458);
nor UO_175 (O_175,N_8082,N_9339);
xnor UO_176 (O_176,N_9813,N_8800);
xor UO_177 (O_177,N_9645,N_9128);
and UO_178 (O_178,N_8795,N_8970);
nor UO_179 (O_179,N_9286,N_8430);
nand UO_180 (O_180,N_8653,N_8472);
xor UO_181 (O_181,N_9232,N_8978);
nand UO_182 (O_182,N_9955,N_9730);
and UO_183 (O_183,N_9592,N_8682);
and UO_184 (O_184,N_8478,N_9325);
and UO_185 (O_185,N_8302,N_8946);
nand UO_186 (O_186,N_8550,N_8818);
or UO_187 (O_187,N_8224,N_8854);
or UO_188 (O_188,N_9662,N_9295);
and UO_189 (O_189,N_9891,N_8619);
nand UO_190 (O_190,N_9860,N_9579);
or UO_191 (O_191,N_8826,N_9515);
or UO_192 (O_192,N_9352,N_9181);
nand UO_193 (O_193,N_9910,N_8892);
nand UO_194 (O_194,N_8517,N_9889);
xnor UO_195 (O_195,N_8518,N_8325);
nand UO_196 (O_196,N_9762,N_9566);
or UO_197 (O_197,N_8320,N_9456);
nand UO_198 (O_198,N_8975,N_8009);
nand UO_199 (O_199,N_8318,N_8249);
or UO_200 (O_200,N_9916,N_9392);
nand UO_201 (O_201,N_8604,N_8631);
nand UO_202 (O_202,N_9111,N_8747);
nand UO_203 (O_203,N_9373,N_9493);
and UO_204 (O_204,N_9229,N_8151);
or UO_205 (O_205,N_8756,N_8264);
and UO_206 (O_206,N_9342,N_9415);
or UO_207 (O_207,N_8221,N_9634);
and UO_208 (O_208,N_8145,N_8623);
nor UO_209 (O_209,N_9678,N_9950);
or UO_210 (O_210,N_8811,N_9516);
or UO_211 (O_211,N_9247,N_8060);
and UO_212 (O_212,N_8489,N_8883);
nand UO_213 (O_213,N_9466,N_9474);
nand UO_214 (O_214,N_9926,N_9193);
and UO_215 (O_215,N_9538,N_8390);
xor UO_216 (O_216,N_8610,N_8986);
or UO_217 (O_217,N_8912,N_8960);
nor UO_218 (O_218,N_8189,N_8690);
or UO_219 (O_219,N_8216,N_9054);
nand UO_220 (O_220,N_9348,N_9925);
nand UO_221 (O_221,N_9414,N_8835);
and UO_222 (O_222,N_9035,N_8701);
nand UO_223 (O_223,N_9585,N_8443);
or UO_224 (O_224,N_9602,N_8042);
xor UO_225 (O_225,N_9022,N_8202);
xor UO_226 (O_226,N_9794,N_8245);
or UO_227 (O_227,N_9141,N_8373);
nor UO_228 (O_228,N_8505,N_9698);
xnor UO_229 (O_229,N_8115,N_9881);
nor UO_230 (O_230,N_8788,N_9313);
or UO_231 (O_231,N_8879,N_9872);
or UO_232 (O_232,N_8869,N_9156);
and UO_233 (O_233,N_8659,N_9750);
xnor UO_234 (O_234,N_9228,N_9019);
or UO_235 (O_235,N_8676,N_9695);
nand UO_236 (O_236,N_8793,N_9347);
xor UO_237 (O_237,N_9576,N_8639);
nor UO_238 (O_238,N_8754,N_9573);
xnor UO_239 (O_239,N_9036,N_8069);
nor UO_240 (O_240,N_8306,N_9007);
and UO_241 (O_241,N_8041,N_9920);
nand UO_242 (O_242,N_9647,N_8219);
and UO_243 (O_243,N_8303,N_8840);
nor UO_244 (O_244,N_8061,N_8680);
xnor UO_245 (O_245,N_9820,N_8874);
nand UO_246 (O_246,N_9208,N_8648);
or UO_247 (O_247,N_9774,N_9554);
nor UO_248 (O_248,N_8093,N_8926);
nor UO_249 (O_249,N_8961,N_8051);
and UO_250 (O_250,N_8901,N_8124);
nor UO_251 (O_251,N_9238,N_9814);
and UO_252 (O_252,N_9088,N_9213);
or UO_253 (O_253,N_8534,N_9665);
nor UO_254 (O_254,N_9283,N_8169);
nor UO_255 (O_255,N_8273,N_9569);
or UO_256 (O_256,N_9321,N_8081);
or UO_257 (O_257,N_9180,N_9905);
and UO_258 (O_258,N_9398,N_9305);
or UO_259 (O_259,N_8310,N_9042);
nor UO_260 (O_260,N_9105,N_9490);
or UO_261 (O_261,N_9811,N_9452);
or UO_262 (O_262,N_9067,N_9432);
nand UO_263 (O_263,N_9998,N_8599);
and UO_264 (O_264,N_9133,N_8052);
nand UO_265 (O_265,N_8324,N_8889);
xor UO_266 (O_266,N_9073,N_8449);
and UO_267 (O_267,N_8474,N_9892);
xor UO_268 (O_268,N_8095,N_8732);
or UO_269 (O_269,N_9858,N_8576);
nor UO_270 (O_270,N_8723,N_8377);
nor UO_271 (O_271,N_9016,N_9039);
xnor UO_272 (O_272,N_8936,N_9720);
nand UO_273 (O_273,N_9158,N_8686);
nand UO_274 (O_274,N_9460,N_9855);
and UO_275 (O_275,N_9402,N_8351);
nor UO_276 (O_276,N_8675,N_9861);
nor UO_277 (O_277,N_9430,N_8342);
nand UO_278 (O_278,N_8580,N_9221);
and UO_279 (O_279,N_9000,N_9962);
xnor UO_280 (O_280,N_9680,N_9847);
and UO_281 (O_281,N_9963,N_8265);
nor UO_282 (O_282,N_9692,N_8241);
and UO_283 (O_283,N_9081,N_8186);
nor UO_284 (O_284,N_8837,N_8594);
xnor UO_285 (O_285,N_8347,N_9854);
xor UO_286 (O_286,N_9069,N_8327);
or UO_287 (O_287,N_9747,N_9358);
nor UO_288 (O_288,N_9808,N_9834);
nand UO_289 (O_289,N_8770,N_8802);
and UO_290 (O_290,N_8053,N_9586);
nor UO_291 (O_291,N_8445,N_9249);
nand UO_292 (O_292,N_8677,N_9131);
and UO_293 (O_293,N_8098,N_8140);
nand UO_294 (O_294,N_8649,N_8029);
and UO_295 (O_295,N_9046,N_9670);
and UO_296 (O_296,N_9696,N_8024);
nor UO_297 (O_297,N_9612,N_9912);
or UO_298 (O_298,N_9688,N_9745);
and UO_299 (O_299,N_8391,N_8644);
nor UO_300 (O_300,N_9594,N_8025);
nand UO_301 (O_301,N_9332,N_8496);
nand UO_302 (O_302,N_9140,N_9377);
and UO_303 (O_303,N_9552,N_9449);
nand UO_304 (O_304,N_9296,N_9494);
and UO_305 (O_305,N_8155,N_8587);
nand UO_306 (O_306,N_8133,N_8720);
nor UO_307 (O_307,N_8557,N_9288);
or UO_308 (O_308,N_9038,N_8481);
or UO_309 (O_309,N_9381,N_8436);
or UO_310 (O_310,N_8158,N_9378);
xor UO_311 (O_311,N_9653,N_9868);
or UO_312 (O_312,N_9190,N_9252);
or UO_313 (O_313,N_8101,N_8441);
nor UO_314 (O_314,N_9772,N_8141);
nor UO_315 (O_315,N_9798,N_9336);
and UO_316 (O_316,N_8708,N_9884);
nand UO_317 (O_317,N_9495,N_9344);
and UO_318 (O_318,N_8692,N_9031);
nand UO_319 (O_319,N_8593,N_8640);
xnor UO_320 (O_320,N_9856,N_8767);
nor UO_321 (O_321,N_9488,N_8156);
nor UO_322 (O_322,N_9240,N_9931);
xnor UO_323 (O_323,N_8323,N_9927);
and UO_324 (O_324,N_9980,N_8192);
or UO_325 (O_325,N_8170,N_8937);
nand UO_326 (O_326,N_8924,N_9061);
or UO_327 (O_327,N_9082,N_8761);
or UO_328 (O_328,N_8954,N_9357);
and UO_329 (O_329,N_9783,N_9650);
nor UO_330 (O_330,N_9239,N_8856);
nand UO_331 (O_331,N_8092,N_8499);
nand UO_332 (O_332,N_8242,N_9721);
and UO_333 (O_333,N_8997,N_9425);
nand UO_334 (O_334,N_9731,N_8482);
nand UO_335 (O_335,N_9646,N_8435);
or UO_336 (O_336,N_9844,N_8437);
nor UO_337 (O_337,N_8178,N_8932);
nand UO_338 (O_338,N_8477,N_8122);
or UO_339 (O_339,N_8762,N_8749);
and UO_340 (O_340,N_9273,N_9735);
or UO_341 (O_341,N_8321,N_8137);
or UO_342 (O_342,N_9399,N_9037);
nand UO_343 (O_343,N_9603,N_9852);
nor UO_344 (O_344,N_9982,N_8262);
nor UO_345 (O_345,N_8319,N_8951);
and UO_346 (O_346,N_8538,N_8378);
nor UO_347 (O_347,N_8357,N_8758);
and UO_348 (O_348,N_9326,N_8113);
nand UO_349 (O_349,N_8697,N_9177);
or UO_350 (O_350,N_8016,N_8707);
and UO_351 (O_351,N_8958,N_8775);
and UO_352 (O_352,N_8583,N_9625);
xnor UO_353 (O_353,N_8058,N_9441);
or UO_354 (O_354,N_9784,N_9214);
and UO_355 (O_355,N_9382,N_8934);
nand UO_356 (O_356,N_9489,N_9829);
or UO_357 (O_357,N_8326,N_9719);
xnor UO_358 (O_358,N_8116,N_9301);
xor UO_359 (O_359,N_9372,N_9959);
nand UO_360 (O_360,N_8279,N_9744);
or UO_361 (O_361,N_8729,N_8218);
nor UO_362 (O_362,N_8969,N_9985);
nand UO_363 (O_363,N_9311,N_9815);
and UO_364 (O_364,N_9504,N_8066);
nand UO_365 (O_365,N_9346,N_8309);
and UO_366 (O_366,N_8974,N_9623);
nor UO_367 (O_367,N_9189,N_8933);
or UO_368 (O_368,N_8714,N_9370);
nand UO_369 (O_369,N_8157,N_9693);
nor UO_370 (O_370,N_8039,N_8067);
and UO_371 (O_371,N_8884,N_9683);
and UO_372 (O_372,N_8750,N_9629);
or UO_373 (O_373,N_8784,N_8737);
or UO_374 (O_374,N_9595,N_8618);
nor UO_375 (O_375,N_9965,N_8847);
nand UO_376 (O_376,N_8510,N_9529);
or UO_377 (O_377,N_9954,N_8080);
nor UO_378 (O_378,N_8004,N_9345);
or UO_379 (O_379,N_9014,N_9063);
nor UO_380 (O_380,N_9002,N_8329);
nand UO_381 (O_381,N_8234,N_8844);
or UO_382 (O_382,N_9198,N_9830);
nand UO_383 (O_383,N_9885,N_8401);
and UO_384 (O_384,N_9976,N_9044);
xor UO_385 (O_385,N_8816,N_8355);
xnor UO_386 (O_386,N_9475,N_9337);
nand UO_387 (O_387,N_8365,N_9655);
xnor UO_388 (O_388,N_8429,N_9101);
and UO_389 (O_389,N_9426,N_9547);
and UO_390 (O_390,N_8923,N_8388);
and UO_391 (O_391,N_9202,N_8915);
nor UO_392 (O_392,N_8394,N_8194);
nand UO_393 (O_393,N_8470,N_8782);
nor UO_394 (O_394,N_8596,N_9997);
nand UO_395 (O_395,N_8566,N_9155);
nand UO_396 (O_396,N_9833,N_8090);
or UO_397 (O_397,N_9324,N_8063);
xnor UO_398 (O_398,N_9258,N_9404);
or UO_399 (O_399,N_8968,N_9702);
xnor UO_400 (O_400,N_8346,N_9395);
and UO_401 (O_401,N_8405,N_9685);
nand UO_402 (O_402,N_8521,N_9694);
and UO_403 (O_403,N_9095,N_9777);
nor UO_404 (O_404,N_9468,N_9224);
nor UO_405 (O_405,N_8740,N_9429);
or UO_406 (O_406,N_8595,N_9331);
and UO_407 (O_407,N_8817,N_8172);
nor UO_408 (O_408,N_9587,N_9179);
or UO_409 (O_409,N_8848,N_9606);
xnor UO_410 (O_410,N_9928,N_9754);
xor UO_411 (O_411,N_8404,N_8403);
or UO_412 (O_412,N_9883,N_9396);
or UO_413 (O_413,N_9899,N_8406);
and UO_414 (O_414,N_9354,N_8700);
nor UO_415 (O_415,N_8425,N_9942);
nand UO_416 (O_416,N_8111,N_8987);
nand UO_417 (O_417,N_8633,N_9098);
and UO_418 (O_418,N_8727,N_9455);
nand UO_419 (O_419,N_8150,N_9072);
and UO_420 (O_420,N_8875,N_9608);
nor UO_421 (O_421,N_8671,N_8803);
and UO_422 (O_422,N_9578,N_9317);
and UO_423 (O_423,N_8331,N_9992);
or UO_424 (O_424,N_9323,N_8198);
nor UO_425 (O_425,N_8182,N_9304);
or UO_426 (O_426,N_9562,N_9314);
or UO_427 (O_427,N_9013,N_8904);
xnor UO_428 (O_428,N_9508,N_9557);
nor UO_429 (O_429,N_8220,N_9701);
and UO_430 (O_430,N_8607,N_8495);
or UO_431 (O_431,N_9284,N_8905);
xor UO_432 (O_432,N_8433,N_8465);
nor UO_433 (O_433,N_9551,N_9435);
nor UO_434 (O_434,N_9677,N_9050);
nand UO_435 (O_435,N_9436,N_9890);
nor UO_436 (O_436,N_9531,N_8684);
xnor UO_437 (O_437,N_8300,N_8371);
and UO_438 (O_438,N_9203,N_9553);
nand UO_439 (O_439,N_8232,N_8919);
nand UO_440 (O_440,N_8337,N_8888);
and UO_441 (O_441,N_8962,N_8246);
nand UO_442 (O_442,N_9851,N_9724);
or UO_443 (O_443,N_8231,N_8999);
or UO_444 (O_444,N_9556,N_8132);
nand UO_445 (O_445,N_8121,N_9903);
nand UO_446 (O_446,N_9433,N_9383);
nor UO_447 (O_447,N_8898,N_8773);
nor UO_448 (O_448,N_8114,N_9267);
nor UO_449 (O_449,N_9064,N_8479);
nor UO_450 (O_450,N_9674,N_8196);
or UO_451 (O_451,N_9930,N_8267);
and UO_452 (O_452,N_9018,N_9671);
nor UO_453 (O_453,N_8948,N_9419);
nand UO_454 (O_454,N_9561,N_9376);
nor UO_455 (O_455,N_8520,N_8392);
xor UO_456 (O_456,N_8467,N_8661);
xor UO_457 (O_457,N_8579,N_9498);
nor UO_458 (O_458,N_8558,N_9497);
nor UO_459 (O_459,N_8483,N_9502);
and UO_460 (O_460,N_8168,N_9349);
nor UO_461 (O_461,N_8230,N_9207);
nor UO_462 (O_462,N_8268,N_8938);
nor UO_463 (O_463,N_9001,N_8598);
nand UO_464 (O_464,N_9666,N_8573);
or UO_465 (O_465,N_9589,N_8089);
or UO_466 (O_466,N_8037,N_9302);
nor UO_467 (O_467,N_9440,N_8537);
and UO_468 (O_468,N_9791,N_9473);
and UO_469 (O_469,N_9405,N_9902);
and UO_470 (O_470,N_8447,N_9096);
or UO_471 (O_471,N_8253,N_8943);
nand UO_472 (O_472,N_8624,N_9041);
nand UO_473 (O_473,N_9026,N_9454);
or UO_474 (O_474,N_8358,N_9628);
nor UO_475 (O_475,N_8953,N_9126);
nor UO_476 (O_476,N_8493,N_9122);
nor UO_477 (O_477,N_9533,N_9341);
or UO_478 (O_478,N_9476,N_9477);
and UO_479 (O_479,N_9684,N_8989);
nor UO_480 (O_480,N_9737,N_8315);
xnor UO_481 (O_481,N_9951,N_9162);
and UO_482 (O_482,N_8745,N_9271);
nor UO_483 (O_483,N_8223,N_8698);
and UO_484 (O_484,N_9049,N_8614);
nand UO_485 (O_485,N_9759,N_8048);
or UO_486 (O_486,N_9004,N_8498);
and UO_487 (O_487,N_8001,N_9149);
nand UO_488 (O_488,N_9713,N_8991);
and UO_489 (O_489,N_8201,N_9280);
and UO_490 (O_490,N_8663,N_8349);
nand UO_491 (O_491,N_8581,N_9770);
nand UO_492 (O_492,N_9599,N_9068);
or UO_493 (O_493,N_8929,N_9509);
and UO_494 (O_494,N_8291,N_9626);
or UO_495 (O_495,N_9307,N_8448);
nor UO_496 (O_496,N_9517,N_8993);
nor UO_497 (O_497,N_8086,N_8733);
or UO_498 (O_498,N_8794,N_8902);
or UO_499 (O_499,N_9824,N_8899);
nand UO_500 (O_500,N_8779,N_9742);
nand UO_501 (O_501,N_8981,N_9661);
and UO_502 (O_502,N_8709,N_8535);
nor UO_503 (O_503,N_8027,N_9279);
and UO_504 (O_504,N_9270,N_8728);
nor UO_505 (O_505,N_8528,N_8380);
nand UO_506 (O_506,N_9781,N_8393);
or UO_507 (O_507,N_8239,N_8385);
nand UO_508 (O_508,N_8353,N_9913);
or UO_509 (O_509,N_9472,N_9114);
nand UO_510 (O_510,N_8731,N_9716);
and UO_511 (O_511,N_9024,N_9617);
and UO_512 (O_512,N_8809,N_9771);
nor UO_513 (O_513,N_9034,N_8200);
and UO_514 (O_514,N_8301,N_8407);
or UO_515 (O_515,N_9544,N_8568);
or UO_516 (O_516,N_8917,N_9151);
nand UO_517 (O_517,N_8621,N_9256);
or UO_518 (O_518,N_8589,N_8939);
and UO_519 (O_519,N_8212,N_8442);
and UO_520 (O_520,N_9079,N_8363);
xnor UO_521 (O_521,N_9921,N_9056);
nor UO_522 (O_522,N_9108,N_8062);
and UO_523 (O_523,N_8928,N_8018);
and UO_524 (O_524,N_9086,N_8079);
or UO_525 (O_525,N_8638,N_9760);
and UO_526 (O_526,N_9871,N_8609);
and UO_527 (O_527,N_8983,N_9896);
nor UO_528 (O_528,N_8977,N_9195);
and UO_529 (O_529,N_8108,N_9215);
or UO_530 (O_530,N_8655,N_8078);
and UO_531 (O_531,N_9259,N_8368);
nand UO_532 (O_532,N_8420,N_8255);
or UO_533 (O_533,N_8908,N_8012);
and UO_534 (O_534,N_8070,N_8608);
and UO_535 (O_535,N_8288,N_9832);
nor UO_536 (O_536,N_8422,N_8451);
or UO_537 (O_537,N_8184,N_9335);
or UO_538 (O_538,N_8772,N_8635);
xor UO_539 (O_539,N_9161,N_9040);
nor UO_540 (O_540,N_9261,N_9292);
nor UO_541 (O_541,N_8164,N_8972);
and UO_542 (O_542,N_9996,N_9722);
nand UO_543 (O_543,N_9597,N_9379);
nand UO_544 (O_544,N_8473,N_9697);
and UO_545 (O_545,N_8641,N_9870);
nor UO_546 (O_546,N_8605,N_9480);
nand UO_547 (O_547,N_9264,N_9333);
nor UO_548 (O_548,N_9387,N_9241);
nor UO_549 (O_549,N_8616,N_9200);
nor UO_550 (O_550,N_9518,N_8492);
or UO_551 (O_551,N_8410,N_9995);
nand UO_552 (O_552,N_9519,N_8428);
nand UO_553 (O_553,N_8742,N_9091);
and UO_554 (O_554,N_8250,N_9150);
and UO_555 (O_555,N_9769,N_8715);
or UO_556 (O_556,N_9875,N_8705);
and UO_557 (O_557,N_9080,N_8480);
nor UO_558 (O_558,N_8862,N_9521);
and UO_559 (O_559,N_9027,N_9755);
xnor UO_560 (O_560,N_8833,N_8755);
or UO_561 (O_561,N_8597,N_9809);
or UO_562 (O_562,N_8440,N_8274);
and UO_563 (O_563,N_8335,N_9938);
or UO_564 (O_564,N_8757,N_8918);
and UO_565 (O_565,N_8555,N_8317);
nand UO_566 (O_566,N_9023,N_9306);
or UO_567 (O_567,N_8672,N_9812);
xor UO_568 (O_568,N_8225,N_8955);
or UO_569 (O_569,N_8167,N_8820);
and UO_570 (O_570,N_8466,N_8841);
xor UO_571 (O_571,N_8668,N_8044);
or UO_572 (O_572,N_9886,N_8781);
nand UO_573 (O_573,N_8871,N_8050);
or UO_574 (O_574,N_9974,N_9243);
or UO_575 (O_575,N_9143,N_9163);
and UO_576 (O_576,N_8135,N_9217);
nor UO_577 (O_577,N_9015,N_9940);
and UO_578 (O_578,N_9482,N_9582);
and UO_579 (O_579,N_8603,N_8459);
and UO_580 (O_580,N_8571,N_9462);
nand UO_581 (O_581,N_8774,N_8965);
nor UO_582 (O_582,N_9756,N_8963);
and UO_583 (O_583,N_9276,N_8452);
and UO_584 (O_584,N_8882,N_9184);
and UO_585 (O_585,N_9192,N_9285);
nand UO_586 (O_586,N_9257,N_9906);
nand UO_587 (O_587,N_9907,N_9074);
nand UO_588 (O_588,N_8990,N_8411);
and UO_589 (O_589,N_9211,N_9469);
nor UO_590 (O_590,N_8810,N_9438);
nand UO_591 (O_591,N_8897,N_8423);
or UO_592 (O_592,N_8413,N_8190);
xor UO_593 (O_593,N_9654,N_8128);
or UO_594 (O_594,N_8147,N_9943);
nand UO_595 (O_595,N_8645,N_9175);
and UO_596 (O_596,N_9804,N_8054);
and UO_597 (O_597,N_9407,N_8881);
and UO_598 (O_598,N_9657,N_9260);
and UO_599 (O_599,N_8504,N_8785);
or UO_600 (O_600,N_9173,N_9715);
nand UO_601 (O_601,N_9363,N_8959);
nand UO_602 (O_602,N_9459,N_9708);
and UO_603 (O_603,N_8525,N_8205);
xnor UO_604 (O_604,N_8464,N_8011);
nor UO_605 (O_605,N_9973,N_9076);
or UO_606 (O_606,N_9581,N_9269);
nand UO_607 (O_607,N_9825,N_9253);
and UO_608 (O_608,N_9277,N_9491);
and UO_609 (O_609,N_9062,N_9879);
nor UO_610 (O_610,N_9659,N_9869);
nand UO_611 (O_611,N_9481,N_9788);
nand UO_612 (O_612,N_8726,N_8426);
nand UO_613 (O_613,N_9417,N_9113);
and UO_614 (O_614,N_9689,N_9590);
or UO_615 (O_615,N_8746,N_9268);
and UO_616 (O_616,N_9511,N_9765);
or UO_617 (O_617,N_8396,N_8204);
or UO_618 (O_618,N_9463,N_8849);
or UO_619 (O_619,N_9077,N_8950);
nor UO_620 (O_620,N_9450,N_8382);
or UO_621 (O_621,N_9525,N_9984);
or UO_622 (O_622,N_9548,N_8276);
nor UO_623 (O_623,N_9549,N_8570);
nand UO_624 (O_624,N_8542,N_9532);
or UO_625 (O_625,N_8896,N_9642);
and UO_626 (O_626,N_9712,N_8828);
and UO_627 (O_627,N_9753,N_8976);
and UO_628 (O_628,N_8462,N_9989);
and UO_629 (O_629,N_9393,N_8088);
nor UO_630 (O_630,N_8439,N_9949);
and UO_631 (O_631,N_9444,N_8161);
nor UO_632 (O_632,N_8836,N_9802);
nand UO_633 (O_633,N_9418,N_8056);
or UO_634 (O_634,N_9318,N_8034);
nand UO_635 (O_635,N_9948,N_8043);
nand UO_636 (O_636,N_8503,N_9672);
nor UO_637 (O_637,N_8711,N_9388);
xor UO_638 (O_638,N_9316,N_8921);
and UO_639 (O_639,N_9961,N_8287);
and UO_640 (O_640,N_9863,N_8359);
and UO_641 (O_641,N_8861,N_8612);
nor UO_642 (O_642,N_9793,N_9028);
nand UO_643 (O_643,N_8724,N_8014);
and UO_644 (O_644,N_8475,N_8446);
nand UO_645 (O_645,N_9743,N_9157);
and UO_646 (O_646,N_8549,N_8316);
nand UO_647 (O_647,N_9673,N_8057);
xor UO_648 (O_648,N_9923,N_8486);
nor UO_649 (O_649,N_9778,N_9312);
or UO_650 (O_650,N_9977,N_8149);
or UO_651 (O_651,N_8177,N_8165);
nand UO_652 (O_652,N_8075,N_8627);
and UO_653 (O_653,N_9539,N_9250);
or UO_654 (O_654,N_9055,N_8033);
xnor UO_655 (O_655,N_8421,N_9527);
xnor UO_656 (O_656,N_8679,N_8290);
and UO_657 (O_657,N_9501,N_8957);
or UO_658 (O_658,N_9386,N_8214);
nor UO_659 (O_659,N_9209,N_8130);
nor UO_660 (O_660,N_9667,N_8613);
nor UO_661 (O_661,N_8490,N_8891);
or UO_662 (O_662,N_8911,N_9758);
nand UO_663 (O_663,N_8536,N_9865);
and UO_664 (O_664,N_8072,N_8988);
nor UO_665 (O_665,N_8669,N_9274);
nor UO_666 (O_666,N_9406,N_8491);
and UO_667 (O_667,N_8509,N_9714);
nor UO_668 (O_668,N_9290,N_8297);
and UO_669 (O_669,N_9479,N_8922);
or UO_670 (O_670,N_8751,N_9664);
or UO_671 (O_671,N_9848,N_8233);
and UO_672 (O_672,N_8362,N_9029);
nor UO_673 (O_673,N_8721,N_9225);
nand UO_674 (O_674,N_8753,N_8444);
and UO_675 (O_675,N_8916,N_9448);
xor UO_676 (O_676,N_9736,N_8615);
and UO_677 (O_677,N_8524,N_8777);
nor UO_678 (O_678,N_8744,N_8281);
or UO_679 (O_679,N_8456,N_9643);
and UO_680 (O_680,N_9152,N_8064);
nand UO_681 (O_681,N_8660,N_8360);
and UO_682 (O_682,N_9236,N_8197);
nand UO_683 (O_683,N_9773,N_9728);
and UO_684 (O_684,N_8685,N_8266);
nand UO_685 (O_685,N_8890,N_8554);
or UO_686 (O_686,N_8188,N_8832);
nand UO_687 (O_687,N_8995,N_9428);
or UO_688 (O_688,N_8665,N_9127);
and UO_689 (O_689,N_8693,N_8419);
nand UO_690 (O_690,N_8552,N_9371);
and UO_691 (O_691,N_9570,N_9185);
and UO_692 (O_692,N_9006,N_8910);
and UO_693 (O_693,N_9281,N_8827);
xnor UO_694 (O_694,N_8112,N_8084);
nand UO_695 (O_695,N_9850,N_9709);
or UO_696 (O_696,N_9584,N_9220);
or UO_697 (O_697,N_8657,N_9568);
or UO_698 (O_698,N_9652,N_9485);
or UO_699 (O_699,N_9424,N_8314);
nor UO_700 (O_700,N_9051,N_9251);
and UO_701 (O_701,N_8632,N_9445);
nor UO_702 (O_702,N_9846,N_8647);
or UO_703 (O_703,N_8211,N_8187);
nor UO_704 (O_704,N_9565,N_8526);
and UO_705 (O_705,N_9648,N_9604);
or UO_706 (O_706,N_8497,N_8650);
or UO_707 (O_707,N_9364,N_9389);
xor UO_708 (O_708,N_8543,N_9766);
and UO_709 (O_709,N_9443,N_9090);
nand UO_710 (O_710,N_8780,N_8944);
nor UO_711 (O_711,N_8654,N_9116);
or UO_712 (O_712,N_9409,N_9607);
nor UO_713 (O_713,N_9789,N_8725);
and UO_714 (O_714,N_8790,N_9353);
nor UO_715 (O_715,N_9968,N_8030);
and UO_716 (O_716,N_9465,N_8895);
xor UO_717 (O_717,N_8244,N_8026);
nand UO_718 (O_718,N_9471,N_8240);
or UO_719 (O_719,N_9059,N_9123);
xor UO_720 (O_720,N_9246,N_9233);
nor UO_721 (O_721,N_9434,N_9102);
nor UO_722 (O_722,N_9191,N_9329);
nand UO_723 (O_723,N_9528,N_9978);
xor UO_724 (O_724,N_9821,N_9144);
or UO_725 (O_725,N_8710,N_8532);
nand UO_726 (O_726,N_8183,N_8453);
xnor UO_727 (O_727,N_9205,N_8369);
or UO_728 (O_728,N_8417,N_9816);
and UO_729 (O_729,N_8338,N_8471);
nand UO_730 (O_730,N_8656,N_8930);
nand UO_731 (O_731,N_9071,N_8578);
nand UO_732 (O_732,N_9641,N_9237);
and UO_733 (O_733,N_8175,N_8144);
nand UO_734 (O_734,N_9422,N_8295);
or UO_735 (O_735,N_9410,N_9663);
xor UO_736 (O_736,N_9638,N_9514);
nor UO_737 (O_737,N_8402,N_8045);
nand UO_738 (O_738,N_9048,N_8176);
nand UO_739 (O_739,N_8361,N_8819);
and UO_740 (O_740,N_9164,N_9795);
nand UO_741 (O_741,N_9580,N_9613);
and UO_742 (O_742,N_9960,N_8125);
nor UO_743 (O_743,N_9622,N_8038);
or UO_744 (O_744,N_8006,N_9952);
nand UO_745 (O_745,N_9857,N_9867);
nor UO_746 (O_746,N_8352,N_9137);
nor UO_747 (O_747,N_9298,N_9165);
xnor UO_748 (O_748,N_8104,N_8887);
nor UO_749 (O_749,N_8506,N_8569);
or UO_750 (O_750,N_9596,N_8031);
nor UO_751 (O_751,N_9803,N_8512);
and UO_752 (O_752,N_8553,N_8107);
nand UO_753 (O_753,N_8015,N_8743);
nor UO_754 (O_754,N_8752,N_9117);
nor UO_755 (O_755,N_8123,N_8808);
nor UO_756 (O_756,N_9843,N_9810);
or UO_757 (O_757,N_8341,N_8625);
nor UO_758 (O_758,N_8257,N_8994);
xnor UO_759 (O_759,N_8813,N_9994);
or UO_760 (O_760,N_9299,N_9362);
nor UO_761 (O_761,N_8935,N_8494);
or UO_762 (O_762,N_8617,N_9204);
or UO_763 (O_763,N_9806,N_8966);
nand UO_764 (O_764,N_9598,N_9524);
or UO_765 (O_765,N_9017,N_9297);
nor UO_766 (O_766,N_8094,N_9255);
nand UO_767 (O_767,N_9679,N_8527);
or UO_768 (O_768,N_9876,N_9403);
nor UO_769 (O_769,N_8865,N_8722);
or UO_770 (O_770,N_8259,N_9859);
or UO_771 (O_771,N_8299,N_8804);
and UO_772 (O_772,N_8821,N_8850);
nand UO_773 (O_773,N_9522,N_9334);
or UO_774 (O_774,N_9222,N_8333);
nor UO_775 (O_775,N_8328,N_9953);
and UO_776 (O_776,N_9446,N_9319);
and UO_777 (O_777,N_9272,N_9725);
nand UO_778 (O_778,N_9842,N_9526);
nand UO_779 (O_779,N_9567,N_8256);
or UO_780 (O_780,N_8611,N_8296);
or UO_781 (O_781,N_8830,N_9615);
or UO_782 (O_782,N_8424,N_9011);
nand UO_783 (O_783,N_9196,N_8040);
nor UO_784 (O_784,N_8488,N_9619);
or UO_785 (O_785,N_9801,N_9300);
and UO_786 (O_786,N_8055,N_9231);
or UO_787 (O_787,N_9154,N_8860);
xnor UO_788 (O_788,N_9717,N_8046);
nand UO_789 (O_789,N_9640,N_8021);
nand UO_790 (O_790,N_8096,N_8925);
or UO_791 (O_791,N_9751,N_8119);
and UO_792 (O_792,N_8823,N_8286);
nor UO_793 (O_793,N_8601,N_8831);
nor UO_794 (O_794,N_8372,N_9136);
and UO_795 (O_795,N_8852,N_9338);
nor UO_796 (O_796,N_8952,N_8091);
and UO_797 (O_797,N_8906,N_9787);
or UO_798 (O_798,N_8866,N_8438);
nand UO_799 (O_799,N_8460,N_9681);
or UO_800 (O_800,N_8049,N_8867);
or UO_801 (O_801,N_8658,N_9874);
xor UO_802 (O_802,N_9070,N_8886);
or UO_803 (O_803,N_9145,N_9124);
or UO_804 (O_804,N_9188,N_8973);
nor UO_805 (O_805,N_9624,N_8017);
and UO_806 (O_806,N_8375,N_8238);
nor UO_807 (O_807,N_9099,N_8606);
or UO_808 (O_808,N_8674,N_8199);
nand UO_809 (O_809,N_9733,N_9169);
xnor UO_810 (O_810,N_9106,N_8461);
nor UO_811 (O_811,N_8967,N_8706);
or UO_812 (O_812,N_8047,N_8222);
xnor UO_813 (O_813,N_9768,N_9411);
nor UO_814 (O_814,N_9397,N_9159);
nor UO_815 (O_815,N_8502,N_9993);
nand UO_816 (O_816,N_8261,N_9112);
nand UO_817 (O_817,N_9366,N_9630);
and UO_818 (O_818,N_8334,N_9287);
xor UO_819 (O_819,N_9427,N_9109);
xor UO_820 (O_820,N_9620,N_8689);
nor UO_821 (O_821,N_9322,N_9374);
and UO_822 (O_822,N_8666,N_8998);
or UO_823 (O_823,N_8843,N_9391);
or UO_824 (O_824,N_8824,N_8185);
nor UO_825 (O_825,N_9464,N_9929);
xnor UO_826 (O_826,N_8148,N_8035);
nand UO_827 (O_827,N_9970,N_8600);
or UO_828 (O_828,N_9384,N_8384);
xnor UO_829 (O_829,N_8400,N_8275);
and UO_830 (O_830,N_9309,N_9616);
and UO_831 (O_831,N_8540,N_9499);
nand UO_832 (O_832,N_9021,N_8389);
or UO_833 (O_833,N_8087,N_9936);
nor UO_834 (O_834,N_9704,N_8292);
nand UO_835 (O_835,N_8642,N_9129);
xor UO_836 (O_836,N_8563,N_8787);
nand UO_837 (O_837,N_8561,N_9831);
and UO_838 (O_838,N_8984,N_8694);
and UO_839 (O_839,N_8894,N_8336);
and UO_840 (O_840,N_8805,N_9780);
or UO_841 (O_841,N_9944,N_8013);
nor UO_842 (O_842,N_8735,N_9900);
and UO_843 (O_843,N_8243,N_8778);
nand UO_844 (O_844,N_8179,N_8541);
and UO_845 (O_845,N_8670,N_9506);
nor UO_846 (O_846,N_9421,N_8739);
and UO_847 (O_847,N_8695,N_9600);
nand UO_848 (O_848,N_8153,N_8846);
and UO_849 (O_849,N_9431,N_8556);
or UO_850 (O_850,N_8293,N_9356);
xor UO_851 (O_851,N_9486,N_9853);
nand UO_852 (O_852,N_9242,N_9045);
nand UO_853 (O_853,N_8367,N_8582);
nor UO_854 (O_854,N_9707,N_9817);
nand UO_855 (O_855,N_9254,N_8529);
nand UO_856 (O_856,N_8878,N_8374);
or UO_857 (O_857,N_9807,N_9265);
nand UO_858 (O_858,N_9206,N_9542);
xnor UO_859 (O_859,N_9636,N_9797);
and UO_860 (O_860,N_9933,N_9457);
nand UO_861 (O_861,N_8945,N_8270);
nor UO_862 (O_862,N_8507,N_9263);
nand UO_863 (O_863,N_9895,N_8643);
nand UO_864 (O_864,N_9218,N_8662);
and UO_865 (O_865,N_9212,N_8964);
nand UO_866 (O_866,N_8409,N_9988);
nor UO_867 (O_867,N_8272,N_9767);
or UO_868 (O_868,N_8893,N_9183);
nor UO_869 (O_869,N_8476,N_9937);
nand UO_870 (O_870,N_8131,N_9560);
nor UO_871 (O_871,N_9609,N_8544);
or UO_872 (O_872,N_8154,N_9703);
nor UO_873 (O_873,N_8636,N_8931);
or UO_874 (O_874,N_8485,N_8408);
xnor UO_875 (O_875,N_9350,N_8768);
nor UO_876 (O_876,N_9644,N_9555);
and UO_877 (O_877,N_9412,N_9065);
nand UO_878 (O_878,N_9461,N_8982);
nand UO_879 (O_879,N_9732,N_8716);
or UO_880 (O_880,N_8381,N_8065);
nand UO_881 (O_881,N_8019,N_8191);
nor UO_882 (O_882,N_9893,N_8248);
or UO_883 (O_883,N_8572,N_9967);
and UO_884 (O_884,N_9327,N_8712);
nand UO_885 (O_885,N_8005,N_8487);
and UO_886 (O_886,N_8741,N_9729);
nand UO_887 (O_887,N_8909,N_8344);
nor UO_888 (O_888,N_9020,N_9043);
nor UO_889 (O_889,N_8354,N_8138);
and UO_890 (O_890,N_9447,N_9142);
and UO_891 (O_891,N_9591,N_9118);
nand UO_892 (O_892,N_9139,N_8602);
and UO_893 (O_893,N_9467,N_8622);
and UO_894 (O_894,N_9888,N_8880);
nand UO_895 (O_895,N_8022,N_9194);
nand UO_896 (O_896,N_9294,N_9915);
nand UO_897 (O_897,N_8687,N_8254);
nand UO_898 (O_898,N_9439,N_8789);
nand UO_899 (O_899,N_9957,N_8434);
and UO_900 (O_900,N_9660,N_9687);
xor UO_901 (O_901,N_8797,N_8469);
nor UO_902 (O_902,N_8171,N_9682);
nand UO_903 (O_903,N_9574,N_8397);
and UO_904 (O_904,N_8237,N_9845);
and UO_905 (O_905,N_8903,N_8907);
nor UO_906 (O_906,N_9174,N_8652);
or UO_907 (O_907,N_8864,N_9003);
or UO_908 (O_908,N_9887,N_9752);
or UO_909 (O_909,N_9132,N_8097);
or UO_910 (O_910,N_8730,N_9877);
or UO_911 (O_911,N_8734,N_9094);
nor UO_912 (O_912,N_9187,N_9805);
xor UO_913 (O_913,N_9782,N_9507);
and UO_914 (O_914,N_8163,N_9827);
xor UO_915 (O_915,N_8345,N_8590);
xnor UO_916 (O_916,N_8522,N_8857);
or UO_917 (O_917,N_8940,N_8313);
or UO_918 (O_918,N_8691,N_8519);
and UO_919 (O_919,N_9505,N_9761);
or UO_920 (O_920,N_8386,N_9983);
and UO_921 (O_921,N_9394,N_9369);
xnor UO_922 (O_922,N_8588,N_9487);
nor UO_923 (O_923,N_9878,N_8251);
or UO_924 (O_924,N_9315,N_8736);
nor UO_925 (O_925,N_9945,N_8523);
xor UO_926 (O_926,N_8129,N_8280);
nor UO_927 (O_927,N_8228,N_8667);
nand UO_928 (O_928,N_8193,N_8143);
and UO_929 (O_929,N_9882,N_8764);
xor UO_930 (O_930,N_9658,N_9060);
xor UO_931 (O_931,N_8941,N_9330);
nor UO_932 (O_932,N_9470,N_8227);
and UO_933 (O_933,N_9201,N_8099);
nand UO_934 (O_934,N_8252,N_9030);
and UO_935 (O_935,N_9130,N_9839);
and UO_936 (O_936,N_8683,N_8545);
or UO_937 (O_937,N_8547,N_8206);
or UO_938 (O_938,N_9289,N_9227);
nand UO_939 (O_939,N_9513,N_8215);
nand UO_940 (O_940,N_9651,N_9822);
nand UO_941 (O_941,N_8226,N_9032);
or UO_942 (O_942,N_8003,N_9451);
or UO_943 (O_943,N_9676,N_8366);
nand UO_944 (O_944,N_8801,N_8139);
nand UO_945 (O_945,N_8551,N_8339);
nand UO_946 (O_946,N_8776,N_8210);
xor UO_947 (O_947,N_8637,N_9649);
nor UO_948 (O_948,N_8340,N_8664);
xnor UO_949 (O_949,N_9981,N_8450);
and UO_950 (O_950,N_9320,N_9934);
and UO_951 (O_951,N_8696,N_9563);
nand UO_952 (O_952,N_8812,N_9503);
nand UO_953 (O_953,N_9360,N_9691);
nand UO_954 (O_954,N_8387,N_9898);
nor UO_955 (O_955,N_9458,N_9245);
nand UO_956 (O_956,N_9104,N_9635);
nand UO_957 (O_957,N_8002,N_9838);
nand UO_958 (O_958,N_9764,N_8160);
or UO_959 (O_959,N_9738,N_8577);
nand UO_960 (O_960,N_9248,N_9705);
nor UO_961 (O_961,N_9535,N_8798);
nand UO_962 (O_962,N_8370,N_9734);
nor UO_963 (O_963,N_9478,N_9632);
and UO_964 (O_964,N_9958,N_8159);
or UO_965 (O_965,N_9262,N_8851);
xor UO_966 (O_966,N_9718,N_9368);
nor UO_967 (O_967,N_8814,N_8628);
nand UO_968 (O_968,N_9799,N_9293);
and UO_969 (O_969,N_8620,N_8992);
and UO_970 (O_970,N_8379,N_9361);
nor UO_971 (O_971,N_8298,N_8463);
nor UO_972 (O_972,N_9841,N_9066);
or UO_973 (O_973,N_9278,N_8284);
or UO_974 (O_974,N_9484,N_9711);
and UO_975 (O_975,N_9559,N_8956);
nor UO_976 (O_976,N_9819,N_9530);
or UO_977 (O_977,N_9575,N_8412);
nor UO_978 (O_978,N_9093,N_8586);
nor UO_979 (O_979,N_8651,N_8626);
or UO_980 (O_980,N_8585,N_9047);
nand UO_981 (O_981,N_9168,N_8565);
nand UO_982 (O_982,N_8364,N_9706);
and UO_983 (O_983,N_9107,N_9757);
and UO_984 (O_984,N_9605,N_8146);
nor UO_985 (O_985,N_9343,N_9775);
nand UO_986 (O_986,N_8786,N_8548);
xor UO_987 (O_987,N_8592,N_8791);
xor UO_988 (O_988,N_8822,N_8271);
and UO_989 (O_989,N_9792,N_8834);
nand UO_990 (O_990,N_9786,N_8681);
nand UO_991 (O_991,N_8704,N_9986);
nand UO_992 (O_992,N_8209,N_9543);
xor UO_993 (O_993,N_8763,N_9135);
nand UO_994 (O_994,N_8028,N_9120);
or UO_995 (O_995,N_9171,N_8876);
and UO_996 (O_996,N_8020,N_9390);
or UO_997 (O_997,N_9919,N_8008);
or UO_998 (O_998,N_9924,N_9053);
or UO_999 (O_999,N_8398,N_8399);
or UO_1000 (O_1000,N_8075,N_8196);
nor UO_1001 (O_1001,N_9615,N_9237);
and UO_1002 (O_1002,N_9003,N_9616);
or UO_1003 (O_1003,N_9735,N_9240);
nor UO_1004 (O_1004,N_8713,N_9188);
and UO_1005 (O_1005,N_8564,N_8871);
nor UO_1006 (O_1006,N_9547,N_9238);
and UO_1007 (O_1007,N_9641,N_8633);
nand UO_1008 (O_1008,N_8702,N_8647);
xor UO_1009 (O_1009,N_9689,N_8883);
or UO_1010 (O_1010,N_9855,N_8999);
nor UO_1011 (O_1011,N_9251,N_9291);
or UO_1012 (O_1012,N_8262,N_8384);
or UO_1013 (O_1013,N_9011,N_9606);
nor UO_1014 (O_1014,N_8805,N_9974);
nand UO_1015 (O_1015,N_8723,N_8681);
or UO_1016 (O_1016,N_9883,N_8772);
or UO_1017 (O_1017,N_8624,N_8962);
nand UO_1018 (O_1018,N_8935,N_8141);
nand UO_1019 (O_1019,N_8931,N_9628);
or UO_1020 (O_1020,N_9136,N_9328);
or UO_1021 (O_1021,N_8662,N_8017);
nor UO_1022 (O_1022,N_9550,N_9991);
and UO_1023 (O_1023,N_9903,N_9853);
or UO_1024 (O_1024,N_9712,N_9136);
nand UO_1025 (O_1025,N_9403,N_8515);
xnor UO_1026 (O_1026,N_8826,N_8722);
or UO_1027 (O_1027,N_9465,N_8533);
nand UO_1028 (O_1028,N_9432,N_8825);
nor UO_1029 (O_1029,N_8518,N_8147);
nand UO_1030 (O_1030,N_9494,N_9669);
or UO_1031 (O_1031,N_9405,N_8587);
nand UO_1032 (O_1032,N_9003,N_9885);
nand UO_1033 (O_1033,N_9004,N_9265);
or UO_1034 (O_1034,N_9109,N_8450);
and UO_1035 (O_1035,N_8169,N_9800);
nand UO_1036 (O_1036,N_9685,N_9933);
and UO_1037 (O_1037,N_8016,N_9892);
or UO_1038 (O_1038,N_9187,N_9533);
and UO_1039 (O_1039,N_8033,N_9185);
nand UO_1040 (O_1040,N_8750,N_9888);
and UO_1041 (O_1041,N_8365,N_9081);
nand UO_1042 (O_1042,N_9984,N_9597);
and UO_1043 (O_1043,N_9409,N_8954);
nand UO_1044 (O_1044,N_9524,N_9910);
or UO_1045 (O_1045,N_9215,N_8501);
and UO_1046 (O_1046,N_8748,N_9905);
and UO_1047 (O_1047,N_8806,N_8919);
and UO_1048 (O_1048,N_9686,N_8127);
nand UO_1049 (O_1049,N_9090,N_8251);
xor UO_1050 (O_1050,N_9525,N_9817);
or UO_1051 (O_1051,N_9735,N_8847);
nor UO_1052 (O_1052,N_8233,N_8154);
nor UO_1053 (O_1053,N_8688,N_8656);
nand UO_1054 (O_1054,N_8546,N_8149);
xor UO_1055 (O_1055,N_9568,N_9831);
nor UO_1056 (O_1056,N_8203,N_9367);
nand UO_1057 (O_1057,N_9587,N_8802);
nor UO_1058 (O_1058,N_9669,N_9368);
and UO_1059 (O_1059,N_8191,N_8106);
and UO_1060 (O_1060,N_8463,N_8442);
or UO_1061 (O_1061,N_8133,N_8552);
or UO_1062 (O_1062,N_9341,N_8289);
nor UO_1063 (O_1063,N_8343,N_9421);
or UO_1064 (O_1064,N_9319,N_8149);
and UO_1065 (O_1065,N_8590,N_8840);
xnor UO_1066 (O_1066,N_8487,N_8183);
nor UO_1067 (O_1067,N_8265,N_9419);
nand UO_1068 (O_1068,N_9694,N_9701);
or UO_1069 (O_1069,N_8811,N_9261);
nor UO_1070 (O_1070,N_8260,N_8401);
and UO_1071 (O_1071,N_8654,N_9701);
or UO_1072 (O_1072,N_9702,N_9627);
nor UO_1073 (O_1073,N_9627,N_9250);
nand UO_1074 (O_1074,N_9640,N_8228);
or UO_1075 (O_1075,N_9574,N_8464);
and UO_1076 (O_1076,N_8148,N_9733);
xnor UO_1077 (O_1077,N_8026,N_9283);
nand UO_1078 (O_1078,N_9617,N_8772);
and UO_1079 (O_1079,N_9425,N_9583);
and UO_1080 (O_1080,N_9674,N_8390);
xnor UO_1081 (O_1081,N_9721,N_9678);
nand UO_1082 (O_1082,N_8912,N_8027);
nor UO_1083 (O_1083,N_9424,N_8243);
nor UO_1084 (O_1084,N_9159,N_8739);
nand UO_1085 (O_1085,N_9282,N_8029);
nand UO_1086 (O_1086,N_8754,N_8694);
and UO_1087 (O_1087,N_9953,N_9639);
or UO_1088 (O_1088,N_9103,N_8384);
nand UO_1089 (O_1089,N_8581,N_8509);
nor UO_1090 (O_1090,N_9813,N_9791);
and UO_1091 (O_1091,N_9248,N_8162);
or UO_1092 (O_1092,N_9776,N_9022);
nand UO_1093 (O_1093,N_9111,N_8100);
and UO_1094 (O_1094,N_8179,N_9590);
nor UO_1095 (O_1095,N_8452,N_9627);
xnor UO_1096 (O_1096,N_9132,N_9055);
or UO_1097 (O_1097,N_9069,N_9984);
xor UO_1098 (O_1098,N_8843,N_9717);
and UO_1099 (O_1099,N_8381,N_8260);
and UO_1100 (O_1100,N_9026,N_8121);
nand UO_1101 (O_1101,N_9777,N_8623);
and UO_1102 (O_1102,N_9807,N_9065);
or UO_1103 (O_1103,N_8617,N_8169);
and UO_1104 (O_1104,N_9492,N_9339);
nor UO_1105 (O_1105,N_9766,N_8176);
xor UO_1106 (O_1106,N_9743,N_8000);
or UO_1107 (O_1107,N_8901,N_9558);
or UO_1108 (O_1108,N_9764,N_9797);
nor UO_1109 (O_1109,N_9288,N_8245);
xnor UO_1110 (O_1110,N_8323,N_8776);
nand UO_1111 (O_1111,N_8945,N_9728);
and UO_1112 (O_1112,N_8566,N_9666);
nand UO_1113 (O_1113,N_9705,N_9103);
xnor UO_1114 (O_1114,N_8084,N_9693);
nor UO_1115 (O_1115,N_8424,N_9205);
nand UO_1116 (O_1116,N_8754,N_8853);
nor UO_1117 (O_1117,N_8847,N_9401);
xnor UO_1118 (O_1118,N_9520,N_9805);
or UO_1119 (O_1119,N_8623,N_9736);
nand UO_1120 (O_1120,N_8403,N_9956);
and UO_1121 (O_1121,N_9766,N_8983);
or UO_1122 (O_1122,N_8871,N_9453);
nor UO_1123 (O_1123,N_9151,N_8542);
or UO_1124 (O_1124,N_8785,N_8959);
nand UO_1125 (O_1125,N_9028,N_8841);
nor UO_1126 (O_1126,N_9137,N_9760);
nor UO_1127 (O_1127,N_8969,N_9852);
nor UO_1128 (O_1128,N_8655,N_9219);
nor UO_1129 (O_1129,N_9025,N_9143);
nand UO_1130 (O_1130,N_9246,N_8752);
or UO_1131 (O_1131,N_8628,N_9341);
nor UO_1132 (O_1132,N_8924,N_8376);
or UO_1133 (O_1133,N_8200,N_8684);
or UO_1134 (O_1134,N_9283,N_8498);
nor UO_1135 (O_1135,N_8982,N_8065);
xor UO_1136 (O_1136,N_9831,N_8420);
nor UO_1137 (O_1137,N_8263,N_8617);
nand UO_1138 (O_1138,N_9663,N_9378);
xnor UO_1139 (O_1139,N_9675,N_8182);
or UO_1140 (O_1140,N_8046,N_9362);
or UO_1141 (O_1141,N_9695,N_8937);
nor UO_1142 (O_1142,N_8224,N_8644);
nor UO_1143 (O_1143,N_8419,N_8004);
and UO_1144 (O_1144,N_9998,N_8628);
nor UO_1145 (O_1145,N_8423,N_8976);
nor UO_1146 (O_1146,N_9116,N_8350);
or UO_1147 (O_1147,N_9556,N_9660);
or UO_1148 (O_1148,N_8808,N_9959);
nor UO_1149 (O_1149,N_9659,N_8919);
and UO_1150 (O_1150,N_8230,N_9376);
and UO_1151 (O_1151,N_9337,N_9477);
nor UO_1152 (O_1152,N_9920,N_9007);
nand UO_1153 (O_1153,N_9811,N_8766);
nand UO_1154 (O_1154,N_8686,N_8529);
or UO_1155 (O_1155,N_9594,N_8193);
xor UO_1156 (O_1156,N_8702,N_9471);
or UO_1157 (O_1157,N_9598,N_8380);
and UO_1158 (O_1158,N_9259,N_9378);
or UO_1159 (O_1159,N_9623,N_9307);
and UO_1160 (O_1160,N_8272,N_9118);
xnor UO_1161 (O_1161,N_8928,N_9469);
or UO_1162 (O_1162,N_9535,N_8519);
and UO_1163 (O_1163,N_9237,N_9089);
and UO_1164 (O_1164,N_8018,N_9077);
or UO_1165 (O_1165,N_8038,N_8966);
xor UO_1166 (O_1166,N_9559,N_8107);
or UO_1167 (O_1167,N_8418,N_8681);
nand UO_1168 (O_1168,N_9868,N_8383);
nand UO_1169 (O_1169,N_8280,N_8821);
nand UO_1170 (O_1170,N_8914,N_8879);
xor UO_1171 (O_1171,N_8910,N_9837);
and UO_1172 (O_1172,N_9516,N_9171);
nand UO_1173 (O_1173,N_8347,N_9822);
or UO_1174 (O_1174,N_8849,N_8106);
and UO_1175 (O_1175,N_9461,N_8121);
or UO_1176 (O_1176,N_9328,N_8351);
or UO_1177 (O_1177,N_8185,N_8342);
or UO_1178 (O_1178,N_8576,N_9489);
nand UO_1179 (O_1179,N_9529,N_9982);
or UO_1180 (O_1180,N_8469,N_8589);
xnor UO_1181 (O_1181,N_9362,N_8614);
nand UO_1182 (O_1182,N_9867,N_9859);
xnor UO_1183 (O_1183,N_9230,N_8268);
and UO_1184 (O_1184,N_9697,N_9935);
nand UO_1185 (O_1185,N_8863,N_9184);
xor UO_1186 (O_1186,N_9361,N_8848);
nand UO_1187 (O_1187,N_9828,N_8564);
nand UO_1188 (O_1188,N_9123,N_9670);
nand UO_1189 (O_1189,N_8478,N_8299);
or UO_1190 (O_1190,N_8257,N_8434);
or UO_1191 (O_1191,N_9046,N_9955);
xor UO_1192 (O_1192,N_9635,N_9848);
nor UO_1193 (O_1193,N_8956,N_9114);
and UO_1194 (O_1194,N_9925,N_9476);
xor UO_1195 (O_1195,N_9045,N_8531);
nor UO_1196 (O_1196,N_9270,N_9672);
xnor UO_1197 (O_1197,N_8453,N_8874);
nand UO_1198 (O_1198,N_9142,N_8799);
and UO_1199 (O_1199,N_9138,N_8467);
xor UO_1200 (O_1200,N_8489,N_8816);
nor UO_1201 (O_1201,N_8692,N_8572);
nor UO_1202 (O_1202,N_8000,N_8661);
xnor UO_1203 (O_1203,N_8961,N_9376);
and UO_1204 (O_1204,N_8156,N_8603);
nand UO_1205 (O_1205,N_8943,N_8164);
nand UO_1206 (O_1206,N_8719,N_8651);
nor UO_1207 (O_1207,N_8481,N_8533);
or UO_1208 (O_1208,N_8550,N_8262);
and UO_1209 (O_1209,N_8913,N_8755);
or UO_1210 (O_1210,N_8511,N_8791);
or UO_1211 (O_1211,N_9790,N_8907);
nand UO_1212 (O_1212,N_8598,N_9629);
or UO_1213 (O_1213,N_9731,N_9859);
nand UO_1214 (O_1214,N_8338,N_8253);
and UO_1215 (O_1215,N_8060,N_8309);
and UO_1216 (O_1216,N_8236,N_9674);
nor UO_1217 (O_1217,N_9844,N_9706);
nand UO_1218 (O_1218,N_8418,N_9478);
nor UO_1219 (O_1219,N_9032,N_9476);
and UO_1220 (O_1220,N_8630,N_8933);
nor UO_1221 (O_1221,N_8770,N_8414);
nor UO_1222 (O_1222,N_8124,N_9147);
nand UO_1223 (O_1223,N_9846,N_8050);
nand UO_1224 (O_1224,N_8798,N_9660);
and UO_1225 (O_1225,N_9171,N_9121);
xor UO_1226 (O_1226,N_9508,N_8194);
and UO_1227 (O_1227,N_9494,N_8098);
or UO_1228 (O_1228,N_9002,N_8136);
nor UO_1229 (O_1229,N_9079,N_8301);
nor UO_1230 (O_1230,N_8787,N_9061);
xnor UO_1231 (O_1231,N_9278,N_8363);
nand UO_1232 (O_1232,N_9653,N_8249);
xnor UO_1233 (O_1233,N_8048,N_9729);
nor UO_1234 (O_1234,N_9599,N_8988);
nor UO_1235 (O_1235,N_9047,N_9909);
nor UO_1236 (O_1236,N_9789,N_9562);
or UO_1237 (O_1237,N_9458,N_9523);
or UO_1238 (O_1238,N_8953,N_9700);
and UO_1239 (O_1239,N_9211,N_9233);
xor UO_1240 (O_1240,N_9602,N_9252);
xor UO_1241 (O_1241,N_8250,N_8590);
or UO_1242 (O_1242,N_8724,N_8982);
xor UO_1243 (O_1243,N_8638,N_9860);
xnor UO_1244 (O_1244,N_8834,N_9584);
and UO_1245 (O_1245,N_9039,N_9892);
nor UO_1246 (O_1246,N_9591,N_9192);
and UO_1247 (O_1247,N_9435,N_9769);
xor UO_1248 (O_1248,N_8044,N_9902);
and UO_1249 (O_1249,N_9131,N_8306);
nand UO_1250 (O_1250,N_8408,N_9358);
or UO_1251 (O_1251,N_8351,N_8593);
and UO_1252 (O_1252,N_8038,N_9018);
nand UO_1253 (O_1253,N_8359,N_8864);
nand UO_1254 (O_1254,N_8655,N_9443);
nand UO_1255 (O_1255,N_8633,N_9642);
or UO_1256 (O_1256,N_9273,N_8941);
and UO_1257 (O_1257,N_9852,N_9436);
nand UO_1258 (O_1258,N_9282,N_9882);
nand UO_1259 (O_1259,N_8096,N_9640);
and UO_1260 (O_1260,N_9699,N_9408);
and UO_1261 (O_1261,N_9025,N_8371);
and UO_1262 (O_1262,N_8501,N_9057);
nand UO_1263 (O_1263,N_9958,N_8633);
and UO_1264 (O_1264,N_8614,N_8356);
xor UO_1265 (O_1265,N_9034,N_9491);
nor UO_1266 (O_1266,N_9320,N_8025);
nor UO_1267 (O_1267,N_9964,N_9842);
nand UO_1268 (O_1268,N_9894,N_9582);
nand UO_1269 (O_1269,N_8315,N_8676);
nor UO_1270 (O_1270,N_9335,N_9995);
nand UO_1271 (O_1271,N_8625,N_8924);
nor UO_1272 (O_1272,N_9674,N_8445);
nand UO_1273 (O_1273,N_8736,N_8546);
nand UO_1274 (O_1274,N_8798,N_9935);
and UO_1275 (O_1275,N_9082,N_8382);
and UO_1276 (O_1276,N_8757,N_8565);
nand UO_1277 (O_1277,N_9800,N_8790);
xnor UO_1278 (O_1278,N_8015,N_8974);
or UO_1279 (O_1279,N_9598,N_8387);
xnor UO_1280 (O_1280,N_9125,N_9480);
or UO_1281 (O_1281,N_8861,N_9713);
or UO_1282 (O_1282,N_8243,N_9436);
or UO_1283 (O_1283,N_9105,N_9166);
and UO_1284 (O_1284,N_9624,N_8813);
and UO_1285 (O_1285,N_8334,N_8977);
and UO_1286 (O_1286,N_8065,N_9411);
nor UO_1287 (O_1287,N_8555,N_9559);
nand UO_1288 (O_1288,N_8724,N_8401);
nand UO_1289 (O_1289,N_9686,N_8488);
or UO_1290 (O_1290,N_9111,N_8106);
xor UO_1291 (O_1291,N_9180,N_9151);
xnor UO_1292 (O_1292,N_9146,N_9234);
or UO_1293 (O_1293,N_8407,N_9101);
nand UO_1294 (O_1294,N_9913,N_9370);
nor UO_1295 (O_1295,N_9656,N_9837);
nand UO_1296 (O_1296,N_8582,N_8356);
and UO_1297 (O_1297,N_9846,N_9847);
or UO_1298 (O_1298,N_9987,N_8158);
nor UO_1299 (O_1299,N_9154,N_9674);
nor UO_1300 (O_1300,N_9766,N_9875);
nor UO_1301 (O_1301,N_9660,N_8639);
nor UO_1302 (O_1302,N_8580,N_9708);
nor UO_1303 (O_1303,N_9742,N_9634);
or UO_1304 (O_1304,N_8724,N_9542);
and UO_1305 (O_1305,N_8447,N_8807);
xor UO_1306 (O_1306,N_8085,N_9054);
or UO_1307 (O_1307,N_9755,N_8316);
nand UO_1308 (O_1308,N_8849,N_8095);
nor UO_1309 (O_1309,N_9700,N_8175);
and UO_1310 (O_1310,N_9621,N_9284);
nor UO_1311 (O_1311,N_8385,N_8563);
nand UO_1312 (O_1312,N_8476,N_9445);
and UO_1313 (O_1313,N_9898,N_9354);
or UO_1314 (O_1314,N_9541,N_8152);
nand UO_1315 (O_1315,N_9389,N_9638);
and UO_1316 (O_1316,N_8766,N_9127);
and UO_1317 (O_1317,N_9088,N_8671);
nor UO_1318 (O_1318,N_8861,N_8592);
xnor UO_1319 (O_1319,N_8530,N_9362);
and UO_1320 (O_1320,N_9793,N_8877);
or UO_1321 (O_1321,N_8553,N_8474);
nor UO_1322 (O_1322,N_9935,N_9830);
nand UO_1323 (O_1323,N_8168,N_9651);
and UO_1324 (O_1324,N_8386,N_8093);
xor UO_1325 (O_1325,N_9035,N_8677);
nor UO_1326 (O_1326,N_8631,N_8262);
or UO_1327 (O_1327,N_8491,N_8390);
or UO_1328 (O_1328,N_8733,N_9460);
nand UO_1329 (O_1329,N_8339,N_9602);
nand UO_1330 (O_1330,N_9520,N_9383);
or UO_1331 (O_1331,N_9000,N_8881);
nand UO_1332 (O_1332,N_8896,N_8303);
or UO_1333 (O_1333,N_8509,N_9737);
nor UO_1334 (O_1334,N_9852,N_8965);
or UO_1335 (O_1335,N_9274,N_9147);
and UO_1336 (O_1336,N_9313,N_9700);
nor UO_1337 (O_1337,N_9682,N_9301);
nor UO_1338 (O_1338,N_8367,N_9848);
xor UO_1339 (O_1339,N_9964,N_8102);
xnor UO_1340 (O_1340,N_9285,N_9928);
or UO_1341 (O_1341,N_8914,N_8413);
nor UO_1342 (O_1342,N_8800,N_8011);
nand UO_1343 (O_1343,N_8030,N_9167);
nor UO_1344 (O_1344,N_9628,N_8132);
and UO_1345 (O_1345,N_8013,N_9755);
or UO_1346 (O_1346,N_8459,N_8016);
nand UO_1347 (O_1347,N_9754,N_8497);
or UO_1348 (O_1348,N_9876,N_8395);
or UO_1349 (O_1349,N_8023,N_9337);
nor UO_1350 (O_1350,N_8263,N_9992);
xnor UO_1351 (O_1351,N_9244,N_9896);
xnor UO_1352 (O_1352,N_8427,N_8447);
and UO_1353 (O_1353,N_8894,N_8852);
nand UO_1354 (O_1354,N_9357,N_9665);
nand UO_1355 (O_1355,N_8107,N_9420);
nor UO_1356 (O_1356,N_9367,N_9802);
and UO_1357 (O_1357,N_8656,N_8360);
nand UO_1358 (O_1358,N_9342,N_8049);
nand UO_1359 (O_1359,N_8611,N_9120);
or UO_1360 (O_1360,N_9837,N_9876);
xnor UO_1361 (O_1361,N_9916,N_9623);
and UO_1362 (O_1362,N_9455,N_8823);
nor UO_1363 (O_1363,N_8093,N_8962);
nor UO_1364 (O_1364,N_8277,N_8319);
or UO_1365 (O_1365,N_9985,N_8579);
nor UO_1366 (O_1366,N_9869,N_9912);
or UO_1367 (O_1367,N_9077,N_9004);
nand UO_1368 (O_1368,N_9110,N_8719);
or UO_1369 (O_1369,N_8440,N_8978);
nor UO_1370 (O_1370,N_8897,N_8134);
nor UO_1371 (O_1371,N_9214,N_9135);
nand UO_1372 (O_1372,N_9082,N_9299);
and UO_1373 (O_1373,N_8195,N_9649);
or UO_1374 (O_1374,N_9684,N_9167);
or UO_1375 (O_1375,N_8825,N_8111);
or UO_1376 (O_1376,N_9023,N_8028);
nand UO_1377 (O_1377,N_9875,N_9361);
xor UO_1378 (O_1378,N_8114,N_8531);
or UO_1379 (O_1379,N_8205,N_8718);
nor UO_1380 (O_1380,N_9673,N_9259);
nand UO_1381 (O_1381,N_8760,N_8144);
nor UO_1382 (O_1382,N_9914,N_9509);
nor UO_1383 (O_1383,N_8824,N_9375);
and UO_1384 (O_1384,N_8440,N_8567);
nor UO_1385 (O_1385,N_8425,N_9870);
nand UO_1386 (O_1386,N_9950,N_9291);
and UO_1387 (O_1387,N_8693,N_8553);
or UO_1388 (O_1388,N_9864,N_8227);
or UO_1389 (O_1389,N_9800,N_8190);
and UO_1390 (O_1390,N_8902,N_9976);
or UO_1391 (O_1391,N_8934,N_8386);
and UO_1392 (O_1392,N_9392,N_8127);
nand UO_1393 (O_1393,N_8821,N_8765);
or UO_1394 (O_1394,N_9202,N_8797);
nor UO_1395 (O_1395,N_8968,N_8463);
and UO_1396 (O_1396,N_9016,N_9181);
or UO_1397 (O_1397,N_9268,N_9189);
nand UO_1398 (O_1398,N_8861,N_9264);
and UO_1399 (O_1399,N_8126,N_9049);
nor UO_1400 (O_1400,N_9063,N_9739);
nand UO_1401 (O_1401,N_9141,N_8280);
and UO_1402 (O_1402,N_8511,N_8239);
nand UO_1403 (O_1403,N_8085,N_9212);
or UO_1404 (O_1404,N_9004,N_8910);
or UO_1405 (O_1405,N_9901,N_8911);
nand UO_1406 (O_1406,N_9045,N_8887);
and UO_1407 (O_1407,N_8035,N_8860);
xor UO_1408 (O_1408,N_9498,N_9586);
and UO_1409 (O_1409,N_9463,N_9121);
nand UO_1410 (O_1410,N_9304,N_9758);
and UO_1411 (O_1411,N_8632,N_8433);
nand UO_1412 (O_1412,N_8107,N_8398);
and UO_1413 (O_1413,N_9829,N_9680);
and UO_1414 (O_1414,N_9121,N_9523);
xnor UO_1415 (O_1415,N_8034,N_8028);
or UO_1416 (O_1416,N_8470,N_8417);
nor UO_1417 (O_1417,N_9442,N_8810);
nor UO_1418 (O_1418,N_8155,N_9586);
nand UO_1419 (O_1419,N_9520,N_9286);
nor UO_1420 (O_1420,N_9028,N_9175);
nand UO_1421 (O_1421,N_8878,N_9555);
nor UO_1422 (O_1422,N_8890,N_9863);
and UO_1423 (O_1423,N_9696,N_8726);
and UO_1424 (O_1424,N_9089,N_9685);
nor UO_1425 (O_1425,N_8497,N_9614);
and UO_1426 (O_1426,N_8009,N_8055);
and UO_1427 (O_1427,N_9964,N_9369);
nor UO_1428 (O_1428,N_9047,N_8813);
and UO_1429 (O_1429,N_9908,N_8237);
and UO_1430 (O_1430,N_8557,N_9196);
nand UO_1431 (O_1431,N_8277,N_9677);
or UO_1432 (O_1432,N_9146,N_8794);
nand UO_1433 (O_1433,N_9587,N_9483);
and UO_1434 (O_1434,N_8671,N_9171);
nand UO_1435 (O_1435,N_8481,N_9057);
and UO_1436 (O_1436,N_8626,N_9871);
nor UO_1437 (O_1437,N_9415,N_8481);
or UO_1438 (O_1438,N_8985,N_9184);
xor UO_1439 (O_1439,N_9665,N_8989);
and UO_1440 (O_1440,N_8267,N_8687);
nand UO_1441 (O_1441,N_8419,N_8147);
and UO_1442 (O_1442,N_9957,N_9094);
nand UO_1443 (O_1443,N_9034,N_9968);
and UO_1444 (O_1444,N_9671,N_8329);
or UO_1445 (O_1445,N_9001,N_8206);
and UO_1446 (O_1446,N_9267,N_8410);
xor UO_1447 (O_1447,N_8703,N_8518);
or UO_1448 (O_1448,N_9330,N_8969);
or UO_1449 (O_1449,N_9661,N_8663);
and UO_1450 (O_1450,N_8598,N_8684);
nor UO_1451 (O_1451,N_9325,N_8393);
nand UO_1452 (O_1452,N_8171,N_9044);
xor UO_1453 (O_1453,N_9076,N_8232);
nor UO_1454 (O_1454,N_9030,N_9873);
nor UO_1455 (O_1455,N_9247,N_9554);
nor UO_1456 (O_1456,N_8030,N_8308);
nand UO_1457 (O_1457,N_9850,N_8018);
nand UO_1458 (O_1458,N_9689,N_9811);
nor UO_1459 (O_1459,N_8880,N_8474);
nor UO_1460 (O_1460,N_8200,N_9373);
and UO_1461 (O_1461,N_9941,N_8797);
nand UO_1462 (O_1462,N_8567,N_8747);
nor UO_1463 (O_1463,N_9032,N_9534);
nor UO_1464 (O_1464,N_8796,N_8471);
nor UO_1465 (O_1465,N_9309,N_8951);
or UO_1466 (O_1466,N_9042,N_9855);
xnor UO_1467 (O_1467,N_9130,N_9164);
and UO_1468 (O_1468,N_9755,N_9899);
nor UO_1469 (O_1469,N_8111,N_9752);
nor UO_1470 (O_1470,N_8435,N_8684);
nor UO_1471 (O_1471,N_9910,N_9812);
nor UO_1472 (O_1472,N_9035,N_9610);
or UO_1473 (O_1473,N_9574,N_9679);
xnor UO_1474 (O_1474,N_8305,N_8146);
xor UO_1475 (O_1475,N_9996,N_9473);
nand UO_1476 (O_1476,N_9860,N_8433);
or UO_1477 (O_1477,N_8451,N_8855);
nand UO_1478 (O_1478,N_9926,N_8254);
nand UO_1479 (O_1479,N_8578,N_8277);
and UO_1480 (O_1480,N_8907,N_8241);
nand UO_1481 (O_1481,N_9772,N_8742);
or UO_1482 (O_1482,N_8344,N_8343);
nand UO_1483 (O_1483,N_9458,N_8743);
nand UO_1484 (O_1484,N_9884,N_9154);
nand UO_1485 (O_1485,N_9929,N_9917);
nand UO_1486 (O_1486,N_9574,N_8824);
or UO_1487 (O_1487,N_8595,N_8384);
nand UO_1488 (O_1488,N_8804,N_9132);
nand UO_1489 (O_1489,N_8480,N_9408);
nor UO_1490 (O_1490,N_9188,N_8345);
or UO_1491 (O_1491,N_9741,N_8779);
and UO_1492 (O_1492,N_9633,N_8453);
nor UO_1493 (O_1493,N_8963,N_8137);
nor UO_1494 (O_1494,N_8591,N_8994);
nor UO_1495 (O_1495,N_8952,N_9381);
xor UO_1496 (O_1496,N_9034,N_8755);
and UO_1497 (O_1497,N_9733,N_9342);
or UO_1498 (O_1498,N_8266,N_8923);
and UO_1499 (O_1499,N_8503,N_9039);
endmodule