module basic_1000_10000_1500_5_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_624,In_323);
xor U1 (N_1,In_539,In_686);
and U2 (N_2,In_788,In_694);
and U3 (N_3,In_571,In_497);
and U4 (N_4,In_358,In_823);
nor U5 (N_5,In_85,In_670);
nand U6 (N_6,In_349,In_715);
or U7 (N_7,In_496,In_545);
nand U8 (N_8,In_92,In_688);
or U9 (N_9,In_508,In_708);
and U10 (N_10,In_998,In_910);
nor U11 (N_11,In_561,In_124);
or U12 (N_12,In_459,In_369);
xor U13 (N_13,In_880,In_86);
and U14 (N_14,In_607,In_639);
or U15 (N_15,In_273,In_113);
nand U16 (N_16,In_490,In_172);
or U17 (N_17,In_696,In_631);
and U18 (N_18,In_598,In_156);
and U19 (N_19,In_507,In_814);
nor U20 (N_20,In_583,In_564);
nand U21 (N_21,In_955,In_640);
and U22 (N_22,In_22,In_858);
or U23 (N_23,In_592,In_39);
and U24 (N_24,In_107,In_372);
and U25 (N_25,In_612,In_572);
or U26 (N_26,In_779,In_438);
or U27 (N_27,In_443,In_57);
nor U28 (N_28,In_799,In_440);
and U29 (N_29,In_394,In_954);
xor U30 (N_30,In_383,In_526);
nor U31 (N_31,In_642,In_802);
xor U32 (N_32,In_519,In_704);
or U33 (N_33,In_214,In_832);
or U34 (N_34,In_155,In_341);
nand U35 (N_35,In_366,In_887);
or U36 (N_36,In_168,In_308);
or U37 (N_37,In_560,In_988);
or U38 (N_38,In_246,In_947);
or U39 (N_39,In_542,In_979);
or U40 (N_40,In_853,In_118);
nor U41 (N_41,In_483,In_337);
nor U42 (N_42,In_744,In_36);
and U43 (N_43,In_651,In_895);
or U44 (N_44,In_252,In_206);
nand U45 (N_45,In_509,In_709);
or U46 (N_46,In_878,In_675);
xor U47 (N_47,In_902,In_233);
and U48 (N_48,In_72,In_790);
xor U49 (N_49,In_112,In_205);
or U50 (N_50,In_740,In_978);
or U51 (N_51,In_837,In_742);
and U52 (N_52,In_711,In_812);
nor U53 (N_53,In_557,In_753);
or U54 (N_54,In_678,In_787);
nor U55 (N_55,In_981,In_730);
nand U56 (N_56,In_75,In_356);
or U57 (N_57,In_136,In_845);
or U58 (N_58,In_284,In_830);
or U59 (N_59,In_807,In_35);
and U60 (N_60,In_319,In_302);
xor U61 (N_61,In_18,In_839);
or U62 (N_62,In_305,In_605);
nor U63 (N_63,In_908,In_444);
nor U64 (N_64,In_140,In_577);
and U65 (N_65,In_520,In_452);
nor U66 (N_66,In_211,In_485);
xnor U67 (N_67,In_946,In_864);
nand U68 (N_68,In_130,In_419);
xnor U69 (N_69,In_149,In_566);
nand U70 (N_70,In_184,In_332);
nor U71 (N_71,In_949,In_238);
and U72 (N_72,In_748,In_403);
and U73 (N_73,In_926,In_404);
or U74 (N_74,In_927,In_276);
and U75 (N_75,In_773,In_568);
nor U76 (N_76,In_277,In_900);
nor U77 (N_77,In_739,In_439);
xor U78 (N_78,In_614,In_396);
or U79 (N_79,In_964,In_856);
nor U80 (N_80,In_78,In_848);
nor U81 (N_81,In_749,In_79);
or U82 (N_82,In_61,In_666);
nor U83 (N_83,In_601,In_693);
nor U84 (N_84,In_153,In_850);
nor U85 (N_85,In_574,In_942);
nor U86 (N_86,In_772,In_762);
or U87 (N_87,In_728,In_227);
and U88 (N_88,In_138,In_881);
nor U89 (N_89,In_258,In_602);
and U90 (N_90,In_585,In_215);
nor U91 (N_91,In_167,In_781);
and U92 (N_92,In_528,In_84);
nand U93 (N_93,In_294,In_83);
or U94 (N_94,In_402,In_93);
and U95 (N_95,In_719,In_523);
and U96 (N_96,In_334,In_108);
nor U97 (N_97,In_25,In_522);
nand U98 (N_98,In_311,In_775);
and U99 (N_99,In_400,In_635);
nor U100 (N_100,In_997,In_662);
xor U101 (N_101,In_27,In_17);
nand U102 (N_102,In_747,In_914);
nand U103 (N_103,In_811,In_549);
or U104 (N_104,In_890,In_906);
or U105 (N_105,In_993,In_985);
nand U106 (N_106,In_892,In_201);
nand U107 (N_107,In_331,In_145);
nor U108 (N_108,In_661,In_296);
or U109 (N_109,In_968,In_875);
or U110 (N_110,In_951,In_865);
or U111 (N_111,In_831,In_2);
nor U112 (N_112,In_795,In_385);
and U113 (N_113,In_267,In_819);
nor U114 (N_114,In_537,In_576);
and U115 (N_115,In_259,In_89);
and U116 (N_116,In_984,In_898);
or U117 (N_117,In_445,In_37);
nand U118 (N_118,In_594,In_120);
nor U119 (N_119,In_553,In_306);
nor U120 (N_120,In_916,In_879);
nor U121 (N_121,In_643,In_973);
or U122 (N_122,In_411,In_854);
and U123 (N_123,In_421,In_745);
nor U124 (N_124,In_114,In_610);
nor U125 (N_125,In_347,In_418);
and U126 (N_126,In_424,In_501);
nor U127 (N_127,In_516,In_46);
or U128 (N_128,In_30,In_533);
xor U129 (N_129,In_453,In_73);
nand U130 (N_130,In_798,In_198);
or U131 (N_131,In_451,In_115);
or U132 (N_132,In_467,In_231);
or U133 (N_133,In_74,In_436);
xor U134 (N_134,In_899,In_959);
nor U135 (N_135,In_518,In_531);
and U136 (N_136,In_464,In_38);
nor U137 (N_137,In_468,In_119);
xnor U138 (N_138,In_558,In_407);
nand U139 (N_139,In_353,In_570);
and U140 (N_140,In_3,In_941);
and U141 (N_141,In_915,In_446);
nand U142 (N_142,In_945,In_230);
xor U143 (N_143,In_345,In_972);
nand U144 (N_144,In_556,In_398);
xnor U145 (N_145,In_471,In_622);
and U146 (N_146,In_187,In_563);
nor U147 (N_147,In_186,In_213);
nor U148 (N_148,In_877,In_203);
or U149 (N_149,In_989,In_660);
nand U150 (N_150,In_283,In_310);
nor U151 (N_151,In_650,In_222);
nor U152 (N_152,In_96,In_503);
or U153 (N_153,In_588,In_499);
and U154 (N_154,In_7,In_293);
or U155 (N_155,In_484,In_101);
or U156 (N_156,In_611,In_554);
and U157 (N_157,In_815,In_532);
and U158 (N_158,In_226,In_94);
or U159 (N_159,In_433,In_32);
nand U160 (N_160,In_913,In_426);
nor U161 (N_161,In_207,In_844);
nor U162 (N_162,In_770,In_106);
nand U163 (N_163,In_876,In_489);
nand U164 (N_164,In_615,In_874);
nor U165 (N_165,In_656,In_741);
nand U166 (N_166,In_548,In_920);
and U167 (N_167,In_559,In_822);
or U168 (N_168,In_194,In_122);
nor U169 (N_169,In_596,In_801);
or U170 (N_170,In_251,In_885);
xnor U171 (N_171,In_434,In_743);
nor U172 (N_172,In_735,In_804);
nor U173 (N_173,In_212,In_986);
nand U174 (N_174,In_768,In_15);
and U175 (N_175,In_161,In_463);
xnor U176 (N_176,In_759,In_47);
nand U177 (N_177,In_692,In_809);
xor U178 (N_178,In_295,In_423);
or U179 (N_179,In_291,In_729);
xor U180 (N_180,In_977,In_0);
nand U181 (N_181,In_150,In_325);
or U182 (N_182,In_966,In_309);
nor U183 (N_183,In_317,In_128);
nand U184 (N_184,In_28,In_725);
or U185 (N_185,In_700,In_943);
nor U186 (N_186,In_912,In_192);
nor U187 (N_187,In_368,In_248);
xnor U188 (N_188,In_689,In_684);
or U189 (N_189,In_657,In_613);
xor U190 (N_190,In_330,In_44);
and U191 (N_191,In_191,In_806);
and U192 (N_192,In_163,In_871);
and U193 (N_193,In_546,In_158);
nor U194 (N_194,In_405,In_617);
or U195 (N_195,In_764,In_506);
nor U196 (N_196,In_384,In_782);
xnor U197 (N_197,In_682,In_838);
nand U198 (N_198,In_491,In_447);
or U199 (N_199,In_975,In_290);
or U200 (N_200,In_808,In_766);
or U201 (N_201,In_458,In_618);
nor U202 (N_202,In_274,In_783);
nand U203 (N_203,In_109,In_415);
nand U204 (N_204,In_278,In_97);
nand U205 (N_205,In_600,In_188);
nand U206 (N_206,In_714,In_91);
and U207 (N_207,In_940,In_166);
and U208 (N_208,In_575,In_71);
nand U209 (N_209,In_282,In_690);
nand U210 (N_210,In_909,In_144);
and U211 (N_211,In_866,In_638);
xnor U212 (N_212,In_843,In_51);
or U213 (N_213,In_751,In_621);
nor U214 (N_214,In_174,In_873);
nor U215 (N_215,In_448,In_774);
nor U216 (N_216,In_703,In_399);
nand U217 (N_217,In_412,In_761);
or U218 (N_218,In_98,In_695);
and U219 (N_219,In_314,In_454);
or U220 (N_220,In_994,In_197);
or U221 (N_221,In_281,In_388);
nor U222 (N_222,In_374,In_250);
and U223 (N_223,In_59,In_182);
nor U224 (N_224,In_377,In_534);
xor U225 (N_225,In_579,In_633);
or U226 (N_226,In_189,In_196);
nand U227 (N_227,In_636,In_100);
or U228 (N_228,In_147,In_886);
xor U229 (N_229,In_970,In_199);
nor U230 (N_230,In_929,In_488);
or U231 (N_231,In_77,In_350);
and U232 (N_232,In_141,In_195);
nand U233 (N_233,In_934,In_237);
and U234 (N_234,In_465,In_375);
and U235 (N_235,In_56,In_363);
or U236 (N_236,In_442,In_235);
and U237 (N_237,In_589,In_313);
nor U238 (N_238,In_272,In_606);
nor U239 (N_239,In_316,In_476);
nand U240 (N_240,In_771,In_724);
and U241 (N_241,In_595,In_584);
and U242 (N_242,In_239,In_6);
and U243 (N_243,In_287,In_225);
nor U244 (N_244,In_521,In_827);
xnor U245 (N_245,In_344,In_181);
nand U246 (N_246,In_364,In_872);
nand U247 (N_247,In_505,In_297);
nand U248 (N_248,In_665,In_386);
and U249 (N_249,In_324,In_301);
xnor U250 (N_250,In_409,In_530);
nand U251 (N_251,In_343,In_604);
or U252 (N_252,In_930,In_637);
or U253 (N_253,In_472,In_234);
and U254 (N_254,In_702,In_710);
or U255 (N_255,In_996,In_65);
xor U256 (N_256,In_387,In_911);
and U257 (N_257,In_907,In_681);
xnor U258 (N_258,In_918,In_544);
nor U259 (N_259,In_190,In_705);
nor U260 (N_260,In_983,In_321);
nor U261 (N_261,In_420,In_133);
nand U262 (N_262,In_517,In_922);
nand U263 (N_263,In_414,In_938);
nor U264 (N_264,In_852,In_470);
and U265 (N_265,In_285,In_591);
and U266 (N_266,In_253,In_132);
or U267 (N_267,In_718,In_990);
xnor U268 (N_268,In_789,In_889);
and U269 (N_269,In_580,In_159);
or U270 (N_270,In_395,In_820);
nand U271 (N_271,In_180,In_373);
nor U272 (N_272,In_732,In_925);
nor U273 (N_273,In_551,In_641);
and U274 (N_274,In_219,In_367);
nand U275 (N_275,In_805,In_683);
or U276 (N_276,In_992,In_70);
nand U277 (N_277,In_66,In_967);
nor U278 (N_278,In_378,In_103);
and U279 (N_279,In_469,In_625);
or U280 (N_280,In_371,In_896);
or U281 (N_281,In_340,In_143);
nand U282 (N_282,In_160,In_50);
nand U283 (N_283,In_179,In_303);
nand U284 (N_284,In_868,In_354);
nand U285 (N_285,In_541,In_220);
nor U286 (N_286,In_137,In_152);
and U287 (N_287,In_401,In_536);
xor U288 (N_288,In_300,In_963);
nor U289 (N_289,In_667,In_723);
or U290 (N_290,In_9,In_34);
nor U291 (N_291,In_578,In_664);
and U292 (N_292,In_720,In_626);
and U293 (N_293,In_339,In_416);
nor U294 (N_294,In_223,In_649);
nand U295 (N_295,In_901,In_826);
or U296 (N_296,In_860,In_193);
and U297 (N_297,In_502,In_142);
and U298 (N_298,In_312,In_49);
nand U299 (N_299,In_738,In_169);
and U300 (N_300,In_221,In_58);
or U301 (N_301,In_746,In_757);
nand U302 (N_302,In_348,In_961);
or U303 (N_303,In_135,In_99);
or U304 (N_304,In_244,In_55);
xnor U305 (N_305,In_413,In_357);
or U306 (N_306,In_264,In_698);
and U307 (N_307,In_699,In_652);
nand U308 (N_308,In_53,In_919);
xor U309 (N_309,In_905,In_841);
nor U310 (N_310,In_478,In_634);
and U311 (N_311,In_824,In_170);
nand U312 (N_312,In_241,In_755);
or U313 (N_313,In_849,In_995);
or U314 (N_314,In_721,In_60);
nand U315 (N_315,In_381,In_261);
and U316 (N_316,In_67,In_380);
nand U317 (N_317,In_177,In_110);
or U318 (N_318,In_165,In_217);
and U319 (N_319,In_62,In_432);
nor U320 (N_320,In_322,In_825);
or U321 (N_321,In_767,In_45);
nand U322 (N_322,In_288,In_209);
or U323 (N_323,In_455,In_847);
nand U324 (N_324,In_888,In_431);
and U325 (N_325,In_645,In_971);
xnor U326 (N_326,In_76,In_410);
nor U327 (N_327,In_8,In_646);
nand U328 (N_328,In_538,In_336);
xor U329 (N_329,In_726,In_632);
xnor U330 (N_330,In_23,In_279);
nand U331 (N_331,In_731,In_500);
or U332 (N_332,In_780,In_792);
or U333 (N_333,In_90,In_701);
and U334 (N_334,In_256,In_26);
and U335 (N_335,In_111,In_462);
nor U336 (N_336,In_857,In_473);
or U337 (N_337,In_449,In_859);
nor U338 (N_338,In_754,In_175);
nand U339 (N_339,In_123,In_543);
nor U340 (N_340,In_48,In_893);
or U341 (N_341,In_178,In_786);
and U342 (N_342,In_619,In_923);
xor U343 (N_343,In_88,In_733);
nand U344 (N_344,In_659,In_224);
xor U345 (N_345,In_525,In_286);
and U346 (N_346,In_917,In_535);
or U347 (N_347,In_833,In_482);
or U348 (N_348,In_836,In_817);
nand U349 (N_349,In_529,In_262);
or U350 (N_350,In_862,In_390);
and U351 (N_351,In_254,In_351);
xnor U352 (N_352,In_430,In_586);
nor U353 (N_353,In_846,In_527);
nand U354 (N_354,In_629,In_894);
nand U355 (N_355,In_391,In_627);
xor U356 (N_356,In_461,In_840);
nand U357 (N_357,In_63,In_329);
and U358 (N_358,In_382,In_102);
and U359 (N_359,In_884,In_33);
nand U360 (N_360,In_569,In_477);
xnor U361 (N_361,In_495,In_355);
and U362 (N_362,In_289,In_280);
nand U363 (N_363,In_987,In_243);
nand U364 (N_364,In_304,In_697);
and U365 (N_365,In_734,In_486);
or U366 (N_366,In_760,In_249);
and U367 (N_367,In_958,In_555);
nand U368 (N_368,In_931,In_957);
and U369 (N_369,In_81,In_104);
and U370 (N_370,In_597,In_31);
nand U371 (N_371,In_376,In_821);
nand U372 (N_372,In_80,In_736);
and U373 (N_373,In_932,In_68);
nor U374 (N_374,In_456,In_722);
and U375 (N_375,In_673,In_512);
xnor U376 (N_376,In_151,In_370);
nor U377 (N_377,In_794,In_352);
nand U378 (N_378,In_752,In_474);
and U379 (N_379,In_183,In_52);
or U380 (N_380,In_552,In_361);
or U381 (N_381,In_457,In_515);
or U382 (N_382,In_204,In_712);
xor U383 (N_383,In_608,In_493);
nand U384 (N_384,In_653,In_342);
nand U385 (N_385,In_164,In_64);
nor U386 (N_386,In_154,In_939);
nand U387 (N_387,In_263,In_674);
nor U388 (N_388,In_437,In_365);
or U389 (N_389,In_573,In_318);
and U390 (N_390,In_524,In_127);
and U391 (N_391,In_691,In_883);
xor U392 (N_392,In_139,In_976);
nand U393 (N_393,In_54,In_320);
or U394 (N_394,In_778,In_679);
and U395 (N_395,In_12,In_565);
nand U396 (N_396,In_924,In_327);
or U397 (N_397,In_750,In_991);
nor U398 (N_398,In_935,In_245);
and U399 (N_399,In_587,In_232);
and U400 (N_400,In_903,In_813);
and U401 (N_401,In_417,In_796);
or U402 (N_402,In_654,In_173);
xor U403 (N_403,In_867,In_216);
or U404 (N_404,In_328,In_897);
and U405 (N_405,In_630,In_359);
and U406 (N_406,In_937,In_668);
and U407 (N_407,In_737,In_540);
or U408 (N_408,In_793,In_863);
and U409 (N_409,In_904,In_504);
and U410 (N_410,In_146,In_389);
nor U411 (N_411,In_861,In_891);
or U412 (N_412,In_427,In_707);
or U413 (N_413,In_777,In_672);
xor U414 (N_414,In_785,In_362);
nand U415 (N_415,In_648,In_335);
nor U416 (N_416,In_948,In_999);
and U417 (N_417,In_628,In_16);
nand U418 (N_418,In_818,In_129);
and U419 (N_419,In_450,In_270);
nand U420 (N_420,In_42,In_481);
xnor U421 (N_421,In_275,In_5);
and U422 (N_422,In_962,In_157);
or U423 (N_423,In_117,In_599);
or U424 (N_424,In_466,In_346);
nand U425 (N_425,In_406,In_265);
and U426 (N_426,In_870,In_593);
or U427 (N_427,In_14,In_933);
nand U428 (N_428,In_228,In_148);
nor U429 (N_429,In_202,In_487);
and U430 (N_430,In_623,In_460);
or U431 (N_431,In_299,In_255);
nor U432 (N_432,In_492,In_271);
or U433 (N_433,In_676,In_965);
or U434 (N_434,In_727,In_247);
or U435 (N_435,In_810,In_428);
nand U436 (N_436,In_1,In_69);
nand U437 (N_437,In_706,In_41);
and U438 (N_438,In_765,In_680);
nor U439 (N_439,In_855,In_562);
or U440 (N_440,In_200,In_208);
nand U441 (N_441,In_763,In_510);
nand U442 (N_442,In_10,In_479);
and U443 (N_443,In_842,In_784);
and U444 (N_444,In_797,In_257);
nor U445 (N_445,In_882,In_269);
or U446 (N_446,In_669,In_980);
and U447 (N_447,In_422,In_658);
nand U448 (N_448,In_717,In_581);
nor U449 (N_449,In_260,In_982);
nand U450 (N_450,In_498,In_835);
and U451 (N_451,In_218,In_338);
nand U452 (N_452,In_511,In_24);
or U453 (N_453,In_121,In_40);
or U454 (N_454,In_928,In_603);
nand U455 (N_455,In_87,In_567);
or U456 (N_456,In_126,In_210);
nand U457 (N_457,In_828,In_663);
or U458 (N_458,In_713,In_974);
nor U459 (N_459,In_834,In_475);
and U460 (N_460,In_514,In_43);
and U461 (N_461,In_758,In_392);
and U462 (N_462,In_307,In_229);
and U463 (N_463,In_236,In_869);
nand U464 (N_464,In_677,In_829);
nor U465 (N_465,In_393,In_19);
or U466 (N_466,In_791,In_240);
nor U467 (N_467,In_547,In_105);
nor U468 (N_468,In_776,In_936);
or U469 (N_469,In_266,In_171);
xnor U470 (N_470,In_4,In_441);
nor U471 (N_471,In_956,In_425);
or U472 (N_472,In_13,In_480);
and U473 (N_473,In_969,In_268);
or U474 (N_474,In_513,In_550);
nand U475 (N_475,In_134,In_125);
or U476 (N_476,In_162,In_326);
and U477 (N_477,In_644,In_816);
and U478 (N_478,In_397,In_582);
nor U479 (N_479,In_11,In_769);
nand U480 (N_480,In_116,In_185);
nor U481 (N_481,In_131,In_408);
nand U482 (N_482,In_756,In_315);
nor U483 (N_483,In_944,In_960);
and U484 (N_484,In_655,In_242);
or U485 (N_485,In_921,In_851);
nor U486 (N_486,In_671,In_620);
nand U487 (N_487,In_953,In_333);
or U488 (N_488,In_685,In_292);
nand U489 (N_489,In_429,In_952);
nand U490 (N_490,In_609,In_716);
nor U491 (N_491,In_800,In_20);
nand U492 (N_492,In_379,In_590);
nor U493 (N_493,In_950,In_21);
nand U494 (N_494,In_435,In_29);
and U495 (N_495,In_803,In_95);
and U496 (N_496,In_647,In_494);
or U497 (N_497,In_616,In_176);
nor U498 (N_498,In_360,In_298);
and U499 (N_499,In_82,In_687);
nand U500 (N_500,In_757,In_668);
xor U501 (N_501,In_50,In_964);
xnor U502 (N_502,In_308,In_383);
and U503 (N_503,In_666,In_878);
and U504 (N_504,In_993,In_663);
nand U505 (N_505,In_414,In_270);
nor U506 (N_506,In_350,In_679);
and U507 (N_507,In_787,In_937);
nand U508 (N_508,In_512,In_243);
nor U509 (N_509,In_947,In_669);
nand U510 (N_510,In_757,In_657);
and U511 (N_511,In_502,In_898);
nand U512 (N_512,In_14,In_411);
xor U513 (N_513,In_22,In_139);
and U514 (N_514,In_594,In_230);
nand U515 (N_515,In_820,In_220);
or U516 (N_516,In_920,In_922);
and U517 (N_517,In_666,In_884);
nand U518 (N_518,In_534,In_567);
nor U519 (N_519,In_296,In_563);
nor U520 (N_520,In_673,In_945);
or U521 (N_521,In_373,In_760);
nand U522 (N_522,In_21,In_875);
xnor U523 (N_523,In_901,In_581);
and U524 (N_524,In_450,In_303);
nor U525 (N_525,In_262,In_326);
xor U526 (N_526,In_683,In_978);
xor U527 (N_527,In_898,In_370);
or U528 (N_528,In_272,In_687);
and U529 (N_529,In_627,In_440);
nand U530 (N_530,In_735,In_96);
and U531 (N_531,In_246,In_77);
and U532 (N_532,In_215,In_237);
nand U533 (N_533,In_747,In_294);
and U534 (N_534,In_903,In_731);
nor U535 (N_535,In_997,In_470);
or U536 (N_536,In_155,In_582);
nor U537 (N_537,In_668,In_388);
nor U538 (N_538,In_7,In_282);
xnor U539 (N_539,In_763,In_402);
nor U540 (N_540,In_60,In_440);
and U541 (N_541,In_749,In_496);
xnor U542 (N_542,In_109,In_617);
and U543 (N_543,In_630,In_801);
nand U544 (N_544,In_188,In_814);
and U545 (N_545,In_609,In_513);
or U546 (N_546,In_918,In_395);
and U547 (N_547,In_573,In_833);
nor U548 (N_548,In_433,In_661);
nand U549 (N_549,In_306,In_210);
and U550 (N_550,In_226,In_95);
nand U551 (N_551,In_109,In_544);
xnor U552 (N_552,In_736,In_135);
nand U553 (N_553,In_23,In_956);
xor U554 (N_554,In_30,In_828);
xor U555 (N_555,In_552,In_631);
nor U556 (N_556,In_174,In_687);
or U557 (N_557,In_288,In_591);
xor U558 (N_558,In_650,In_826);
nand U559 (N_559,In_701,In_234);
or U560 (N_560,In_735,In_644);
nor U561 (N_561,In_503,In_864);
or U562 (N_562,In_640,In_807);
nor U563 (N_563,In_365,In_933);
and U564 (N_564,In_834,In_297);
xnor U565 (N_565,In_127,In_33);
and U566 (N_566,In_564,In_290);
nand U567 (N_567,In_733,In_202);
and U568 (N_568,In_600,In_658);
nor U569 (N_569,In_152,In_332);
and U570 (N_570,In_542,In_613);
and U571 (N_571,In_12,In_415);
nand U572 (N_572,In_864,In_751);
nor U573 (N_573,In_216,In_233);
nand U574 (N_574,In_320,In_835);
nor U575 (N_575,In_345,In_45);
or U576 (N_576,In_869,In_652);
xnor U577 (N_577,In_166,In_758);
nor U578 (N_578,In_115,In_355);
nand U579 (N_579,In_289,In_119);
nor U580 (N_580,In_772,In_267);
nand U581 (N_581,In_474,In_510);
nand U582 (N_582,In_975,In_30);
and U583 (N_583,In_258,In_382);
nand U584 (N_584,In_168,In_730);
nor U585 (N_585,In_8,In_941);
nor U586 (N_586,In_300,In_276);
or U587 (N_587,In_23,In_437);
nand U588 (N_588,In_494,In_886);
xnor U589 (N_589,In_230,In_768);
nand U590 (N_590,In_376,In_293);
nor U591 (N_591,In_318,In_615);
and U592 (N_592,In_780,In_285);
or U593 (N_593,In_143,In_300);
nand U594 (N_594,In_740,In_568);
xor U595 (N_595,In_818,In_107);
and U596 (N_596,In_820,In_320);
or U597 (N_597,In_871,In_98);
nand U598 (N_598,In_192,In_639);
or U599 (N_599,In_447,In_300);
xnor U600 (N_600,In_522,In_751);
and U601 (N_601,In_323,In_646);
nor U602 (N_602,In_654,In_319);
nand U603 (N_603,In_943,In_386);
nor U604 (N_604,In_760,In_134);
or U605 (N_605,In_647,In_279);
and U606 (N_606,In_786,In_974);
and U607 (N_607,In_533,In_704);
nand U608 (N_608,In_273,In_45);
nor U609 (N_609,In_544,In_477);
or U610 (N_610,In_340,In_679);
nand U611 (N_611,In_619,In_277);
xor U612 (N_612,In_341,In_770);
or U613 (N_613,In_470,In_509);
and U614 (N_614,In_202,In_765);
and U615 (N_615,In_783,In_819);
or U616 (N_616,In_21,In_929);
nand U617 (N_617,In_915,In_538);
and U618 (N_618,In_121,In_794);
and U619 (N_619,In_834,In_73);
or U620 (N_620,In_200,In_301);
nor U621 (N_621,In_209,In_296);
and U622 (N_622,In_999,In_64);
or U623 (N_623,In_326,In_676);
nor U624 (N_624,In_691,In_788);
and U625 (N_625,In_479,In_730);
and U626 (N_626,In_646,In_743);
nand U627 (N_627,In_316,In_658);
and U628 (N_628,In_518,In_127);
nor U629 (N_629,In_374,In_567);
and U630 (N_630,In_758,In_40);
nand U631 (N_631,In_460,In_748);
and U632 (N_632,In_355,In_908);
nor U633 (N_633,In_833,In_144);
nor U634 (N_634,In_569,In_257);
nor U635 (N_635,In_925,In_361);
and U636 (N_636,In_983,In_666);
nor U637 (N_637,In_882,In_142);
or U638 (N_638,In_264,In_334);
nor U639 (N_639,In_739,In_495);
nor U640 (N_640,In_333,In_922);
and U641 (N_641,In_191,In_407);
nand U642 (N_642,In_228,In_326);
nor U643 (N_643,In_612,In_439);
and U644 (N_644,In_332,In_591);
xor U645 (N_645,In_71,In_865);
and U646 (N_646,In_104,In_77);
nor U647 (N_647,In_628,In_444);
or U648 (N_648,In_977,In_392);
nand U649 (N_649,In_523,In_813);
or U650 (N_650,In_465,In_991);
or U651 (N_651,In_648,In_226);
nor U652 (N_652,In_308,In_277);
xnor U653 (N_653,In_460,In_450);
nand U654 (N_654,In_403,In_222);
and U655 (N_655,In_668,In_116);
nand U656 (N_656,In_946,In_242);
or U657 (N_657,In_5,In_600);
or U658 (N_658,In_762,In_93);
or U659 (N_659,In_188,In_628);
or U660 (N_660,In_937,In_264);
nor U661 (N_661,In_51,In_669);
and U662 (N_662,In_383,In_107);
or U663 (N_663,In_988,In_964);
and U664 (N_664,In_95,In_654);
nor U665 (N_665,In_903,In_44);
nand U666 (N_666,In_949,In_377);
nand U667 (N_667,In_874,In_148);
nand U668 (N_668,In_373,In_101);
nor U669 (N_669,In_212,In_557);
xor U670 (N_670,In_728,In_818);
nor U671 (N_671,In_179,In_27);
and U672 (N_672,In_221,In_600);
nand U673 (N_673,In_325,In_761);
nor U674 (N_674,In_953,In_350);
or U675 (N_675,In_811,In_842);
nor U676 (N_676,In_82,In_317);
and U677 (N_677,In_686,In_755);
and U678 (N_678,In_89,In_608);
or U679 (N_679,In_9,In_353);
nand U680 (N_680,In_101,In_562);
xor U681 (N_681,In_700,In_433);
nand U682 (N_682,In_778,In_495);
and U683 (N_683,In_374,In_313);
nor U684 (N_684,In_581,In_595);
nor U685 (N_685,In_963,In_243);
nor U686 (N_686,In_215,In_57);
or U687 (N_687,In_893,In_803);
nor U688 (N_688,In_382,In_348);
nand U689 (N_689,In_948,In_191);
xnor U690 (N_690,In_711,In_19);
and U691 (N_691,In_364,In_211);
xor U692 (N_692,In_278,In_285);
nand U693 (N_693,In_658,In_769);
nand U694 (N_694,In_772,In_15);
or U695 (N_695,In_882,In_120);
nand U696 (N_696,In_677,In_623);
xor U697 (N_697,In_780,In_743);
nor U698 (N_698,In_159,In_747);
and U699 (N_699,In_51,In_238);
or U700 (N_700,In_472,In_484);
and U701 (N_701,In_966,In_265);
or U702 (N_702,In_845,In_594);
or U703 (N_703,In_208,In_40);
or U704 (N_704,In_849,In_531);
xor U705 (N_705,In_770,In_663);
nor U706 (N_706,In_399,In_616);
or U707 (N_707,In_356,In_38);
or U708 (N_708,In_672,In_440);
or U709 (N_709,In_765,In_127);
or U710 (N_710,In_21,In_690);
and U711 (N_711,In_416,In_422);
nor U712 (N_712,In_592,In_171);
nor U713 (N_713,In_65,In_957);
or U714 (N_714,In_99,In_337);
or U715 (N_715,In_869,In_821);
nand U716 (N_716,In_863,In_281);
nor U717 (N_717,In_968,In_768);
and U718 (N_718,In_137,In_270);
or U719 (N_719,In_972,In_679);
nor U720 (N_720,In_960,In_6);
or U721 (N_721,In_895,In_460);
xnor U722 (N_722,In_656,In_949);
nor U723 (N_723,In_93,In_405);
and U724 (N_724,In_835,In_258);
nand U725 (N_725,In_877,In_48);
nor U726 (N_726,In_335,In_902);
and U727 (N_727,In_989,In_551);
and U728 (N_728,In_192,In_598);
and U729 (N_729,In_902,In_170);
nor U730 (N_730,In_945,In_656);
nor U731 (N_731,In_956,In_721);
nand U732 (N_732,In_137,In_0);
nor U733 (N_733,In_942,In_888);
nand U734 (N_734,In_477,In_438);
nor U735 (N_735,In_283,In_830);
nand U736 (N_736,In_432,In_428);
or U737 (N_737,In_756,In_425);
or U738 (N_738,In_727,In_617);
xnor U739 (N_739,In_790,In_417);
and U740 (N_740,In_781,In_235);
and U741 (N_741,In_228,In_931);
nor U742 (N_742,In_787,In_165);
nand U743 (N_743,In_443,In_347);
xor U744 (N_744,In_25,In_317);
and U745 (N_745,In_743,In_416);
nor U746 (N_746,In_512,In_690);
and U747 (N_747,In_582,In_825);
or U748 (N_748,In_699,In_708);
and U749 (N_749,In_530,In_996);
and U750 (N_750,In_85,In_450);
xor U751 (N_751,In_496,In_451);
and U752 (N_752,In_896,In_960);
and U753 (N_753,In_254,In_953);
nor U754 (N_754,In_89,In_822);
nand U755 (N_755,In_863,In_937);
and U756 (N_756,In_94,In_732);
or U757 (N_757,In_732,In_610);
nor U758 (N_758,In_682,In_520);
nor U759 (N_759,In_725,In_728);
xnor U760 (N_760,In_202,In_978);
nand U761 (N_761,In_3,In_998);
or U762 (N_762,In_606,In_427);
or U763 (N_763,In_492,In_807);
xnor U764 (N_764,In_936,In_930);
xor U765 (N_765,In_347,In_658);
and U766 (N_766,In_730,In_676);
or U767 (N_767,In_863,In_737);
and U768 (N_768,In_698,In_862);
nand U769 (N_769,In_655,In_462);
nand U770 (N_770,In_193,In_387);
and U771 (N_771,In_390,In_288);
nand U772 (N_772,In_755,In_620);
nand U773 (N_773,In_240,In_377);
nand U774 (N_774,In_713,In_806);
nor U775 (N_775,In_467,In_680);
nor U776 (N_776,In_576,In_108);
or U777 (N_777,In_991,In_883);
and U778 (N_778,In_106,In_459);
nand U779 (N_779,In_641,In_554);
and U780 (N_780,In_516,In_794);
nor U781 (N_781,In_142,In_780);
nor U782 (N_782,In_534,In_873);
and U783 (N_783,In_421,In_600);
or U784 (N_784,In_405,In_802);
nand U785 (N_785,In_316,In_43);
or U786 (N_786,In_484,In_284);
or U787 (N_787,In_418,In_509);
or U788 (N_788,In_740,In_537);
or U789 (N_789,In_914,In_549);
and U790 (N_790,In_237,In_678);
nor U791 (N_791,In_899,In_337);
nor U792 (N_792,In_263,In_594);
and U793 (N_793,In_544,In_332);
nand U794 (N_794,In_973,In_487);
or U795 (N_795,In_123,In_182);
or U796 (N_796,In_135,In_69);
and U797 (N_797,In_497,In_174);
nor U798 (N_798,In_619,In_341);
or U799 (N_799,In_470,In_736);
nand U800 (N_800,In_895,In_157);
nand U801 (N_801,In_318,In_134);
nor U802 (N_802,In_594,In_555);
and U803 (N_803,In_257,In_560);
nor U804 (N_804,In_581,In_470);
nor U805 (N_805,In_253,In_371);
nor U806 (N_806,In_596,In_692);
and U807 (N_807,In_517,In_384);
or U808 (N_808,In_692,In_434);
or U809 (N_809,In_181,In_316);
xor U810 (N_810,In_836,In_975);
nor U811 (N_811,In_475,In_677);
nand U812 (N_812,In_207,In_774);
nand U813 (N_813,In_826,In_358);
and U814 (N_814,In_305,In_237);
and U815 (N_815,In_184,In_531);
nand U816 (N_816,In_751,In_796);
nor U817 (N_817,In_33,In_535);
or U818 (N_818,In_801,In_994);
nand U819 (N_819,In_784,In_428);
nor U820 (N_820,In_942,In_622);
or U821 (N_821,In_502,In_777);
xor U822 (N_822,In_54,In_676);
and U823 (N_823,In_635,In_174);
and U824 (N_824,In_389,In_458);
nand U825 (N_825,In_990,In_624);
and U826 (N_826,In_301,In_146);
nor U827 (N_827,In_524,In_715);
nand U828 (N_828,In_447,In_264);
and U829 (N_829,In_864,In_625);
nand U830 (N_830,In_317,In_566);
or U831 (N_831,In_161,In_349);
xor U832 (N_832,In_491,In_707);
xnor U833 (N_833,In_592,In_288);
and U834 (N_834,In_930,In_67);
nor U835 (N_835,In_172,In_608);
nand U836 (N_836,In_952,In_319);
or U837 (N_837,In_149,In_45);
nand U838 (N_838,In_501,In_80);
and U839 (N_839,In_945,In_506);
nor U840 (N_840,In_531,In_328);
xnor U841 (N_841,In_728,In_982);
and U842 (N_842,In_312,In_682);
or U843 (N_843,In_781,In_906);
nand U844 (N_844,In_679,In_659);
nand U845 (N_845,In_548,In_940);
nand U846 (N_846,In_348,In_64);
nor U847 (N_847,In_112,In_272);
and U848 (N_848,In_235,In_109);
nand U849 (N_849,In_871,In_419);
nor U850 (N_850,In_842,In_564);
and U851 (N_851,In_473,In_467);
or U852 (N_852,In_779,In_65);
or U853 (N_853,In_377,In_159);
and U854 (N_854,In_292,In_53);
and U855 (N_855,In_267,In_32);
nor U856 (N_856,In_893,In_179);
or U857 (N_857,In_893,In_972);
nor U858 (N_858,In_333,In_441);
or U859 (N_859,In_737,In_807);
or U860 (N_860,In_563,In_547);
xnor U861 (N_861,In_804,In_481);
nor U862 (N_862,In_263,In_230);
or U863 (N_863,In_773,In_964);
or U864 (N_864,In_494,In_701);
and U865 (N_865,In_517,In_888);
nor U866 (N_866,In_192,In_700);
nor U867 (N_867,In_18,In_877);
and U868 (N_868,In_237,In_528);
or U869 (N_869,In_20,In_928);
nor U870 (N_870,In_599,In_305);
nor U871 (N_871,In_281,In_598);
or U872 (N_872,In_786,In_260);
nor U873 (N_873,In_402,In_516);
xnor U874 (N_874,In_72,In_50);
and U875 (N_875,In_740,In_583);
nand U876 (N_876,In_993,In_415);
nand U877 (N_877,In_917,In_688);
nand U878 (N_878,In_683,In_35);
nand U879 (N_879,In_440,In_521);
nor U880 (N_880,In_857,In_69);
nor U881 (N_881,In_67,In_467);
or U882 (N_882,In_815,In_973);
nand U883 (N_883,In_117,In_572);
or U884 (N_884,In_355,In_913);
nor U885 (N_885,In_178,In_868);
or U886 (N_886,In_985,In_784);
and U887 (N_887,In_672,In_283);
nand U888 (N_888,In_823,In_632);
or U889 (N_889,In_935,In_394);
and U890 (N_890,In_257,In_492);
xnor U891 (N_891,In_998,In_704);
nor U892 (N_892,In_969,In_552);
and U893 (N_893,In_437,In_775);
xor U894 (N_894,In_681,In_548);
nand U895 (N_895,In_749,In_601);
nand U896 (N_896,In_543,In_653);
or U897 (N_897,In_424,In_618);
nand U898 (N_898,In_21,In_724);
nor U899 (N_899,In_367,In_446);
or U900 (N_900,In_25,In_806);
nand U901 (N_901,In_429,In_365);
nand U902 (N_902,In_875,In_417);
or U903 (N_903,In_158,In_925);
nand U904 (N_904,In_327,In_808);
or U905 (N_905,In_637,In_154);
or U906 (N_906,In_332,In_616);
nand U907 (N_907,In_891,In_232);
nor U908 (N_908,In_421,In_408);
nor U909 (N_909,In_517,In_220);
nand U910 (N_910,In_802,In_145);
xor U911 (N_911,In_402,In_932);
nand U912 (N_912,In_655,In_912);
nand U913 (N_913,In_232,In_215);
or U914 (N_914,In_743,In_98);
nand U915 (N_915,In_281,In_687);
nor U916 (N_916,In_183,In_884);
and U917 (N_917,In_335,In_580);
and U918 (N_918,In_100,In_739);
and U919 (N_919,In_864,In_11);
nor U920 (N_920,In_691,In_100);
nor U921 (N_921,In_789,In_525);
nand U922 (N_922,In_67,In_358);
nand U923 (N_923,In_969,In_860);
nor U924 (N_924,In_291,In_228);
nand U925 (N_925,In_725,In_587);
nand U926 (N_926,In_194,In_366);
nor U927 (N_927,In_383,In_930);
or U928 (N_928,In_377,In_958);
nand U929 (N_929,In_642,In_553);
nor U930 (N_930,In_295,In_360);
nand U931 (N_931,In_155,In_324);
and U932 (N_932,In_826,In_870);
nor U933 (N_933,In_255,In_411);
xor U934 (N_934,In_679,In_475);
nor U935 (N_935,In_165,In_702);
or U936 (N_936,In_572,In_345);
or U937 (N_937,In_906,In_74);
or U938 (N_938,In_814,In_542);
nor U939 (N_939,In_894,In_542);
nor U940 (N_940,In_32,In_296);
and U941 (N_941,In_839,In_20);
nor U942 (N_942,In_564,In_879);
and U943 (N_943,In_352,In_612);
and U944 (N_944,In_15,In_850);
or U945 (N_945,In_91,In_901);
nand U946 (N_946,In_417,In_869);
or U947 (N_947,In_473,In_823);
or U948 (N_948,In_370,In_323);
or U949 (N_949,In_122,In_678);
or U950 (N_950,In_788,In_225);
or U951 (N_951,In_307,In_537);
nand U952 (N_952,In_858,In_515);
nor U953 (N_953,In_740,In_193);
and U954 (N_954,In_257,In_245);
and U955 (N_955,In_730,In_84);
and U956 (N_956,In_601,In_504);
nor U957 (N_957,In_774,In_173);
nand U958 (N_958,In_861,In_136);
or U959 (N_959,In_672,In_144);
nor U960 (N_960,In_714,In_653);
nor U961 (N_961,In_448,In_898);
and U962 (N_962,In_207,In_553);
or U963 (N_963,In_493,In_611);
and U964 (N_964,In_682,In_821);
and U965 (N_965,In_726,In_98);
nand U966 (N_966,In_171,In_716);
and U967 (N_967,In_641,In_38);
xor U968 (N_968,In_878,In_363);
nand U969 (N_969,In_905,In_645);
or U970 (N_970,In_828,In_138);
and U971 (N_971,In_875,In_737);
and U972 (N_972,In_502,In_738);
or U973 (N_973,In_366,In_234);
or U974 (N_974,In_132,In_613);
xor U975 (N_975,In_642,In_220);
or U976 (N_976,In_743,In_323);
and U977 (N_977,In_930,In_120);
nor U978 (N_978,In_104,In_328);
nor U979 (N_979,In_719,In_449);
nor U980 (N_980,In_474,In_385);
xor U981 (N_981,In_620,In_253);
xnor U982 (N_982,In_285,In_934);
nor U983 (N_983,In_631,In_255);
and U984 (N_984,In_476,In_589);
nand U985 (N_985,In_989,In_683);
nand U986 (N_986,In_342,In_324);
or U987 (N_987,In_254,In_205);
and U988 (N_988,In_570,In_872);
nor U989 (N_989,In_400,In_267);
xnor U990 (N_990,In_792,In_898);
or U991 (N_991,In_786,In_213);
or U992 (N_992,In_22,In_836);
nor U993 (N_993,In_237,In_947);
and U994 (N_994,In_380,In_870);
nor U995 (N_995,In_813,In_264);
or U996 (N_996,In_759,In_117);
and U997 (N_997,In_865,In_613);
nor U998 (N_998,In_445,In_510);
and U999 (N_999,In_326,In_511);
or U1000 (N_1000,In_305,In_184);
and U1001 (N_1001,In_629,In_858);
or U1002 (N_1002,In_78,In_598);
or U1003 (N_1003,In_865,In_479);
and U1004 (N_1004,In_858,In_632);
nor U1005 (N_1005,In_429,In_519);
nand U1006 (N_1006,In_670,In_68);
nor U1007 (N_1007,In_236,In_581);
or U1008 (N_1008,In_669,In_696);
nor U1009 (N_1009,In_800,In_792);
nor U1010 (N_1010,In_106,In_491);
nor U1011 (N_1011,In_582,In_446);
and U1012 (N_1012,In_706,In_238);
or U1013 (N_1013,In_467,In_888);
xnor U1014 (N_1014,In_187,In_185);
nor U1015 (N_1015,In_115,In_256);
or U1016 (N_1016,In_220,In_781);
and U1017 (N_1017,In_108,In_291);
nand U1018 (N_1018,In_319,In_786);
nand U1019 (N_1019,In_19,In_950);
nand U1020 (N_1020,In_81,In_58);
xnor U1021 (N_1021,In_422,In_120);
nand U1022 (N_1022,In_771,In_817);
xor U1023 (N_1023,In_455,In_666);
nor U1024 (N_1024,In_868,In_81);
nor U1025 (N_1025,In_711,In_303);
and U1026 (N_1026,In_276,In_349);
or U1027 (N_1027,In_284,In_914);
nand U1028 (N_1028,In_489,In_518);
nand U1029 (N_1029,In_225,In_984);
or U1030 (N_1030,In_824,In_234);
or U1031 (N_1031,In_943,In_812);
xnor U1032 (N_1032,In_851,In_696);
nand U1033 (N_1033,In_494,In_242);
nand U1034 (N_1034,In_465,In_546);
xnor U1035 (N_1035,In_600,In_601);
or U1036 (N_1036,In_281,In_798);
nor U1037 (N_1037,In_39,In_868);
nor U1038 (N_1038,In_15,In_172);
nand U1039 (N_1039,In_655,In_137);
nor U1040 (N_1040,In_881,In_216);
and U1041 (N_1041,In_289,In_954);
nor U1042 (N_1042,In_977,In_891);
and U1043 (N_1043,In_228,In_667);
and U1044 (N_1044,In_543,In_394);
nor U1045 (N_1045,In_255,In_529);
xnor U1046 (N_1046,In_603,In_45);
nand U1047 (N_1047,In_340,In_389);
nand U1048 (N_1048,In_300,In_637);
and U1049 (N_1049,In_690,In_601);
or U1050 (N_1050,In_345,In_651);
nand U1051 (N_1051,In_596,In_817);
xnor U1052 (N_1052,In_607,In_272);
xor U1053 (N_1053,In_804,In_139);
and U1054 (N_1054,In_544,In_206);
or U1055 (N_1055,In_47,In_459);
nand U1056 (N_1056,In_999,In_183);
nand U1057 (N_1057,In_730,In_65);
nand U1058 (N_1058,In_536,In_313);
xnor U1059 (N_1059,In_577,In_163);
xor U1060 (N_1060,In_788,In_922);
or U1061 (N_1061,In_167,In_372);
or U1062 (N_1062,In_213,In_403);
or U1063 (N_1063,In_278,In_766);
and U1064 (N_1064,In_68,In_32);
and U1065 (N_1065,In_901,In_123);
and U1066 (N_1066,In_852,In_991);
nor U1067 (N_1067,In_618,In_469);
nand U1068 (N_1068,In_414,In_975);
and U1069 (N_1069,In_153,In_87);
and U1070 (N_1070,In_277,In_524);
xor U1071 (N_1071,In_244,In_8);
or U1072 (N_1072,In_491,In_506);
xnor U1073 (N_1073,In_174,In_265);
nor U1074 (N_1074,In_570,In_323);
nor U1075 (N_1075,In_403,In_538);
nor U1076 (N_1076,In_944,In_137);
and U1077 (N_1077,In_503,In_562);
nand U1078 (N_1078,In_324,In_343);
and U1079 (N_1079,In_219,In_105);
nor U1080 (N_1080,In_57,In_209);
nor U1081 (N_1081,In_322,In_199);
and U1082 (N_1082,In_290,In_430);
and U1083 (N_1083,In_139,In_870);
nor U1084 (N_1084,In_33,In_415);
or U1085 (N_1085,In_514,In_246);
nand U1086 (N_1086,In_54,In_485);
xnor U1087 (N_1087,In_151,In_834);
and U1088 (N_1088,In_404,In_453);
nor U1089 (N_1089,In_643,In_787);
or U1090 (N_1090,In_974,In_719);
nor U1091 (N_1091,In_617,In_107);
nor U1092 (N_1092,In_383,In_111);
nand U1093 (N_1093,In_336,In_476);
nand U1094 (N_1094,In_982,In_76);
nand U1095 (N_1095,In_150,In_723);
or U1096 (N_1096,In_861,In_463);
xor U1097 (N_1097,In_434,In_395);
nor U1098 (N_1098,In_834,In_827);
and U1099 (N_1099,In_589,In_543);
nor U1100 (N_1100,In_172,In_607);
xnor U1101 (N_1101,In_508,In_859);
nand U1102 (N_1102,In_641,In_106);
and U1103 (N_1103,In_673,In_541);
or U1104 (N_1104,In_374,In_505);
and U1105 (N_1105,In_820,In_680);
and U1106 (N_1106,In_297,In_703);
or U1107 (N_1107,In_692,In_632);
or U1108 (N_1108,In_387,In_777);
or U1109 (N_1109,In_663,In_261);
and U1110 (N_1110,In_682,In_145);
and U1111 (N_1111,In_19,In_94);
and U1112 (N_1112,In_506,In_19);
and U1113 (N_1113,In_774,In_416);
and U1114 (N_1114,In_553,In_758);
nor U1115 (N_1115,In_737,In_695);
nor U1116 (N_1116,In_662,In_672);
nor U1117 (N_1117,In_849,In_425);
nor U1118 (N_1118,In_846,In_913);
or U1119 (N_1119,In_413,In_584);
or U1120 (N_1120,In_276,In_529);
and U1121 (N_1121,In_625,In_841);
or U1122 (N_1122,In_81,In_963);
nand U1123 (N_1123,In_682,In_562);
or U1124 (N_1124,In_391,In_610);
and U1125 (N_1125,In_920,In_444);
or U1126 (N_1126,In_545,In_543);
or U1127 (N_1127,In_36,In_993);
nand U1128 (N_1128,In_867,In_210);
and U1129 (N_1129,In_801,In_490);
and U1130 (N_1130,In_958,In_774);
xor U1131 (N_1131,In_18,In_405);
and U1132 (N_1132,In_187,In_152);
nand U1133 (N_1133,In_75,In_314);
nor U1134 (N_1134,In_548,In_942);
nor U1135 (N_1135,In_931,In_831);
or U1136 (N_1136,In_787,In_897);
nand U1137 (N_1137,In_935,In_752);
xor U1138 (N_1138,In_771,In_996);
xnor U1139 (N_1139,In_677,In_846);
and U1140 (N_1140,In_613,In_939);
nor U1141 (N_1141,In_749,In_879);
or U1142 (N_1142,In_245,In_217);
xor U1143 (N_1143,In_92,In_577);
xor U1144 (N_1144,In_853,In_106);
xor U1145 (N_1145,In_977,In_401);
nor U1146 (N_1146,In_4,In_52);
nor U1147 (N_1147,In_884,In_711);
and U1148 (N_1148,In_579,In_239);
nor U1149 (N_1149,In_18,In_633);
or U1150 (N_1150,In_105,In_802);
or U1151 (N_1151,In_940,In_276);
nand U1152 (N_1152,In_723,In_988);
or U1153 (N_1153,In_562,In_749);
xor U1154 (N_1154,In_335,In_597);
and U1155 (N_1155,In_520,In_459);
or U1156 (N_1156,In_923,In_598);
nand U1157 (N_1157,In_217,In_16);
or U1158 (N_1158,In_811,In_642);
nor U1159 (N_1159,In_757,In_323);
and U1160 (N_1160,In_967,In_957);
nand U1161 (N_1161,In_484,In_801);
nand U1162 (N_1162,In_786,In_376);
nor U1163 (N_1163,In_64,In_645);
xnor U1164 (N_1164,In_555,In_879);
or U1165 (N_1165,In_963,In_866);
and U1166 (N_1166,In_792,In_777);
or U1167 (N_1167,In_307,In_282);
and U1168 (N_1168,In_396,In_573);
nor U1169 (N_1169,In_783,In_581);
and U1170 (N_1170,In_836,In_587);
nor U1171 (N_1171,In_552,In_851);
xor U1172 (N_1172,In_297,In_702);
nand U1173 (N_1173,In_878,In_253);
and U1174 (N_1174,In_275,In_222);
or U1175 (N_1175,In_671,In_96);
nor U1176 (N_1176,In_834,In_513);
xnor U1177 (N_1177,In_758,In_678);
nand U1178 (N_1178,In_624,In_60);
xnor U1179 (N_1179,In_496,In_272);
nor U1180 (N_1180,In_689,In_552);
or U1181 (N_1181,In_100,In_723);
or U1182 (N_1182,In_93,In_508);
or U1183 (N_1183,In_473,In_273);
nand U1184 (N_1184,In_741,In_489);
nor U1185 (N_1185,In_375,In_68);
nand U1186 (N_1186,In_408,In_487);
nor U1187 (N_1187,In_965,In_223);
nor U1188 (N_1188,In_279,In_209);
nand U1189 (N_1189,In_193,In_912);
nand U1190 (N_1190,In_697,In_320);
nor U1191 (N_1191,In_626,In_929);
or U1192 (N_1192,In_248,In_784);
xor U1193 (N_1193,In_131,In_912);
nand U1194 (N_1194,In_217,In_37);
nand U1195 (N_1195,In_431,In_973);
nand U1196 (N_1196,In_744,In_284);
and U1197 (N_1197,In_663,In_957);
nand U1198 (N_1198,In_259,In_640);
or U1199 (N_1199,In_60,In_47);
nand U1200 (N_1200,In_113,In_112);
nand U1201 (N_1201,In_699,In_662);
and U1202 (N_1202,In_92,In_207);
xor U1203 (N_1203,In_449,In_595);
nor U1204 (N_1204,In_350,In_370);
xor U1205 (N_1205,In_104,In_682);
nand U1206 (N_1206,In_842,In_304);
xor U1207 (N_1207,In_151,In_558);
and U1208 (N_1208,In_48,In_902);
and U1209 (N_1209,In_73,In_150);
nor U1210 (N_1210,In_278,In_833);
and U1211 (N_1211,In_936,In_931);
or U1212 (N_1212,In_155,In_245);
and U1213 (N_1213,In_966,In_276);
nor U1214 (N_1214,In_889,In_588);
xnor U1215 (N_1215,In_824,In_215);
nand U1216 (N_1216,In_114,In_699);
or U1217 (N_1217,In_629,In_420);
nand U1218 (N_1218,In_77,In_352);
nor U1219 (N_1219,In_153,In_575);
and U1220 (N_1220,In_637,In_964);
nor U1221 (N_1221,In_430,In_551);
nor U1222 (N_1222,In_153,In_984);
xor U1223 (N_1223,In_117,In_112);
or U1224 (N_1224,In_610,In_31);
or U1225 (N_1225,In_579,In_92);
xnor U1226 (N_1226,In_628,In_503);
or U1227 (N_1227,In_459,In_680);
or U1228 (N_1228,In_776,In_613);
nor U1229 (N_1229,In_714,In_253);
xnor U1230 (N_1230,In_491,In_748);
or U1231 (N_1231,In_682,In_908);
or U1232 (N_1232,In_270,In_7);
or U1233 (N_1233,In_15,In_314);
xor U1234 (N_1234,In_245,In_428);
or U1235 (N_1235,In_839,In_560);
or U1236 (N_1236,In_850,In_135);
or U1237 (N_1237,In_750,In_580);
or U1238 (N_1238,In_161,In_776);
and U1239 (N_1239,In_64,In_436);
and U1240 (N_1240,In_126,In_199);
nor U1241 (N_1241,In_436,In_804);
or U1242 (N_1242,In_479,In_375);
nand U1243 (N_1243,In_277,In_197);
and U1244 (N_1244,In_821,In_928);
nand U1245 (N_1245,In_434,In_732);
nand U1246 (N_1246,In_812,In_947);
nand U1247 (N_1247,In_577,In_558);
nor U1248 (N_1248,In_600,In_886);
and U1249 (N_1249,In_698,In_596);
nor U1250 (N_1250,In_320,In_876);
or U1251 (N_1251,In_253,In_534);
or U1252 (N_1252,In_308,In_682);
nor U1253 (N_1253,In_290,In_674);
nor U1254 (N_1254,In_694,In_887);
nand U1255 (N_1255,In_689,In_908);
and U1256 (N_1256,In_631,In_606);
and U1257 (N_1257,In_685,In_968);
nor U1258 (N_1258,In_727,In_473);
nand U1259 (N_1259,In_665,In_907);
and U1260 (N_1260,In_987,In_443);
xor U1261 (N_1261,In_830,In_34);
nor U1262 (N_1262,In_753,In_797);
nor U1263 (N_1263,In_123,In_663);
nand U1264 (N_1264,In_468,In_331);
or U1265 (N_1265,In_162,In_934);
and U1266 (N_1266,In_494,In_802);
xor U1267 (N_1267,In_395,In_563);
nor U1268 (N_1268,In_916,In_926);
and U1269 (N_1269,In_43,In_562);
nor U1270 (N_1270,In_635,In_966);
or U1271 (N_1271,In_110,In_658);
or U1272 (N_1272,In_957,In_886);
and U1273 (N_1273,In_970,In_241);
nor U1274 (N_1274,In_233,In_101);
and U1275 (N_1275,In_680,In_733);
nand U1276 (N_1276,In_25,In_769);
nand U1277 (N_1277,In_628,In_617);
or U1278 (N_1278,In_549,In_590);
nor U1279 (N_1279,In_130,In_777);
or U1280 (N_1280,In_846,In_226);
xnor U1281 (N_1281,In_643,In_715);
nand U1282 (N_1282,In_472,In_462);
and U1283 (N_1283,In_150,In_384);
nor U1284 (N_1284,In_30,In_190);
xnor U1285 (N_1285,In_789,In_886);
and U1286 (N_1286,In_946,In_858);
and U1287 (N_1287,In_141,In_119);
xnor U1288 (N_1288,In_714,In_246);
and U1289 (N_1289,In_474,In_773);
xor U1290 (N_1290,In_68,In_317);
and U1291 (N_1291,In_781,In_178);
nand U1292 (N_1292,In_558,In_792);
nor U1293 (N_1293,In_684,In_986);
nor U1294 (N_1294,In_340,In_622);
or U1295 (N_1295,In_909,In_326);
xor U1296 (N_1296,In_812,In_836);
or U1297 (N_1297,In_568,In_97);
and U1298 (N_1298,In_626,In_605);
and U1299 (N_1299,In_528,In_958);
nand U1300 (N_1300,In_675,In_829);
nor U1301 (N_1301,In_797,In_854);
or U1302 (N_1302,In_46,In_332);
or U1303 (N_1303,In_369,In_26);
and U1304 (N_1304,In_234,In_542);
and U1305 (N_1305,In_502,In_91);
or U1306 (N_1306,In_430,In_690);
or U1307 (N_1307,In_34,In_229);
and U1308 (N_1308,In_776,In_387);
nor U1309 (N_1309,In_496,In_49);
and U1310 (N_1310,In_574,In_565);
nand U1311 (N_1311,In_993,In_234);
or U1312 (N_1312,In_297,In_283);
and U1313 (N_1313,In_985,In_888);
nor U1314 (N_1314,In_57,In_659);
and U1315 (N_1315,In_737,In_450);
nand U1316 (N_1316,In_436,In_681);
xnor U1317 (N_1317,In_749,In_271);
nor U1318 (N_1318,In_67,In_263);
and U1319 (N_1319,In_302,In_515);
and U1320 (N_1320,In_402,In_969);
nor U1321 (N_1321,In_784,In_33);
nor U1322 (N_1322,In_175,In_851);
nor U1323 (N_1323,In_705,In_506);
or U1324 (N_1324,In_471,In_791);
xor U1325 (N_1325,In_470,In_514);
and U1326 (N_1326,In_71,In_649);
xnor U1327 (N_1327,In_538,In_95);
nor U1328 (N_1328,In_103,In_652);
nor U1329 (N_1329,In_115,In_897);
or U1330 (N_1330,In_141,In_803);
or U1331 (N_1331,In_162,In_125);
nor U1332 (N_1332,In_696,In_346);
and U1333 (N_1333,In_399,In_187);
nand U1334 (N_1334,In_74,In_606);
or U1335 (N_1335,In_173,In_935);
or U1336 (N_1336,In_400,In_414);
or U1337 (N_1337,In_707,In_201);
and U1338 (N_1338,In_672,In_348);
nand U1339 (N_1339,In_340,In_381);
nand U1340 (N_1340,In_789,In_952);
and U1341 (N_1341,In_710,In_765);
or U1342 (N_1342,In_801,In_745);
or U1343 (N_1343,In_41,In_732);
nor U1344 (N_1344,In_745,In_608);
and U1345 (N_1345,In_457,In_977);
xor U1346 (N_1346,In_592,In_724);
nor U1347 (N_1347,In_386,In_895);
and U1348 (N_1348,In_196,In_823);
xnor U1349 (N_1349,In_124,In_667);
xor U1350 (N_1350,In_503,In_423);
nor U1351 (N_1351,In_610,In_125);
nand U1352 (N_1352,In_295,In_458);
or U1353 (N_1353,In_277,In_125);
and U1354 (N_1354,In_268,In_354);
and U1355 (N_1355,In_946,In_819);
xor U1356 (N_1356,In_100,In_825);
nand U1357 (N_1357,In_480,In_127);
nor U1358 (N_1358,In_561,In_837);
and U1359 (N_1359,In_303,In_517);
nand U1360 (N_1360,In_541,In_580);
or U1361 (N_1361,In_374,In_174);
or U1362 (N_1362,In_634,In_159);
or U1363 (N_1363,In_517,In_457);
and U1364 (N_1364,In_0,In_494);
and U1365 (N_1365,In_775,In_155);
nor U1366 (N_1366,In_791,In_982);
or U1367 (N_1367,In_448,In_644);
xnor U1368 (N_1368,In_837,In_92);
and U1369 (N_1369,In_53,In_609);
nand U1370 (N_1370,In_902,In_320);
nor U1371 (N_1371,In_440,In_928);
or U1372 (N_1372,In_50,In_447);
nor U1373 (N_1373,In_425,In_258);
nor U1374 (N_1374,In_883,In_648);
xnor U1375 (N_1375,In_941,In_142);
nor U1376 (N_1376,In_320,In_172);
nor U1377 (N_1377,In_294,In_112);
nand U1378 (N_1378,In_440,In_626);
or U1379 (N_1379,In_799,In_577);
nor U1380 (N_1380,In_391,In_741);
nand U1381 (N_1381,In_52,In_446);
or U1382 (N_1382,In_968,In_973);
nand U1383 (N_1383,In_799,In_511);
nand U1384 (N_1384,In_198,In_683);
or U1385 (N_1385,In_490,In_279);
nor U1386 (N_1386,In_663,In_766);
xor U1387 (N_1387,In_638,In_117);
nor U1388 (N_1388,In_950,In_697);
nor U1389 (N_1389,In_170,In_622);
or U1390 (N_1390,In_270,In_762);
and U1391 (N_1391,In_864,In_2);
or U1392 (N_1392,In_844,In_343);
and U1393 (N_1393,In_753,In_735);
nor U1394 (N_1394,In_8,In_669);
nand U1395 (N_1395,In_275,In_605);
or U1396 (N_1396,In_389,In_554);
or U1397 (N_1397,In_773,In_311);
nor U1398 (N_1398,In_701,In_138);
or U1399 (N_1399,In_27,In_25);
and U1400 (N_1400,In_247,In_522);
and U1401 (N_1401,In_987,In_4);
and U1402 (N_1402,In_990,In_506);
nand U1403 (N_1403,In_842,In_915);
nor U1404 (N_1404,In_667,In_484);
nand U1405 (N_1405,In_848,In_903);
nand U1406 (N_1406,In_434,In_842);
nor U1407 (N_1407,In_713,In_964);
nand U1408 (N_1408,In_206,In_205);
and U1409 (N_1409,In_899,In_1);
xnor U1410 (N_1410,In_477,In_497);
and U1411 (N_1411,In_666,In_132);
or U1412 (N_1412,In_654,In_30);
or U1413 (N_1413,In_279,In_627);
or U1414 (N_1414,In_970,In_704);
or U1415 (N_1415,In_824,In_403);
or U1416 (N_1416,In_256,In_208);
and U1417 (N_1417,In_172,In_209);
nor U1418 (N_1418,In_505,In_335);
or U1419 (N_1419,In_697,In_337);
nor U1420 (N_1420,In_849,In_356);
xnor U1421 (N_1421,In_235,In_428);
nand U1422 (N_1422,In_319,In_334);
and U1423 (N_1423,In_993,In_137);
or U1424 (N_1424,In_937,In_580);
and U1425 (N_1425,In_157,In_112);
nand U1426 (N_1426,In_585,In_388);
xor U1427 (N_1427,In_923,In_858);
nand U1428 (N_1428,In_720,In_195);
and U1429 (N_1429,In_29,In_356);
nor U1430 (N_1430,In_360,In_109);
and U1431 (N_1431,In_621,In_594);
nor U1432 (N_1432,In_589,In_692);
nor U1433 (N_1433,In_545,In_656);
xor U1434 (N_1434,In_40,In_858);
and U1435 (N_1435,In_50,In_707);
and U1436 (N_1436,In_953,In_593);
nor U1437 (N_1437,In_257,In_700);
xnor U1438 (N_1438,In_440,In_574);
and U1439 (N_1439,In_820,In_869);
nand U1440 (N_1440,In_964,In_736);
nor U1441 (N_1441,In_190,In_257);
or U1442 (N_1442,In_649,In_542);
or U1443 (N_1443,In_724,In_805);
nand U1444 (N_1444,In_281,In_302);
and U1445 (N_1445,In_551,In_642);
or U1446 (N_1446,In_696,In_293);
nand U1447 (N_1447,In_342,In_112);
and U1448 (N_1448,In_844,In_213);
nand U1449 (N_1449,In_531,In_863);
or U1450 (N_1450,In_642,In_450);
and U1451 (N_1451,In_161,In_184);
nand U1452 (N_1452,In_262,In_750);
nand U1453 (N_1453,In_377,In_472);
nand U1454 (N_1454,In_46,In_976);
and U1455 (N_1455,In_171,In_918);
and U1456 (N_1456,In_28,In_281);
and U1457 (N_1457,In_33,In_794);
xnor U1458 (N_1458,In_625,In_867);
nor U1459 (N_1459,In_902,In_846);
nor U1460 (N_1460,In_864,In_203);
nor U1461 (N_1461,In_703,In_66);
or U1462 (N_1462,In_198,In_516);
nor U1463 (N_1463,In_225,In_0);
or U1464 (N_1464,In_882,In_865);
and U1465 (N_1465,In_861,In_864);
nor U1466 (N_1466,In_755,In_391);
nand U1467 (N_1467,In_429,In_3);
nor U1468 (N_1468,In_225,In_412);
or U1469 (N_1469,In_280,In_888);
and U1470 (N_1470,In_798,In_337);
or U1471 (N_1471,In_311,In_604);
and U1472 (N_1472,In_270,In_476);
nor U1473 (N_1473,In_257,In_449);
nand U1474 (N_1474,In_45,In_164);
and U1475 (N_1475,In_314,In_272);
or U1476 (N_1476,In_474,In_209);
or U1477 (N_1477,In_76,In_934);
and U1478 (N_1478,In_246,In_556);
and U1479 (N_1479,In_424,In_194);
nor U1480 (N_1480,In_123,In_155);
or U1481 (N_1481,In_227,In_861);
nor U1482 (N_1482,In_162,In_267);
nor U1483 (N_1483,In_197,In_588);
and U1484 (N_1484,In_966,In_621);
xor U1485 (N_1485,In_901,In_833);
and U1486 (N_1486,In_426,In_620);
or U1487 (N_1487,In_867,In_873);
nor U1488 (N_1488,In_85,In_673);
nand U1489 (N_1489,In_827,In_328);
and U1490 (N_1490,In_218,In_207);
or U1491 (N_1491,In_391,In_961);
nor U1492 (N_1492,In_913,In_299);
and U1493 (N_1493,In_196,In_768);
or U1494 (N_1494,In_183,In_312);
xnor U1495 (N_1495,In_994,In_977);
and U1496 (N_1496,In_518,In_530);
nand U1497 (N_1497,In_761,In_677);
or U1498 (N_1498,In_156,In_436);
nor U1499 (N_1499,In_162,In_221);
nand U1500 (N_1500,In_330,In_126);
or U1501 (N_1501,In_317,In_552);
and U1502 (N_1502,In_102,In_134);
nor U1503 (N_1503,In_661,In_897);
and U1504 (N_1504,In_655,In_333);
or U1505 (N_1505,In_314,In_644);
xor U1506 (N_1506,In_243,In_932);
nand U1507 (N_1507,In_784,In_915);
nor U1508 (N_1508,In_518,In_803);
and U1509 (N_1509,In_534,In_577);
nand U1510 (N_1510,In_471,In_611);
and U1511 (N_1511,In_587,In_813);
and U1512 (N_1512,In_986,In_647);
nor U1513 (N_1513,In_28,In_952);
xor U1514 (N_1514,In_236,In_198);
and U1515 (N_1515,In_748,In_395);
and U1516 (N_1516,In_347,In_185);
and U1517 (N_1517,In_540,In_19);
or U1518 (N_1518,In_698,In_827);
or U1519 (N_1519,In_241,In_250);
and U1520 (N_1520,In_336,In_641);
nor U1521 (N_1521,In_334,In_737);
and U1522 (N_1522,In_867,In_870);
nor U1523 (N_1523,In_151,In_411);
xor U1524 (N_1524,In_548,In_747);
or U1525 (N_1525,In_292,In_626);
or U1526 (N_1526,In_264,In_290);
and U1527 (N_1527,In_4,In_586);
and U1528 (N_1528,In_338,In_673);
or U1529 (N_1529,In_335,In_616);
and U1530 (N_1530,In_270,In_860);
nor U1531 (N_1531,In_962,In_43);
nand U1532 (N_1532,In_17,In_108);
nand U1533 (N_1533,In_787,In_120);
and U1534 (N_1534,In_851,In_172);
nand U1535 (N_1535,In_769,In_100);
nand U1536 (N_1536,In_141,In_94);
nor U1537 (N_1537,In_309,In_943);
or U1538 (N_1538,In_549,In_995);
and U1539 (N_1539,In_799,In_395);
nor U1540 (N_1540,In_897,In_256);
nand U1541 (N_1541,In_600,In_488);
and U1542 (N_1542,In_472,In_436);
nand U1543 (N_1543,In_651,In_890);
and U1544 (N_1544,In_4,In_231);
and U1545 (N_1545,In_640,In_597);
and U1546 (N_1546,In_715,In_178);
nand U1547 (N_1547,In_713,In_912);
or U1548 (N_1548,In_527,In_379);
nand U1549 (N_1549,In_912,In_456);
nor U1550 (N_1550,In_587,In_811);
xnor U1551 (N_1551,In_578,In_713);
nand U1552 (N_1552,In_823,In_22);
nor U1553 (N_1553,In_532,In_427);
xnor U1554 (N_1554,In_453,In_342);
and U1555 (N_1555,In_584,In_193);
nand U1556 (N_1556,In_918,In_826);
nor U1557 (N_1557,In_176,In_685);
xnor U1558 (N_1558,In_643,In_745);
or U1559 (N_1559,In_343,In_712);
nor U1560 (N_1560,In_615,In_345);
and U1561 (N_1561,In_263,In_482);
nand U1562 (N_1562,In_666,In_470);
nand U1563 (N_1563,In_651,In_351);
xor U1564 (N_1564,In_286,In_768);
xnor U1565 (N_1565,In_550,In_859);
and U1566 (N_1566,In_351,In_934);
xor U1567 (N_1567,In_415,In_763);
and U1568 (N_1568,In_444,In_969);
xnor U1569 (N_1569,In_884,In_988);
nor U1570 (N_1570,In_559,In_878);
xnor U1571 (N_1571,In_463,In_320);
nand U1572 (N_1572,In_686,In_377);
nand U1573 (N_1573,In_216,In_777);
or U1574 (N_1574,In_74,In_212);
nand U1575 (N_1575,In_183,In_745);
nand U1576 (N_1576,In_758,In_724);
and U1577 (N_1577,In_328,In_489);
or U1578 (N_1578,In_832,In_776);
nand U1579 (N_1579,In_740,In_223);
or U1580 (N_1580,In_447,In_51);
nand U1581 (N_1581,In_909,In_199);
and U1582 (N_1582,In_23,In_88);
or U1583 (N_1583,In_42,In_296);
nand U1584 (N_1584,In_842,In_548);
nor U1585 (N_1585,In_886,In_161);
nand U1586 (N_1586,In_291,In_616);
nor U1587 (N_1587,In_600,In_743);
or U1588 (N_1588,In_14,In_206);
nor U1589 (N_1589,In_749,In_839);
or U1590 (N_1590,In_895,In_757);
xor U1591 (N_1591,In_760,In_578);
and U1592 (N_1592,In_336,In_102);
nand U1593 (N_1593,In_433,In_889);
xnor U1594 (N_1594,In_569,In_343);
nor U1595 (N_1595,In_289,In_297);
nor U1596 (N_1596,In_450,In_495);
or U1597 (N_1597,In_839,In_247);
xor U1598 (N_1598,In_800,In_493);
nor U1599 (N_1599,In_26,In_482);
xor U1600 (N_1600,In_469,In_461);
nand U1601 (N_1601,In_418,In_158);
nor U1602 (N_1602,In_569,In_55);
or U1603 (N_1603,In_179,In_634);
and U1604 (N_1604,In_994,In_854);
xnor U1605 (N_1605,In_832,In_709);
nand U1606 (N_1606,In_106,In_644);
xnor U1607 (N_1607,In_819,In_461);
and U1608 (N_1608,In_168,In_299);
and U1609 (N_1609,In_725,In_849);
xnor U1610 (N_1610,In_431,In_80);
nand U1611 (N_1611,In_398,In_366);
or U1612 (N_1612,In_79,In_996);
or U1613 (N_1613,In_850,In_223);
nor U1614 (N_1614,In_93,In_675);
nand U1615 (N_1615,In_135,In_321);
nor U1616 (N_1616,In_804,In_2);
or U1617 (N_1617,In_76,In_344);
nand U1618 (N_1618,In_741,In_84);
nor U1619 (N_1619,In_676,In_85);
nor U1620 (N_1620,In_635,In_710);
and U1621 (N_1621,In_633,In_598);
and U1622 (N_1622,In_802,In_854);
or U1623 (N_1623,In_180,In_513);
or U1624 (N_1624,In_715,In_782);
nand U1625 (N_1625,In_311,In_914);
nand U1626 (N_1626,In_401,In_266);
nand U1627 (N_1627,In_64,In_717);
and U1628 (N_1628,In_553,In_613);
nor U1629 (N_1629,In_459,In_265);
xnor U1630 (N_1630,In_120,In_885);
nor U1631 (N_1631,In_350,In_545);
xor U1632 (N_1632,In_509,In_475);
nor U1633 (N_1633,In_120,In_897);
nor U1634 (N_1634,In_691,In_402);
nand U1635 (N_1635,In_466,In_370);
nor U1636 (N_1636,In_423,In_521);
nor U1637 (N_1637,In_46,In_251);
nor U1638 (N_1638,In_558,In_704);
and U1639 (N_1639,In_716,In_196);
nor U1640 (N_1640,In_206,In_422);
xor U1641 (N_1641,In_75,In_82);
and U1642 (N_1642,In_219,In_589);
or U1643 (N_1643,In_615,In_937);
and U1644 (N_1644,In_317,In_394);
nor U1645 (N_1645,In_142,In_731);
or U1646 (N_1646,In_872,In_187);
xnor U1647 (N_1647,In_390,In_74);
xor U1648 (N_1648,In_592,In_900);
nor U1649 (N_1649,In_654,In_432);
nand U1650 (N_1650,In_715,In_621);
xnor U1651 (N_1651,In_507,In_495);
nand U1652 (N_1652,In_244,In_608);
nand U1653 (N_1653,In_633,In_730);
nand U1654 (N_1654,In_97,In_221);
or U1655 (N_1655,In_305,In_744);
xnor U1656 (N_1656,In_0,In_457);
xnor U1657 (N_1657,In_459,In_941);
or U1658 (N_1658,In_871,In_91);
and U1659 (N_1659,In_618,In_83);
nor U1660 (N_1660,In_185,In_734);
nand U1661 (N_1661,In_320,In_360);
xor U1662 (N_1662,In_279,In_289);
or U1663 (N_1663,In_454,In_598);
nand U1664 (N_1664,In_49,In_859);
or U1665 (N_1665,In_752,In_339);
and U1666 (N_1666,In_922,In_783);
or U1667 (N_1667,In_429,In_167);
nor U1668 (N_1668,In_935,In_226);
and U1669 (N_1669,In_783,In_190);
nand U1670 (N_1670,In_702,In_43);
and U1671 (N_1671,In_316,In_775);
or U1672 (N_1672,In_930,In_273);
nor U1673 (N_1673,In_346,In_12);
xor U1674 (N_1674,In_332,In_513);
nor U1675 (N_1675,In_707,In_673);
and U1676 (N_1676,In_87,In_180);
nand U1677 (N_1677,In_610,In_718);
xnor U1678 (N_1678,In_371,In_133);
nor U1679 (N_1679,In_344,In_302);
or U1680 (N_1680,In_549,In_374);
nor U1681 (N_1681,In_656,In_797);
nor U1682 (N_1682,In_951,In_813);
and U1683 (N_1683,In_539,In_338);
nor U1684 (N_1684,In_216,In_463);
nor U1685 (N_1685,In_6,In_293);
or U1686 (N_1686,In_8,In_975);
and U1687 (N_1687,In_31,In_892);
xnor U1688 (N_1688,In_972,In_312);
and U1689 (N_1689,In_264,In_203);
nand U1690 (N_1690,In_902,In_563);
and U1691 (N_1691,In_507,In_16);
xnor U1692 (N_1692,In_763,In_105);
or U1693 (N_1693,In_190,In_996);
or U1694 (N_1694,In_274,In_958);
or U1695 (N_1695,In_837,In_175);
nor U1696 (N_1696,In_888,In_959);
or U1697 (N_1697,In_535,In_791);
and U1698 (N_1698,In_270,In_858);
nor U1699 (N_1699,In_61,In_879);
and U1700 (N_1700,In_126,In_749);
xnor U1701 (N_1701,In_427,In_46);
nor U1702 (N_1702,In_34,In_98);
xor U1703 (N_1703,In_505,In_53);
and U1704 (N_1704,In_211,In_978);
nor U1705 (N_1705,In_954,In_814);
nand U1706 (N_1706,In_157,In_24);
nor U1707 (N_1707,In_226,In_10);
or U1708 (N_1708,In_895,In_337);
nand U1709 (N_1709,In_995,In_373);
or U1710 (N_1710,In_327,In_293);
nor U1711 (N_1711,In_78,In_929);
nor U1712 (N_1712,In_636,In_166);
and U1713 (N_1713,In_724,In_306);
or U1714 (N_1714,In_472,In_973);
and U1715 (N_1715,In_794,In_340);
nand U1716 (N_1716,In_109,In_364);
and U1717 (N_1717,In_378,In_925);
and U1718 (N_1718,In_786,In_160);
nor U1719 (N_1719,In_71,In_736);
and U1720 (N_1720,In_159,In_666);
and U1721 (N_1721,In_142,In_444);
nand U1722 (N_1722,In_14,In_705);
or U1723 (N_1723,In_942,In_573);
and U1724 (N_1724,In_430,In_458);
xor U1725 (N_1725,In_279,In_373);
nor U1726 (N_1726,In_719,In_953);
nand U1727 (N_1727,In_448,In_181);
nand U1728 (N_1728,In_622,In_881);
nand U1729 (N_1729,In_316,In_879);
or U1730 (N_1730,In_169,In_572);
or U1731 (N_1731,In_365,In_559);
nor U1732 (N_1732,In_483,In_49);
and U1733 (N_1733,In_944,In_866);
or U1734 (N_1734,In_405,In_304);
and U1735 (N_1735,In_284,In_92);
nand U1736 (N_1736,In_35,In_787);
or U1737 (N_1737,In_329,In_621);
nor U1738 (N_1738,In_849,In_235);
xor U1739 (N_1739,In_815,In_929);
nand U1740 (N_1740,In_523,In_297);
nand U1741 (N_1741,In_64,In_7);
nand U1742 (N_1742,In_402,In_886);
and U1743 (N_1743,In_253,In_539);
nand U1744 (N_1744,In_367,In_586);
nand U1745 (N_1745,In_225,In_32);
or U1746 (N_1746,In_763,In_103);
and U1747 (N_1747,In_569,In_858);
nor U1748 (N_1748,In_534,In_203);
nand U1749 (N_1749,In_55,In_898);
xor U1750 (N_1750,In_205,In_456);
xor U1751 (N_1751,In_792,In_697);
nor U1752 (N_1752,In_881,In_625);
nor U1753 (N_1753,In_319,In_215);
nor U1754 (N_1754,In_947,In_953);
or U1755 (N_1755,In_308,In_305);
nor U1756 (N_1756,In_108,In_800);
or U1757 (N_1757,In_19,In_778);
xor U1758 (N_1758,In_105,In_9);
xnor U1759 (N_1759,In_175,In_863);
or U1760 (N_1760,In_361,In_32);
nand U1761 (N_1761,In_772,In_79);
xor U1762 (N_1762,In_727,In_720);
nand U1763 (N_1763,In_417,In_351);
nor U1764 (N_1764,In_224,In_161);
and U1765 (N_1765,In_613,In_107);
or U1766 (N_1766,In_637,In_884);
xnor U1767 (N_1767,In_136,In_455);
or U1768 (N_1768,In_212,In_151);
nor U1769 (N_1769,In_722,In_956);
and U1770 (N_1770,In_207,In_727);
nand U1771 (N_1771,In_981,In_809);
and U1772 (N_1772,In_427,In_360);
or U1773 (N_1773,In_807,In_652);
and U1774 (N_1774,In_558,In_965);
nand U1775 (N_1775,In_184,In_543);
or U1776 (N_1776,In_886,In_603);
xor U1777 (N_1777,In_11,In_835);
nand U1778 (N_1778,In_158,In_191);
nand U1779 (N_1779,In_358,In_596);
and U1780 (N_1780,In_81,In_832);
and U1781 (N_1781,In_243,In_631);
or U1782 (N_1782,In_166,In_723);
nor U1783 (N_1783,In_21,In_694);
or U1784 (N_1784,In_749,In_596);
xor U1785 (N_1785,In_378,In_598);
or U1786 (N_1786,In_378,In_894);
xor U1787 (N_1787,In_591,In_400);
and U1788 (N_1788,In_138,In_291);
nand U1789 (N_1789,In_849,In_726);
or U1790 (N_1790,In_262,In_140);
nand U1791 (N_1791,In_834,In_939);
nand U1792 (N_1792,In_30,In_782);
nor U1793 (N_1793,In_716,In_740);
nand U1794 (N_1794,In_704,In_778);
or U1795 (N_1795,In_774,In_468);
nand U1796 (N_1796,In_844,In_570);
or U1797 (N_1797,In_271,In_295);
and U1798 (N_1798,In_996,In_707);
nand U1799 (N_1799,In_58,In_532);
or U1800 (N_1800,In_61,In_863);
nor U1801 (N_1801,In_463,In_439);
or U1802 (N_1802,In_171,In_809);
and U1803 (N_1803,In_982,In_674);
xor U1804 (N_1804,In_219,In_740);
and U1805 (N_1805,In_47,In_253);
nor U1806 (N_1806,In_50,In_269);
nand U1807 (N_1807,In_739,In_367);
nand U1808 (N_1808,In_380,In_199);
and U1809 (N_1809,In_897,In_678);
nand U1810 (N_1810,In_327,In_587);
nor U1811 (N_1811,In_884,In_47);
xor U1812 (N_1812,In_431,In_886);
nand U1813 (N_1813,In_696,In_58);
and U1814 (N_1814,In_201,In_951);
and U1815 (N_1815,In_345,In_18);
nor U1816 (N_1816,In_294,In_167);
nand U1817 (N_1817,In_888,In_904);
and U1818 (N_1818,In_406,In_531);
nand U1819 (N_1819,In_124,In_373);
nor U1820 (N_1820,In_484,In_777);
xor U1821 (N_1821,In_292,In_570);
and U1822 (N_1822,In_412,In_636);
nand U1823 (N_1823,In_697,In_249);
nor U1824 (N_1824,In_590,In_781);
xor U1825 (N_1825,In_206,In_37);
xnor U1826 (N_1826,In_494,In_279);
and U1827 (N_1827,In_33,In_630);
or U1828 (N_1828,In_198,In_935);
or U1829 (N_1829,In_710,In_146);
and U1830 (N_1830,In_352,In_940);
and U1831 (N_1831,In_617,In_498);
or U1832 (N_1832,In_67,In_630);
nand U1833 (N_1833,In_359,In_784);
nand U1834 (N_1834,In_371,In_402);
nand U1835 (N_1835,In_829,In_678);
and U1836 (N_1836,In_395,In_849);
nand U1837 (N_1837,In_300,In_434);
nor U1838 (N_1838,In_732,In_741);
or U1839 (N_1839,In_403,In_717);
xnor U1840 (N_1840,In_328,In_915);
or U1841 (N_1841,In_560,In_466);
or U1842 (N_1842,In_220,In_398);
nand U1843 (N_1843,In_29,In_704);
or U1844 (N_1844,In_517,In_954);
nor U1845 (N_1845,In_894,In_332);
nand U1846 (N_1846,In_213,In_815);
nand U1847 (N_1847,In_439,In_291);
and U1848 (N_1848,In_51,In_636);
and U1849 (N_1849,In_708,In_813);
nand U1850 (N_1850,In_863,In_455);
xor U1851 (N_1851,In_818,In_622);
and U1852 (N_1852,In_563,In_821);
nor U1853 (N_1853,In_45,In_790);
nor U1854 (N_1854,In_683,In_27);
nand U1855 (N_1855,In_412,In_957);
nand U1856 (N_1856,In_506,In_70);
and U1857 (N_1857,In_229,In_139);
nand U1858 (N_1858,In_270,In_679);
or U1859 (N_1859,In_68,In_457);
nor U1860 (N_1860,In_433,In_342);
or U1861 (N_1861,In_295,In_128);
nor U1862 (N_1862,In_916,In_587);
and U1863 (N_1863,In_377,In_160);
nand U1864 (N_1864,In_389,In_830);
nor U1865 (N_1865,In_673,In_783);
or U1866 (N_1866,In_659,In_487);
nor U1867 (N_1867,In_982,In_649);
and U1868 (N_1868,In_388,In_486);
nand U1869 (N_1869,In_785,In_759);
and U1870 (N_1870,In_662,In_785);
or U1871 (N_1871,In_234,In_666);
nand U1872 (N_1872,In_657,In_512);
or U1873 (N_1873,In_238,In_137);
nor U1874 (N_1874,In_153,In_942);
or U1875 (N_1875,In_66,In_841);
and U1876 (N_1876,In_547,In_826);
or U1877 (N_1877,In_1,In_786);
xor U1878 (N_1878,In_746,In_69);
nand U1879 (N_1879,In_363,In_614);
and U1880 (N_1880,In_102,In_292);
nor U1881 (N_1881,In_720,In_104);
xor U1882 (N_1882,In_483,In_446);
or U1883 (N_1883,In_481,In_145);
or U1884 (N_1884,In_890,In_622);
and U1885 (N_1885,In_415,In_681);
nand U1886 (N_1886,In_845,In_914);
or U1887 (N_1887,In_961,In_259);
xor U1888 (N_1888,In_205,In_774);
nand U1889 (N_1889,In_419,In_633);
nand U1890 (N_1890,In_896,In_713);
and U1891 (N_1891,In_394,In_964);
and U1892 (N_1892,In_213,In_264);
nor U1893 (N_1893,In_644,In_574);
or U1894 (N_1894,In_975,In_434);
or U1895 (N_1895,In_637,In_861);
or U1896 (N_1896,In_922,In_227);
xor U1897 (N_1897,In_386,In_403);
or U1898 (N_1898,In_632,In_904);
or U1899 (N_1899,In_458,In_836);
or U1900 (N_1900,In_112,In_778);
or U1901 (N_1901,In_482,In_265);
nor U1902 (N_1902,In_190,In_674);
nand U1903 (N_1903,In_695,In_544);
xor U1904 (N_1904,In_834,In_414);
xnor U1905 (N_1905,In_264,In_970);
nand U1906 (N_1906,In_218,In_808);
or U1907 (N_1907,In_402,In_458);
and U1908 (N_1908,In_498,In_744);
or U1909 (N_1909,In_5,In_221);
nand U1910 (N_1910,In_805,In_116);
nand U1911 (N_1911,In_14,In_589);
or U1912 (N_1912,In_532,In_594);
or U1913 (N_1913,In_569,In_38);
nand U1914 (N_1914,In_881,In_400);
and U1915 (N_1915,In_317,In_877);
and U1916 (N_1916,In_688,In_818);
or U1917 (N_1917,In_870,In_351);
nor U1918 (N_1918,In_192,In_384);
or U1919 (N_1919,In_677,In_613);
nor U1920 (N_1920,In_56,In_655);
nand U1921 (N_1921,In_322,In_850);
nand U1922 (N_1922,In_303,In_938);
and U1923 (N_1923,In_429,In_615);
or U1924 (N_1924,In_244,In_319);
nand U1925 (N_1925,In_632,In_326);
nand U1926 (N_1926,In_146,In_757);
nor U1927 (N_1927,In_259,In_558);
nand U1928 (N_1928,In_575,In_931);
nor U1929 (N_1929,In_282,In_179);
nor U1930 (N_1930,In_555,In_324);
nand U1931 (N_1931,In_746,In_395);
and U1932 (N_1932,In_858,In_821);
or U1933 (N_1933,In_825,In_66);
nor U1934 (N_1934,In_763,In_347);
nand U1935 (N_1935,In_17,In_146);
and U1936 (N_1936,In_522,In_295);
or U1937 (N_1937,In_251,In_417);
and U1938 (N_1938,In_92,In_724);
nand U1939 (N_1939,In_617,In_50);
nor U1940 (N_1940,In_557,In_585);
and U1941 (N_1941,In_636,In_157);
nor U1942 (N_1942,In_728,In_930);
or U1943 (N_1943,In_811,In_679);
and U1944 (N_1944,In_209,In_146);
nand U1945 (N_1945,In_596,In_840);
nor U1946 (N_1946,In_316,In_450);
xor U1947 (N_1947,In_276,In_113);
nor U1948 (N_1948,In_916,In_501);
and U1949 (N_1949,In_91,In_900);
xor U1950 (N_1950,In_291,In_417);
and U1951 (N_1951,In_6,In_18);
or U1952 (N_1952,In_557,In_989);
and U1953 (N_1953,In_196,In_289);
nand U1954 (N_1954,In_698,In_732);
and U1955 (N_1955,In_7,In_279);
or U1956 (N_1956,In_767,In_112);
or U1957 (N_1957,In_583,In_512);
xor U1958 (N_1958,In_940,In_89);
nand U1959 (N_1959,In_700,In_526);
nor U1960 (N_1960,In_975,In_339);
nor U1961 (N_1961,In_168,In_230);
xor U1962 (N_1962,In_372,In_199);
or U1963 (N_1963,In_46,In_301);
nor U1964 (N_1964,In_858,In_345);
or U1965 (N_1965,In_812,In_261);
or U1966 (N_1966,In_290,In_539);
and U1967 (N_1967,In_794,In_380);
or U1968 (N_1968,In_113,In_209);
nor U1969 (N_1969,In_82,In_987);
or U1970 (N_1970,In_689,In_621);
nor U1971 (N_1971,In_625,In_222);
or U1972 (N_1972,In_636,In_21);
or U1973 (N_1973,In_555,In_73);
and U1974 (N_1974,In_948,In_550);
nand U1975 (N_1975,In_230,In_645);
nor U1976 (N_1976,In_571,In_446);
or U1977 (N_1977,In_884,In_615);
or U1978 (N_1978,In_5,In_932);
or U1979 (N_1979,In_725,In_654);
nand U1980 (N_1980,In_726,In_787);
nand U1981 (N_1981,In_265,In_199);
nor U1982 (N_1982,In_106,In_873);
nand U1983 (N_1983,In_396,In_37);
or U1984 (N_1984,In_29,In_80);
nand U1985 (N_1985,In_87,In_704);
or U1986 (N_1986,In_421,In_483);
or U1987 (N_1987,In_932,In_584);
or U1988 (N_1988,In_202,In_586);
or U1989 (N_1989,In_753,In_902);
nand U1990 (N_1990,In_364,In_3);
and U1991 (N_1991,In_394,In_527);
or U1992 (N_1992,In_589,In_450);
nor U1993 (N_1993,In_566,In_302);
xnor U1994 (N_1994,In_83,In_468);
xor U1995 (N_1995,In_350,In_536);
and U1996 (N_1996,In_373,In_833);
xor U1997 (N_1997,In_4,In_813);
and U1998 (N_1998,In_523,In_509);
or U1999 (N_1999,In_121,In_390);
or U2000 (N_2000,N_1282,N_1505);
nor U2001 (N_2001,N_870,N_1931);
and U2002 (N_2002,N_1059,N_1401);
xor U2003 (N_2003,N_790,N_1810);
nand U2004 (N_2004,N_1247,N_1574);
or U2005 (N_2005,N_42,N_581);
nand U2006 (N_2006,N_1051,N_1591);
nand U2007 (N_2007,N_378,N_1891);
or U2008 (N_2008,N_31,N_148);
and U2009 (N_2009,N_24,N_1892);
or U2010 (N_2010,N_449,N_191);
nand U2011 (N_2011,N_1695,N_713);
nand U2012 (N_2012,N_642,N_891);
nor U2013 (N_2013,N_1728,N_1765);
nand U2014 (N_2014,N_1182,N_785);
or U2015 (N_2015,N_1467,N_569);
and U2016 (N_2016,N_1339,N_1229);
nor U2017 (N_2017,N_533,N_528);
or U2018 (N_2018,N_927,N_1409);
xor U2019 (N_2019,N_1763,N_56);
or U2020 (N_2020,N_621,N_1469);
or U2021 (N_2021,N_956,N_821);
or U2022 (N_2022,N_1704,N_206);
nor U2023 (N_2023,N_1048,N_1329);
nand U2024 (N_2024,N_249,N_1534);
and U2025 (N_2025,N_1203,N_981);
nor U2026 (N_2026,N_1290,N_1402);
nand U2027 (N_2027,N_1159,N_273);
and U2028 (N_2028,N_407,N_1184);
or U2029 (N_2029,N_872,N_1672);
or U2030 (N_2030,N_1733,N_1817);
or U2031 (N_2031,N_1821,N_301);
nor U2032 (N_2032,N_1877,N_375);
nand U2033 (N_2033,N_1601,N_1418);
nand U2034 (N_2034,N_547,N_1355);
nand U2035 (N_2035,N_93,N_110);
and U2036 (N_2036,N_1894,N_1304);
nand U2037 (N_2037,N_550,N_1538);
or U2038 (N_2038,N_915,N_1648);
nor U2039 (N_2039,N_1364,N_117);
or U2040 (N_2040,N_1980,N_304);
nor U2041 (N_2041,N_539,N_1729);
nor U2042 (N_2042,N_950,N_668);
nor U2043 (N_2043,N_201,N_1326);
or U2044 (N_2044,N_32,N_1767);
nor U2045 (N_2045,N_1983,N_1450);
or U2046 (N_2046,N_59,N_1676);
nand U2047 (N_2047,N_438,N_847);
xor U2048 (N_2048,N_101,N_1639);
nor U2049 (N_2049,N_267,N_11);
and U2050 (N_2050,N_510,N_1793);
nor U2051 (N_2051,N_168,N_1617);
nor U2052 (N_2052,N_1598,N_1301);
nand U2053 (N_2053,N_1239,N_1558);
and U2054 (N_2054,N_1726,N_1270);
nand U2055 (N_2055,N_740,N_1794);
and U2056 (N_2056,N_819,N_1691);
xor U2057 (N_2057,N_1963,N_1047);
nor U2058 (N_2058,N_1531,N_1820);
nor U2059 (N_2059,N_1634,N_1619);
and U2060 (N_2060,N_1626,N_1719);
nand U2061 (N_2061,N_1010,N_8);
or U2062 (N_2062,N_1214,N_34);
nor U2063 (N_2063,N_1019,N_1008);
and U2064 (N_2064,N_905,N_1310);
and U2065 (N_2065,N_76,N_430);
nor U2066 (N_2066,N_1426,N_1782);
or U2067 (N_2067,N_925,N_685);
and U2068 (N_2068,N_823,N_262);
nand U2069 (N_2069,N_321,N_1692);
nand U2070 (N_2070,N_937,N_1910);
nand U2071 (N_2071,N_170,N_220);
xnor U2072 (N_2072,N_1572,N_1445);
and U2073 (N_2073,N_1712,N_254);
or U2074 (N_2074,N_1466,N_1515);
nand U2075 (N_2075,N_1775,N_627);
xnor U2076 (N_2076,N_1786,N_496);
and U2077 (N_2077,N_1623,N_1074);
and U2078 (N_2078,N_734,N_898);
nor U2079 (N_2079,N_1559,N_1707);
and U2080 (N_2080,N_1438,N_224);
and U2081 (N_2081,N_1528,N_291);
nor U2082 (N_2082,N_1783,N_43);
nor U2083 (N_2083,N_1813,N_39);
nor U2084 (N_2084,N_1705,N_1385);
nor U2085 (N_2085,N_238,N_638);
nor U2086 (N_2086,N_1237,N_1493);
or U2087 (N_2087,N_347,N_230);
and U2088 (N_2088,N_1555,N_1399);
nand U2089 (N_2089,N_312,N_839);
or U2090 (N_2090,N_1573,N_838);
or U2091 (N_2091,N_876,N_1193);
nand U2092 (N_2092,N_1388,N_279);
nand U2093 (N_2093,N_1777,N_520);
nor U2094 (N_2094,N_748,N_1302);
nand U2095 (N_2095,N_1348,N_830);
or U2096 (N_2096,N_145,N_1525);
nand U2097 (N_2097,N_1485,N_406);
and U2098 (N_2098,N_508,N_13);
and U2099 (N_2099,N_657,N_91);
xor U2100 (N_2100,N_530,N_473);
nor U2101 (N_2101,N_270,N_55);
and U2102 (N_2102,N_1678,N_1622);
and U2103 (N_2103,N_1213,N_402);
nor U2104 (N_2104,N_1742,N_1846);
and U2105 (N_2105,N_648,N_1442);
nor U2106 (N_2106,N_74,N_1296);
nor U2107 (N_2107,N_1447,N_65);
nand U2108 (N_2108,N_422,N_1834);
xnor U2109 (N_2109,N_1036,N_104);
and U2110 (N_2110,N_1333,N_1138);
nand U2111 (N_2111,N_672,N_1962);
or U2112 (N_2112,N_590,N_1003);
nand U2113 (N_2113,N_793,N_196);
nor U2114 (N_2114,N_240,N_909);
and U2115 (N_2115,N_243,N_1780);
or U2116 (N_2116,N_1123,N_666);
and U2117 (N_2117,N_1584,N_755);
nand U2118 (N_2118,N_150,N_1795);
nor U2119 (N_2119,N_1377,N_1608);
nor U2120 (N_2120,N_667,N_722);
xor U2121 (N_2121,N_883,N_1907);
and U2122 (N_2122,N_1413,N_1243);
or U2123 (N_2123,N_746,N_1909);
or U2124 (N_2124,N_255,N_1071);
nor U2125 (N_2125,N_1318,N_1057);
and U2126 (N_2126,N_182,N_1933);
nor U2127 (N_2127,N_1044,N_380);
nand U2128 (N_2128,N_1665,N_998);
nor U2129 (N_2129,N_1365,N_1112);
or U2130 (N_2130,N_322,N_1249);
nand U2131 (N_2131,N_1224,N_1353);
or U2132 (N_2132,N_779,N_505);
and U2133 (N_2133,N_1391,N_237);
or U2134 (N_2134,N_1700,N_678);
or U2135 (N_2135,N_922,N_565);
and U2136 (N_2136,N_741,N_857);
or U2137 (N_2137,N_22,N_163);
and U2138 (N_2138,N_176,N_419);
nor U2139 (N_2139,N_1839,N_1088);
and U2140 (N_2140,N_160,N_1972);
nand U2141 (N_2141,N_865,N_1679);
or U2142 (N_2142,N_733,N_1953);
nand U2143 (N_2143,N_271,N_427);
and U2144 (N_2144,N_608,N_357);
nor U2145 (N_2145,N_1336,N_641);
xor U2146 (N_2146,N_1058,N_417);
xor U2147 (N_2147,N_1052,N_335);
and U2148 (N_2148,N_1373,N_1993);
and U2149 (N_2149,N_828,N_1444);
and U2150 (N_2150,N_1487,N_868);
and U2151 (N_2151,N_63,N_374);
xor U2152 (N_2152,N_560,N_1830);
nor U2153 (N_2153,N_1702,N_1836);
nand U2154 (N_2154,N_1039,N_1424);
nand U2155 (N_2155,N_345,N_1108);
nor U2156 (N_2156,N_1870,N_78);
nor U2157 (N_2157,N_948,N_1666);
nor U2158 (N_2158,N_251,N_1197);
or U2159 (N_2159,N_578,N_1343);
and U2160 (N_2160,N_146,N_1151);
nor U2161 (N_2161,N_1616,N_1754);
nand U2162 (N_2162,N_1300,N_1292);
nand U2163 (N_2163,N_618,N_1107);
xnor U2164 (N_2164,N_1756,N_1271);
or U2165 (N_2165,N_226,N_1849);
or U2166 (N_2166,N_719,N_1536);
and U2167 (N_2167,N_1784,N_1285);
and U2168 (N_2168,N_1518,N_1737);
and U2169 (N_2169,N_193,N_650);
or U2170 (N_2170,N_1670,N_863);
or U2171 (N_2171,N_1699,N_624);
and U2172 (N_2172,N_323,N_1750);
xor U2173 (N_2173,N_390,N_124);
and U2174 (N_2174,N_1186,N_1211);
xor U2175 (N_2175,N_1319,N_120);
nand U2176 (N_2176,N_774,N_48);
nor U2177 (N_2177,N_1139,N_920);
or U2178 (N_2178,N_771,N_526);
and U2179 (N_2179,N_1183,N_1260);
nand U2180 (N_2180,N_1419,N_57);
nor U2181 (N_2181,N_1772,N_385);
or U2182 (N_2182,N_669,N_1740);
and U2183 (N_2183,N_366,N_1609);
or U2184 (N_2184,N_328,N_947);
or U2185 (N_2185,N_664,N_1092);
nand U2186 (N_2186,N_67,N_278);
nand U2187 (N_2187,N_1287,N_919);
and U2188 (N_2188,N_1994,N_944);
nand U2189 (N_2189,N_571,N_1252);
and U2190 (N_2190,N_645,N_1553);
nor U2191 (N_2191,N_1878,N_825);
nor U2192 (N_2192,N_171,N_404);
xor U2193 (N_2193,N_613,N_831);
nand U2194 (N_2194,N_1654,N_940);
nor U2195 (N_2195,N_1068,N_836);
and U2196 (N_2196,N_1232,N_619);
nor U2197 (N_2197,N_235,N_461);
xor U2198 (N_2198,N_1664,N_691);
nor U2199 (N_2199,N_568,N_1504);
and U2200 (N_2200,N_367,N_245);
xor U2201 (N_2201,N_714,N_1165);
or U2202 (N_2202,N_487,N_786);
and U2203 (N_2203,N_1317,N_396);
nor U2204 (N_2204,N_1513,N_344);
xor U2205 (N_2205,N_1884,N_1250);
nor U2206 (N_2206,N_1779,N_1567);
nor U2207 (N_2207,N_1338,N_1647);
or U2208 (N_2208,N_595,N_478);
or U2209 (N_2209,N_1768,N_1412);
nand U2210 (N_2210,N_83,N_1236);
nand U2211 (N_2211,N_739,N_178);
and U2212 (N_2212,N_1337,N_1129);
and U2213 (N_2213,N_356,N_504);
nand U2214 (N_2214,N_1991,N_695);
nand U2215 (N_2215,N_1792,N_1833);
or U2216 (N_2216,N_1625,N_1200);
nor U2217 (N_2217,N_125,N_1050);
or U2218 (N_2218,N_1741,N_1638);
or U2219 (N_2219,N_363,N_1462);
and U2220 (N_2220,N_1581,N_218);
nor U2221 (N_2221,N_319,N_141);
nor U2222 (N_2222,N_123,N_1630);
nor U2223 (N_2223,N_303,N_598);
and U2224 (N_2224,N_1807,N_269);
or U2225 (N_2225,N_1565,N_1069);
nor U2226 (N_2226,N_1172,N_896);
or U2227 (N_2227,N_309,N_1471);
xnor U2228 (N_2228,N_631,N_1913);
and U2229 (N_2229,N_1483,N_1307);
or U2230 (N_2230,N_346,N_1620);
and U2231 (N_2231,N_551,N_503);
or U2232 (N_2232,N_1605,N_759);
nand U2233 (N_2233,N_1421,N_1921);
or U2234 (N_2234,N_1761,N_706);
xor U2235 (N_2235,N_369,N_1356);
xor U2236 (N_2236,N_990,N_1441);
nor U2237 (N_2237,N_1005,N_1927);
nor U2238 (N_2238,N_1137,N_1788);
nand U2239 (N_2239,N_425,N_1323);
nor U2240 (N_2240,N_29,N_890);
and U2241 (N_2241,N_1420,N_559);
or U2242 (N_2242,N_377,N_189);
and U2243 (N_2243,N_250,N_21);
nand U2244 (N_2244,N_1669,N_928);
nor U2245 (N_2245,N_1856,N_1073);
and U2246 (N_2246,N_681,N_986);
or U2247 (N_2247,N_1109,N_953);
nor U2248 (N_2248,N_1130,N_874);
and U2249 (N_2249,N_1724,N_1818);
or U2250 (N_2250,N_263,N_1579);
and U2251 (N_2251,N_878,N_654);
xnor U2252 (N_2252,N_38,N_1956);
and U2253 (N_2253,N_1562,N_1860);
and U2254 (N_2254,N_1379,N_454);
or U2255 (N_2255,N_1357,N_1967);
xnor U2256 (N_2256,N_1597,N_995);
and U2257 (N_2257,N_1557,N_481);
nand U2258 (N_2258,N_597,N_310);
nor U2259 (N_2259,N_1110,N_1455);
xnor U2260 (N_2260,N_463,N_1998);
and U2261 (N_2261,N_579,N_1629);
and U2262 (N_2262,N_812,N_1481);
nor U2263 (N_2263,N_1014,N_517);
nor U2264 (N_2264,N_983,N_1946);
nand U2265 (N_2265,N_1906,N_128);
nor U2266 (N_2266,N_1033,N_1354);
nand U2267 (N_2267,N_1334,N_1407);
nor U2268 (N_2268,N_161,N_1847);
nor U2269 (N_2269,N_835,N_916);
nand U2270 (N_2270,N_829,N_1537);
or U2271 (N_2271,N_1519,N_386);
xor U2272 (N_2272,N_1686,N_745);
nor U2273 (N_2273,N_1066,N_147);
nand U2274 (N_2274,N_1376,N_929);
nand U2275 (N_2275,N_1857,N_1230);
and U2276 (N_2276,N_1613,N_105);
or U2277 (N_2277,N_127,N_381);
xnor U2278 (N_2278,N_1762,N_361);
and U2279 (N_2279,N_817,N_1038);
and U2280 (N_2280,N_116,N_429);
nand U2281 (N_2281,N_77,N_456);
nor U2282 (N_2282,N_1470,N_203);
or U2283 (N_2283,N_1217,N_1134);
and U2284 (N_2284,N_1098,N_211);
or U2285 (N_2285,N_867,N_1721);
or U2286 (N_2286,N_1627,N_1206);
and U2287 (N_2287,N_1231,N_1416);
and U2288 (N_2288,N_1945,N_999);
xnor U2289 (N_2289,N_1175,N_1263);
and U2290 (N_2290,N_783,N_1541);
and U2291 (N_2291,N_708,N_1486);
and U2292 (N_2292,N_736,N_442);
nor U2293 (N_2293,N_1935,N_1035);
nor U2294 (N_2294,N_181,N_16);
nor U2295 (N_2295,N_1293,N_1570);
nor U2296 (N_2296,N_1883,N_1411);
and U2297 (N_2297,N_985,N_1090);
nand U2298 (N_2298,N_1852,N_675);
and U2299 (N_2299,N_1361,N_1873);
and U2300 (N_2300,N_180,N_215);
and U2301 (N_2301,N_26,N_862);
nand U2302 (N_2302,N_1841,N_1031);
nor U2303 (N_2303,N_1636,N_100);
nand U2304 (N_2304,N_1291,N_1312);
nor U2305 (N_2305,N_801,N_605);
nor U2306 (N_2306,N_738,N_1898);
nand U2307 (N_2307,N_1022,N_1596);
and U2308 (N_2308,N_1164,N_721);
nor U2309 (N_2309,N_1615,N_1132);
and U2310 (N_2310,N_1770,N_207);
and U2311 (N_2311,N_900,N_292);
and U2312 (N_2312,N_90,N_1328);
nand U2313 (N_2313,N_1899,N_12);
xnor U2314 (N_2314,N_432,N_1716);
or U2315 (N_2315,N_1097,N_40);
or U2316 (N_2316,N_371,N_1053);
xnor U2317 (N_2317,N_644,N_1812);
nand U2318 (N_2318,N_1111,N_527);
or U2319 (N_2319,N_700,N_866);
or U2320 (N_2320,N_894,N_744);
nand U2321 (N_2321,N_1578,N_846);
nand U2322 (N_2322,N_917,N_754);
or U2323 (N_2323,N_295,N_389);
nand U2324 (N_2324,N_1947,N_280);
and U2325 (N_2325,N_1517,N_975);
nor U2326 (N_2326,N_99,N_1248);
and U2327 (N_2327,N_1785,N_1815);
nand U2328 (N_2328,N_532,N_1769);
and U2329 (N_2329,N_966,N_1589);
or U2330 (N_2330,N_911,N_852);
nor U2331 (N_2331,N_1932,N_564);
nand U2332 (N_2332,N_1173,N_987);
xor U2333 (N_2333,N_1673,N_247);
or U2334 (N_2334,N_1595,N_1226);
or U2335 (N_2335,N_459,N_694);
or U2336 (N_2336,N_431,N_1168);
xor U2337 (N_2337,N_239,N_534);
nand U2338 (N_2338,N_1734,N_317);
xor U2339 (N_2339,N_1844,N_1453);
nor U2340 (N_2340,N_364,N_1196);
nand U2341 (N_2341,N_573,N_1494);
nor U2342 (N_2342,N_1372,N_1922);
nand U2343 (N_2343,N_1273,N_484);
nor U2344 (N_2344,N_1276,N_1593);
xnor U2345 (N_2345,N_223,N_1222);
and U2346 (N_2346,N_1162,N_932);
nor U2347 (N_2347,N_1403,N_1332);
and U2348 (N_2348,N_167,N_490);
nor U2349 (N_2349,N_1408,N_1509);
nor U2350 (N_2350,N_1602,N_1103);
xnor U2351 (N_2351,N_633,N_1545);
and U2352 (N_2352,N_807,N_274);
nor U2353 (N_2353,N_1133,N_804);
and U2354 (N_2354,N_996,N_1662);
nor U2355 (N_2355,N_1244,N_913);
nand U2356 (N_2356,N_318,N_525);
nor U2357 (N_2357,N_227,N_1503);
nor U2358 (N_2358,N_1116,N_1124);
or U2359 (N_2359,N_717,N_643);
xnor U2360 (N_2360,N_1394,N_1392);
nand U2361 (N_2361,N_1422,N_516);
nand U2362 (N_2362,N_1136,N_80);
and U2363 (N_2363,N_462,N_1314);
nand U2364 (N_2364,N_955,N_540);
nor U2365 (N_2365,N_582,N_1127);
and U2366 (N_2366,N_1286,N_1521);
nor U2367 (N_2367,N_1923,N_1997);
or U2368 (N_2368,N_1649,N_1439);
xnor U2369 (N_2369,N_1027,N_1976);
or U2370 (N_2370,N_244,N_612);
xor U2371 (N_2371,N_6,N_1212);
or U2372 (N_2372,N_538,N_1245);
nor U2373 (N_2373,N_855,N_885);
nand U2374 (N_2374,N_475,N_546);
and U2375 (N_2375,N_690,N_1640);
and U2376 (N_2376,N_735,N_938);
nand U2377 (N_2377,N_1207,N_200);
or U2378 (N_2378,N_358,N_513);
or U2379 (N_2379,N_458,N_229);
nand U2380 (N_2380,N_1095,N_1984);
xor U2381 (N_2381,N_446,N_1903);
xnor U2382 (N_2382,N_777,N_136);
nand U2383 (N_2383,N_1979,N_1952);
nor U2384 (N_2384,N_555,N_709);
and U2385 (N_2385,N_455,N_1085);
or U2386 (N_2386,N_860,N_311);
nor U2387 (N_2387,N_594,N_626);
or U2388 (N_2388,N_1800,N_1738);
nor U2389 (N_2389,N_1524,N_1170);
nand U2390 (N_2390,N_584,N_1942);
nand U2391 (N_2391,N_1937,N_810);
nor U2392 (N_2392,N_1791,N_1614);
and U2393 (N_2393,N_1757,N_994);
or U2394 (N_2394,N_886,N_320);
or U2395 (N_2395,N_1826,N_1556);
nor U2396 (N_2396,N_1081,N_1653);
and U2397 (N_2397,N_172,N_984);
or U2398 (N_2398,N_1266,N_1056);
and U2399 (N_2399,N_854,N_1461);
nor U2400 (N_2400,N_96,N_73);
and U2401 (N_2401,N_285,N_1720);
or U2402 (N_2402,N_0,N_1167);
xor U2403 (N_2403,N_1020,N_253);
nand U2404 (N_2404,N_1215,N_1482);
nand U2405 (N_2405,N_1275,N_1703);
and U2406 (N_2406,N_325,N_1683);
nor U2407 (N_2407,N_1925,N_1034);
and U2408 (N_2408,N_166,N_1688);
and U2409 (N_2409,N_972,N_1280);
nor U2410 (N_2410,N_1369,N_33);
and U2411 (N_2411,N_187,N_660);
and U2412 (N_2412,N_699,N_1018);
nor U2413 (N_2413,N_712,N_1859);
or U2414 (N_2414,N_1100,N_766);
or U2415 (N_2415,N_1971,N_1837);
and U2416 (N_2416,N_416,N_1886);
nand U2417 (N_2417,N_762,N_1028);
or U2418 (N_2418,N_1701,N_188);
xnor U2419 (N_2419,N_365,N_1105);
nand U2420 (N_2420,N_1948,N_1660);
nor U2421 (N_2421,N_1759,N_1747);
nand U2422 (N_2422,N_1939,N_606);
nor U2423 (N_2423,N_1241,N_1397);
nand U2424 (N_2424,N_1201,N_1987);
nor U2425 (N_2425,N_493,N_842);
and U2426 (N_2426,N_770,N_1543);
or U2427 (N_2427,N_1753,N_1722);
or U2428 (N_2428,N_282,N_1764);
and U2429 (N_2429,N_1468,N_901);
nand U2430 (N_2430,N_499,N_1690);
nand U2431 (N_2431,N_199,N_1867);
nor U2432 (N_2432,N_337,N_1163);
nor U2433 (N_2433,N_742,N_281);
and U2434 (N_2434,N_1969,N_1571);
and U2435 (N_2435,N_1564,N_1457);
and U2436 (N_2436,N_97,N_1599);
nand U2437 (N_2437,N_287,N_1911);
nand U2438 (N_2438,N_1067,N_843);
nand U2439 (N_2439,N_617,N_382);
and U2440 (N_2440,N_1375,N_1350);
nor U2441 (N_2441,N_1324,N_28);
and U2442 (N_2442,N_570,N_1781);
and U2443 (N_2443,N_252,N_1806);
and U2444 (N_2444,N_302,N_683);
nand U2445 (N_2445,N_1309,N_1011);
nor U2446 (N_2446,N_701,N_1472);
and U2447 (N_2447,N_789,N_453);
and U2448 (N_2448,N_376,N_542);
nand U2449 (N_2449,N_1055,N_1588);
nor U2450 (N_2450,N_173,N_1996);
nor U2451 (N_2451,N_1363,N_236);
nor U2452 (N_2452,N_776,N_1644);
nand U2453 (N_2453,N_632,N_1508);
and U2454 (N_2454,N_1985,N_769);
or U2455 (N_2455,N_1154,N_1828);
or U2456 (N_2456,N_1208,N_1727);
and U2457 (N_2457,N_869,N_1089);
or U2458 (N_2458,N_307,N_543);
nand U2459 (N_2459,N_949,N_1436);
nand U2460 (N_2460,N_1776,N_368);
xnor U2461 (N_2461,N_297,N_1002);
nand U2462 (N_2462,N_17,N_306);
and U2463 (N_2463,N_1577,N_635);
nand U2464 (N_2464,N_1,N_715);
or U2465 (N_2465,N_859,N_408);
xnor U2466 (N_2466,N_511,N_1966);
xor U2467 (N_2467,N_1344,N_1443);
or U2468 (N_2468,N_1840,N_46);
nor U2469 (N_2469,N_1233,N_1065);
and U2470 (N_2470,N_609,N_1185);
nand U2471 (N_2471,N_1887,N_483);
nor U2472 (N_2472,N_492,N_1272);
nor U2473 (N_2473,N_435,N_294);
nor U2474 (N_2474,N_1009,N_348);
nand U2475 (N_2475,N_1115,N_1973);
nor U2476 (N_2476,N_1456,N_276);
nand U2477 (N_2477,N_818,N_512);
nand U2478 (N_2478,N_1851,N_1677);
xor U2479 (N_2479,N_1289,N_314);
and U2480 (N_2480,N_1934,N_1256);
nand U2481 (N_2481,N_775,N_1888);
nand U2482 (N_2482,N_1989,N_387);
or U2483 (N_2483,N_958,N_142);
nand U2484 (N_2484,N_327,N_1015);
and U2485 (N_2485,N_440,N_155);
nand U2486 (N_2486,N_1658,N_554);
and U2487 (N_2487,N_799,N_1084);
and U2488 (N_2488,N_1417,N_765);
and U2489 (N_2489,N_72,N_576);
nand U2490 (N_2490,N_509,N_1853);
nor U2491 (N_2491,N_135,N_602);
nand U2492 (N_2492,N_151,N_557);
nor U2493 (N_2493,N_198,N_433);
nand U2494 (N_2494,N_1507,N_840);
or U2495 (N_2495,N_305,N_1501);
nand U2496 (N_2496,N_1970,N_780);
or U2497 (N_2497,N_787,N_283);
or U2498 (N_2498,N_1893,N_1930);
and U2499 (N_2499,N_1778,N_1195);
or U2500 (N_2500,N_85,N_122);
and U2501 (N_2501,N_1001,N_1446);
nor U2502 (N_2502,N_1227,N_1798);
nor U2503 (N_2503,N_1079,N_60);
nor U2504 (N_2504,N_849,N_1140);
nand U2505 (N_2505,N_952,N_718);
or U2506 (N_2506,N_791,N_1264);
nor U2507 (N_2507,N_1076,N_284);
nor U2508 (N_2508,N_175,N_1495);
or U2509 (N_2509,N_1267,N_1492);
nand U2510 (N_2510,N_339,N_1816);
and U2511 (N_2511,N_1706,N_1992);
nor U2512 (N_2512,N_51,N_340);
and U2513 (N_2513,N_1671,N_1122);
and U2514 (N_2514,N_464,N_871);
nand U2515 (N_2515,N_1876,N_680);
nand U2516 (N_2516,N_333,N_1434);
nor U2517 (N_2517,N_164,N_1606);
or U2518 (N_2518,N_1862,N_1575);
nor U2519 (N_2519,N_1205,N_98);
and U2520 (N_2520,N_1512,N_805);
nand U2521 (N_2521,N_980,N_214);
xor U2522 (N_2522,N_231,N_9);
and U2523 (N_2523,N_1158,N_1773);
or U2524 (N_2524,N_684,N_1316);
nor U2525 (N_2525,N_1835,N_476);
and U2526 (N_2526,N_1030,N_1752);
and U2527 (N_2527,N_1179,N_1760);
or U2528 (N_2528,N_1101,N_697);
and U2529 (N_2529,N_1255,N_1362);
xnor U2530 (N_2530,N_964,N_313);
nand U2531 (N_2531,N_1281,N_1811);
nor U2532 (N_2532,N_1150,N_1511);
and U2533 (N_2533,N_501,N_903);
nand U2534 (N_2534,N_1396,N_822);
and U2535 (N_2535,N_845,N_257);
or U2536 (N_2536,N_1974,N_795);
xor U2537 (N_2537,N_912,N_585);
nor U2538 (N_2538,N_1335,N_1360);
xnor U2539 (N_2539,N_782,N_979);
nor U2540 (N_2540,N_784,N_809);
or U2541 (N_2541,N_1061,N_758);
and U2542 (N_2542,N_1113,N_138);
and U2543 (N_2543,N_655,N_1743);
nand U2544 (N_2544,N_904,N_1382);
nor U2545 (N_2545,N_359,N_1919);
xor U2546 (N_2546,N_592,N_1174);
nand U2547 (N_2547,N_1526,N_1060);
or U2548 (N_2548,N_1268,N_1072);
nor U2549 (N_2549,N_82,N_1687);
nor U2550 (N_2550,N_1410,N_1476);
and U2551 (N_2551,N_1554,N_1879);
or U2552 (N_2552,N_935,N_1221);
xor U2553 (N_2553,N_157,N_1610);
nand U2554 (N_2554,N_1094,N_974);
and U2555 (N_2555,N_1464,N_1460);
nor U2556 (N_2556,N_1012,N_58);
nand U2557 (N_2557,N_963,N_796);
and U2558 (N_2558,N_445,N_1083);
nand U2559 (N_2559,N_88,N_951);
nand U2560 (N_2560,N_66,N_1077);
nand U2561 (N_2561,N_1251,N_628);
xor U2562 (N_2562,N_1498,N_1550);
xnor U2563 (N_2563,N_190,N_1400);
or U2564 (N_2564,N_1656,N_1751);
and U2565 (N_2565,N_452,N_601);
nor U2566 (N_2566,N_27,N_556);
and U2567 (N_2567,N_811,N_130);
nand U2568 (N_2568,N_1126,N_1929);
nand U2569 (N_2569,N_1313,N_682);
and U2570 (N_2570,N_1961,N_1725);
and U2571 (N_2571,N_1981,N_1171);
xnor U2572 (N_2572,N_233,N_500);
nor U2573 (N_2573,N_1995,N_1041);
nand U2574 (N_2574,N_1790,N_106);
nand U2575 (N_2575,N_1191,N_737);
nand U2576 (N_2576,N_162,N_1358);
nand U2577 (N_2577,N_1474,N_521);
nand U2578 (N_2578,N_68,N_931);
and U2579 (N_2579,N_781,N_1583);
or U2580 (N_2580,N_1771,N_209);
nand U2581 (N_2581,N_1386,N_676);
nor U2582 (N_2582,N_329,N_892);
xor U2583 (N_2583,N_1042,N_698);
and U2584 (N_2584,N_720,N_414);
nor U2585 (N_2585,N_808,N_729);
nand U2586 (N_2586,N_139,N_1850);
nand U2587 (N_2587,N_1540,N_1585);
xor U2588 (N_2588,N_1143,N_600);
or U2589 (N_2589,N_1954,N_992);
nor U2590 (N_2590,N_1188,N_558);
nor U2591 (N_2591,N_1674,N_880);
and U2592 (N_2592,N_1624,N_62);
and U2593 (N_2593,N_391,N_651);
nand U2594 (N_2594,N_1730,N_259);
and U2595 (N_2595,N_562,N_877);
xnor U2596 (N_2596,N_997,N_1516);
and U2597 (N_2597,N_1148,N_1529);
or U2598 (N_2598,N_1955,N_89);
or U2599 (N_2599,N_1383,N_1454);
or U2600 (N_2600,N_1958,N_388);
nand U2601 (N_2601,N_192,N_184);
nand U2602 (N_2602,N_205,N_1711);
nand U2603 (N_2603,N_930,N_1819);
and U2604 (N_2604,N_1091,N_10);
and U2605 (N_2605,N_967,N_1822);
nor U2606 (N_2606,N_1548,N_1723);
or U2607 (N_2607,N_126,N_1160);
nand U2608 (N_2608,N_502,N_1219);
nand U2609 (N_2609,N_300,N_1149);
and U2610 (N_2610,N_1693,N_1535);
or U2611 (N_2611,N_217,N_54);
nor U2612 (N_2612,N_1938,N_1189);
or U2613 (N_2613,N_649,N_918);
nand U2614 (N_2614,N_1587,N_768);
and U2615 (N_2615,N_1904,N_1390);
nand U2616 (N_2616,N_677,N_1315);
and U2617 (N_2617,N_1990,N_399);
nor U2618 (N_2618,N_225,N_1135);
or U2619 (N_2619,N_1238,N_1327);
or U2620 (N_2620,N_577,N_1890);
nor U2621 (N_2621,N_338,N_316);
nand U2622 (N_2622,N_1560,N_1299);
nor U2623 (N_2623,N_514,N_596);
nand U2624 (N_2624,N_861,N_7);
or U2625 (N_2625,N_1240,N_647);
or U2626 (N_2626,N_1523,N_465);
or U2627 (N_2627,N_580,N_272);
or U2628 (N_2628,N_1477,N_25);
nand U2629 (N_2629,N_1568,N_794);
nor U2630 (N_2630,N_837,N_1261);
or U2631 (N_2631,N_1199,N_757);
xor U2632 (N_2632,N_234,N_1459);
or U2633 (N_2633,N_806,N_658);
or U2634 (N_2634,N_289,N_723);
nand U2635 (N_2635,N_1566,N_506);
and U2636 (N_2636,N_696,N_583);
xor U2637 (N_2637,N_485,N_1988);
or U2638 (N_2638,N_1257,N_724);
nor U2639 (N_2639,N_750,N_1187);
and U2640 (N_2640,N_611,N_1746);
nor U2641 (N_2641,N_336,N_760);
nor U2642 (N_2642,N_1037,N_833);
nor U2643 (N_2643,N_1539,N_332);
nor U2644 (N_2644,N_1440,N_1650);
or U2645 (N_2645,N_824,N_489);
nor U2646 (N_2646,N_424,N_725);
or U2647 (N_2647,N_92,N_946);
or U2648 (N_2648,N_1117,N_474);
nand U2649 (N_2649,N_1977,N_1978);
xnor U2650 (N_2650,N_1604,N_1594);
or U2651 (N_2651,N_971,N_405);
or U2652 (N_2652,N_299,N_942);
nand U2653 (N_2653,N_394,N_1114);
nand U2654 (N_2654,N_119,N_152);
nor U2655 (N_2655,N_541,N_349);
nand U2656 (N_2656,N_1437,N_471);
nand U2657 (N_2657,N_523,N_418);
and U2658 (N_2658,N_1398,N_1965);
or U2659 (N_2659,N_507,N_1864);
nand U2660 (N_2660,N_1075,N_1552);
nand U2661 (N_2661,N_488,N_140);
nand U2662 (N_2662,N_1607,N_1082);
or U2663 (N_2663,N_434,N_1941);
nor U2664 (N_2664,N_674,N_298);
nand U2665 (N_2665,N_50,N_960);
and U2666 (N_2666,N_1875,N_79);
and U2667 (N_2667,N_107,N_1352);
or U2668 (N_2668,N_118,N_1713);
or U2669 (N_2669,N_1889,N_1387);
nor U2670 (N_2670,N_826,N_1530);
xnor U2671 (N_2671,N_1749,N_1311);
or U2672 (N_2672,N_330,N_1544);
nor U2673 (N_2673,N_216,N_1774);
nand U2674 (N_2674,N_1803,N_1885);
and U2675 (N_2675,N_1863,N_841);
and U2676 (N_2676,N_625,N_1960);
and U2677 (N_2677,N_1374,N_1448);
nand U2678 (N_2678,N_1128,N_246);
nor U2679 (N_2679,N_355,N_977);
nand U2680 (N_2680,N_84,N_242);
nor U2681 (N_2681,N_1533,N_1147);
or U2682 (N_2682,N_1510,N_1914);
xnor U2683 (N_2683,N_1986,N_1435);
nand U2684 (N_2684,N_1882,N_1582);
or U2685 (N_2685,N_174,N_395);
nand U2686 (N_2686,N_524,N_1298);
or U2687 (N_2687,N_673,N_797);
nand U2688 (N_2688,N_1652,N_544);
nor U2689 (N_2689,N_1106,N_49);
or U2690 (N_2690,N_934,N_1406);
or U2691 (N_2691,N_1957,N_1119);
or U2692 (N_2692,N_1586,N_112);
nand U2693 (N_2693,N_1789,N_1641);
and U2694 (N_2694,N_1062,N_1320);
and U2695 (N_2695,N_881,N_288);
xor U2696 (N_2696,N_1415,N_1542);
or U2697 (N_2697,N_773,N_1569);
nor U2698 (N_2698,N_661,N_467);
and U2699 (N_2699,N_1367,N_1680);
xor U2700 (N_2700,N_1936,N_256);
or U2701 (N_2701,N_392,N_1499);
or U2702 (N_2702,N_1141,N_468);
or U2703 (N_2703,N_591,N_315);
or U2704 (N_2704,N_772,N_1659);
or U2705 (N_2705,N_277,N_1180);
nor U2706 (N_2706,N_132,N_1643);
and U2707 (N_2707,N_1169,N_1698);
or U2708 (N_2708,N_308,N_159);
or U2709 (N_2709,N_1359,N_149);
or U2710 (N_2710,N_1999,N_536);
nand U2711 (N_2711,N_94,N_1854);
nor U2712 (N_2712,N_933,N_704);
nand U2713 (N_2713,N_1799,N_352);
nor U2714 (N_2714,N_1430,N_1384);
nor U2715 (N_2715,N_888,N_1475);
and U2716 (N_2716,N_1216,N_707);
and U2717 (N_2717,N_204,N_902);
or U2718 (N_2718,N_410,N_572);
nand U2719 (N_2719,N_910,N_1433);
and U2720 (N_2720,N_924,N_535);
or U2721 (N_2721,N_1824,N_1121);
xnor U2722 (N_2722,N_1322,N_884);
nand U2723 (N_2723,N_1796,N_943);
and U2724 (N_2724,N_1234,N_1026);
nand U2725 (N_2725,N_1908,N_756);
nor U2726 (N_2726,N_1046,N_450);
nor U2727 (N_2727,N_1900,N_515);
nor U2728 (N_2728,N_858,N_194);
nand U2729 (N_2729,N_61,N_529);
and U2730 (N_2730,N_71,N_1684);
nor U2731 (N_2731,N_1178,N_87);
nor U2732 (N_2732,N_1177,N_1940);
nand U2733 (N_2733,N_753,N_653);
nor U2734 (N_2734,N_102,N_370);
or U2735 (N_2735,N_290,N_241);
or U2736 (N_2736,N_411,N_803);
nor U2737 (N_2737,N_383,N_457);
xnor U2738 (N_2738,N_914,N_1425);
and U2739 (N_2739,N_443,N_814);
nand U2740 (N_2740,N_144,N_1943);
nor U2741 (N_2741,N_957,N_561);
nor U2742 (N_2742,N_324,N_604);
xor U2743 (N_2743,N_1736,N_1488);
nor U2744 (N_2744,N_472,N_1120);
nor U2745 (N_2745,N_1655,N_401);
or U2746 (N_2746,N_623,N_202);
nand U2747 (N_2747,N_1479,N_45);
or U2748 (N_2748,N_1345,N_1242);
nand U2749 (N_2749,N_908,N_637);
or U2750 (N_2750,N_1532,N_1351);
or U2751 (N_2751,N_1592,N_137);
or U2752 (N_2752,N_1802,N_4);
and U2753 (N_2753,N_815,N_5);
or U2754 (N_2754,N_1428,N_1497);
or U2755 (N_2755,N_679,N_716);
or U2756 (N_2756,N_730,N_1845);
or U2757 (N_2757,N_397,N_656);
nand U2758 (N_2758,N_111,N_1023);
nand U2759 (N_2759,N_616,N_400);
or U2760 (N_2760,N_553,N_688);
or U2761 (N_2761,N_1228,N_1748);
nor U2762 (N_2762,N_1745,N_1370);
xor U2763 (N_2763,N_195,N_1848);
nor U2764 (N_2764,N_1070,N_1869);
nor U2765 (N_2765,N_1006,N_882);
nand U2766 (N_2766,N_1580,N_1118);
nor U2767 (N_2767,N_109,N_1078);
xnor U2768 (N_2768,N_1209,N_409);
and U2769 (N_2769,N_379,N_1731);
nor U2770 (N_2770,N_15,N_351);
nor U2771 (N_2771,N_761,N_1277);
and U2772 (N_2772,N_1561,N_1855);
nand U2773 (N_2773,N_751,N_1717);
nand U2774 (N_2774,N_1920,N_1004);
nor U2775 (N_2775,N_959,N_1710);
or U2776 (N_2776,N_1758,N_342);
nand U2777 (N_2777,N_498,N_1871);
nand U2778 (N_2778,N_659,N_1087);
and U2779 (N_2779,N_343,N_887);
and U2780 (N_2780,N_726,N_326);
and U2781 (N_2781,N_1262,N_491);
or U2782 (N_2782,N_1284,N_1389);
nor U2783 (N_2783,N_1831,N_1645);
xnor U2784 (N_2784,N_183,N_179);
and U2785 (N_2785,N_1040,N_1928);
nand U2786 (N_2786,N_1801,N_477);
and U2787 (N_2787,N_296,N_567);
and U2788 (N_2788,N_1696,N_221);
xnor U2789 (N_2789,N_143,N_1013);
and U2790 (N_2790,N_470,N_1657);
nand U2791 (N_2791,N_899,N_1024);
or U2792 (N_2792,N_1347,N_1895);
and U2793 (N_2793,N_1744,N_1125);
and U2794 (N_2794,N_1017,N_398);
nand U2795 (N_2795,N_1288,N_1866);
or U2796 (N_2796,N_210,N_670);
and U2797 (N_2797,N_86,N_14);
or U2798 (N_2798,N_1480,N_1192);
or U2799 (N_2799,N_1917,N_1194);
or U2800 (N_2800,N_1295,N_1331);
or U2801 (N_2801,N_451,N_652);
or U2802 (N_2802,N_35,N_1681);
and U2803 (N_2803,N_1366,N_646);
or U2804 (N_2804,N_1661,N_1804);
nand U2805 (N_2805,N_75,N_970);
xnor U2806 (N_2806,N_731,N_778);
xor U2807 (N_2807,N_703,N_537);
nor U2808 (N_2808,N_1667,N_1253);
and U2809 (N_2809,N_69,N_767);
or U2810 (N_2810,N_563,N_1825);
nand U2811 (N_2811,N_1016,N_1093);
nor U2812 (N_2812,N_1342,N_549);
or U2813 (N_2813,N_1235,N_921);
or U2814 (N_2814,N_800,N_1915);
nor U2815 (N_2815,N_372,N_44);
nand U2816 (N_2816,N_460,N_607);
nand U2817 (N_2817,N_1708,N_945);
nor U2818 (N_2818,N_1766,N_610);
nand U2819 (N_2819,N_1086,N_978);
or U2820 (N_2820,N_177,N_1600);
and U2821 (N_2821,N_693,N_1489);
and U2822 (N_2822,N_362,N_1395);
xnor U2823 (N_2823,N_1404,N_1633);
or U2824 (N_2824,N_373,N_1522);
and U2825 (N_2825,N_1043,N_1675);
nor U2826 (N_2826,N_1896,N_689);
nor U2827 (N_2827,N_788,N_1861);
nand U2828 (N_2828,N_1912,N_436);
nor U2829 (N_2829,N_1340,N_965);
or U2830 (N_2830,N_437,N_1709);
nor U2831 (N_2831,N_1305,N_763);
or U2832 (N_2832,N_728,N_853);
or U2833 (N_2833,N_1637,N_423);
nand U2834 (N_2834,N_1157,N_941);
nor U2835 (N_2835,N_1631,N_1218);
xnor U2836 (N_2836,N_1805,N_1924);
xnor U2837 (N_2837,N_133,N_640);
and U2838 (N_2838,N_848,N_154);
xor U2839 (N_2839,N_1689,N_1063);
nor U2840 (N_2840,N_1181,N_851);
nor U2841 (N_2841,N_1918,N_1491);
nand U2842 (N_2842,N_212,N_64);
or U2843 (N_2843,N_587,N_662);
nand U2844 (N_2844,N_1330,N_134);
nor U2845 (N_2845,N_1210,N_1797);
nor U2846 (N_2846,N_448,N_350);
or U2847 (N_2847,N_832,N_261);
and U2848 (N_2848,N_131,N_614);
nor U2849 (N_2849,N_705,N_1490);
nor U2850 (N_2850,N_1651,N_620);
nand U2851 (N_2851,N_906,N_1809);
or U2852 (N_2852,N_354,N_1827);
and U2853 (N_2853,N_1901,N_466);
nor U2854 (N_2854,N_1563,N_1427);
nor U2855 (N_2855,N_1142,N_1321);
xnor U2856 (N_2856,N_1452,N_973);
or U2857 (N_2857,N_615,N_495);
nor U2858 (N_2858,N_792,N_1449);
nand U2859 (N_2859,N_1872,N_1858);
nand U2860 (N_2860,N_1968,N_1663);
nand U2861 (N_2861,N_519,N_566);
and U2862 (N_2862,N_1926,N_421);
or U2863 (N_2863,N_636,N_426);
nor U2864 (N_2864,N_816,N_873);
nor U2865 (N_2865,N_1303,N_692);
nand U2866 (N_2866,N_480,N_1735);
and U2867 (N_2867,N_213,N_266);
and U2868 (N_2868,N_531,N_258);
nand U2869 (N_2869,N_747,N_260);
nand U2870 (N_2870,N_1429,N_1520);
nor U2871 (N_2871,N_497,N_41);
nand U2872 (N_2872,N_228,N_634);
nor U2873 (N_2873,N_622,N_1393);
or U2874 (N_2874,N_1611,N_1590);
nand U2875 (N_2875,N_1032,N_1714);
or U2876 (N_2876,N_798,N_1368);
nor U2877 (N_2877,N_1950,N_1612);
or U2878 (N_2878,N_844,N_856);
xor U2879 (N_2879,N_1152,N_1951);
and U2880 (N_2880,N_265,N_1668);
or U2881 (N_2881,N_420,N_293);
xor U2882 (N_2882,N_982,N_991);
and U2883 (N_2883,N_103,N_95);
nand U2884 (N_2884,N_665,N_3);
nor U2885 (N_2885,N_926,N_1258);
nor U2886 (N_2886,N_114,N_575);
nor U2887 (N_2887,N_1306,N_1381);
nor U2888 (N_2888,N_248,N_121);
nor U2889 (N_2889,N_962,N_439);
or U2890 (N_2890,N_19,N_599);
nor U2891 (N_2891,N_1204,N_895);
and U2892 (N_2892,N_1814,N_586);
nor U2893 (N_2893,N_820,N_1897);
nor U2894 (N_2894,N_968,N_1144);
or U2895 (N_2895,N_52,N_1635);
and U2896 (N_2896,N_702,N_1099);
or U2897 (N_2897,N_802,N_1975);
and U2898 (N_2898,N_1269,N_545);
nand U2899 (N_2899,N_574,N_360);
or U2900 (N_2900,N_53,N_1380);
nand U2901 (N_2901,N_1202,N_486);
and U2902 (N_2902,N_2,N_1064);
and U2903 (N_2903,N_393,N_1096);
nand U2904 (N_2904,N_1378,N_1732);
nand U2905 (N_2905,N_156,N_1325);
and U2906 (N_2906,N_1451,N_1294);
or U2907 (N_2907,N_20,N_444);
xnor U2908 (N_2908,N_850,N_1131);
nand U2909 (N_2909,N_1838,N_47);
or U2910 (N_2910,N_413,N_1755);
nand U2911 (N_2911,N_1049,N_518);
nand U2912 (N_2912,N_23,N_671);
and U2913 (N_2913,N_732,N_961);
and U2914 (N_2914,N_889,N_1308);
nand U2915 (N_2915,N_1832,N_1484);
nor U2916 (N_2916,N_1551,N_1496);
and U2917 (N_2917,N_81,N_1220);
or U2918 (N_2918,N_923,N_353);
nor U2919 (N_2919,N_1465,N_1514);
or U2920 (N_2920,N_1225,N_939);
and U2921 (N_2921,N_1682,N_1506);
nand U2922 (N_2922,N_1349,N_1628);
xor U2923 (N_2923,N_1473,N_1274);
or U2924 (N_2924,N_764,N_603);
nand U2925 (N_2925,N_1715,N_1341);
xor U2926 (N_2926,N_264,N_158);
nand U2927 (N_2927,N_1916,N_1500);
nand U2928 (N_2928,N_639,N_522);
and U2929 (N_2929,N_428,N_1259);
nand U2930 (N_2930,N_1223,N_153);
and U2931 (N_2931,N_969,N_1823);
nor U2932 (N_2932,N_907,N_1787);
nor U2933 (N_2933,N_1054,N_1829);
nor U2934 (N_2934,N_1371,N_1478);
or U2935 (N_2935,N_993,N_1959);
nand U2936 (N_2936,N_1104,N_1982);
nand U2937 (N_2937,N_1279,N_1549);
nand U2938 (N_2938,N_1156,N_711);
and U2939 (N_2939,N_1007,N_286);
and U2940 (N_2940,N_1145,N_331);
and U2941 (N_2941,N_1718,N_827);
and U2942 (N_2942,N_384,N_1576);
nand U2943 (N_2943,N_1246,N_1902);
or U2944 (N_2944,N_494,N_1176);
and U2945 (N_2945,N_976,N_1868);
nand U2946 (N_2946,N_727,N_275);
nand U2947 (N_2947,N_1283,N_1502);
nor U2948 (N_2948,N_875,N_268);
and U2949 (N_2949,N_834,N_108);
nand U2950 (N_2950,N_403,N_18);
and U2951 (N_2951,N_1527,N_1843);
nor U2952 (N_2952,N_232,N_1842);
and U2953 (N_2953,N_1414,N_1964);
xnor U2954 (N_2954,N_552,N_1155);
nand U2955 (N_2955,N_208,N_469);
and U2956 (N_2956,N_1346,N_30);
nor U2957 (N_2957,N_593,N_1405);
nand U2958 (N_2958,N_589,N_879);
xor U2959 (N_2959,N_897,N_185);
nor U2960 (N_2960,N_169,N_752);
nor U2961 (N_2961,N_113,N_1297);
and U2962 (N_2962,N_1278,N_186);
and U2963 (N_2963,N_1949,N_115);
nor U2964 (N_2964,N_222,N_1458);
xor U2965 (N_2965,N_629,N_1905);
xor U2966 (N_2966,N_165,N_1944);
or U2967 (N_2967,N_1463,N_936);
or U2968 (N_2968,N_1166,N_1025);
xor U2969 (N_2969,N_1880,N_1546);
nor U2970 (N_2970,N_1000,N_893);
and U2971 (N_2971,N_1021,N_1618);
or U2972 (N_2972,N_482,N_1423);
or U2973 (N_2973,N_954,N_1697);
or U2974 (N_2974,N_1146,N_1161);
or U2975 (N_2975,N_341,N_1694);
nor U2976 (N_2976,N_813,N_1190);
nor U2977 (N_2977,N_1153,N_1739);
nand U2978 (N_2978,N_412,N_1808);
nor U2979 (N_2979,N_1547,N_1865);
nand U2980 (N_2980,N_686,N_1102);
nand U2981 (N_2981,N_710,N_1874);
and U2982 (N_2982,N_988,N_334);
nor U2983 (N_2983,N_1685,N_1431);
nor U2984 (N_2984,N_37,N_1642);
or U2985 (N_2985,N_749,N_415);
and U2986 (N_2986,N_197,N_1432);
xor U2987 (N_2987,N_1603,N_1646);
or U2988 (N_2988,N_70,N_479);
nand U2989 (N_2989,N_1265,N_1621);
nor U2990 (N_2990,N_441,N_1632);
or U2991 (N_2991,N_1045,N_447);
and U2992 (N_2992,N_219,N_1881);
and U2993 (N_2993,N_588,N_548);
and U2994 (N_2994,N_864,N_989);
nor U2995 (N_2995,N_1254,N_1080);
and U2996 (N_2996,N_1198,N_743);
and U2997 (N_2997,N_129,N_1029);
or U2998 (N_2998,N_687,N_630);
xnor U2999 (N_2999,N_663,N_36);
xnor U3000 (N_3000,N_16,N_790);
nand U3001 (N_3001,N_1566,N_1367);
or U3002 (N_3002,N_1308,N_167);
nand U3003 (N_3003,N_1480,N_732);
nand U3004 (N_3004,N_810,N_693);
xor U3005 (N_3005,N_1850,N_187);
or U3006 (N_3006,N_1412,N_346);
nor U3007 (N_3007,N_1410,N_1084);
xor U3008 (N_3008,N_590,N_831);
or U3009 (N_3009,N_418,N_1104);
nand U3010 (N_3010,N_1361,N_519);
and U3011 (N_3011,N_1494,N_1022);
nand U3012 (N_3012,N_489,N_1628);
or U3013 (N_3013,N_661,N_1028);
nor U3014 (N_3014,N_608,N_1092);
nor U3015 (N_3015,N_1376,N_59);
nand U3016 (N_3016,N_1928,N_693);
xnor U3017 (N_3017,N_1428,N_1321);
nor U3018 (N_3018,N_1658,N_1127);
or U3019 (N_3019,N_975,N_1931);
and U3020 (N_3020,N_1911,N_1902);
or U3021 (N_3021,N_1393,N_802);
xor U3022 (N_3022,N_370,N_1747);
xor U3023 (N_3023,N_1651,N_324);
or U3024 (N_3024,N_1212,N_497);
and U3025 (N_3025,N_320,N_1313);
nand U3026 (N_3026,N_126,N_178);
or U3027 (N_3027,N_1947,N_219);
nor U3028 (N_3028,N_1425,N_1727);
nand U3029 (N_3029,N_1844,N_1143);
and U3030 (N_3030,N_154,N_720);
nor U3031 (N_3031,N_1363,N_1548);
or U3032 (N_3032,N_927,N_1949);
or U3033 (N_3033,N_1298,N_453);
and U3034 (N_3034,N_1491,N_55);
and U3035 (N_3035,N_1229,N_844);
nor U3036 (N_3036,N_500,N_1153);
nor U3037 (N_3037,N_323,N_1694);
xnor U3038 (N_3038,N_82,N_1395);
or U3039 (N_3039,N_689,N_917);
or U3040 (N_3040,N_19,N_1086);
or U3041 (N_3041,N_1536,N_979);
and U3042 (N_3042,N_1705,N_712);
and U3043 (N_3043,N_924,N_1145);
nor U3044 (N_3044,N_881,N_1429);
nor U3045 (N_3045,N_734,N_212);
nor U3046 (N_3046,N_923,N_1380);
nand U3047 (N_3047,N_1053,N_345);
and U3048 (N_3048,N_1077,N_1579);
and U3049 (N_3049,N_700,N_735);
and U3050 (N_3050,N_67,N_1664);
and U3051 (N_3051,N_1343,N_100);
xor U3052 (N_3052,N_249,N_567);
nor U3053 (N_3053,N_1018,N_406);
and U3054 (N_3054,N_920,N_32);
nor U3055 (N_3055,N_778,N_1745);
nor U3056 (N_3056,N_849,N_60);
nor U3057 (N_3057,N_1759,N_1442);
nor U3058 (N_3058,N_1360,N_1996);
nand U3059 (N_3059,N_40,N_1935);
and U3060 (N_3060,N_194,N_1319);
and U3061 (N_3061,N_1362,N_1695);
and U3062 (N_3062,N_313,N_1761);
and U3063 (N_3063,N_1064,N_88);
nor U3064 (N_3064,N_347,N_449);
or U3065 (N_3065,N_1872,N_541);
and U3066 (N_3066,N_1239,N_2);
or U3067 (N_3067,N_552,N_1826);
nor U3068 (N_3068,N_1506,N_740);
and U3069 (N_3069,N_203,N_1633);
and U3070 (N_3070,N_465,N_1294);
nand U3071 (N_3071,N_490,N_1782);
nand U3072 (N_3072,N_1072,N_165);
and U3073 (N_3073,N_29,N_782);
or U3074 (N_3074,N_771,N_1168);
nor U3075 (N_3075,N_1274,N_1562);
or U3076 (N_3076,N_1072,N_367);
and U3077 (N_3077,N_1150,N_93);
nor U3078 (N_3078,N_1129,N_1902);
or U3079 (N_3079,N_13,N_590);
nor U3080 (N_3080,N_1852,N_1665);
nand U3081 (N_3081,N_411,N_936);
xnor U3082 (N_3082,N_1865,N_1804);
or U3083 (N_3083,N_1499,N_1231);
nand U3084 (N_3084,N_1301,N_704);
nand U3085 (N_3085,N_358,N_208);
nor U3086 (N_3086,N_1302,N_1015);
nand U3087 (N_3087,N_1816,N_850);
nor U3088 (N_3088,N_835,N_1797);
and U3089 (N_3089,N_535,N_285);
nor U3090 (N_3090,N_1137,N_657);
nand U3091 (N_3091,N_337,N_1077);
nand U3092 (N_3092,N_1758,N_1174);
xor U3093 (N_3093,N_1646,N_327);
and U3094 (N_3094,N_1557,N_1835);
and U3095 (N_3095,N_1760,N_1019);
nor U3096 (N_3096,N_993,N_1930);
and U3097 (N_3097,N_886,N_36);
and U3098 (N_3098,N_193,N_1896);
xnor U3099 (N_3099,N_1054,N_387);
xor U3100 (N_3100,N_1463,N_999);
nand U3101 (N_3101,N_1271,N_1990);
nand U3102 (N_3102,N_1128,N_1002);
or U3103 (N_3103,N_1069,N_181);
nand U3104 (N_3104,N_1863,N_495);
and U3105 (N_3105,N_1197,N_1390);
nand U3106 (N_3106,N_57,N_1229);
or U3107 (N_3107,N_733,N_732);
nand U3108 (N_3108,N_180,N_269);
or U3109 (N_3109,N_319,N_93);
and U3110 (N_3110,N_404,N_456);
or U3111 (N_3111,N_1249,N_1681);
and U3112 (N_3112,N_1433,N_607);
and U3113 (N_3113,N_1687,N_808);
and U3114 (N_3114,N_1633,N_267);
nor U3115 (N_3115,N_918,N_1552);
and U3116 (N_3116,N_1115,N_1478);
xor U3117 (N_3117,N_1708,N_1906);
and U3118 (N_3118,N_1432,N_1134);
nor U3119 (N_3119,N_705,N_1731);
nand U3120 (N_3120,N_488,N_45);
and U3121 (N_3121,N_94,N_1725);
xnor U3122 (N_3122,N_298,N_122);
nand U3123 (N_3123,N_1525,N_1527);
or U3124 (N_3124,N_1952,N_1350);
nor U3125 (N_3125,N_659,N_1099);
or U3126 (N_3126,N_113,N_147);
nor U3127 (N_3127,N_1189,N_1234);
or U3128 (N_3128,N_968,N_1921);
or U3129 (N_3129,N_1144,N_1574);
and U3130 (N_3130,N_1054,N_1242);
nor U3131 (N_3131,N_964,N_675);
or U3132 (N_3132,N_681,N_139);
and U3133 (N_3133,N_1002,N_1283);
xnor U3134 (N_3134,N_1672,N_409);
or U3135 (N_3135,N_143,N_1451);
nor U3136 (N_3136,N_45,N_1427);
or U3137 (N_3137,N_209,N_930);
or U3138 (N_3138,N_1507,N_1641);
nand U3139 (N_3139,N_1613,N_11);
xnor U3140 (N_3140,N_1142,N_549);
and U3141 (N_3141,N_203,N_1994);
and U3142 (N_3142,N_332,N_1910);
nor U3143 (N_3143,N_1178,N_1337);
nand U3144 (N_3144,N_883,N_277);
and U3145 (N_3145,N_1960,N_1005);
xnor U3146 (N_3146,N_136,N_345);
and U3147 (N_3147,N_1843,N_15);
nand U3148 (N_3148,N_235,N_18);
or U3149 (N_3149,N_464,N_659);
and U3150 (N_3150,N_1866,N_151);
and U3151 (N_3151,N_1742,N_910);
or U3152 (N_3152,N_1054,N_468);
and U3153 (N_3153,N_255,N_1434);
nor U3154 (N_3154,N_1925,N_301);
nand U3155 (N_3155,N_799,N_320);
xnor U3156 (N_3156,N_1758,N_78);
or U3157 (N_3157,N_1987,N_230);
nand U3158 (N_3158,N_1527,N_1212);
or U3159 (N_3159,N_1493,N_240);
and U3160 (N_3160,N_1546,N_701);
and U3161 (N_3161,N_666,N_1249);
and U3162 (N_3162,N_745,N_757);
nor U3163 (N_3163,N_372,N_1246);
nand U3164 (N_3164,N_1873,N_7);
or U3165 (N_3165,N_463,N_1418);
and U3166 (N_3166,N_169,N_1318);
nor U3167 (N_3167,N_1425,N_314);
or U3168 (N_3168,N_54,N_11);
nor U3169 (N_3169,N_431,N_88);
nor U3170 (N_3170,N_1129,N_1652);
and U3171 (N_3171,N_76,N_1309);
nand U3172 (N_3172,N_1948,N_806);
or U3173 (N_3173,N_606,N_658);
and U3174 (N_3174,N_681,N_724);
and U3175 (N_3175,N_1224,N_352);
and U3176 (N_3176,N_283,N_84);
nand U3177 (N_3177,N_1085,N_1073);
and U3178 (N_3178,N_458,N_578);
nand U3179 (N_3179,N_1818,N_1713);
and U3180 (N_3180,N_1165,N_98);
nand U3181 (N_3181,N_507,N_128);
nand U3182 (N_3182,N_1519,N_1939);
or U3183 (N_3183,N_370,N_1247);
and U3184 (N_3184,N_1821,N_1022);
nor U3185 (N_3185,N_1233,N_750);
xor U3186 (N_3186,N_1433,N_275);
nor U3187 (N_3187,N_1988,N_1330);
and U3188 (N_3188,N_887,N_1048);
nand U3189 (N_3189,N_993,N_1941);
or U3190 (N_3190,N_985,N_473);
or U3191 (N_3191,N_310,N_1917);
and U3192 (N_3192,N_1841,N_830);
nor U3193 (N_3193,N_637,N_1122);
or U3194 (N_3194,N_286,N_1267);
nor U3195 (N_3195,N_931,N_333);
or U3196 (N_3196,N_551,N_1091);
nor U3197 (N_3197,N_1018,N_11);
nor U3198 (N_3198,N_1111,N_737);
or U3199 (N_3199,N_316,N_1845);
and U3200 (N_3200,N_1878,N_1720);
nand U3201 (N_3201,N_626,N_1855);
nand U3202 (N_3202,N_1230,N_89);
xor U3203 (N_3203,N_231,N_431);
nand U3204 (N_3204,N_607,N_1023);
nor U3205 (N_3205,N_1324,N_1572);
or U3206 (N_3206,N_106,N_604);
or U3207 (N_3207,N_360,N_483);
nor U3208 (N_3208,N_388,N_673);
xor U3209 (N_3209,N_63,N_1130);
nand U3210 (N_3210,N_1653,N_842);
nor U3211 (N_3211,N_320,N_794);
and U3212 (N_3212,N_532,N_334);
xnor U3213 (N_3213,N_1775,N_1013);
xnor U3214 (N_3214,N_1643,N_108);
xnor U3215 (N_3215,N_634,N_1157);
nor U3216 (N_3216,N_1786,N_1352);
nand U3217 (N_3217,N_1251,N_1146);
xor U3218 (N_3218,N_213,N_138);
xnor U3219 (N_3219,N_465,N_233);
nor U3220 (N_3220,N_725,N_454);
nand U3221 (N_3221,N_187,N_1541);
xor U3222 (N_3222,N_1575,N_1932);
nor U3223 (N_3223,N_1981,N_1162);
and U3224 (N_3224,N_260,N_177);
nand U3225 (N_3225,N_1782,N_1430);
or U3226 (N_3226,N_1979,N_533);
or U3227 (N_3227,N_1721,N_775);
xnor U3228 (N_3228,N_176,N_625);
nand U3229 (N_3229,N_17,N_454);
nand U3230 (N_3230,N_61,N_180);
and U3231 (N_3231,N_1509,N_710);
or U3232 (N_3232,N_483,N_351);
and U3233 (N_3233,N_750,N_1195);
nand U3234 (N_3234,N_1341,N_883);
nor U3235 (N_3235,N_818,N_915);
xnor U3236 (N_3236,N_276,N_787);
and U3237 (N_3237,N_874,N_1786);
or U3238 (N_3238,N_1745,N_90);
and U3239 (N_3239,N_901,N_127);
or U3240 (N_3240,N_196,N_1297);
or U3241 (N_3241,N_518,N_1834);
or U3242 (N_3242,N_486,N_1200);
or U3243 (N_3243,N_1135,N_1160);
or U3244 (N_3244,N_1451,N_1705);
and U3245 (N_3245,N_1077,N_349);
nor U3246 (N_3246,N_1620,N_837);
nor U3247 (N_3247,N_802,N_1966);
and U3248 (N_3248,N_1659,N_423);
xor U3249 (N_3249,N_1912,N_486);
and U3250 (N_3250,N_713,N_1616);
or U3251 (N_3251,N_976,N_1418);
nor U3252 (N_3252,N_547,N_384);
nor U3253 (N_3253,N_423,N_559);
nor U3254 (N_3254,N_682,N_1757);
nor U3255 (N_3255,N_1379,N_452);
or U3256 (N_3256,N_1955,N_1401);
nand U3257 (N_3257,N_1675,N_675);
or U3258 (N_3258,N_848,N_698);
nor U3259 (N_3259,N_1395,N_989);
nor U3260 (N_3260,N_1039,N_843);
or U3261 (N_3261,N_1483,N_713);
or U3262 (N_3262,N_115,N_1879);
nand U3263 (N_3263,N_1436,N_310);
xor U3264 (N_3264,N_1528,N_1504);
and U3265 (N_3265,N_746,N_715);
nand U3266 (N_3266,N_1511,N_1578);
nor U3267 (N_3267,N_1487,N_1206);
nand U3268 (N_3268,N_1747,N_577);
nand U3269 (N_3269,N_394,N_729);
or U3270 (N_3270,N_1649,N_1180);
or U3271 (N_3271,N_39,N_1781);
and U3272 (N_3272,N_1849,N_565);
nand U3273 (N_3273,N_1959,N_973);
and U3274 (N_3274,N_859,N_871);
nand U3275 (N_3275,N_1297,N_1511);
or U3276 (N_3276,N_1494,N_1391);
nand U3277 (N_3277,N_727,N_711);
nand U3278 (N_3278,N_193,N_1769);
and U3279 (N_3279,N_29,N_757);
or U3280 (N_3280,N_1305,N_1211);
nor U3281 (N_3281,N_803,N_1167);
nor U3282 (N_3282,N_927,N_469);
and U3283 (N_3283,N_1260,N_1951);
and U3284 (N_3284,N_1167,N_1467);
nor U3285 (N_3285,N_933,N_686);
or U3286 (N_3286,N_227,N_1831);
nand U3287 (N_3287,N_296,N_13);
xor U3288 (N_3288,N_1759,N_1698);
nor U3289 (N_3289,N_25,N_606);
and U3290 (N_3290,N_1745,N_446);
nor U3291 (N_3291,N_76,N_866);
or U3292 (N_3292,N_935,N_1184);
or U3293 (N_3293,N_998,N_1581);
xnor U3294 (N_3294,N_1136,N_1090);
or U3295 (N_3295,N_1298,N_331);
nor U3296 (N_3296,N_1068,N_1749);
nor U3297 (N_3297,N_1450,N_571);
or U3298 (N_3298,N_986,N_1170);
and U3299 (N_3299,N_886,N_1354);
or U3300 (N_3300,N_167,N_1371);
xor U3301 (N_3301,N_983,N_1495);
nand U3302 (N_3302,N_873,N_310);
or U3303 (N_3303,N_124,N_609);
or U3304 (N_3304,N_1266,N_647);
nand U3305 (N_3305,N_1926,N_761);
nand U3306 (N_3306,N_511,N_1633);
nor U3307 (N_3307,N_1189,N_782);
or U3308 (N_3308,N_1502,N_1647);
nand U3309 (N_3309,N_1753,N_607);
and U3310 (N_3310,N_307,N_1704);
and U3311 (N_3311,N_201,N_1213);
or U3312 (N_3312,N_481,N_1600);
nor U3313 (N_3313,N_1313,N_880);
nand U3314 (N_3314,N_414,N_5);
nor U3315 (N_3315,N_415,N_1760);
and U3316 (N_3316,N_1022,N_557);
and U3317 (N_3317,N_487,N_1449);
nor U3318 (N_3318,N_322,N_965);
and U3319 (N_3319,N_228,N_616);
and U3320 (N_3320,N_1913,N_801);
nor U3321 (N_3321,N_1688,N_498);
nor U3322 (N_3322,N_972,N_1917);
and U3323 (N_3323,N_1531,N_1643);
nor U3324 (N_3324,N_1951,N_1184);
nand U3325 (N_3325,N_1185,N_768);
or U3326 (N_3326,N_691,N_335);
xnor U3327 (N_3327,N_526,N_355);
nor U3328 (N_3328,N_511,N_1255);
and U3329 (N_3329,N_103,N_1905);
nand U3330 (N_3330,N_366,N_1640);
and U3331 (N_3331,N_1751,N_448);
or U3332 (N_3332,N_500,N_1627);
and U3333 (N_3333,N_794,N_642);
and U3334 (N_3334,N_398,N_772);
or U3335 (N_3335,N_1698,N_731);
xnor U3336 (N_3336,N_1772,N_205);
nor U3337 (N_3337,N_92,N_377);
nand U3338 (N_3338,N_1604,N_420);
nand U3339 (N_3339,N_1939,N_1029);
nand U3340 (N_3340,N_250,N_1298);
xnor U3341 (N_3341,N_1971,N_765);
xor U3342 (N_3342,N_1043,N_438);
nor U3343 (N_3343,N_1492,N_1312);
xnor U3344 (N_3344,N_1792,N_132);
and U3345 (N_3345,N_32,N_555);
and U3346 (N_3346,N_1140,N_1797);
nand U3347 (N_3347,N_783,N_647);
nand U3348 (N_3348,N_1292,N_427);
nand U3349 (N_3349,N_1900,N_1113);
and U3350 (N_3350,N_457,N_1104);
and U3351 (N_3351,N_139,N_1852);
or U3352 (N_3352,N_501,N_1279);
and U3353 (N_3353,N_929,N_1131);
and U3354 (N_3354,N_1882,N_1699);
and U3355 (N_3355,N_161,N_220);
nand U3356 (N_3356,N_1492,N_1265);
and U3357 (N_3357,N_587,N_1962);
or U3358 (N_3358,N_1864,N_1319);
or U3359 (N_3359,N_773,N_1470);
and U3360 (N_3360,N_52,N_699);
nor U3361 (N_3361,N_1869,N_516);
nor U3362 (N_3362,N_877,N_1978);
and U3363 (N_3363,N_1958,N_1573);
xor U3364 (N_3364,N_308,N_1739);
and U3365 (N_3365,N_550,N_285);
and U3366 (N_3366,N_1736,N_1383);
or U3367 (N_3367,N_1234,N_1509);
and U3368 (N_3368,N_1700,N_3);
nand U3369 (N_3369,N_196,N_628);
nor U3370 (N_3370,N_74,N_1466);
or U3371 (N_3371,N_1425,N_113);
and U3372 (N_3372,N_283,N_553);
or U3373 (N_3373,N_1272,N_818);
nor U3374 (N_3374,N_1638,N_247);
or U3375 (N_3375,N_1219,N_764);
and U3376 (N_3376,N_1862,N_657);
and U3377 (N_3377,N_679,N_72);
nand U3378 (N_3378,N_1236,N_685);
nand U3379 (N_3379,N_1946,N_231);
nand U3380 (N_3380,N_1611,N_1896);
nor U3381 (N_3381,N_1496,N_840);
nor U3382 (N_3382,N_1455,N_1959);
nand U3383 (N_3383,N_1244,N_1);
and U3384 (N_3384,N_1719,N_48);
or U3385 (N_3385,N_851,N_1610);
nand U3386 (N_3386,N_1412,N_1770);
nor U3387 (N_3387,N_41,N_1745);
nand U3388 (N_3388,N_1743,N_1155);
nor U3389 (N_3389,N_202,N_1171);
and U3390 (N_3390,N_1022,N_1765);
nand U3391 (N_3391,N_1920,N_44);
xnor U3392 (N_3392,N_1533,N_1158);
nor U3393 (N_3393,N_1253,N_311);
nand U3394 (N_3394,N_824,N_1895);
or U3395 (N_3395,N_1072,N_154);
and U3396 (N_3396,N_1051,N_1440);
and U3397 (N_3397,N_1470,N_1416);
nand U3398 (N_3398,N_22,N_694);
and U3399 (N_3399,N_26,N_635);
and U3400 (N_3400,N_1879,N_359);
or U3401 (N_3401,N_553,N_565);
nand U3402 (N_3402,N_545,N_1260);
or U3403 (N_3403,N_1147,N_323);
and U3404 (N_3404,N_1654,N_849);
nor U3405 (N_3405,N_773,N_1189);
xnor U3406 (N_3406,N_1734,N_179);
or U3407 (N_3407,N_1312,N_444);
nor U3408 (N_3408,N_657,N_1901);
nor U3409 (N_3409,N_315,N_1000);
nand U3410 (N_3410,N_527,N_1906);
or U3411 (N_3411,N_1554,N_1523);
nor U3412 (N_3412,N_993,N_204);
xnor U3413 (N_3413,N_387,N_880);
xor U3414 (N_3414,N_1239,N_1403);
and U3415 (N_3415,N_1541,N_1359);
xnor U3416 (N_3416,N_385,N_967);
or U3417 (N_3417,N_992,N_1018);
or U3418 (N_3418,N_1818,N_168);
nor U3419 (N_3419,N_1088,N_1091);
nor U3420 (N_3420,N_268,N_171);
and U3421 (N_3421,N_1822,N_1794);
and U3422 (N_3422,N_1206,N_179);
xnor U3423 (N_3423,N_1193,N_1508);
nor U3424 (N_3424,N_538,N_1761);
or U3425 (N_3425,N_937,N_1344);
nand U3426 (N_3426,N_88,N_86);
nor U3427 (N_3427,N_130,N_271);
and U3428 (N_3428,N_1183,N_266);
or U3429 (N_3429,N_610,N_1466);
or U3430 (N_3430,N_1914,N_1836);
and U3431 (N_3431,N_1414,N_1954);
and U3432 (N_3432,N_905,N_1851);
nand U3433 (N_3433,N_822,N_959);
or U3434 (N_3434,N_1799,N_141);
and U3435 (N_3435,N_1023,N_1836);
and U3436 (N_3436,N_133,N_52);
nor U3437 (N_3437,N_981,N_958);
nor U3438 (N_3438,N_1814,N_776);
and U3439 (N_3439,N_1356,N_795);
or U3440 (N_3440,N_1960,N_1423);
or U3441 (N_3441,N_1284,N_772);
nor U3442 (N_3442,N_572,N_1469);
or U3443 (N_3443,N_1874,N_1389);
nor U3444 (N_3444,N_651,N_521);
nand U3445 (N_3445,N_1398,N_533);
or U3446 (N_3446,N_746,N_152);
nor U3447 (N_3447,N_781,N_1928);
or U3448 (N_3448,N_1718,N_1005);
or U3449 (N_3449,N_1177,N_1584);
nor U3450 (N_3450,N_1940,N_849);
nand U3451 (N_3451,N_626,N_884);
nand U3452 (N_3452,N_679,N_351);
nand U3453 (N_3453,N_85,N_427);
and U3454 (N_3454,N_880,N_1767);
xor U3455 (N_3455,N_1007,N_998);
nand U3456 (N_3456,N_592,N_497);
xnor U3457 (N_3457,N_1622,N_549);
and U3458 (N_3458,N_1775,N_843);
xor U3459 (N_3459,N_549,N_1848);
nor U3460 (N_3460,N_363,N_756);
and U3461 (N_3461,N_1600,N_609);
nand U3462 (N_3462,N_920,N_465);
nand U3463 (N_3463,N_1486,N_1649);
and U3464 (N_3464,N_1566,N_503);
nor U3465 (N_3465,N_819,N_1341);
and U3466 (N_3466,N_361,N_176);
nor U3467 (N_3467,N_213,N_410);
nand U3468 (N_3468,N_1570,N_565);
or U3469 (N_3469,N_469,N_1020);
nand U3470 (N_3470,N_1221,N_920);
nor U3471 (N_3471,N_1263,N_758);
nor U3472 (N_3472,N_1013,N_1668);
and U3473 (N_3473,N_1778,N_1004);
or U3474 (N_3474,N_356,N_292);
xnor U3475 (N_3475,N_211,N_309);
nand U3476 (N_3476,N_1041,N_482);
nor U3477 (N_3477,N_1208,N_649);
nand U3478 (N_3478,N_646,N_278);
nand U3479 (N_3479,N_798,N_1739);
nor U3480 (N_3480,N_365,N_1193);
nand U3481 (N_3481,N_1236,N_1682);
nand U3482 (N_3482,N_1518,N_1497);
and U3483 (N_3483,N_578,N_978);
xnor U3484 (N_3484,N_811,N_906);
nand U3485 (N_3485,N_892,N_1444);
nor U3486 (N_3486,N_1073,N_1961);
and U3487 (N_3487,N_1562,N_1066);
nor U3488 (N_3488,N_407,N_1259);
and U3489 (N_3489,N_1289,N_7);
xnor U3490 (N_3490,N_347,N_1082);
xnor U3491 (N_3491,N_1623,N_1743);
nand U3492 (N_3492,N_1951,N_154);
nand U3493 (N_3493,N_1891,N_880);
and U3494 (N_3494,N_169,N_1199);
and U3495 (N_3495,N_95,N_1307);
xnor U3496 (N_3496,N_297,N_601);
xor U3497 (N_3497,N_235,N_985);
nor U3498 (N_3498,N_1731,N_1932);
nor U3499 (N_3499,N_312,N_1736);
and U3500 (N_3500,N_1317,N_456);
nor U3501 (N_3501,N_1129,N_113);
or U3502 (N_3502,N_201,N_411);
or U3503 (N_3503,N_1137,N_1657);
and U3504 (N_3504,N_1641,N_300);
and U3505 (N_3505,N_1984,N_406);
nor U3506 (N_3506,N_1192,N_1146);
and U3507 (N_3507,N_1086,N_390);
nand U3508 (N_3508,N_1218,N_957);
and U3509 (N_3509,N_1779,N_987);
nor U3510 (N_3510,N_704,N_369);
nor U3511 (N_3511,N_354,N_1537);
xnor U3512 (N_3512,N_1849,N_199);
nor U3513 (N_3513,N_314,N_1643);
nand U3514 (N_3514,N_855,N_266);
xnor U3515 (N_3515,N_189,N_1821);
nand U3516 (N_3516,N_1266,N_1267);
nand U3517 (N_3517,N_1027,N_1551);
and U3518 (N_3518,N_20,N_898);
and U3519 (N_3519,N_1385,N_1283);
and U3520 (N_3520,N_444,N_275);
nor U3521 (N_3521,N_860,N_286);
and U3522 (N_3522,N_1751,N_1834);
and U3523 (N_3523,N_1607,N_1327);
or U3524 (N_3524,N_658,N_260);
nand U3525 (N_3525,N_3,N_483);
nor U3526 (N_3526,N_1078,N_684);
and U3527 (N_3527,N_1024,N_1770);
nand U3528 (N_3528,N_1285,N_1050);
and U3529 (N_3529,N_789,N_246);
nand U3530 (N_3530,N_428,N_1875);
and U3531 (N_3531,N_295,N_675);
nand U3532 (N_3532,N_1523,N_1526);
and U3533 (N_3533,N_1932,N_641);
or U3534 (N_3534,N_1352,N_184);
nor U3535 (N_3535,N_391,N_50);
and U3536 (N_3536,N_1865,N_1471);
nor U3537 (N_3537,N_9,N_981);
nor U3538 (N_3538,N_1179,N_1160);
nand U3539 (N_3539,N_478,N_1614);
nand U3540 (N_3540,N_554,N_1755);
xor U3541 (N_3541,N_1637,N_1050);
nor U3542 (N_3542,N_1998,N_664);
or U3543 (N_3543,N_1425,N_754);
or U3544 (N_3544,N_796,N_1695);
or U3545 (N_3545,N_1280,N_230);
nand U3546 (N_3546,N_997,N_1910);
nor U3547 (N_3547,N_1148,N_1015);
nor U3548 (N_3548,N_1861,N_1280);
and U3549 (N_3549,N_377,N_853);
or U3550 (N_3550,N_886,N_281);
xor U3551 (N_3551,N_1595,N_1646);
or U3552 (N_3552,N_262,N_570);
nor U3553 (N_3553,N_1118,N_1416);
or U3554 (N_3554,N_447,N_665);
or U3555 (N_3555,N_1673,N_1050);
and U3556 (N_3556,N_1073,N_1737);
nor U3557 (N_3557,N_1815,N_1517);
and U3558 (N_3558,N_1513,N_19);
or U3559 (N_3559,N_1722,N_660);
and U3560 (N_3560,N_1991,N_646);
nand U3561 (N_3561,N_1506,N_1296);
or U3562 (N_3562,N_188,N_331);
nor U3563 (N_3563,N_1419,N_548);
and U3564 (N_3564,N_171,N_1249);
or U3565 (N_3565,N_813,N_883);
nand U3566 (N_3566,N_339,N_480);
or U3567 (N_3567,N_553,N_891);
nor U3568 (N_3568,N_1002,N_263);
nand U3569 (N_3569,N_1433,N_21);
nand U3570 (N_3570,N_1033,N_1961);
and U3571 (N_3571,N_1173,N_1112);
and U3572 (N_3572,N_668,N_740);
and U3573 (N_3573,N_1530,N_1567);
or U3574 (N_3574,N_1995,N_918);
xor U3575 (N_3575,N_668,N_1093);
nand U3576 (N_3576,N_372,N_61);
nand U3577 (N_3577,N_356,N_1933);
and U3578 (N_3578,N_1766,N_310);
and U3579 (N_3579,N_135,N_1446);
and U3580 (N_3580,N_925,N_1871);
or U3581 (N_3581,N_1348,N_887);
nor U3582 (N_3582,N_1490,N_1644);
and U3583 (N_3583,N_116,N_1430);
nor U3584 (N_3584,N_272,N_1776);
nor U3585 (N_3585,N_1037,N_59);
nor U3586 (N_3586,N_732,N_1977);
and U3587 (N_3587,N_573,N_723);
xor U3588 (N_3588,N_1581,N_1345);
nand U3589 (N_3589,N_1441,N_1206);
xnor U3590 (N_3590,N_1737,N_664);
xnor U3591 (N_3591,N_1653,N_1018);
and U3592 (N_3592,N_648,N_1172);
and U3593 (N_3593,N_1060,N_594);
and U3594 (N_3594,N_188,N_1277);
and U3595 (N_3595,N_1790,N_194);
nand U3596 (N_3596,N_1275,N_952);
and U3597 (N_3597,N_1875,N_1223);
nor U3598 (N_3598,N_1213,N_1613);
and U3599 (N_3599,N_1248,N_652);
and U3600 (N_3600,N_1189,N_1867);
nor U3601 (N_3601,N_1123,N_38);
nand U3602 (N_3602,N_1845,N_46);
nand U3603 (N_3603,N_1496,N_1899);
nor U3604 (N_3604,N_922,N_1653);
and U3605 (N_3605,N_372,N_604);
nand U3606 (N_3606,N_775,N_1559);
nor U3607 (N_3607,N_63,N_1028);
and U3608 (N_3608,N_1888,N_1513);
nand U3609 (N_3609,N_1590,N_467);
or U3610 (N_3610,N_118,N_550);
nand U3611 (N_3611,N_1067,N_20);
or U3612 (N_3612,N_1895,N_1924);
or U3613 (N_3613,N_704,N_1411);
and U3614 (N_3614,N_247,N_444);
nand U3615 (N_3615,N_1427,N_1394);
nand U3616 (N_3616,N_1189,N_951);
or U3617 (N_3617,N_352,N_770);
and U3618 (N_3618,N_1906,N_1297);
xnor U3619 (N_3619,N_1740,N_760);
or U3620 (N_3620,N_1594,N_1520);
or U3621 (N_3621,N_903,N_364);
or U3622 (N_3622,N_77,N_1563);
nand U3623 (N_3623,N_729,N_61);
and U3624 (N_3624,N_404,N_1848);
or U3625 (N_3625,N_1192,N_1696);
and U3626 (N_3626,N_179,N_1789);
xor U3627 (N_3627,N_1894,N_37);
and U3628 (N_3628,N_23,N_1057);
nand U3629 (N_3629,N_1955,N_1276);
nand U3630 (N_3630,N_1423,N_1613);
and U3631 (N_3631,N_546,N_417);
and U3632 (N_3632,N_293,N_511);
or U3633 (N_3633,N_1497,N_1120);
nand U3634 (N_3634,N_1105,N_1242);
and U3635 (N_3635,N_799,N_1269);
or U3636 (N_3636,N_1867,N_30);
and U3637 (N_3637,N_1484,N_535);
or U3638 (N_3638,N_522,N_1834);
nand U3639 (N_3639,N_315,N_34);
or U3640 (N_3640,N_1610,N_1981);
or U3641 (N_3641,N_959,N_315);
and U3642 (N_3642,N_1160,N_1352);
nor U3643 (N_3643,N_17,N_1003);
nor U3644 (N_3644,N_1937,N_1418);
nor U3645 (N_3645,N_1810,N_867);
and U3646 (N_3646,N_1935,N_353);
and U3647 (N_3647,N_639,N_450);
nor U3648 (N_3648,N_139,N_1156);
xnor U3649 (N_3649,N_1580,N_1718);
nor U3650 (N_3650,N_809,N_1384);
xor U3651 (N_3651,N_297,N_763);
nor U3652 (N_3652,N_1114,N_1794);
xor U3653 (N_3653,N_115,N_1782);
xor U3654 (N_3654,N_1431,N_1893);
nand U3655 (N_3655,N_844,N_218);
or U3656 (N_3656,N_434,N_219);
nand U3657 (N_3657,N_188,N_1505);
nor U3658 (N_3658,N_1238,N_118);
or U3659 (N_3659,N_973,N_1251);
or U3660 (N_3660,N_913,N_1572);
or U3661 (N_3661,N_586,N_1545);
or U3662 (N_3662,N_1041,N_167);
and U3663 (N_3663,N_1128,N_380);
nor U3664 (N_3664,N_364,N_812);
and U3665 (N_3665,N_19,N_970);
or U3666 (N_3666,N_931,N_1552);
nor U3667 (N_3667,N_1535,N_591);
nor U3668 (N_3668,N_781,N_1762);
nand U3669 (N_3669,N_952,N_1643);
and U3670 (N_3670,N_609,N_86);
or U3671 (N_3671,N_1039,N_1556);
nor U3672 (N_3672,N_1930,N_1117);
nor U3673 (N_3673,N_217,N_939);
and U3674 (N_3674,N_1055,N_376);
nor U3675 (N_3675,N_167,N_832);
or U3676 (N_3676,N_279,N_337);
nand U3677 (N_3677,N_1705,N_1120);
nor U3678 (N_3678,N_299,N_1833);
and U3679 (N_3679,N_560,N_1075);
and U3680 (N_3680,N_481,N_1073);
xnor U3681 (N_3681,N_846,N_8);
or U3682 (N_3682,N_939,N_527);
and U3683 (N_3683,N_1531,N_1176);
nor U3684 (N_3684,N_377,N_395);
or U3685 (N_3685,N_233,N_1422);
nor U3686 (N_3686,N_343,N_1024);
nand U3687 (N_3687,N_1598,N_654);
nor U3688 (N_3688,N_104,N_834);
nand U3689 (N_3689,N_1963,N_1108);
and U3690 (N_3690,N_1346,N_603);
or U3691 (N_3691,N_1903,N_132);
nand U3692 (N_3692,N_0,N_573);
and U3693 (N_3693,N_1262,N_1951);
nor U3694 (N_3694,N_593,N_1837);
and U3695 (N_3695,N_1822,N_361);
xnor U3696 (N_3696,N_1846,N_1732);
and U3697 (N_3697,N_1623,N_560);
nor U3698 (N_3698,N_937,N_765);
nand U3699 (N_3699,N_1599,N_1483);
or U3700 (N_3700,N_307,N_446);
and U3701 (N_3701,N_498,N_290);
and U3702 (N_3702,N_1908,N_1975);
nor U3703 (N_3703,N_31,N_556);
or U3704 (N_3704,N_1578,N_1679);
or U3705 (N_3705,N_81,N_885);
and U3706 (N_3706,N_364,N_964);
nand U3707 (N_3707,N_1490,N_1353);
and U3708 (N_3708,N_373,N_802);
and U3709 (N_3709,N_1922,N_1687);
nor U3710 (N_3710,N_520,N_1834);
and U3711 (N_3711,N_1583,N_646);
nand U3712 (N_3712,N_33,N_1721);
or U3713 (N_3713,N_1882,N_1356);
and U3714 (N_3714,N_1006,N_461);
nand U3715 (N_3715,N_1806,N_677);
nor U3716 (N_3716,N_289,N_429);
and U3717 (N_3717,N_1101,N_388);
xor U3718 (N_3718,N_1004,N_1719);
nor U3719 (N_3719,N_1807,N_475);
nor U3720 (N_3720,N_845,N_872);
xor U3721 (N_3721,N_1328,N_545);
nand U3722 (N_3722,N_1217,N_911);
xor U3723 (N_3723,N_1250,N_1767);
nand U3724 (N_3724,N_322,N_1990);
nand U3725 (N_3725,N_1979,N_859);
nand U3726 (N_3726,N_1390,N_998);
nor U3727 (N_3727,N_1232,N_60);
and U3728 (N_3728,N_450,N_989);
or U3729 (N_3729,N_569,N_286);
nand U3730 (N_3730,N_30,N_1040);
and U3731 (N_3731,N_1585,N_444);
nand U3732 (N_3732,N_168,N_1015);
or U3733 (N_3733,N_748,N_237);
or U3734 (N_3734,N_371,N_1678);
nor U3735 (N_3735,N_421,N_1835);
xor U3736 (N_3736,N_164,N_1763);
nand U3737 (N_3737,N_1970,N_1689);
nand U3738 (N_3738,N_903,N_239);
nor U3739 (N_3739,N_418,N_837);
nor U3740 (N_3740,N_5,N_1661);
nand U3741 (N_3741,N_1670,N_1165);
and U3742 (N_3742,N_175,N_541);
nand U3743 (N_3743,N_980,N_1352);
nand U3744 (N_3744,N_1904,N_1783);
or U3745 (N_3745,N_381,N_1743);
nor U3746 (N_3746,N_1274,N_833);
or U3747 (N_3747,N_1272,N_561);
or U3748 (N_3748,N_1824,N_859);
or U3749 (N_3749,N_1009,N_852);
or U3750 (N_3750,N_10,N_1754);
and U3751 (N_3751,N_1597,N_684);
and U3752 (N_3752,N_1724,N_1740);
and U3753 (N_3753,N_493,N_1225);
nand U3754 (N_3754,N_162,N_589);
or U3755 (N_3755,N_239,N_684);
xnor U3756 (N_3756,N_141,N_24);
or U3757 (N_3757,N_1236,N_1728);
nor U3758 (N_3758,N_51,N_846);
xnor U3759 (N_3759,N_382,N_1263);
and U3760 (N_3760,N_1704,N_1871);
nand U3761 (N_3761,N_963,N_1617);
and U3762 (N_3762,N_1712,N_1226);
xor U3763 (N_3763,N_1009,N_112);
or U3764 (N_3764,N_1936,N_1078);
nor U3765 (N_3765,N_1406,N_555);
and U3766 (N_3766,N_1478,N_1250);
nor U3767 (N_3767,N_1496,N_785);
xor U3768 (N_3768,N_538,N_964);
nor U3769 (N_3769,N_1659,N_1816);
nand U3770 (N_3770,N_270,N_1646);
or U3771 (N_3771,N_892,N_1727);
nand U3772 (N_3772,N_1427,N_1283);
nor U3773 (N_3773,N_234,N_1958);
nand U3774 (N_3774,N_335,N_34);
or U3775 (N_3775,N_1515,N_258);
nor U3776 (N_3776,N_108,N_1458);
nand U3777 (N_3777,N_742,N_1778);
or U3778 (N_3778,N_9,N_409);
nor U3779 (N_3779,N_158,N_1690);
and U3780 (N_3780,N_1099,N_479);
nor U3781 (N_3781,N_778,N_594);
nand U3782 (N_3782,N_1722,N_76);
nand U3783 (N_3783,N_1055,N_180);
nand U3784 (N_3784,N_818,N_1020);
xnor U3785 (N_3785,N_1552,N_464);
or U3786 (N_3786,N_719,N_1541);
and U3787 (N_3787,N_220,N_921);
nor U3788 (N_3788,N_1468,N_130);
or U3789 (N_3789,N_1990,N_438);
nor U3790 (N_3790,N_976,N_991);
nor U3791 (N_3791,N_135,N_1897);
or U3792 (N_3792,N_1130,N_706);
nor U3793 (N_3793,N_1261,N_524);
xnor U3794 (N_3794,N_1320,N_1121);
and U3795 (N_3795,N_1165,N_1608);
nand U3796 (N_3796,N_87,N_327);
and U3797 (N_3797,N_859,N_1104);
and U3798 (N_3798,N_282,N_269);
and U3799 (N_3799,N_1530,N_460);
nand U3800 (N_3800,N_1876,N_1051);
nand U3801 (N_3801,N_1873,N_305);
or U3802 (N_3802,N_968,N_1599);
nand U3803 (N_3803,N_849,N_697);
nand U3804 (N_3804,N_1711,N_731);
or U3805 (N_3805,N_969,N_1150);
and U3806 (N_3806,N_466,N_1270);
nand U3807 (N_3807,N_285,N_459);
nand U3808 (N_3808,N_667,N_1064);
or U3809 (N_3809,N_1161,N_175);
and U3810 (N_3810,N_1582,N_844);
and U3811 (N_3811,N_856,N_738);
nand U3812 (N_3812,N_1769,N_1525);
xnor U3813 (N_3813,N_508,N_1195);
nor U3814 (N_3814,N_1736,N_741);
and U3815 (N_3815,N_1687,N_634);
nand U3816 (N_3816,N_1306,N_837);
or U3817 (N_3817,N_985,N_1816);
nor U3818 (N_3818,N_1616,N_780);
or U3819 (N_3819,N_610,N_1746);
nand U3820 (N_3820,N_1199,N_37);
and U3821 (N_3821,N_1276,N_874);
nand U3822 (N_3822,N_1351,N_1327);
nand U3823 (N_3823,N_60,N_364);
nor U3824 (N_3824,N_1336,N_1279);
and U3825 (N_3825,N_380,N_1054);
nand U3826 (N_3826,N_1881,N_1306);
and U3827 (N_3827,N_1934,N_1889);
nor U3828 (N_3828,N_74,N_232);
nor U3829 (N_3829,N_1182,N_771);
nor U3830 (N_3830,N_1938,N_1789);
xor U3831 (N_3831,N_116,N_807);
and U3832 (N_3832,N_1117,N_256);
nand U3833 (N_3833,N_764,N_459);
or U3834 (N_3834,N_1500,N_699);
nor U3835 (N_3835,N_25,N_402);
or U3836 (N_3836,N_1747,N_1011);
or U3837 (N_3837,N_143,N_1677);
nor U3838 (N_3838,N_1949,N_1988);
or U3839 (N_3839,N_1628,N_1702);
and U3840 (N_3840,N_1291,N_1825);
nor U3841 (N_3841,N_513,N_1627);
or U3842 (N_3842,N_509,N_1162);
and U3843 (N_3843,N_1081,N_519);
and U3844 (N_3844,N_750,N_674);
or U3845 (N_3845,N_1548,N_1296);
or U3846 (N_3846,N_91,N_1884);
xnor U3847 (N_3847,N_1666,N_194);
nor U3848 (N_3848,N_1112,N_1009);
nor U3849 (N_3849,N_868,N_776);
nand U3850 (N_3850,N_1329,N_1445);
or U3851 (N_3851,N_52,N_536);
nand U3852 (N_3852,N_605,N_1766);
or U3853 (N_3853,N_723,N_832);
nand U3854 (N_3854,N_198,N_1218);
nand U3855 (N_3855,N_982,N_180);
nand U3856 (N_3856,N_1866,N_17);
xnor U3857 (N_3857,N_1047,N_395);
nand U3858 (N_3858,N_819,N_1868);
nor U3859 (N_3859,N_1540,N_1297);
nor U3860 (N_3860,N_135,N_1427);
nand U3861 (N_3861,N_1724,N_1701);
or U3862 (N_3862,N_417,N_537);
or U3863 (N_3863,N_1208,N_1136);
nand U3864 (N_3864,N_1595,N_548);
nand U3865 (N_3865,N_550,N_461);
and U3866 (N_3866,N_1055,N_1234);
nand U3867 (N_3867,N_1452,N_856);
or U3868 (N_3868,N_1146,N_1836);
nor U3869 (N_3869,N_1688,N_105);
or U3870 (N_3870,N_534,N_1028);
and U3871 (N_3871,N_1777,N_1656);
nor U3872 (N_3872,N_537,N_1719);
nor U3873 (N_3873,N_291,N_1713);
nand U3874 (N_3874,N_543,N_985);
nand U3875 (N_3875,N_955,N_391);
nor U3876 (N_3876,N_1068,N_1953);
or U3877 (N_3877,N_1535,N_1999);
and U3878 (N_3878,N_1802,N_620);
nor U3879 (N_3879,N_1799,N_1780);
and U3880 (N_3880,N_1800,N_784);
and U3881 (N_3881,N_764,N_1929);
nor U3882 (N_3882,N_368,N_1384);
or U3883 (N_3883,N_8,N_303);
and U3884 (N_3884,N_1230,N_266);
nor U3885 (N_3885,N_234,N_573);
nand U3886 (N_3886,N_944,N_549);
nand U3887 (N_3887,N_574,N_1946);
nand U3888 (N_3888,N_1640,N_182);
or U3889 (N_3889,N_1818,N_1987);
or U3890 (N_3890,N_1255,N_600);
or U3891 (N_3891,N_1965,N_180);
nand U3892 (N_3892,N_730,N_1400);
nor U3893 (N_3893,N_1796,N_667);
nor U3894 (N_3894,N_1034,N_693);
xnor U3895 (N_3895,N_1357,N_1641);
nand U3896 (N_3896,N_1118,N_7);
or U3897 (N_3897,N_1939,N_1512);
nor U3898 (N_3898,N_462,N_1906);
nor U3899 (N_3899,N_1248,N_1027);
nand U3900 (N_3900,N_1434,N_1126);
nor U3901 (N_3901,N_486,N_1643);
xnor U3902 (N_3902,N_165,N_1190);
or U3903 (N_3903,N_630,N_1707);
or U3904 (N_3904,N_8,N_776);
xnor U3905 (N_3905,N_1409,N_376);
nand U3906 (N_3906,N_550,N_732);
nand U3907 (N_3907,N_402,N_1800);
and U3908 (N_3908,N_299,N_1083);
nand U3909 (N_3909,N_694,N_895);
and U3910 (N_3910,N_517,N_1693);
and U3911 (N_3911,N_1996,N_835);
xnor U3912 (N_3912,N_579,N_1604);
nand U3913 (N_3913,N_667,N_56);
nand U3914 (N_3914,N_1958,N_1170);
or U3915 (N_3915,N_1171,N_608);
xor U3916 (N_3916,N_1464,N_581);
nor U3917 (N_3917,N_181,N_1749);
or U3918 (N_3918,N_1841,N_927);
nand U3919 (N_3919,N_1067,N_1568);
nor U3920 (N_3920,N_1801,N_829);
xor U3921 (N_3921,N_777,N_1713);
and U3922 (N_3922,N_1980,N_286);
or U3923 (N_3923,N_851,N_988);
and U3924 (N_3924,N_1208,N_83);
or U3925 (N_3925,N_1735,N_27);
and U3926 (N_3926,N_38,N_1478);
and U3927 (N_3927,N_520,N_1558);
nor U3928 (N_3928,N_371,N_103);
and U3929 (N_3929,N_599,N_1611);
or U3930 (N_3930,N_944,N_1919);
nand U3931 (N_3931,N_1126,N_1982);
nor U3932 (N_3932,N_775,N_1942);
nand U3933 (N_3933,N_363,N_566);
nor U3934 (N_3934,N_667,N_850);
and U3935 (N_3935,N_1260,N_123);
and U3936 (N_3936,N_1810,N_321);
or U3937 (N_3937,N_1654,N_1864);
and U3938 (N_3938,N_1437,N_80);
nand U3939 (N_3939,N_586,N_1557);
nand U3940 (N_3940,N_403,N_1247);
and U3941 (N_3941,N_38,N_1502);
nand U3942 (N_3942,N_758,N_1103);
xor U3943 (N_3943,N_908,N_409);
xor U3944 (N_3944,N_1241,N_1080);
or U3945 (N_3945,N_838,N_1364);
nand U3946 (N_3946,N_534,N_505);
nor U3947 (N_3947,N_1642,N_304);
nor U3948 (N_3948,N_1667,N_1094);
or U3949 (N_3949,N_1802,N_711);
xor U3950 (N_3950,N_1058,N_789);
nand U3951 (N_3951,N_1773,N_1342);
nor U3952 (N_3952,N_1463,N_1187);
xnor U3953 (N_3953,N_22,N_135);
and U3954 (N_3954,N_595,N_1849);
nand U3955 (N_3955,N_788,N_1736);
nand U3956 (N_3956,N_632,N_386);
and U3957 (N_3957,N_548,N_1315);
xor U3958 (N_3958,N_1053,N_1492);
and U3959 (N_3959,N_116,N_22);
nand U3960 (N_3960,N_1836,N_138);
or U3961 (N_3961,N_1601,N_1211);
and U3962 (N_3962,N_1327,N_1848);
and U3963 (N_3963,N_823,N_1516);
nand U3964 (N_3964,N_1031,N_319);
xor U3965 (N_3965,N_1361,N_219);
or U3966 (N_3966,N_1624,N_567);
nor U3967 (N_3967,N_800,N_475);
nor U3968 (N_3968,N_786,N_1911);
and U3969 (N_3969,N_274,N_1942);
nor U3970 (N_3970,N_492,N_1736);
or U3971 (N_3971,N_1490,N_1706);
and U3972 (N_3972,N_1333,N_492);
xor U3973 (N_3973,N_1189,N_289);
nand U3974 (N_3974,N_1614,N_1528);
nor U3975 (N_3975,N_814,N_319);
or U3976 (N_3976,N_241,N_1308);
and U3977 (N_3977,N_1772,N_610);
nor U3978 (N_3978,N_878,N_1891);
or U3979 (N_3979,N_992,N_861);
or U3980 (N_3980,N_1977,N_776);
or U3981 (N_3981,N_1249,N_573);
nor U3982 (N_3982,N_817,N_1559);
and U3983 (N_3983,N_882,N_299);
xnor U3984 (N_3984,N_960,N_1292);
xor U3985 (N_3985,N_1008,N_65);
nor U3986 (N_3986,N_1438,N_1894);
and U3987 (N_3987,N_1426,N_944);
and U3988 (N_3988,N_1938,N_148);
nor U3989 (N_3989,N_1614,N_1594);
and U3990 (N_3990,N_118,N_1919);
and U3991 (N_3991,N_1540,N_1923);
or U3992 (N_3992,N_577,N_728);
and U3993 (N_3993,N_199,N_361);
xnor U3994 (N_3994,N_1676,N_1240);
nand U3995 (N_3995,N_1590,N_1196);
nand U3996 (N_3996,N_1742,N_494);
nand U3997 (N_3997,N_871,N_884);
nor U3998 (N_3998,N_905,N_1053);
nor U3999 (N_3999,N_1092,N_983);
nand U4000 (N_4000,N_2061,N_2762);
nand U4001 (N_4001,N_3962,N_2535);
xor U4002 (N_4002,N_2462,N_3744);
nand U4003 (N_4003,N_3582,N_3325);
or U4004 (N_4004,N_2139,N_3292);
or U4005 (N_4005,N_2500,N_3863);
or U4006 (N_4006,N_3546,N_3491);
xor U4007 (N_4007,N_2408,N_2340);
xor U4008 (N_4008,N_2419,N_2414);
nand U4009 (N_4009,N_3144,N_3284);
and U4010 (N_4010,N_2632,N_3643);
nor U4011 (N_4011,N_3571,N_3404);
nand U4012 (N_4012,N_3667,N_3456);
xor U4013 (N_4013,N_3206,N_2895);
or U4014 (N_4014,N_2696,N_2910);
nand U4015 (N_4015,N_2147,N_3652);
nor U4016 (N_4016,N_2357,N_3311);
and U4017 (N_4017,N_2600,N_3992);
or U4018 (N_4018,N_2562,N_2608);
or U4019 (N_4019,N_2598,N_2431);
nand U4020 (N_4020,N_3376,N_2889);
nand U4021 (N_4021,N_2993,N_2890);
nand U4022 (N_4022,N_3415,N_2132);
nor U4023 (N_4023,N_3893,N_3225);
nand U4024 (N_4024,N_3087,N_3921);
or U4025 (N_4025,N_2222,N_3909);
or U4026 (N_4026,N_2808,N_3705);
or U4027 (N_4027,N_2013,N_3003);
nor U4028 (N_4028,N_2700,N_3094);
nand U4029 (N_4029,N_3021,N_2255);
or U4030 (N_4030,N_2536,N_2878);
or U4031 (N_4031,N_2292,N_2131);
or U4032 (N_4032,N_2763,N_2706);
nor U4033 (N_4033,N_3857,N_3572);
nor U4034 (N_4034,N_3825,N_2741);
nand U4035 (N_4035,N_3031,N_2621);
or U4036 (N_4036,N_2786,N_3259);
nor U4037 (N_4037,N_2393,N_3700);
nor U4038 (N_4038,N_3357,N_2454);
and U4039 (N_4039,N_3540,N_2363);
or U4040 (N_4040,N_2160,N_2827);
xnor U4041 (N_4041,N_2217,N_3648);
and U4042 (N_4042,N_2892,N_3855);
nand U4043 (N_4043,N_2218,N_3627);
or U4044 (N_4044,N_3786,N_2877);
nand U4045 (N_4045,N_3459,N_2410);
nand U4046 (N_4046,N_2100,N_3645);
and U4047 (N_4047,N_3812,N_3304);
and U4048 (N_4048,N_3661,N_2617);
nand U4049 (N_4049,N_3473,N_3635);
xor U4050 (N_4050,N_2815,N_3166);
nand U4051 (N_4051,N_3019,N_2656);
or U4052 (N_4052,N_3498,N_3506);
xnor U4053 (N_4053,N_2845,N_2926);
nand U4054 (N_4054,N_3137,N_3447);
nand U4055 (N_4055,N_3297,N_3011);
and U4056 (N_4056,N_2451,N_2436);
and U4057 (N_4057,N_3853,N_2407);
nor U4058 (N_4058,N_2113,N_2011);
nand U4059 (N_4059,N_2425,N_3324);
and U4060 (N_4060,N_3906,N_2273);
and U4061 (N_4061,N_2070,N_3566);
nor U4062 (N_4062,N_3056,N_2901);
or U4063 (N_4063,N_3027,N_3753);
or U4064 (N_4064,N_3622,N_3760);
nor U4065 (N_4065,N_3783,N_3043);
nand U4066 (N_4066,N_3560,N_2166);
nor U4067 (N_4067,N_2007,N_3406);
nand U4068 (N_4068,N_3053,N_2293);
and U4069 (N_4069,N_3923,N_2884);
nand U4070 (N_4070,N_3086,N_3435);
nand U4071 (N_4071,N_3826,N_2261);
and U4072 (N_4072,N_3486,N_3973);
and U4073 (N_4073,N_2221,N_3776);
xnor U4074 (N_4074,N_3696,N_3949);
and U4075 (N_4075,N_3051,N_3028);
nand U4076 (N_4076,N_3122,N_3879);
or U4077 (N_4077,N_3055,N_2981);
nor U4078 (N_4078,N_3308,N_2494);
and U4079 (N_4079,N_3544,N_3749);
or U4080 (N_4080,N_2580,N_2365);
nand U4081 (N_4081,N_2597,N_3090);
nor U4082 (N_4082,N_3139,N_3547);
or U4083 (N_4083,N_2846,N_2213);
nand U4084 (N_4084,N_3332,N_2093);
and U4085 (N_4085,N_3837,N_3203);
xor U4086 (N_4086,N_2917,N_3590);
or U4087 (N_4087,N_2920,N_3610);
and U4088 (N_4088,N_3537,N_2944);
or U4089 (N_4089,N_3690,N_3132);
or U4090 (N_4090,N_2144,N_2380);
xnor U4091 (N_4091,N_3639,N_2039);
xnor U4092 (N_4092,N_3687,N_2599);
nand U4093 (N_4093,N_2125,N_3271);
nand U4094 (N_4094,N_3410,N_3649);
xor U4095 (N_4095,N_2933,N_2238);
or U4096 (N_4096,N_2409,N_2278);
or U4097 (N_4097,N_2969,N_2711);
nor U4098 (N_4098,N_2888,N_3561);
nand U4099 (N_4099,N_3101,N_2539);
and U4100 (N_4100,N_2383,N_2760);
and U4101 (N_4101,N_2818,N_2992);
and U4102 (N_4102,N_2973,N_2157);
and U4103 (N_4103,N_2082,N_2275);
and U4104 (N_4104,N_2504,N_3396);
nand U4105 (N_4105,N_3482,N_2382);
and U4106 (N_4106,N_3497,N_2122);
nand U4107 (N_4107,N_2483,N_2914);
nor U4108 (N_4108,N_3769,N_2886);
and U4109 (N_4109,N_2831,N_2753);
or U4110 (N_4110,N_2282,N_3875);
and U4111 (N_4111,N_2778,N_2162);
nor U4112 (N_4112,N_2868,N_2294);
nand U4113 (N_4113,N_3197,N_3465);
or U4114 (N_4114,N_3301,N_2077);
and U4115 (N_4115,N_2894,N_2349);
or U4116 (N_4116,N_3626,N_2306);
or U4117 (N_4117,N_3836,N_2675);
nand U4118 (N_4118,N_3545,N_2523);
xnor U4119 (N_4119,N_3298,N_3955);
and U4120 (N_4120,N_2676,N_2102);
and U4121 (N_4121,N_2479,N_2487);
nand U4122 (N_4122,N_2552,N_2809);
and U4123 (N_4123,N_2618,N_2976);
or U4124 (N_4124,N_2524,N_2189);
xnor U4125 (N_4125,N_3978,N_2574);
nand U4126 (N_4126,N_3142,N_3337);
nor U4127 (N_4127,N_2634,N_2528);
or U4128 (N_4128,N_2283,N_2505);
or U4129 (N_4129,N_2545,N_3468);
and U4130 (N_4130,N_2076,N_3095);
and U4131 (N_4131,N_2657,N_3559);
xnor U4132 (N_4132,N_3001,N_3780);
and U4133 (N_4133,N_3444,N_2610);
and U4134 (N_4134,N_2605,N_3300);
nand U4135 (N_4135,N_3047,N_2876);
nand U4136 (N_4136,N_2241,N_2647);
or U4137 (N_4137,N_2925,N_2736);
or U4138 (N_4138,N_2072,N_2949);
and U4139 (N_4139,N_3887,N_3599);
xor U4140 (N_4140,N_2210,N_2399);
and U4141 (N_4141,N_3367,N_2701);
and U4142 (N_4142,N_3516,N_3107);
nand U4143 (N_4143,N_2206,N_2905);
nand U4144 (N_4144,N_3928,N_2946);
nand U4145 (N_4145,N_3806,N_3264);
or U4146 (N_4146,N_2502,N_3767);
nor U4147 (N_4147,N_3905,N_3691);
and U4148 (N_4148,N_2604,N_3196);
nand U4149 (N_4149,N_3071,N_3959);
and U4150 (N_4150,N_3596,N_2937);
nand U4151 (N_4151,N_2947,N_2900);
nor U4152 (N_4152,N_3052,N_3088);
and U4153 (N_4153,N_2152,N_2127);
nand U4154 (N_4154,N_3405,N_3219);
nor U4155 (N_4155,N_3430,N_3771);
or U4156 (N_4156,N_3778,N_2685);
nor U4157 (N_4157,N_2743,N_2134);
and U4158 (N_4158,N_2176,N_3674);
and U4159 (N_4159,N_2126,N_2650);
or U4160 (N_4160,N_2033,N_2682);
and U4161 (N_4161,N_3215,N_2475);
and U4162 (N_4162,N_3568,N_3530);
or U4163 (N_4163,N_3490,N_3676);
or U4164 (N_4164,N_2923,N_2522);
nor U4165 (N_4165,N_3589,N_2641);
nand U4166 (N_4166,N_3323,N_2246);
or U4167 (N_4167,N_2046,N_3218);
nand U4168 (N_4168,N_3570,N_2034);
nand U4169 (N_4169,N_2887,N_3424);
and U4170 (N_4170,N_3333,N_2795);
nand U4171 (N_4171,N_3952,N_3161);
or U4172 (N_4172,N_3188,N_3105);
or U4173 (N_4173,N_2154,N_3654);
and U4174 (N_4174,N_3126,N_3556);
nor U4175 (N_4175,N_2765,N_2554);
nor U4176 (N_4176,N_2514,N_3838);
or U4177 (N_4177,N_3427,N_2994);
nor U4178 (N_4178,N_2195,N_2744);
or U4179 (N_4179,N_3385,N_2774);
nor U4180 (N_4180,N_3069,N_2354);
or U4181 (N_4181,N_3348,N_2049);
nand U4182 (N_4182,N_3081,N_3179);
or U4183 (N_4183,N_2427,N_3791);
nor U4184 (N_4184,N_3703,N_3035);
nand U4185 (N_4185,N_2314,N_2151);
nor U4186 (N_4186,N_2968,N_3869);
or U4187 (N_4187,N_2509,N_2153);
nand U4188 (N_4188,N_3967,N_2821);
nor U4189 (N_4189,N_3951,N_2432);
nor U4190 (N_4190,N_2421,N_3555);
nor U4191 (N_4191,N_3452,N_3725);
nand U4192 (N_4192,N_3680,N_2777);
nor U4193 (N_4193,N_2798,N_2582);
and U4194 (N_4194,N_2956,N_2406);
nand U4195 (N_4195,N_3241,N_2236);
nand U4196 (N_4196,N_3508,N_2655);
xnor U4197 (N_4197,N_3002,N_2304);
and U4198 (N_4198,N_2342,N_3723);
nand U4199 (N_4199,N_3664,N_3818);
xnor U4200 (N_4200,N_3233,N_3612);
or U4201 (N_4201,N_3079,N_3975);
or U4202 (N_4202,N_3658,N_3143);
nand U4203 (N_4203,N_2540,N_3672);
and U4204 (N_4204,N_3010,N_2167);
nand U4205 (N_4205,N_2053,N_3554);
nor U4206 (N_4206,N_3880,N_3721);
nand U4207 (N_4207,N_2026,N_3026);
and U4208 (N_4208,N_2679,N_3147);
and U4209 (N_4209,N_3469,N_3697);
nor U4210 (N_4210,N_2587,N_3195);
nand U4211 (N_4211,N_3029,N_2603);
nand U4212 (N_4212,N_3476,N_3379);
xor U4213 (N_4213,N_3784,N_3266);
nand U4214 (N_4214,N_2224,N_3252);
and U4215 (N_4215,N_2503,N_2577);
nor U4216 (N_4216,N_2654,N_2196);
nand U4217 (N_4217,N_2187,N_3866);
nor U4218 (N_4218,N_2561,N_3922);
nor U4219 (N_4219,N_2424,N_2541);
or U4220 (N_4220,N_2315,N_2099);
or U4221 (N_4221,N_3030,N_2975);
nor U4222 (N_4222,N_2005,N_3462);
xor U4223 (N_4223,N_3970,N_2704);
nand U4224 (N_4224,N_2857,N_2435);
nor U4225 (N_4225,N_2300,N_2271);
nand U4226 (N_4226,N_3316,N_3140);
and U4227 (N_4227,N_2705,N_2334);
xnor U4228 (N_4228,N_3881,N_3223);
nand U4229 (N_4229,N_2220,N_3461);
and U4230 (N_4230,N_2974,N_3719);
nor U4231 (N_4231,N_2103,N_3231);
or U4232 (N_4232,N_2557,N_2867);
or U4233 (N_4233,N_2727,N_3865);
and U4234 (N_4234,N_2193,N_3014);
and U4235 (N_4235,N_3229,N_2909);
nor U4236 (N_4236,N_3351,N_3135);
nor U4237 (N_4237,N_3979,N_3209);
nor U4238 (N_4238,N_2040,N_3150);
nor U4239 (N_4239,N_3045,N_3202);
nor U4240 (N_4240,N_3739,N_3637);
or U4241 (N_4241,N_2995,N_3609);
or U4242 (N_4242,N_2287,N_2385);
nor U4243 (N_4243,N_3904,N_2757);
nor U4244 (N_4244,N_2405,N_3213);
xor U4245 (N_4245,N_2086,N_3466);
or U4246 (N_4246,N_2836,N_2112);
nor U4247 (N_4247,N_3581,N_3686);
or U4248 (N_4248,N_2515,N_3724);
xor U4249 (N_4249,N_2227,N_3670);
nor U4250 (N_4250,N_2932,N_2563);
or U4251 (N_4251,N_3743,N_2138);
nor U4252 (N_4252,N_3123,N_3699);
or U4253 (N_4253,N_2341,N_3382);
and U4254 (N_4254,N_2308,N_2434);
nor U4255 (N_4255,N_3102,N_2806);
nor U4256 (N_4256,N_2172,N_3080);
nand U4257 (N_4257,N_2477,N_3873);
nand U4258 (N_4258,N_3835,N_2398);
and U4259 (N_4259,N_2239,N_2672);
and U4260 (N_4260,N_2457,N_3200);
and U4261 (N_4261,N_2761,N_2066);
nand U4262 (N_4262,N_3020,N_2096);
nand U4263 (N_4263,N_2602,N_3457);
nor U4264 (N_4264,N_3623,N_3205);
and U4265 (N_4265,N_3034,N_2547);
nand U4266 (N_4266,N_3551,N_3387);
or U4267 (N_4267,N_2056,N_3248);
or U4268 (N_4268,N_2359,N_2623);
nor U4269 (N_4269,N_2724,N_3945);
or U4270 (N_4270,N_3016,N_3334);
and U4271 (N_4271,N_2594,N_3173);
and U4272 (N_4272,N_2411,N_2165);
nor U4273 (N_4273,N_3824,N_2447);
or U4274 (N_4274,N_2396,N_3965);
nand U4275 (N_4275,N_3008,N_3756);
nor U4276 (N_4276,N_3931,N_2871);
nand U4277 (N_4277,N_3280,N_3024);
xnor U4278 (N_4278,N_2358,N_3941);
and U4279 (N_4279,N_2337,N_2756);
xnor U4280 (N_4280,N_3860,N_3493);
or U4281 (N_4281,N_3897,N_2529);
and U4282 (N_4282,N_3341,N_2109);
nand U4283 (N_4283,N_3526,N_3303);
and U4284 (N_4284,N_3985,N_2532);
and U4285 (N_4285,N_3996,N_2781);
nor U4286 (N_4286,N_2107,N_3238);
and U4287 (N_4287,N_3247,N_2525);
or U4288 (N_4288,N_2027,N_2829);
or U4289 (N_4289,N_3841,N_3710);
and U4290 (N_4290,N_2170,N_3160);
nor U4291 (N_4291,N_2546,N_2615);
or U4292 (N_4292,N_3892,N_3854);
and U4293 (N_4293,N_3124,N_3840);
nand U4294 (N_4294,N_2813,N_3244);
and U4295 (N_4295,N_2402,N_3414);
or U4296 (N_4296,N_2197,N_2560);
and U4297 (N_4297,N_3453,N_2356);
xor U4298 (N_4298,N_2714,N_2216);
nor U4299 (N_4299,N_3651,N_2361);
or U4300 (N_4300,N_3063,N_3671);
or U4301 (N_4301,N_2404,N_3458);
nand U4302 (N_4302,N_3317,N_2247);
nand U4303 (N_4303,N_3103,N_3309);
and U4304 (N_4304,N_2473,N_3242);
and U4305 (N_4305,N_2175,N_3155);
nand U4306 (N_4306,N_3089,N_3846);
nor U4307 (N_4307,N_3182,N_3372);
nor U4308 (N_4308,N_3982,N_2145);
nand U4309 (N_4309,N_2942,N_2355);
nand U4310 (N_4310,N_2012,N_2028);
nand U4311 (N_4311,N_3023,N_2572);
nor U4312 (N_4312,N_3679,N_3594);
or U4313 (N_4313,N_2695,N_2542);
nor U4314 (N_4314,N_2799,N_2970);
nand U4315 (N_4315,N_2038,N_3895);
nor U4316 (N_4316,N_3629,N_3330);
or U4317 (N_4317,N_3956,N_2254);
or U4318 (N_4318,N_2498,N_3092);
or U4319 (N_4319,N_2842,N_3810);
or U4320 (N_4320,N_2448,N_2286);
nor U4321 (N_4321,N_2652,N_2052);
nand U4322 (N_4322,N_3606,N_2928);
nor U4323 (N_4323,N_2873,N_3733);
nor U4324 (N_4324,N_3918,N_2787);
nand U4325 (N_4325,N_2938,N_2804);
or U4326 (N_4326,N_2377,N_3113);
nor U4327 (N_4327,N_2050,N_2601);
or U4328 (N_4328,N_2630,N_3802);
or U4329 (N_4329,N_3129,N_2149);
and U4330 (N_4330,N_3575,N_3577);
and U4331 (N_4331,N_3843,N_2029);
nor U4332 (N_4332,N_2309,N_3750);
or U4333 (N_4333,N_2268,N_2180);
or U4334 (N_4334,N_2158,N_3184);
and U4335 (N_4335,N_3842,N_2759);
nand U4336 (N_4336,N_2228,N_2506);
nor U4337 (N_4337,N_2110,N_2793);
nand U4338 (N_4338,N_3175,N_3258);
nand U4339 (N_4339,N_3888,N_2150);
and U4340 (N_4340,N_2609,N_3618);
nand U4341 (N_4341,N_2025,N_3717);
nor U4342 (N_4342,N_2130,N_2872);
and U4343 (N_4343,N_3673,N_3402);
xnor U4344 (N_4344,N_2595,N_2305);
nand U4345 (N_4345,N_2573,N_3017);
nor U4346 (N_4346,N_3039,N_3522);
and U4347 (N_4347,N_2856,N_2137);
and U4348 (N_4348,N_3022,N_2171);
and U4349 (N_4349,N_2392,N_2075);
or U4350 (N_4350,N_3167,N_3119);
nand U4351 (N_4351,N_2474,N_2371);
nor U4352 (N_4352,N_2834,N_3764);
and U4353 (N_4353,N_3240,N_3060);
or U4354 (N_4354,N_3910,N_2186);
or U4355 (N_4355,N_2629,N_3958);
nand U4356 (N_4356,N_2990,N_3156);
and U4357 (N_4357,N_2098,N_2775);
nor U4358 (N_4358,N_3374,N_2468);
nand U4359 (N_4359,N_3726,N_2715);
nor U4360 (N_4360,N_2260,N_3711);
and U4361 (N_4361,N_2902,N_3270);
and U4362 (N_4362,N_2586,N_3442);
and U4363 (N_4363,N_2530,N_3944);
nand U4364 (N_4364,N_3220,N_3595);
nand U4365 (N_4365,N_2919,N_3816);
nand U4366 (N_4366,N_2088,N_3600);
and U4367 (N_4367,N_2833,N_2350);
nand U4368 (N_4368,N_2148,N_2692);
nand U4369 (N_4369,N_3883,N_2094);
xnor U4370 (N_4370,N_3634,N_2664);
nor U4371 (N_4371,N_3646,N_2472);
or U4372 (N_4372,N_3210,N_2703);
or U4373 (N_4373,N_3328,N_2381);
xor U4374 (N_4374,N_2140,N_3138);
or U4375 (N_4375,N_2329,N_3698);
nor U4376 (N_4376,N_2119,N_3722);
nor U4377 (N_4377,N_2327,N_3278);
nand U4378 (N_4378,N_2658,N_2687);
nor U4379 (N_4379,N_3187,N_3692);
or U4380 (N_4380,N_2467,N_3641);
nand U4381 (N_4381,N_2510,N_3499);
and U4382 (N_4382,N_2980,N_2333);
nand U4383 (N_4383,N_3236,N_3552);
nand U4384 (N_4384,N_3272,N_2348);
xor U4385 (N_4385,N_3386,N_3714);
nand U4386 (N_4386,N_3432,N_3246);
or U4387 (N_4387,N_3800,N_3742);
nand U4388 (N_4388,N_2003,N_2512);
and U4389 (N_4389,N_3449,N_3400);
nor U4390 (N_4390,N_2812,N_2810);
nor U4391 (N_4391,N_2607,N_2688);
nor U4392 (N_4392,N_2559,N_3429);
nand U4393 (N_4393,N_3265,N_2875);
nor U4394 (N_4394,N_2129,N_3127);
nor U4395 (N_4395,N_2250,N_3625);
and U4396 (N_4396,N_3408,N_2588);
nor U4397 (N_4397,N_2486,N_3657);
nor U4398 (N_4398,N_3250,N_2667);
or U4399 (N_4399,N_2370,N_2362);
nor U4400 (N_4400,N_2670,N_3208);
nand U4401 (N_4401,N_2986,N_3913);
or U4402 (N_4402,N_3740,N_2754);
nand U4403 (N_4403,N_2177,N_2079);
or U4404 (N_4404,N_2459,N_3141);
nand U4405 (N_4405,N_2784,N_3758);
nand U4406 (N_4406,N_2764,N_3773);
nand U4407 (N_4407,N_3709,N_2345);
and U4408 (N_4408,N_3098,N_3267);
nand U4409 (N_4409,N_3520,N_2493);
or U4410 (N_4410,N_2678,N_3084);
and U4411 (N_4411,N_2972,N_3312);
nand U4412 (N_4412,N_2032,N_3077);
and U4413 (N_4413,N_2517,N_2665);
or U4414 (N_4414,N_3932,N_2814);
and U4415 (N_4415,N_3578,N_3974);
or U4416 (N_4416,N_3377,N_3314);
nor U4417 (N_4417,N_3291,N_3586);
and U4418 (N_4418,N_3583,N_2495);
or U4419 (N_4419,N_2527,N_3503);
and U4420 (N_4420,N_3689,N_3799);
nand U4421 (N_4421,N_3823,N_3104);
and U4422 (N_4422,N_2668,N_3867);
or U4423 (N_4423,N_3957,N_3287);
nor U4424 (N_4424,N_2006,N_3917);
nor U4425 (N_4425,N_3186,N_3889);
nor U4426 (N_4426,N_3603,N_3075);
nor U4427 (N_4427,N_3536,N_3216);
nor U4428 (N_4428,N_3484,N_2281);
and U4429 (N_4429,N_2870,N_3048);
xnor U4430 (N_4430,N_3748,N_2551);
nor U4431 (N_4431,N_3523,N_2584);
and U4432 (N_4432,N_2780,N_3381);
nand U4433 (N_4433,N_2533,N_3777);
nand U4434 (N_4434,N_3683,N_3347);
and U4435 (N_4435,N_3025,N_3929);
or U4436 (N_4436,N_2779,N_2897);
or U4437 (N_4437,N_2859,N_3640);
nand U4438 (N_4438,N_3798,N_3116);
nor U4439 (N_4439,N_3145,N_3796);
or U4440 (N_4440,N_3994,N_2936);
and U4441 (N_4441,N_2214,N_2063);
nor U4442 (N_4442,N_2624,N_2095);
nor U4443 (N_4443,N_2299,N_2484);
nor U4444 (N_4444,N_3797,N_3878);
xnor U4445 (N_4445,N_2924,N_2478);
or U4446 (N_4446,N_3384,N_2360);
nand U4447 (N_4447,N_3302,N_3434);
nor U4448 (N_4448,N_3318,N_2142);
nand U4449 (N_4449,N_3870,N_2373);
and U4450 (N_4450,N_2939,N_2430);
xor U4451 (N_4451,N_2482,N_2497);
nand U4452 (N_4452,N_2200,N_3392);
xnor U4453 (N_4453,N_3305,N_3423);
nand U4454 (N_4454,N_2782,N_2323);
nor U4455 (N_4455,N_2596,N_2883);
or U4456 (N_4456,N_2252,N_3227);
nand U4457 (N_4457,N_2750,N_3194);
nand U4458 (N_4458,N_2412,N_3428);
nor U4459 (N_4459,N_2089,N_3190);
xnor U4460 (N_4460,N_3380,N_2344);
and U4461 (N_4461,N_2415,N_3630);
and U4462 (N_4462,N_3774,N_3820);
nand U4463 (N_4463,N_3787,N_3057);
or U4464 (N_4464,N_3693,N_3704);
and U4465 (N_4465,N_2458,N_2449);
nor U4466 (N_4466,N_2499,N_2017);
or U4467 (N_4467,N_3033,N_3938);
or U4468 (N_4468,N_3356,N_2031);
and U4469 (N_4469,N_3900,N_3488);
nand U4470 (N_4470,N_2712,N_2576);
xor U4471 (N_4471,N_3919,N_2916);
and U4472 (N_4472,N_3966,N_3631);
or U4473 (N_4473,N_2401,N_2861);
nor U4474 (N_4474,N_3728,N_3849);
xor U4475 (N_4475,N_3276,N_2863);
nor U4476 (N_4476,N_3808,N_2234);
nor U4477 (N_4477,N_3005,N_2997);
nor U4478 (N_4478,N_2291,N_3009);
and U4479 (N_4479,N_3065,N_2740);
or U4480 (N_4480,N_3567,N_3833);
xor U4481 (N_4481,N_2043,N_2606);
nor U4482 (N_4482,N_3040,N_3814);
and U4483 (N_4483,N_2826,N_3668);
and U4484 (N_4484,N_3411,N_2862);
xnor U4485 (N_4485,N_3548,N_2248);
xor U4486 (N_4486,N_2376,N_2469);
or U4487 (N_4487,N_3793,N_3997);
and U4488 (N_4488,N_2651,N_3322);
and U4489 (N_4489,N_3489,N_2721);
nor U4490 (N_4490,N_2316,N_2440);
nor U4491 (N_4491,N_3085,N_3154);
nor U4492 (N_4492,N_3193,N_3707);
nand U4493 (N_4493,N_2881,N_2792);
nor U4494 (N_4494,N_3557,N_2556);
or U4495 (N_4495,N_3789,N_3514);
nor U4496 (N_4496,N_2716,N_2243);
xor U4497 (N_4497,N_2183,N_2748);
or U4498 (N_4498,N_2830,N_2805);
or U4499 (N_4499,N_3364,N_3759);
nand U4500 (N_4500,N_2274,N_3954);
nor U4501 (N_4501,N_2637,N_2908);
nand U4502 (N_4502,N_3443,N_2702);
xnor U4503 (N_4503,N_2796,N_2069);
and U4504 (N_4504,N_2375,N_3983);
nor U4505 (N_4505,N_3616,N_2689);
nand U4506 (N_4506,N_3871,N_2934);
nor U4507 (N_4507,N_2693,N_3934);
xnor U4508 (N_4508,N_3779,N_3925);
nor U4509 (N_4509,N_2788,N_3282);
or U4510 (N_4510,N_2335,N_2828);
xor U4511 (N_4511,N_2416,N_3390);
or U4512 (N_4512,N_2369,N_2520);
xor U4513 (N_4513,N_2627,N_2683);
or U4514 (N_4514,N_2133,N_3827);
and U4515 (N_4515,N_2090,N_2708);
nor U4516 (N_4516,N_3100,N_2644);
and U4517 (N_4517,N_2906,N_2544);
nor U4518 (N_4518,N_2019,N_3315);
nand U4519 (N_4519,N_3354,N_3339);
xnor U4520 (N_4520,N_3914,N_3481);
and U4521 (N_4521,N_3212,N_2347);
or U4522 (N_4522,N_2611,N_2789);
nand U4523 (N_4523,N_3734,N_3074);
and U4524 (N_4524,N_2747,N_3948);
or U4525 (N_4525,N_2209,N_3862);
or U4526 (N_4526,N_2844,N_2092);
nor U4527 (N_4527,N_3662,N_2521);
or U4528 (N_4528,N_3562,N_3781);
or U4529 (N_4529,N_3527,N_3159);
and U4530 (N_4530,N_3647,N_3500);
nand U4531 (N_4531,N_2619,N_2639);
nor U4532 (N_4532,N_2581,N_3257);
nand U4533 (N_4533,N_3587,N_3851);
and U4534 (N_4534,N_3279,N_2280);
or U4535 (N_4535,N_2951,N_3702);
nor U4536 (N_4536,N_3253,N_3507);
and U4537 (N_4537,N_2583,N_3108);
or U4538 (N_4538,N_3650,N_3968);
xnor U4539 (N_4539,N_2124,N_3986);
xor U4540 (N_4540,N_2625,N_3737);
nand U4541 (N_4541,N_2461,N_3450);
xnor U4542 (N_4542,N_3908,N_2164);
xor U4543 (N_4543,N_3856,N_2680);
xor U4544 (N_4544,N_2659,N_3602);
nor U4545 (N_4545,N_2749,N_2083);
and U4546 (N_4546,N_2940,N_2204);
or U4547 (N_4547,N_2135,N_3448);
xnor U4548 (N_4548,N_2198,N_3588);
or U4549 (N_4549,N_3891,N_2453);
or U4550 (N_4550,N_2684,N_3117);
or U4551 (N_4551,N_2681,N_3902);
or U4552 (N_4552,N_2879,N_2492);
nor U4553 (N_4553,N_2568,N_2346);
or U4554 (N_4554,N_3226,N_2979);
xor U4555 (N_4555,N_2330,N_2874);
and U4556 (N_4556,N_3655,N_3727);
or U4557 (N_4557,N_2394,N_3953);
xnor U4558 (N_4558,N_2015,N_2108);
and U4559 (N_4559,N_2470,N_3576);
and U4560 (N_4560,N_2643,N_3701);
nand U4561 (N_4561,N_3128,N_2232);
nand U4562 (N_4562,N_3199,N_2265);
xnor U4563 (N_4563,N_3401,N_2009);
or U4564 (N_4564,N_2686,N_2303);
and U4565 (N_4565,N_3882,N_3677);
nor U4566 (N_4566,N_3565,N_3999);
xnor U4567 (N_4567,N_2450,N_2593);
nand U4568 (N_4568,N_2123,N_2065);
or U4569 (N_4569,N_2378,N_3006);
xor U4570 (N_4570,N_2297,N_2825);
and U4571 (N_4571,N_2044,N_3950);
or U4572 (N_4572,N_2097,N_3694);
nor U4573 (N_4573,N_3534,N_2731);
nor U4574 (N_4574,N_3636,N_2384);
nand U4575 (N_4575,N_3352,N_2231);
nand U4576 (N_4576,N_2037,N_3494);
xnor U4577 (N_4577,N_3180,N_2985);
xnor U4578 (N_4578,N_3393,N_2054);
nand U4579 (N_4579,N_2913,N_2852);
xor U4580 (N_4580,N_3483,N_3426);
xor U4581 (N_4581,N_3281,N_3930);
xnor U4582 (N_4582,N_3653,N_3732);
and U4583 (N_4583,N_2677,N_2045);
or U4584 (N_4584,N_2071,N_2725);
nand U4585 (N_4585,N_2136,N_2445);
nor U4586 (N_4586,N_2797,N_3815);
and U4587 (N_4587,N_2242,N_3416);
nand U4588 (N_4588,N_2948,N_3148);
nor U4589 (N_4589,N_3501,N_3136);
nor U4590 (N_4590,N_2640,N_2785);
nand U4591 (N_4591,N_3505,N_3288);
and U4592 (N_4592,N_3340,N_2379);
xor U4593 (N_4593,N_3296,N_3924);
or U4594 (N_4594,N_3042,N_2891);
or U4595 (N_4595,N_3964,N_2752);
or U4596 (N_4596,N_2988,N_2548);
and U4597 (N_4597,N_2965,N_3407);
and U4598 (N_4598,N_2790,N_3715);
xor U4599 (N_4599,N_2203,N_2730);
nor U4600 (N_4600,N_3511,N_2225);
or U4601 (N_4601,N_3512,N_3998);
or U4602 (N_4602,N_3822,N_3532);
and U4603 (N_4603,N_2735,N_3149);
nor U4604 (N_4604,N_3419,N_3937);
and U4605 (N_4605,N_2041,N_3395);
nor U4606 (N_4606,N_2391,N_3936);
or U4607 (N_4607,N_2104,N_3942);
or U4608 (N_4608,N_2996,N_2163);
and U4609 (N_4609,N_3307,N_3884);
nand U4610 (N_4610,N_3162,N_2987);
nand U4611 (N_4611,N_2155,N_3663);
xnor U4612 (N_4612,N_3821,N_2463);
nand U4613 (N_4613,N_3736,N_2922);
or U4614 (N_4614,N_3477,N_3585);
or U4615 (N_4615,N_3363,N_2628);
xor U4616 (N_4616,N_3366,N_3441);
and U4617 (N_4617,N_3656,N_2169);
nand U4618 (N_4618,N_3681,N_2531);
and U4619 (N_4619,N_2114,N_3358);
and U4620 (N_4620,N_3605,N_3972);
or U4621 (N_4621,N_3336,N_2352);
xor U4622 (N_4622,N_2320,N_3438);
or U4623 (N_4623,N_2935,N_3189);
xnor U4624 (N_4624,N_2770,N_3976);
nor U4625 (N_4625,N_3845,N_2000);
nor U4626 (N_4626,N_3378,N_2783);
nand U4627 (N_4627,N_3874,N_3614);
nor U4628 (N_4628,N_3059,N_2374);
nor U4629 (N_4629,N_3133,N_2885);
nor U4630 (N_4630,N_2253,N_3070);
nor U4631 (N_4631,N_2794,N_2964);
or U4632 (N_4632,N_2507,N_2156);
nor U4633 (N_4633,N_3943,N_2417);
nand U4634 (N_4634,N_3886,N_3260);
nand U4635 (N_4635,N_3529,N_3805);
and U4636 (N_4636,N_2694,N_3487);
xnor U4637 (N_4637,N_3608,N_2589);
and U4638 (N_4638,N_3172,N_2439);
xor U4639 (N_4639,N_3290,N_2386);
nor U4640 (N_4640,N_2751,N_2322);
nand U4641 (N_4641,N_2277,N_2565);
and U4642 (N_4642,N_2722,N_3479);
nand U4643 (N_4643,N_2691,N_3920);
or U4644 (N_4644,N_2413,N_2898);
and U4645 (N_4645,N_3121,N_2443);
nand U4646 (N_4646,N_3598,N_3531);
xor U4647 (N_4647,N_2418,N_3062);
nor U4648 (N_4648,N_3607,N_2929);
or U4649 (N_4649,N_3170,N_2513);
nand U4650 (N_4650,N_3746,N_3169);
nor U4651 (N_4651,N_3399,N_2087);
nor U4652 (N_4652,N_3644,N_3584);
or U4653 (N_4653,N_2613,N_2543);
or U4654 (N_4654,N_3359,N_2566);
or U4655 (N_4655,N_2626,N_3361);
xnor U4656 (N_4656,N_3695,N_2592);
and U4657 (N_4657,N_2508,N_3464);
nand U4658 (N_4658,N_3437,N_2237);
nor U4659 (N_4659,N_3961,N_3898);
nand U4660 (N_4660,N_3365,N_3178);
nand U4661 (N_4661,N_3454,N_2837);
nand U4662 (N_4662,N_2055,N_2555);
nor U4663 (N_4663,N_2907,N_3417);
xnor U4664 (N_4664,N_2403,N_3369);
xor U4665 (N_4665,N_3243,N_3096);
nor U4666 (N_4666,N_2428,N_3064);
nand U4667 (N_4667,N_2848,N_3539);
and U4668 (N_4668,N_2420,N_2128);
or U4669 (N_4669,N_2481,N_3890);
and U4670 (N_4670,N_2635,N_3518);
nor U4671 (N_4671,N_2918,N_3872);
and U4672 (N_4672,N_2207,N_3114);
or U4673 (N_4673,N_3642,N_2899);
nand U4674 (N_4674,N_2553,N_2324);
nor U4675 (N_4675,N_2850,N_2738);
xor U4676 (N_4676,N_3158,N_3068);
nand U4677 (N_4677,N_2276,N_2726);
nand U4678 (N_4678,N_2190,N_2105);
nand U4679 (N_4679,N_3176,N_2511);
or U4680 (N_4680,N_3593,N_3110);
or U4681 (N_4681,N_2538,N_2967);
or U4682 (N_4682,N_3632,N_2219);
and U4683 (N_4683,N_3335,N_2016);
nor U4684 (N_4684,N_3112,N_3751);
nand U4685 (N_4685,N_2851,N_3370);
nand U4686 (N_4686,N_2064,N_3067);
and U4687 (N_4687,N_3817,N_3896);
nand U4688 (N_4688,N_3903,N_2422);
nand U4689 (N_4689,N_3012,N_3072);
and U4690 (N_4690,N_3804,N_3097);
or U4691 (N_4691,N_3550,N_3519);
nor U4692 (N_4692,N_2262,N_2719);
nor U4693 (N_4693,N_2591,N_3885);
or U4694 (N_4694,N_3713,N_3295);
and U4695 (N_4695,N_2460,N_3790);
and U4696 (N_4696,N_3201,N_3597);
xor U4697 (N_4697,N_3451,N_3362);
nand U4698 (N_4698,N_3475,N_3111);
nor U4699 (N_4699,N_3988,N_2115);
nor U4700 (N_4700,N_3757,N_2244);
or U4701 (N_4701,N_2991,N_2230);
or U4702 (N_4702,N_3174,N_2866);
nor U4703 (N_4703,N_3058,N_2245);
xor U4704 (N_4704,N_2820,N_2622);
or U4705 (N_4705,N_2663,N_2208);
nor U4706 (N_4706,N_2084,N_2769);
nand U4707 (N_4707,N_3007,N_2042);
and U4708 (N_4708,N_2771,N_2811);
or U4709 (N_4709,N_2389,N_3394);
and U4710 (N_4710,N_3706,N_3478);
nor U4711 (N_4711,N_2982,N_2710);
and U4712 (N_4712,N_2023,N_2896);
and U4713 (N_4713,N_3099,N_3752);
nand U4714 (N_4714,N_2387,N_2057);
nor U4715 (N_4715,N_2737,N_2091);
nor U4716 (N_4716,N_2179,N_2960);
nand U4717 (N_4717,N_3041,N_3852);
and U4718 (N_4718,N_2073,N_2317);
nor U4719 (N_4719,N_2945,N_3185);
and U4720 (N_4720,N_2817,N_2564);
nor U4721 (N_4721,N_3230,N_2390);
xnor U4722 (N_4722,N_2791,N_2847);
nor U4723 (N_4723,N_3355,N_3558);
nand U4724 (N_4724,N_2698,N_3061);
nor U4725 (N_4725,N_3542,N_3807);
or U4726 (N_4726,N_3289,N_3249);
and U4727 (N_4727,N_3331,N_2835);
nor U4728 (N_4728,N_3346,N_2256);
nand U4729 (N_4729,N_2674,N_3214);
nand U4730 (N_4730,N_2441,N_3344);
nor U4731 (N_4731,N_3850,N_3621);
or U4732 (N_4732,N_3682,N_2911);
or U4733 (N_4733,N_3788,N_3073);
xnor U4734 (N_4734,N_2022,N_2661);
or U4735 (N_4735,N_2807,N_3198);
and U4736 (N_4736,N_3735,N_2030);
and U4737 (N_4737,N_2950,N_3708);
xor U4738 (N_4738,N_3222,N_3939);
xnor U4739 (N_4739,N_3830,N_3947);
xnor U4740 (N_4740,N_2002,N_2058);
and U4741 (N_4741,N_3165,N_2372);
or U4742 (N_4742,N_3251,N_2638);
nor U4743 (N_4743,N_2295,N_3502);
nor U4744 (N_4744,N_3440,N_2021);
and U4745 (N_4745,N_3375,N_2266);
or U4746 (N_4746,N_3991,N_2259);
nor U4747 (N_4747,N_2288,N_2279);
nand U4748 (N_4748,N_3373,N_2534);
and U4749 (N_4749,N_2931,N_2035);
and U4750 (N_4750,N_2860,N_3911);
nand U4751 (N_4751,N_2464,N_2010);
and U4752 (N_4752,N_2174,N_3293);
or U4753 (N_4753,N_3433,N_3775);
and U4754 (N_4754,N_2575,N_3015);
or U4755 (N_4755,N_3446,N_3660);
nand U4756 (N_4756,N_2739,N_3217);
or U4757 (N_4757,N_3659,N_2310);
or U4758 (N_4758,N_2018,N_2893);
and U4759 (N_4759,N_2120,N_3183);
nor U4760 (N_4760,N_3720,N_3765);
nor U4761 (N_4761,N_2366,N_3963);
and U4762 (N_4762,N_3899,N_3125);
or U4763 (N_4763,N_2014,N_3345);
nor U4764 (N_4764,N_2307,N_2958);
nand U4765 (N_4765,N_3803,N_3485);
and U4766 (N_4766,N_3989,N_3839);
nand U4767 (N_4767,N_3977,N_2671);
and U4768 (N_4768,N_3940,N_3960);
or U4769 (N_4769,N_3263,N_3146);
nor U4770 (N_4770,N_3004,N_2971);
and U4771 (N_4771,N_2117,N_3741);
and U4772 (N_4772,N_3754,N_3013);
and U4773 (N_4773,N_2353,N_3834);
and U4774 (N_4774,N_2733,N_2321);
and U4775 (N_4775,N_2840,N_2465);
xor U4776 (N_4776,N_3460,N_2351);
nand U4777 (N_4777,N_3245,N_2212);
xor U4778 (N_4778,N_3971,N_3801);
or U4779 (N_4779,N_2311,N_3993);
nor U4780 (N_4780,N_2168,N_2205);
or U4781 (N_4781,N_2616,N_2776);
nand U4782 (N_4782,N_2496,N_2802);
nor U4783 (N_4783,N_2822,N_3794);
and U4784 (N_4784,N_3504,N_2388);
nor U4785 (N_4785,N_2537,N_2912);
xnor U4786 (N_4786,N_3601,N_2192);
nor U4787 (N_4787,N_2476,N_2301);
or U4788 (N_4788,N_3350,N_3549);
and U4789 (N_4789,N_2062,N_3981);
or U4790 (N_4790,N_3038,N_2338);
xor U4791 (N_4791,N_2116,N_3036);
and U4792 (N_4792,N_3747,N_3844);
or U4793 (N_4793,N_3234,N_3471);
or U4794 (N_4794,N_2233,N_3969);
and U4795 (N_4795,N_3403,N_2631);
xor U4796 (N_4796,N_3613,N_3083);
or U4797 (N_4797,N_2767,N_3269);
and U4798 (N_4798,N_2660,N_2111);
nor U4799 (N_4799,N_3360,N_2312);
nor U4800 (N_4800,N_2569,N_2364);
or U4801 (N_4801,N_3738,N_3412);
and U4802 (N_4802,N_2526,N_2646);
nand U4803 (N_4803,N_2426,N_2669);
and U4804 (N_4804,N_2201,N_3078);
and U4805 (N_4805,N_3617,N_2318);
nor U4806 (N_4806,N_2709,N_3191);
and U4807 (N_4807,N_2466,N_3755);
and U4808 (N_4808,N_3018,N_2485);
nor U4809 (N_4809,N_2249,N_2433);
nand U4810 (N_4810,N_3688,N_3299);
or U4811 (N_4811,N_3177,N_3995);
nand U4812 (N_4812,N_2957,N_2161);
xor U4813 (N_4813,N_3543,N_2325);
or U4814 (N_4814,N_3811,N_3912);
nand U4815 (N_4815,N_3861,N_3368);
nor U4816 (N_4816,N_2800,N_2284);
and U4817 (N_4817,N_3730,N_3513);
or U4818 (N_4818,N_2336,N_2620);
nor U4819 (N_4819,N_3525,N_3391);
nand U4820 (N_4820,N_2746,N_3353);
and U4821 (N_4821,N_2954,N_2326);
xor U4822 (N_4822,N_3894,N_2258);
or U4823 (N_4823,N_2118,N_2903);
xnor U4824 (N_4824,N_2296,N_2059);
nor U4825 (N_4825,N_3980,N_3809);
or U4826 (N_4826,N_2745,N_2865);
nand U4827 (N_4827,N_2267,N_3731);
and U4828 (N_4828,N_3772,N_3604);
nand U4829 (N_4829,N_2653,N_2614);
nand U4830 (N_4830,N_2673,N_3320);
nand U4831 (N_4831,N_2047,N_2880);
nand U4832 (N_4832,N_2185,N_2717);
and U4833 (N_4833,N_2961,N_2983);
nor U4834 (N_4834,N_3868,N_2943);
nand U4835 (N_4835,N_2194,N_2343);
nor U4836 (N_4836,N_3573,N_3848);
and U4837 (N_4837,N_2713,N_3580);
nand U4838 (N_4838,N_3901,N_2229);
nor U4839 (N_4839,N_3768,N_2930);
and U4840 (N_4840,N_2008,N_2080);
nand U4841 (N_4841,N_2853,N_2178);
nor U4842 (N_4842,N_2036,N_3927);
nand U4843 (N_4843,N_2832,N_3037);
nor U4844 (N_4844,N_3569,N_3745);
nand U4845 (N_4845,N_3564,N_2636);
nand U4846 (N_4846,N_3164,N_3915);
xnor U4847 (N_4847,N_2839,N_3044);
nor U4848 (N_4848,N_2882,N_2302);
nand U4849 (N_4849,N_3049,N_3876);
nor U4850 (N_4850,N_2331,N_3371);
or U4851 (N_4851,N_3611,N_2984);
xnor U4852 (N_4852,N_2772,N_3528);
or U4853 (N_4853,N_3859,N_3261);
xor U4854 (N_4854,N_3716,N_2452);
and U4855 (N_4855,N_3832,N_3684);
nor U4856 (N_4856,N_3907,N_2758);
nor U4857 (N_4857,N_2211,N_3262);
and U4858 (N_4858,N_3046,N_2732);
and U4859 (N_4859,N_3256,N_3211);
or U4860 (N_4860,N_3134,N_3524);
nor U4861 (N_4861,N_3847,N_3192);
nor U4862 (N_4862,N_3120,N_3495);
nor U4863 (N_4863,N_2141,N_2855);
and U4864 (N_4864,N_2742,N_3455);
nand U4865 (N_4865,N_3467,N_3761);
nor U4866 (N_4866,N_3349,N_2226);
xor U4867 (N_4867,N_3538,N_3286);
or U4868 (N_4868,N_2567,N_2838);
nor U4869 (N_4869,N_3050,N_2819);
xor U4870 (N_4870,N_3157,N_2718);
nand U4871 (N_4871,N_3306,N_3678);
and U4872 (N_4872,N_3268,N_2173);
or U4873 (N_4873,N_2191,N_3093);
and U4874 (N_4874,N_2423,N_3115);
and U4875 (N_4875,N_2633,N_2471);
and U4876 (N_4876,N_3343,N_2339);
and U4877 (N_4877,N_3151,N_3397);
nand U4878 (N_4878,N_2146,N_2690);
nand U4879 (N_4879,N_3420,N_3254);
nor U4880 (N_4880,N_3987,N_3926);
nand U4881 (N_4881,N_2697,N_3984);
and U4882 (N_4882,N_2550,N_2298);
or U4883 (N_4883,N_3235,N_2579);
nor U4884 (N_4884,N_2182,N_3712);
and U4885 (N_4885,N_2488,N_3338);
nor U4886 (N_4886,N_3492,N_2723);
nor U4887 (N_4887,N_3445,N_2869);
or U4888 (N_4888,N_3933,N_3321);
or U4889 (N_4889,N_3000,N_2854);
nand U4890 (N_4890,N_3275,N_3541);
nor U4891 (N_4891,N_3782,N_3329);
xnor U4892 (N_4892,N_3828,N_3592);
nand U4893 (N_4893,N_3421,N_3628);
nor U4894 (N_4894,N_2858,N_3054);
nor U4895 (N_4895,N_3813,N_3436);
or U4896 (N_4896,N_2766,N_3131);
and U4897 (N_4897,N_2501,N_2328);
or U4898 (N_4898,N_2962,N_3521);
nor U4899 (N_4899,N_3666,N_2289);
xnor U4900 (N_4900,N_2444,N_2367);
and U4901 (N_4901,N_3207,N_3327);
or U4902 (N_4902,N_3574,N_2490);
xnor U4903 (N_4903,N_2319,N_3792);
and U4904 (N_4904,N_3472,N_2803);
nor U4905 (N_4905,N_2060,N_3109);
nand U4906 (N_4906,N_2313,N_2666);
nand U4907 (N_4907,N_2269,N_2734);
nor U4908 (N_4908,N_3294,N_3729);
and U4909 (N_4909,N_2489,N_2518);
or U4910 (N_4910,N_3082,N_2078);
nor U4911 (N_4911,N_3342,N_2101);
and U4912 (N_4912,N_2085,N_2181);
xor U4913 (N_4913,N_3237,N_2519);
and U4914 (N_4914,N_2020,N_3619);
nor U4915 (N_4915,N_3633,N_3470);
nor U4916 (N_4916,N_3510,N_2904);
or U4917 (N_4917,N_2202,N_3221);
and U4918 (N_4918,N_2251,N_2998);
nor U4919 (N_4919,N_3763,N_3831);
and U4920 (N_4920,N_2823,N_2395);
and U4921 (N_4921,N_2121,N_3066);
nand U4922 (N_4922,N_3171,N_2051);
or U4923 (N_4923,N_3463,N_3669);
nand U4924 (N_4924,N_2953,N_2004);
nand U4925 (N_4925,N_2999,N_2001);
nand U4926 (N_4926,N_2455,N_3615);
xor U4927 (N_4927,N_3277,N_2921);
nand U4928 (N_4928,N_3389,N_2645);
and U4929 (N_4929,N_2989,N_2397);
or U4930 (N_4930,N_3591,N_2024);
or U4931 (N_4931,N_2729,N_3422);
nor U4932 (N_4932,N_3563,N_3665);
nor U4933 (N_4933,N_2915,N_3313);
or U4934 (N_4934,N_2442,N_2068);
nor U4935 (N_4935,N_3388,N_3474);
nor U4936 (N_4936,N_3232,N_3480);
nand U4937 (N_4937,N_2662,N_2081);
or U4938 (N_4938,N_3032,N_2491);
or U4939 (N_4939,N_2978,N_2768);
nor U4940 (N_4940,N_2184,N_2235);
and U4941 (N_4941,N_2590,N_2223);
and U4942 (N_4942,N_2570,N_2270);
nand U4943 (N_4943,N_3439,N_3118);
and U4944 (N_4944,N_2963,N_3152);
nand U4945 (N_4945,N_2446,N_2106);
or U4946 (N_4946,N_3935,N_3285);
nor U4947 (N_4947,N_2755,N_3515);
or U4948 (N_4948,N_2959,N_3181);
xnor U4949 (N_4949,N_3425,N_2927);
nor U4950 (N_4950,N_2642,N_3163);
and U4951 (N_4951,N_3168,N_2849);
xor U4952 (N_4952,N_3228,N_3638);
xnor U4953 (N_4953,N_2480,N_3409);
and U4954 (N_4954,N_2159,N_3496);
xor U4955 (N_4955,N_2549,N_2400);
nor U4956 (N_4956,N_3509,N_3770);
nand U4957 (N_4957,N_3553,N_3624);
xnor U4958 (N_4958,N_2263,N_2240);
nand U4959 (N_4959,N_2290,N_3319);
and U4960 (N_4960,N_2977,N_3431);
nor U4961 (N_4961,N_3310,N_2585);
or U4962 (N_4962,N_3130,N_2648);
or U4963 (N_4963,N_2801,N_2728);
or U4964 (N_4964,N_2966,N_2824);
and U4965 (N_4965,N_3106,N_3675);
nor U4966 (N_4966,N_3274,N_2188);
and U4967 (N_4967,N_3239,N_2067);
or U4968 (N_4968,N_2864,N_3383);
xnor U4969 (N_4969,N_2516,N_3990);
nand U4970 (N_4970,N_2720,N_2429);
xnor U4971 (N_4971,N_3819,N_3418);
or U4972 (N_4972,N_2368,N_3829);
or U4973 (N_4973,N_2285,N_3864);
or U4974 (N_4974,N_2707,N_3273);
or U4975 (N_4975,N_3091,N_2558);
xnor U4976 (N_4976,N_2456,N_3579);
and U4977 (N_4977,N_3076,N_2332);
nor U4978 (N_4978,N_3762,N_3877);
nand U4979 (N_4979,N_3533,N_3718);
or U4980 (N_4980,N_2955,N_2612);
nor U4981 (N_4981,N_3224,N_3795);
nand U4982 (N_4982,N_2437,N_2941);
nor U4983 (N_4983,N_3535,N_3685);
nand U4984 (N_4984,N_3858,N_2272);
nand U4985 (N_4985,N_2264,N_2578);
nand U4986 (N_4986,N_2816,N_3398);
nand U4987 (N_4987,N_3413,N_3785);
or U4988 (N_4988,N_3517,N_3153);
nand U4989 (N_4989,N_3255,N_3326);
or U4990 (N_4990,N_2074,N_2571);
or U4991 (N_4991,N_2143,N_2215);
and U4992 (N_4992,N_2257,N_3204);
nor U4993 (N_4993,N_2773,N_3946);
or U4994 (N_4994,N_2199,N_2438);
nand U4995 (N_4995,N_2843,N_2649);
and U4996 (N_4996,N_2048,N_3916);
or U4997 (N_4997,N_2699,N_3620);
or U4998 (N_4998,N_3766,N_2841);
and U4999 (N_4999,N_2952,N_3283);
xor U5000 (N_5000,N_2354,N_2454);
nand U5001 (N_5001,N_2898,N_3065);
xnor U5002 (N_5002,N_2154,N_2763);
nand U5003 (N_5003,N_2635,N_2325);
and U5004 (N_5004,N_3326,N_2718);
nor U5005 (N_5005,N_3047,N_3358);
and U5006 (N_5006,N_3980,N_3581);
nand U5007 (N_5007,N_2757,N_2434);
and U5008 (N_5008,N_3076,N_3664);
or U5009 (N_5009,N_3304,N_2087);
nor U5010 (N_5010,N_3118,N_2277);
nor U5011 (N_5011,N_3318,N_2539);
or U5012 (N_5012,N_2198,N_3662);
nor U5013 (N_5013,N_2173,N_3849);
or U5014 (N_5014,N_3897,N_3701);
and U5015 (N_5015,N_3776,N_2012);
nor U5016 (N_5016,N_3836,N_3999);
nor U5017 (N_5017,N_3313,N_2914);
or U5018 (N_5018,N_3937,N_3659);
xnor U5019 (N_5019,N_3262,N_2176);
nand U5020 (N_5020,N_2900,N_2566);
nand U5021 (N_5021,N_2338,N_2154);
and U5022 (N_5022,N_3337,N_3574);
and U5023 (N_5023,N_2380,N_3157);
or U5024 (N_5024,N_2798,N_2688);
or U5025 (N_5025,N_3571,N_2849);
and U5026 (N_5026,N_3032,N_3193);
xor U5027 (N_5027,N_3763,N_3263);
nor U5028 (N_5028,N_3017,N_2968);
nand U5029 (N_5029,N_3496,N_2504);
nand U5030 (N_5030,N_2349,N_3742);
xnor U5031 (N_5031,N_3756,N_3918);
xor U5032 (N_5032,N_3265,N_3585);
nand U5033 (N_5033,N_2395,N_2504);
nand U5034 (N_5034,N_2569,N_2725);
nand U5035 (N_5035,N_2874,N_2154);
nor U5036 (N_5036,N_2922,N_3433);
or U5037 (N_5037,N_2046,N_2631);
and U5038 (N_5038,N_2572,N_2201);
nor U5039 (N_5039,N_2038,N_3927);
nand U5040 (N_5040,N_2544,N_3598);
nor U5041 (N_5041,N_2599,N_2626);
nand U5042 (N_5042,N_2074,N_2529);
nand U5043 (N_5043,N_3425,N_3555);
nand U5044 (N_5044,N_2070,N_3046);
and U5045 (N_5045,N_3237,N_3154);
nand U5046 (N_5046,N_2661,N_3872);
nand U5047 (N_5047,N_3575,N_2217);
or U5048 (N_5048,N_3309,N_3868);
or U5049 (N_5049,N_2045,N_2208);
or U5050 (N_5050,N_3501,N_2344);
nand U5051 (N_5051,N_3026,N_3707);
nor U5052 (N_5052,N_3930,N_2976);
xnor U5053 (N_5053,N_2633,N_3674);
or U5054 (N_5054,N_2449,N_2689);
and U5055 (N_5055,N_2954,N_3139);
xor U5056 (N_5056,N_3360,N_2332);
and U5057 (N_5057,N_2975,N_3980);
and U5058 (N_5058,N_2277,N_3442);
nor U5059 (N_5059,N_3676,N_2845);
nand U5060 (N_5060,N_3240,N_3036);
nand U5061 (N_5061,N_2272,N_3970);
nor U5062 (N_5062,N_3962,N_3522);
or U5063 (N_5063,N_2635,N_3464);
or U5064 (N_5064,N_2218,N_3009);
nor U5065 (N_5065,N_3196,N_2489);
nor U5066 (N_5066,N_3987,N_3886);
and U5067 (N_5067,N_2432,N_3506);
nand U5068 (N_5068,N_3241,N_3507);
nand U5069 (N_5069,N_2777,N_2328);
nand U5070 (N_5070,N_3823,N_3155);
and U5071 (N_5071,N_3807,N_3587);
nor U5072 (N_5072,N_3619,N_3541);
and U5073 (N_5073,N_2956,N_3974);
nand U5074 (N_5074,N_3234,N_3443);
nor U5075 (N_5075,N_3193,N_2678);
or U5076 (N_5076,N_2656,N_3745);
xor U5077 (N_5077,N_3140,N_3565);
nor U5078 (N_5078,N_3325,N_3249);
nor U5079 (N_5079,N_3051,N_2674);
and U5080 (N_5080,N_3937,N_3932);
xor U5081 (N_5081,N_2632,N_3628);
nand U5082 (N_5082,N_2701,N_2118);
or U5083 (N_5083,N_2059,N_3374);
nor U5084 (N_5084,N_2366,N_2552);
xnor U5085 (N_5085,N_3386,N_3510);
and U5086 (N_5086,N_2528,N_3997);
nand U5087 (N_5087,N_3967,N_3348);
or U5088 (N_5088,N_2270,N_2387);
or U5089 (N_5089,N_2006,N_3453);
nand U5090 (N_5090,N_3355,N_2433);
xnor U5091 (N_5091,N_2278,N_3255);
and U5092 (N_5092,N_3347,N_2230);
nor U5093 (N_5093,N_2292,N_3711);
and U5094 (N_5094,N_3004,N_3054);
nor U5095 (N_5095,N_3114,N_2317);
nand U5096 (N_5096,N_3973,N_3653);
nor U5097 (N_5097,N_2041,N_2492);
nor U5098 (N_5098,N_2026,N_2988);
nor U5099 (N_5099,N_2692,N_2200);
and U5100 (N_5100,N_2832,N_3739);
nand U5101 (N_5101,N_2072,N_3286);
or U5102 (N_5102,N_3057,N_2868);
nor U5103 (N_5103,N_3088,N_3905);
and U5104 (N_5104,N_2010,N_3159);
nor U5105 (N_5105,N_2484,N_2470);
xnor U5106 (N_5106,N_3911,N_2952);
nor U5107 (N_5107,N_3709,N_3584);
xnor U5108 (N_5108,N_2727,N_3105);
and U5109 (N_5109,N_2710,N_3284);
or U5110 (N_5110,N_2177,N_2767);
nor U5111 (N_5111,N_2372,N_2221);
nor U5112 (N_5112,N_2261,N_3525);
and U5113 (N_5113,N_3696,N_3019);
or U5114 (N_5114,N_2523,N_3265);
nand U5115 (N_5115,N_2519,N_3260);
or U5116 (N_5116,N_3177,N_2405);
or U5117 (N_5117,N_2128,N_3971);
or U5118 (N_5118,N_3974,N_3549);
or U5119 (N_5119,N_3234,N_3066);
xnor U5120 (N_5120,N_2863,N_3024);
and U5121 (N_5121,N_3954,N_2087);
nand U5122 (N_5122,N_3753,N_3109);
nand U5123 (N_5123,N_2737,N_3740);
nand U5124 (N_5124,N_3436,N_3073);
and U5125 (N_5125,N_3563,N_2975);
nand U5126 (N_5126,N_3132,N_2391);
or U5127 (N_5127,N_3319,N_2636);
and U5128 (N_5128,N_2350,N_3517);
xnor U5129 (N_5129,N_2438,N_2671);
nor U5130 (N_5130,N_2367,N_3689);
nor U5131 (N_5131,N_3445,N_3294);
nand U5132 (N_5132,N_2548,N_3966);
nand U5133 (N_5133,N_2251,N_3079);
nor U5134 (N_5134,N_3890,N_2811);
nand U5135 (N_5135,N_2703,N_3371);
or U5136 (N_5136,N_2073,N_2443);
nand U5137 (N_5137,N_2868,N_3271);
or U5138 (N_5138,N_3415,N_3428);
nor U5139 (N_5139,N_2160,N_3842);
nor U5140 (N_5140,N_2082,N_2950);
and U5141 (N_5141,N_2564,N_3295);
xor U5142 (N_5142,N_3735,N_3185);
nor U5143 (N_5143,N_2050,N_3242);
nand U5144 (N_5144,N_2976,N_3470);
xnor U5145 (N_5145,N_3917,N_3982);
and U5146 (N_5146,N_2115,N_2273);
or U5147 (N_5147,N_2983,N_2030);
xnor U5148 (N_5148,N_3049,N_3028);
and U5149 (N_5149,N_3946,N_2013);
nand U5150 (N_5150,N_3180,N_2947);
nand U5151 (N_5151,N_3335,N_2981);
or U5152 (N_5152,N_2848,N_3827);
nand U5153 (N_5153,N_3963,N_3474);
and U5154 (N_5154,N_3752,N_2291);
nand U5155 (N_5155,N_3146,N_2634);
nor U5156 (N_5156,N_3882,N_2728);
and U5157 (N_5157,N_2258,N_2635);
nor U5158 (N_5158,N_3115,N_2906);
nand U5159 (N_5159,N_2992,N_2613);
nand U5160 (N_5160,N_2969,N_2734);
nor U5161 (N_5161,N_2324,N_3508);
xnor U5162 (N_5162,N_3604,N_3080);
or U5163 (N_5163,N_3075,N_2645);
and U5164 (N_5164,N_2313,N_3280);
nor U5165 (N_5165,N_3985,N_2195);
nand U5166 (N_5166,N_2880,N_2608);
or U5167 (N_5167,N_3238,N_2090);
and U5168 (N_5168,N_2413,N_3057);
and U5169 (N_5169,N_2789,N_2791);
or U5170 (N_5170,N_3657,N_2675);
nor U5171 (N_5171,N_3751,N_2993);
nor U5172 (N_5172,N_3216,N_2674);
xnor U5173 (N_5173,N_2255,N_2310);
nand U5174 (N_5174,N_3572,N_2257);
nor U5175 (N_5175,N_2584,N_3625);
nor U5176 (N_5176,N_2213,N_3871);
or U5177 (N_5177,N_3972,N_2875);
nand U5178 (N_5178,N_3256,N_3678);
nor U5179 (N_5179,N_3454,N_2458);
and U5180 (N_5180,N_3359,N_3046);
and U5181 (N_5181,N_3176,N_2395);
nand U5182 (N_5182,N_2906,N_2322);
xnor U5183 (N_5183,N_3405,N_3727);
or U5184 (N_5184,N_2793,N_2278);
nand U5185 (N_5185,N_3180,N_2574);
nand U5186 (N_5186,N_3409,N_3324);
and U5187 (N_5187,N_2296,N_3377);
and U5188 (N_5188,N_3699,N_3080);
nor U5189 (N_5189,N_3070,N_2135);
and U5190 (N_5190,N_2286,N_2504);
and U5191 (N_5191,N_3972,N_2008);
or U5192 (N_5192,N_2606,N_3414);
xor U5193 (N_5193,N_2252,N_3839);
and U5194 (N_5194,N_3131,N_3233);
or U5195 (N_5195,N_2714,N_3931);
or U5196 (N_5196,N_3694,N_2090);
nand U5197 (N_5197,N_3040,N_3113);
and U5198 (N_5198,N_2285,N_3852);
or U5199 (N_5199,N_2129,N_3844);
nor U5200 (N_5200,N_3039,N_3535);
xnor U5201 (N_5201,N_3105,N_3166);
xor U5202 (N_5202,N_3320,N_2303);
or U5203 (N_5203,N_3611,N_2808);
nand U5204 (N_5204,N_2042,N_2037);
nand U5205 (N_5205,N_2580,N_2385);
and U5206 (N_5206,N_2557,N_3977);
or U5207 (N_5207,N_2677,N_3898);
or U5208 (N_5208,N_3704,N_3221);
and U5209 (N_5209,N_2996,N_2095);
nor U5210 (N_5210,N_2346,N_2710);
nor U5211 (N_5211,N_3847,N_2244);
xor U5212 (N_5212,N_2807,N_2792);
nor U5213 (N_5213,N_2289,N_2786);
nand U5214 (N_5214,N_2620,N_3002);
and U5215 (N_5215,N_2994,N_3173);
nor U5216 (N_5216,N_3590,N_2892);
nand U5217 (N_5217,N_2866,N_2036);
nor U5218 (N_5218,N_3086,N_2887);
or U5219 (N_5219,N_3835,N_3378);
and U5220 (N_5220,N_3262,N_3564);
nand U5221 (N_5221,N_2649,N_3251);
or U5222 (N_5222,N_3051,N_2875);
and U5223 (N_5223,N_2037,N_3690);
and U5224 (N_5224,N_3609,N_3952);
nor U5225 (N_5225,N_3812,N_3200);
nand U5226 (N_5226,N_2627,N_3745);
or U5227 (N_5227,N_3301,N_2280);
and U5228 (N_5228,N_3762,N_3576);
nor U5229 (N_5229,N_3275,N_2398);
and U5230 (N_5230,N_3807,N_2813);
nand U5231 (N_5231,N_3378,N_3907);
nor U5232 (N_5232,N_2736,N_3224);
nor U5233 (N_5233,N_2333,N_3971);
or U5234 (N_5234,N_2341,N_3016);
or U5235 (N_5235,N_2308,N_3519);
nand U5236 (N_5236,N_2126,N_2988);
nor U5237 (N_5237,N_2202,N_3591);
nor U5238 (N_5238,N_2025,N_2154);
nand U5239 (N_5239,N_2169,N_2156);
or U5240 (N_5240,N_3384,N_2337);
nor U5241 (N_5241,N_2635,N_2575);
nand U5242 (N_5242,N_3973,N_2638);
and U5243 (N_5243,N_2750,N_2806);
and U5244 (N_5244,N_2530,N_2076);
or U5245 (N_5245,N_3855,N_3587);
nand U5246 (N_5246,N_3561,N_2252);
and U5247 (N_5247,N_3487,N_3829);
or U5248 (N_5248,N_2652,N_3848);
nor U5249 (N_5249,N_3228,N_2824);
nand U5250 (N_5250,N_2356,N_3253);
and U5251 (N_5251,N_2626,N_3942);
and U5252 (N_5252,N_2552,N_3960);
and U5253 (N_5253,N_3553,N_3653);
or U5254 (N_5254,N_2519,N_3972);
nand U5255 (N_5255,N_2909,N_3076);
or U5256 (N_5256,N_3951,N_2279);
and U5257 (N_5257,N_2776,N_2907);
or U5258 (N_5258,N_3576,N_2298);
nor U5259 (N_5259,N_3287,N_2225);
and U5260 (N_5260,N_3067,N_3912);
nor U5261 (N_5261,N_3770,N_3608);
and U5262 (N_5262,N_2762,N_2065);
or U5263 (N_5263,N_3707,N_2585);
nor U5264 (N_5264,N_2418,N_2296);
and U5265 (N_5265,N_3887,N_3540);
nand U5266 (N_5266,N_3385,N_2890);
or U5267 (N_5267,N_2253,N_2288);
or U5268 (N_5268,N_2474,N_2208);
xor U5269 (N_5269,N_3747,N_2956);
and U5270 (N_5270,N_3689,N_2055);
nor U5271 (N_5271,N_3054,N_3373);
or U5272 (N_5272,N_2496,N_3119);
or U5273 (N_5273,N_3793,N_3425);
nor U5274 (N_5274,N_2513,N_3572);
nor U5275 (N_5275,N_2523,N_2018);
xor U5276 (N_5276,N_3374,N_2693);
or U5277 (N_5277,N_3437,N_3388);
or U5278 (N_5278,N_2871,N_3112);
nor U5279 (N_5279,N_2387,N_2673);
nor U5280 (N_5280,N_2793,N_2073);
xnor U5281 (N_5281,N_3549,N_2513);
and U5282 (N_5282,N_3467,N_3766);
nor U5283 (N_5283,N_3149,N_3898);
and U5284 (N_5284,N_2777,N_3935);
nand U5285 (N_5285,N_2527,N_3137);
nand U5286 (N_5286,N_3859,N_3440);
and U5287 (N_5287,N_2758,N_2580);
nor U5288 (N_5288,N_3845,N_2856);
nand U5289 (N_5289,N_3004,N_3508);
xor U5290 (N_5290,N_3219,N_2607);
or U5291 (N_5291,N_3319,N_2381);
or U5292 (N_5292,N_2917,N_2343);
xnor U5293 (N_5293,N_2099,N_2612);
xor U5294 (N_5294,N_2035,N_3307);
nand U5295 (N_5295,N_3485,N_3910);
and U5296 (N_5296,N_3040,N_2506);
nor U5297 (N_5297,N_3297,N_2350);
and U5298 (N_5298,N_2616,N_3821);
nand U5299 (N_5299,N_2680,N_3494);
nor U5300 (N_5300,N_2987,N_3605);
xnor U5301 (N_5301,N_2988,N_2334);
and U5302 (N_5302,N_2294,N_2056);
nor U5303 (N_5303,N_3495,N_3149);
xor U5304 (N_5304,N_3764,N_3048);
nand U5305 (N_5305,N_3476,N_3318);
and U5306 (N_5306,N_2305,N_3119);
or U5307 (N_5307,N_2523,N_2901);
nand U5308 (N_5308,N_3068,N_2717);
or U5309 (N_5309,N_2557,N_3246);
or U5310 (N_5310,N_2191,N_2650);
nand U5311 (N_5311,N_3788,N_2592);
or U5312 (N_5312,N_2767,N_2142);
nand U5313 (N_5313,N_2451,N_3276);
and U5314 (N_5314,N_2518,N_3205);
or U5315 (N_5315,N_2098,N_2418);
nand U5316 (N_5316,N_2754,N_3475);
or U5317 (N_5317,N_3961,N_3685);
nand U5318 (N_5318,N_3574,N_3066);
xnor U5319 (N_5319,N_3470,N_3794);
nand U5320 (N_5320,N_2454,N_2468);
and U5321 (N_5321,N_3202,N_3777);
nand U5322 (N_5322,N_3055,N_3090);
nand U5323 (N_5323,N_3226,N_2673);
nor U5324 (N_5324,N_3511,N_2672);
and U5325 (N_5325,N_3598,N_3962);
nand U5326 (N_5326,N_3760,N_2592);
and U5327 (N_5327,N_3233,N_2276);
or U5328 (N_5328,N_3092,N_3048);
or U5329 (N_5329,N_3783,N_3778);
and U5330 (N_5330,N_3474,N_3797);
nand U5331 (N_5331,N_3675,N_3900);
and U5332 (N_5332,N_3743,N_2824);
nor U5333 (N_5333,N_3296,N_3580);
xor U5334 (N_5334,N_2988,N_3124);
nand U5335 (N_5335,N_2053,N_3832);
nor U5336 (N_5336,N_3105,N_2537);
and U5337 (N_5337,N_3818,N_2925);
nand U5338 (N_5338,N_2781,N_3370);
nor U5339 (N_5339,N_3203,N_3497);
nand U5340 (N_5340,N_2832,N_3433);
or U5341 (N_5341,N_2626,N_3595);
or U5342 (N_5342,N_3396,N_2355);
xor U5343 (N_5343,N_2649,N_2930);
and U5344 (N_5344,N_3261,N_3997);
or U5345 (N_5345,N_2571,N_2358);
and U5346 (N_5346,N_2351,N_2487);
nor U5347 (N_5347,N_3320,N_2208);
nand U5348 (N_5348,N_3098,N_2570);
xnor U5349 (N_5349,N_2481,N_2042);
or U5350 (N_5350,N_2271,N_3986);
or U5351 (N_5351,N_2247,N_2564);
or U5352 (N_5352,N_2526,N_3823);
nand U5353 (N_5353,N_3058,N_3359);
xor U5354 (N_5354,N_3978,N_2030);
nor U5355 (N_5355,N_3198,N_3749);
or U5356 (N_5356,N_2319,N_3643);
or U5357 (N_5357,N_3139,N_3779);
and U5358 (N_5358,N_3788,N_3684);
xnor U5359 (N_5359,N_3587,N_3788);
nand U5360 (N_5360,N_3739,N_3008);
nor U5361 (N_5361,N_3095,N_2819);
or U5362 (N_5362,N_3811,N_2051);
and U5363 (N_5363,N_3700,N_2520);
nor U5364 (N_5364,N_2148,N_3052);
nand U5365 (N_5365,N_3090,N_2325);
and U5366 (N_5366,N_3453,N_2179);
nor U5367 (N_5367,N_2633,N_2984);
nor U5368 (N_5368,N_3394,N_3725);
or U5369 (N_5369,N_2582,N_3997);
nand U5370 (N_5370,N_2913,N_3062);
and U5371 (N_5371,N_2111,N_2802);
nor U5372 (N_5372,N_3608,N_2444);
nand U5373 (N_5373,N_2174,N_2538);
nor U5374 (N_5374,N_3301,N_2269);
nor U5375 (N_5375,N_3050,N_2602);
nand U5376 (N_5376,N_2555,N_2127);
nand U5377 (N_5377,N_2836,N_3172);
xnor U5378 (N_5378,N_3389,N_2677);
nand U5379 (N_5379,N_2343,N_2828);
or U5380 (N_5380,N_3864,N_3488);
xnor U5381 (N_5381,N_3742,N_2381);
nand U5382 (N_5382,N_3356,N_2923);
and U5383 (N_5383,N_2972,N_2462);
nand U5384 (N_5384,N_3344,N_3251);
or U5385 (N_5385,N_2859,N_2509);
xor U5386 (N_5386,N_3831,N_2584);
xnor U5387 (N_5387,N_3193,N_3063);
and U5388 (N_5388,N_3741,N_2787);
nor U5389 (N_5389,N_3578,N_3804);
and U5390 (N_5390,N_3052,N_2641);
nor U5391 (N_5391,N_2803,N_2636);
nor U5392 (N_5392,N_2789,N_3702);
or U5393 (N_5393,N_2579,N_3187);
and U5394 (N_5394,N_3526,N_2323);
xnor U5395 (N_5395,N_2625,N_2855);
nand U5396 (N_5396,N_3057,N_2349);
nand U5397 (N_5397,N_2451,N_2111);
xnor U5398 (N_5398,N_3602,N_2825);
nor U5399 (N_5399,N_3476,N_2105);
nor U5400 (N_5400,N_3722,N_3240);
and U5401 (N_5401,N_3221,N_3346);
and U5402 (N_5402,N_3829,N_3983);
nor U5403 (N_5403,N_2149,N_3167);
or U5404 (N_5404,N_2647,N_2913);
nor U5405 (N_5405,N_3546,N_3438);
nand U5406 (N_5406,N_2112,N_3447);
or U5407 (N_5407,N_3504,N_2475);
or U5408 (N_5408,N_3512,N_2460);
or U5409 (N_5409,N_2755,N_3745);
xnor U5410 (N_5410,N_3478,N_2369);
or U5411 (N_5411,N_3205,N_3616);
nand U5412 (N_5412,N_2771,N_3799);
nor U5413 (N_5413,N_2404,N_3094);
and U5414 (N_5414,N_3210,N_3285);
nand U5415 (N_5415,N_2262,N_2841);
and U5416 (N_5416,N_3302,N_3545);
or U5417 (N_5417,N_2985,N_3705);
and U5418 (N_5418,N_2925,N_2350);
nor U5419 (N_5419,N_3690,N_2122);
or U5420 (N_5420,N_3970,N_3327);
nand U5421 (N_5421,N_2285,N_3074);
nand U5422 (N_5422,N_3125,N_3856);
nand U5423 (N_5423,N_2786,N_3934);
nand U5424 (N_5424,N_3226,N_3855);
nor U5425 (N_5425,N_3482,N_3182);
and U5426 (N_5426,N_3964,N_2912);
nand U5427 (N_5427,N_3938,N_3706);
nor U5428 (N_5428,N_3590,N_3637);
nand U5429 (N_5429,N_2631,N_2270);
xor U5430 (N_5430,N_2473,N_2772);
or U5431 (N_5431,N_2288,N_2190);
nand U5432 (N_5432,N_2471,N_2744);
xnor U5433 (N_5433,N_2249,N_2411);
nand U5434 (N_5434,N_2166,N_2945);
nor U5435 (N_5435,N_2055,N_2164);
nand U5436 (N_5436,N_2032,N_3156);
and U5437 (N_5437,N_2880,N_2454);
nor U5438 (N_5438,N_3967,N_2145);
xor U5439 (N_5439,N_3994,N_3115);
xnor U5440 (N_5440,N_2757,N_3824);
or U5441 (N_5441,N_3960,N_2954);
nor U5442 (N_5442,N_3917,N_3935);
nand U5443 (N_5443,N_3365,N_2234);
and U5444 (N_5444,N_3246,N_2234);
xor U5445 (N_5445,N_3376,N_3021);
or U5446 (N_5446,N_3018,N_3984);
nand U5447 (N_5447,N_3873,N_3357);
and U5448 (N_5448,N_3270,N_2093);
or U5449 (N_5449,N_3383,N_2504);
and U5450 (N_5450,N_3043,N_2991);
xnor U5451 (N_5451,N_2312,N_3662);
or U5452 (N_5452,N_2886,N_2479);
nand U5453 (N_5453,N_3262,N_3749);
nand U5454 (N_5454,N_3568,N_2925);
and U5455 (N_5455,N_2506,N_2982);
xor U5456 (N_5456,N_2751,N_3413);
or U5457 (N_5457,N_2376,N_3370);
nand U5458 (N_5458,N_3760,N_3389);
xnor U5459 (N_5459,N_2451,N_2068);
nor U5460 (N_5460,N_2165,N_2924);
and U5461 (N_5461,N_3141,N_3963);
nor U5462 (N_5462,N_2148,N_3895);
nor U5463 (N_5463,N_3162,N_2839);
nand U5464 (N_5464,N_2109,N_2361);
nor U5465 (N_5465,N_3412,N_2346);
and U5466 (N_5466,N_3591,N_2868);
and U5467 (N_5467,N_2882,N_3271);
xnor U5468 (N_5468,N_3267,N_2213);
or U5469 (N_5469,N_3414,N_3280);
xnor U5470 (N_5470,N_2091,N_2023);
nor U5471 (N_5471,N_2034,N_2287);
nor U5472 (N_5472,N_2636,N_2276);
xnor U5473 (N_5473,N_3319,N_2101);
and U5474 (N_5474,N_2273,N_2566);
nor U5475 (N_5475,N_2373,N_2060);
nor U5476 (N_5476,N_2779,N_2178);
xor U5477 (N_5477,N_2166,N_3743);
or U5478 (N_5478,N_3634,N_3537);
and U5479 (N_5479,N_3571,N_2455);
and U5480 (N_5480,N_2851,N_2158);
and U5481 (N_5481,N_3237,N_2763);
and U5482 (N_5482,N_2384,N_2447);
nor U5483 (N_5483,N_3405,N_3722);
or U5484 (N_5484,N_3900,N_2856);
nand U5485 (N_5485,N_2845,N_3246);
nand U5486 (N_5486,N_2360,N_2042);
or U5487 (N_5487,N_2632,N_3680);
and U5488 (N_5488,N_2551,N_3947);
and U5489 (N_5489,N_2127,N_2783);
and U5490 (N_5490,N_3693,N_2464);
or U5491 (N_5491,N_3330,N_3369);
xor U5492 (N_5492,N_2629,N_3615);
and U5493 (N_5493,N_2538,N_2550);
or U5494 (N_5494,N_2723,N_3419);
or U5495 (N_5495,N_3699,N_2205);
and U5496 (N_5496,N_3761,N_3513);
xor U5497 (N_5497,N_3271,N_3118);
nor U5498 (N_5498,N_3010,N_3826);
or U5499 (N_5499,N_2873,N_3361);
or U5500 (N_5500,N_3877,N_3247);
or U5501 (N_5501,N_3034,N_2796);
and U5502 (N_5502,N_3550,N_3483);
and U5503 (N_5503,N_2498,N_2463);
nand U5504 (N_5504,N_2135,N_3833);
or U5505 (N_5505,N_3204,N_3247);
xor U5506 (N_5506,N_3744,N_3195);
or U5507 (N_5507,N_3988,N_2026);
xor U5508 (N_5508,N_3712,N_3914);
nand U5509 (N_5509,N_2004,N_2159);
nand U5510 (N_5510,N_2844,N_3006);
and U5511 (N_5511,N_2881,N_2687);
or U5512 (N_5512,N_2601,N_3654);
or U5513 (N_5513,N_3229,N_2367);
nand U5514 (N_5514,N_2516,N_2762);
or U5515 (N_5515,N_2978,N_3583);
nor U5516 (N_5516,N_3281,N_2504);
xor U5517 (N_5517,N_2876,N_3271);
and U5518 (N_5518,N_3065,N_2263);
nand U5519 (N_5519,N_3622,N_3116);
nand U5520 (N_5520,N_2067,N_2058);
or U5521 (N_5521,N_2051,N_2189);
or U5522 (N_5522,N_3274,N_2529);
and U5523 (N_5523,N_2173,N_3543);
and U5524 (N_5524,N_3857,N_3917);
nand U5525 (N_5525,N_3366,N_2110);
or U5526 (N_5526,N_3232,N_3114);
nor U5527 (N_5527,N_3273,N_2533);
or U5528 (N_5528,N_2072,N_3614);
and U5529 (N_5529,N_2996,N_2189);
nor U5530 (N_5530,N_2903,N_2386);
nand U5531 (N_5531,N_2319,N_3235);
and U5532 (N_5532,N_2605,N_2009);
or U5533 (N_5533,N_2824,N_3020);
or U5534 (N_5534,N_2680,N_3357);
and U5535 (N_5535,N_2112,N_3057);
nand U5536 (N_5536,N_2586,N_3888);
nand U5537 (N_5537,N_2212,N_2334);
xnor U5538 (N_5538,N_3162,N_2380);
or U5539 (N_5539,N_3331,N_2283);
and U5540 (N_5540,N_2540,N_3852);
or U5541 (N_5541,N_3915,N_2352);
xnor U5542 (N_5542,N_2012,N_3125);
and U5543 (N_5543,N_3512,N_3469);
nor U5544 (N_5544,N_2456,N_2896);
and U5545 (N_5545,N_3185,N_2218);
nand U5546 (N_5546,N_2854,N_3374);
nor U5547 (N_5547,N_3604,N_3841);
and U5548 (N_5548,N_2188,N_2094);
nand U5549 (N_5549,N_3633,N_2361);
or U5550 (N_5550,N_2163,N_2007);
and U5551 (N_5551,N_2264,N_3823);
and U5552 (N_5552,N_3235,N_2790);
and U5553 (N_5553,N_3589,N_2511);
nor U5554 (N_5554,N_2794,N_2739);
xnor U5555 (N_5555,N_2127,N_2106);
nor U5556 (N_5556,N_3614,N_3967);
and U5557 (N_5557,N_3466,N_2454);
xor U5558 (N_5558,N_2954,N_2172);
or U5559 (N_5559,N_2016,N_3518);
or U5560 (N_5560,N_3522,N_3013);
and U5561 (N_5561,N_3547,N_2481);
or U5562 (N_5562,N_3465,N_2082);
and U5563 (N_5563,N_2543,N_2299);
or U5564 (N_5564,N_3155,N_2050);
nor U5565 (N_5565,N_3836,N_3591);
nor U5566 (N_5566,N_2411,N_3769);
or U5567 (N_5567,N_3468,N_3216);
or U5568 (N_5568,N_3039,N_2361);
nor U5569 (N_5569,N_3168,N_2142);
and U5570 (N_5570,N_2291,N_2290);
or U5571 (N_5571,N_3202,N_2526);
nand U5572 (N_5572,N_2358,N_3060);
xnor U5573 (N_5573,N_2789,N_2817);
and U5574 (N_5574,N_3433,N_3012);
xnor U5575 (N_5575,N_2716,N_3306);
nor U5576 (N_5576,N_3540,N_2795);
or U5577 (N_5577,N_3313,N_3710);
nand U5578 (N_5578,N_2877,N_3297);
nor U5579 (N_5579,N_3498,N_2499);
and U5580 (N_5580,N_3283,N_3632);
or U5581 (N_5581,N_2481,N_2835);
nand U5582 (N_5582,N_2853,N_3156);
nand U5583 (N_5583,N_3079,N_3009);
nor U5584 (N_5584,N_3831,N_2624);
or U5585 (N_5585,N_3081,N_2354);
and U5586 (N_5586,N_3449,N_2923);
nand U5587 (N_5587,N_3255,N_2295);
and U5588 (N_5588,N_2391,N_2051);
xnor U5589 (N_5589,N_2506,N_3252);
and U5590 (N_5590,N_2595,N_2327);
and U5591 (N_5591,N_2093,N_3947);
and U5592 (N_5592,N_3848,N_2380);
nand U5593 (N_5593,N_3866,N_2326);
or U5594 (N_5594,N_3799,N_3088);
or U5595 (N_5595,N_2583,N_2910);
nand U5596 (N_5596,N_2458,N_3924);
nand U5597 (N_5597,N_2527,N_3246);
xor U5598 (N_5598,N_3307,N_2522);
nor U5599 (N_5599,N_3547,N_3867);
and U5600 (N_5600,N_3157,N_3163);
or U5601 (N_5601,N_2258,N_3537);
or U5602 (N_5602,N_2501,N_2253);
xor U5603 (N_5603,N_3042,N_3139);
xnor U5604 (N_5604,N_2706,N_3309);
nand U5605 (N_5605,N_3272,N_2355);
nor U5606 (N_5606,N_3187,N_2952);
nor U5607 (N_5607,N_2796,N_2568);
xor U5608 (N_5608,N_2950,N_3582);
nand U5609 (N_5609,N_3104,N_2685);
nor U5610 (N_5610,N_2625,N_2022);
or U5611 (N_5611,N_2170,N_3509);
or U5612 (N_5612,N_2070,N_3128);
and U5613 (N_5613,N_3236,N_2340);
nor U5614 (N_5614,N_3230,N_3868);
xnor U5615 (N_5615,N_3065,N_2480);
or U5616 (N_5616,N_2060,N_3309);
or U5617 (N_5617,N_2870,N_3274);
and U5618 (N_5618,N_3272,N_2154);
nand U5619 (N_5619,N_2293,N_3868);
nand U5620 (N_5620,N_3756,N_2649);
xnor U5621 (N_5621,N_3914,N_2273);
xnor U5622 (N_5622,N_2353,N_3436);
and U5623 (N_5623,N_3464,N_3136);
nand U5624 (N_5624,N_3836,N_2937);
nand U5625 (N_5625,N_2732,N_2022);
nor U5626 (N_5626,N_2303,N_2755);
xor U5627 (N_5627,N_3435,N_3147);
nand U5628 (N_5628,N_3361,N_2570);
and U5629 (N_5629,N_2136,N_3343);
nand U5630 (N_5630,N_3192,N_2452);
and U5631 (N_5631,N_2147,N_3430);
or U5632 (N_5632,N_3428,N_2425);
xor U5633 (N_5633,N_3674,N_3538);
nand U5634 (N_5634,N_2213,N_2459);
nand U5635 (N_5635,N_2821,N_2521);
nand U5636 (N_5636,N_2245,N_2496);
or U5637 (N_5637,N_2713,N_3650);
nand U5638 (N_5638,N_2604,N_3327);
nor U5639 (N_5639,N_3907,N_2121);
and U5640 (N_5640,N_3554,N_2438);
nand U5641 (N_5641,N_2282,N_3744);
or U5642 (N_5642,N_2823,N_3910);
or U5643 (N_5643,N_2326,N_2463);
and U5644 (N_5644,N_2753,N_2190);
nor U5645 (N_5645,N_3765,N_3242);
nand U5646 (N_5646,N_3557,N_3537);
xnor U5647 (N_5647,N_3176,N_2477);
or U5648 (N_5648,N_2695,N_2570);
or U5649 (N_5649,N_3623,N_3637);
nand U5650 (N_5650,N_2048,N_3322);
and U5651 (N_5651,N_3262,N_3962);
or U5652 (N_5652,N_3029,N_2794);
nor U5653 (N_5653,N_3370,N_3477);
nand U5654 (N_5654,N_3124,N_3528);
nand U5655 (N_5655,N_2023,N_3215);
and U5656 (N_5656,N_2901,N_3747);
or U5657 (N_5657,N_3280,N_3764);
or U5658 (N_5658,N_2230,N_2837);
xnor U5659 (N_5659,N_2968,N_2815);
nor U5660 (N_5660,N_3382,N_3794);
and U5661 (N_5661,N_3160,N_2718);
nor U5662 (N_5662,N_2956,N_2710);
nand U5663 (N_5663,N_2022,N_3681);
nand U5664 (N_5664,N_2987,N_3717);
or U5665 (N_5665,N_2179,N_3177);
nor U5666 (N_5666,N_3990,N_3513);
and U5667 (N_5667,N_2353,N_2670);
or U5668 (N_5668,N_3745,N_2104);
nor U5669 (N_5669,N_3056,N_2990);
nor U5670 (N_5670,N_2948,N_3775);
and U5671 (N_5671,N_3140,N_2816);
nor U5672 (N_5672,N_3088,N_2320);
or U5673 (N_5673,N_3416,N_2217);
nand U5674 (N_5674,N_2343,N_2735);
xnor U5675 (N_5675,N_3373,N_3922);
nor U5676 (N_5676,N_2274,N_3595);
and U5677 (N_5677,N_3247,N_3044);
nor U5678 (N_5678,N_3657,N_3519);
and U5679 (N_5679,N_2059,N_3644);
and U5680 (N_5680,N_3999,N_3361);
or U5681 (N_5681,N_2295,N_2998);
and U5682 (N_5682,N_3277,N_2820);
and U5683 (N_5683,N_2168,N_3178);
and U5684 (N_5684,N_3009,N_3922);
xor U5685 (N_5685,N_3479,N_2679);
nor U5686 (N_5686,N_3901,N_3125);
xor U5687 (N_5687,N_2417,N_2677);
or U5688 (N_5688,N_3265,N_3171);
or U5689 (N_5689,N_3582,N_3301);
or U5690 (N_5690,N_3452,N_3033);
nand U5691 (N_5691,N_2675,N_3227);
nand U5692 (N_5692,N_2668,N_2201);
nor U5693 (N_5693,N_3478,N_2076);
and U5694 (N_5694,N_2790,N_3635);
nand U5695 (N_5695,N_2354,N_2018);
or U5696 (N_5696,N_3906,N_3600);
or U5697 (N_5697,N_2459,N_3918);
and U5698 (N_5698,N_3690,N_3330);
nor U5699 (N_5699,N_3112,N_2205);
and U5700 (N_5700,N_2674,N_3039);
and U5701 (N_5701,N_2737,N_2568);
or U5702 (N_5702,N_3488,N_3292);
and U5703 (N_5703,N_3206,N_3812);
nor U5704 (N_5704,N_3801,N_3510);
or U5705 (N_5705,N_3038,N_2057);
nor U5706 (N_5706,N_2505,N_2588);
or U5707 (N_5707,N_2371,N_3130);
or U5708 (N_5708,N_2568,N_2996);
nor U5709 (N_5709,N_3641,N_3990);
nor U5710 (N_5710,N_2026,N_2809);
xor U5711 (N_5711,N_3566,N_3927);
nand U5712 (N_5712,N_2548,N_3946);
and U5713 (N_5713,N_2283,N_2226);
and U5714 (N_5714,N_2940,N_3940);
nor U5715 (N_5715,N_2548,N_3303);
or U5716 (N_5716,N_2874,N_3677);
or U5717 (N_5717,N_2926,N_2662);
and U5718 (N_5718,N_2119,N_2632);
xor U5719 (N_5719,N_3932,N_3723);
nor U5720 (N_5720,N_3485,N_2954);
or U5721 (N_5721,N_3791,N_2057);
xnor U5722 (N_5722,N_2741,N_2637);
and U5723 (N_5723,N_2117,N_2871);
and U5724 (N_5724,N_2741,N_3656);
and U5725 (N_5725,N_3157,N_3274);
and U5726 (N_5726,N_2571,N_2601);
nand U5727 (N_5727,N_3257,N_2570);
nor U5728 (N_5728,N_2011,N_2965);
and U5729 (N_5729,N_3602,N_2988);
and U5730 (N_5730,N_3818,N_2753);
or U5731 (N_5731,N_3914,N_2869);
or U5732 (N_5732,N_2695,N_3683);
or U5733 (N_5733,N_2025,N_3438);
and U5734 (N_5734,N_2625,N_3467);
nand U5735 (N_5735,N_3654,N_2161);
nor U5736 (N_5736,N_3053,N_3589);
and U5737 (N_5737,N_2112,N_2981);
or U5738 (N_5738,N_3761,N_3697);
nor U5739 (N_5739,N_3776,N_3834);
nor U5740 (N_5740,N_2276,N_2529);
or U5741 (N_5741,N_3601,N_3123);
nor U5742 (N_5742,N_2785,N_3224);
and U5743 (N_5743,N_2658,N_3670);
and U5744 (N_5744,N_3857,N_2453);
nand U5745 (N_5745,N_3229,N_3521);
nor U5746 (N_5746,N_2090,N_3376);
xor U5747 (N_5747,N_3032,N_2347);
nand U5748 (N_5748,N_2397,N_3091);
nand U5749 (N_5749,N_3028,N_3551);
nor U5750 (N_5750,N_2507,N_3889);
xnor U5751 (N_5751,N_3885,N_3171);
or U5752 (N_5752,N_2931,N_2856);
nor U5753 (N_5753,N_3918,N_3525);
or U5754 (N_5754,N_3735,N_2307);
or U5755 (N_5755,N_2744,N_2230);
or U5756 (N_5756,N_2471,N_2580);
nand U5757 (N_5757,N_3604,N_3171);
and U5758 (N_5758,N_2991,N_3775);
or U5759 (N_5759,N_3647,N_2733);
or U5760 (N_5760,N_3890,N_2100);
and U5761 (N_5761,N_2304,N_2861);
or U5762 (N_5762,N_3204,N_3704);
nand U5763 (N_5763,N_3162,N_3835);
xor U5764 (N_5764,N_3373,N_2156);
or U5765 (N_5765,N_3241,N_2108);
or U5766 (N_5766,N_3999,N_2864);
and U5767 (N_5767,N_3842,N_2217);
nand U5768 (N_5768,N_3273,N_3189);
nor U5769 (N_5769,N_3611,N_2035);
nor U5770 (N_5770,N_3450,N_3263);
and U5771 (N_5771,N_3479,N_3156);
and U5772 (N_5772,N_2031,N_2817);
and U5773 (N_5773,N_2783,N_2505);
nand U5774 (N_5774,N_2610,N_3367);
and U5775 (N_5775,N_3887,N_3353);
xor U5776 (N_5776,N_2798,N_2548);
and U5777 (N_5777,N_2908,N_2488);
nor U5778 (N_5778,N_3445,N_3565);
and U5779 (N_5779,N_2030,N_3831);
xnor U5780 (N_5780,N_2316,N_2807);
nor U5781 (N_5781,N_3495,N_3317);
nor U5782 (N_5782,N_2240,N_2107);
nand U5783 (N_5783,N_3570,N_2075);
xor U5784 (N_5784,N_3083,N_3108);
and U5785 (N_5785,N_2127,N_3479);
nand U5786 (N_5786,N_2034,N_2265);
or U5787 (N_5787,N_2158,N_3066);
nand U5788 (N_5788,N_2105,N_3511);
nor U5789 (N_5789,N_2722,N_2627);
nor U5790 (N_5790,N_2757,N_2231);
nand U5791 (N_5791,N_3824,N_2673);
nand U5792 (N_5792,N_3723,N_2780);
nor U5793 (N_5793,N_2724,N_2420);
or U5794 (N_5794,N_3199,N_2936);
and U5795 (N_5795,N_3460,N_2279);
xnor U5796 (N_5796,N_3955,N_2243);
or U5797 (N_5797,N_3727,N_2070);
and U5798 (N_5798,N_2363,N_2947);
or U5799 (N_5799,N_3872,N_2394);
xnor U5800 (N_5800,N_3196,N_3653);
and U5801 (N_5801,N_2784,N_2400);
nand U5802 (N_5802,N_3103,N_3240);
or U5803 (N_5803,N_3912,N_2090);
and U5804 (N_5804,N_2368,N_3824);
nand U5805 (N_5805,N_3088,N_3588);
or U5806 (N_5806,N_2222,N_3691);
and U5807 (N_5807,N_3581,N_3700);
and U5808 (N_5808,N_2678,N_2613);
or U5809 (N_5809,N_3390,N_2528);
or U5810 (N_5810,N_3362,N_3096);
or U5811 (N_5811,N_3800,N_3114);
and U5812 (N_5812,N_3094,N_2539);
or U5813 (N_5813,N_3801,N_2376);
nor U5814 (N_5814,N_3553,N_2101);
and U5815 (N_5815,N_2714,N_2793);
or U5816 (N_5816,N_2909,N_2018);
nor U5817 (N_5817,N_2554,N_3958);
or U5818 (N_5818,N_2376,N_2919);
nor U5819 (N_5819,N_2740,N_3944);
nor U5820 (N_5820,N_3927,N_3140);
and U5821 (N_5821,N_2327,N_2412);
nand U5822 (N_5822,N_3289,N_2463);
and U5823 (N_5823,N_3275,N_3893);
and U5824 (N_5824,N_3799,N_2575);
or U5825 (N_5825,N_3890,N_2533);
nor U5826 (N_5826,N_3499,N_2906);
nand U5827 (N_5827,N_2753,N_2948);
nand U5828 (N_5828,N_2530,N_2264);
xor U5829 (N_5829,N_3829,N_2945);
nand U5830 (N_5830,N_3792,N_2210);
or U5831 (N_5831,N_2200,N_2629);
and U5832 (N_5832,N_2391,N_3823);
and U5833 (N_5833,N_2978,N_3622);
or U5834 (N_5834,N_3650,N_3976);
nand U5835 (N_5835,N_2117,N_2559);
nor U5836 (N_5836,N_3016,N_3659);
nor U5837 (N_5837,N_3867,N_3058);
and U5838 (N_5838,N_2998,N_2529);
or U5839 (N_5839,N_2198,N_2594);
or U5840 (N_5840,N_2680,N_2404);
xor U5841 (N_5841,N_3117,N_3094);
nand U5842 (N_5842,N_3619,N_3342);
and U5843 (N_5843,N_2409,N_2659);
nor U5844 (N_5844,N_3295,N_2309);
xnor U5845 (N_5845,N_3917,N_2075);
and U5846 (N_5846,N_3519,N_2287);
xor U5847 (N_5847,N_3150,N_3491);
and U5848 (N_5848,N_2169,N_3931);
and U5849 (N_5849,N_3325,N_3091);
or U5850 (N_5850,N_2803,N_3568);
or U5851 (N_5851,N_2381,N_2641);
nor U5852 (N_5852,N_3993,N_2984);
nand U5853 (N_5853,N_2139,N_2634);
and U5854 (N_5854,N_3171,N_2371);
and U5855 (N_5855,N_2582,N_2649);
nand U5856 (N_5856,N_2288,N_3841);
nand U5857 (N_5857,N_2972,N_3711);
and U5858 (N_5858,N_3434,N_3714);
xor U5859 (N_5859,N_2425,N_3249);
nand U5860 (N_5860,N_3048,N_3760);
nand U5861 (N_5861,N_3844,N_2259);
nor U5862 (N_5862,N_2204,N_2316);
or U5863 (N_5863,N_3699,N_3725);
and U5864 (N_5864,N_2162,N_3672);
nand U5865 (N_5865,N_2831,N_2030);
xnor U5866 (N_5866,N_2020,N_3347);
and U5867 (N_5867,N_2039,N_2188);
or U5868 (N_5868,N_3377,N_2711);
nor U5869 (N_5869,N_3327,N_3296);
nor U5870 (N_5870,N_3670,N_3702);
xor U5871 (N_5871,N_2364,N_3941);
nand U5872 (N_5872,N_2399,N_2179);
or U5873 (N_5873,N_2877,N_3648);
and U5874 (N_5874,N_3382,N_2953);
nand U5875 (N_5875,N_2215,N_3567);
xor U5876 (N_5876,N_3911,N_3922);
xor U5877 (N_5877,N_2886,N_3734);
or U5878 (N_5878,N_3288,N_2215);
nand U5879 (N_5879,N_3050,N_2240);
nor U5880 (N_5880,N_3090,N_2830);
and U5881 (N_5881,N_2981,N_3415);
and U5882 (N_5882,N_3265,N_2348);
or U5883 (N_5883,N_3643,N_2768);
nand U5884 (N_5884,N_3648,N_3630);
nor U5885 (N_5885,N_2795,N_2126);
and U5886 (N_5886,N_2336,N_2144);
or U5887 (N_5887,N_2630,N_2813);
nor U5888 (N_5888,N_2117,N_3971);
nor U5889 (N_5889,N_3457,N_3981);
and U5890 (N_5890,N_2561,N_2045);
or U5891 (N_5891,N_2279,N_2692);
nor U5892 (N_5892,N_2866,N_3790);
nor U5893 (N_5893,N_3003,N_2734);
nand U5894 (N_5894,N_2690,N_2199);
and U5895 (N_5895,N_3459,N_2578);
and U5896 (N_5896,N_2841,N_2486);
nor U5897 (N_5897,N_2650,N_3215);
nor U5898 (N_5898,N_2819,N_3959);
nand U5899 (N_5899,N_2387,N_3189);
nor U5900 (N_5900,N_3418,N_2594);
nor U5901 (N_5901,N_3885,N_3112);
nand U5902 (N_5902,N_2452,N_2199);
or U5903 (N_5903,N_2444,N_3794);
and U5904 (N_5904,N_2227,N_2651);
nand U5905 (N_5905,N_3588,N_3468);
and U5906 (N_5906,N_2774,N_2706);
nor U5907 (N_5907,N_3098,N_3135);
or U5908 (N_5908,N_3680,N_3632);
or U5909 (N_5909,N_2736,N_3907);
nand U5910 (N_5910,N_2455,N_2110);
or U5911 (N_5911,N_3144,N_2032);
nor U5912 (N_5912,N_2375,N_2890);
nor U5913 (N_5913,N_2003,N_3733);
nand U5914 (N_5914,N_2101,N_2685);
or U5915 (N_5915,N_3815,N_2298);
nand U5916 (N_5916,N_3798,N_3405);
and U5917 (N_5917,N_3655,N_3800);
nor U5918 (N_5918,N_2831,N_2518);
nor U5919 (N_5919,N_3424,N_3336);
and U5920 (N_5920,N_2302,N_2844);
or U5921 (N_5921,N_3870,N_2073);
and U5922 (N_5922,N_2203,N_2760);
nor U5923 (N_5923,N_3108,N_3465);
and U5924 (N_5924,N_3193,N_2579);
nand U5925 (N_5925,N_2492,N_3582);
nor U5926 (N_5926,N_2715,N_2737);
and U5927 (N_5927,N_3348,N_2448);
nor U5928 (N_5928,N_2349,N_2094);
nor U5929 (N_5929,N_3540,N_2977);
nor U5930 (N_5930,N_3458,N_3828);
and U5931 (N_5931,N_3221,N_2553);
or U5932 (N_5932,N_3575,N_3900);
and U5933 (N_5933,N_3035,N_2274);
nand U5934 (N_5934,N_3254,N_3625);
nor U5935 (N_5935,N_2887,N_3969);
xor U5936 (N_5936,N_2264,N_3584);
and U5937 (N_5937,N_2384,N_3088);
nor U5938 (N_5938,N_2310,N_3574);
nand U5939 (N_5939,N_3407,N_3210);
xor U5940 (N_5940,N_2351,N_3761);
nand U5941 (N_5941,N_3202,N_3908);
or U5942 (N_5942,N_3000,N_2900);
nand U5943 (N_5943,N_2070,N_2164);
or U5944 (N_5944,N_3142,N_3855);
and U5945 (N_5945,N_2983,N_2622);
nor U5946 (N_5946,N_3228,N_3962);
or U5947 (N_5947,N_3104,N_2905);
or U5948 (N_5948,N_2790,N_2767);
xnor U5949 (N_5949,N_2646,N_2068);
or U5950 (N_5950,N_2922,N_3492);
nand U5951 (N_5951,N_3103,N_3081);
or U5952 (N_5952,N_3735,N_3024);
nor U5953 (N_5953,N_3849,N_2937);
nand U5954 (N_5954,N_2967,N_2811);
nand U5955 (N_5955,N_3331,N_2335);
nand U5956 (N_5956,N_3039,N_3392);
and U5957 (N_5957,N_3077,N_3483);
nand U5958 (N_5958,N_3154,N_2492);
or U5959 (N_5959,N_2485,N_2049);
or U5960 (N_5960,N_2947,N_3491);
nand U5961 (N_5961,N_3219,N_3978);
nand U5962 (N_5962,N_2327,N_3880);
nand U5963 (N_5963,N_3835,N_3996);
nor U5964 (N_5964,N_3933,N_2947);
xor U5965 (N_5965,N_3208,N_3472);
nor U5966 (N_5966,N_2977,N_3315);
nand U5967 (N_5967,N_3466,N_3873);
nand U5968 (N_5968,N_3813,N_2726);
and U5969 (N_5969,N_3153,N_2784);
nand U5970 (N_5970,N_3611,N_3336);
xnor U5971 (N_5971,N_3366,N_3046);
nor U5972 (N_5972,N_2588,N_3485);
or U5973 (N_5973,N_3222,N_3985);
nand U5974 (N_5974,N_3176,N_2720);
nor U5975 (N_5975,N_2629,N_3785);
or U5976 (N_5976,N_2656,N_2520);
nor U5977 (N_5977,N_2942,N_2266);
and U5978 (N_5978,N_3714,N_3735);
or U5979 (N_5979,N_2313,N_2667);
and U5980 (N_5980,N_3073,N_2207);
xnor U5981 (N_5981,N_3629,N_2053);
and U5982 (N_5982,N_2622,N_2564);
nor U5983 (N_5983,N_3087,N_3778);
nor U5984 (N_5984,N_2351,N_3369);
or U5985 (N_5985,N_3772,N_2170);
and U5986 (N_5986,N_2570,N_3525);
and U5987 (N_5987,N_3671,N_2709);
xor U5988 (N_5988,N_2837,N_3963);
xor U5989 (N_5989,N_3516,N_2150);
xnor U5990 (N_5990,N_2711,N_3814);
nor U5991 (N_5991,N_3971,N_2631);
or U5992 (N_5992,N_3961,N_2854);
and U5993 (N_5993,N_2286,N_2351);
and U5994 (N_5994,N_3013,N_3511);
and U5995 (N_5995,N_3682,N_3577);
or U5996 (N_5996,N_2024,N_3495);
and U5997 (N_5997,N_2267,N_2470);
nand U5998 (N_5998,N_3927,N_3997);
and U5999 (N_5999,N_2991,N_2423);
nor U6000 (N_6000,N_4985,N_5928);
and U6001 (N_6001,N_4163,N_5493);
and U6002 (N_6002,N_4045,N_5284);
nand U6003 (N_6003,N_4334,N_4039);
xnor U6004 (N_6004,N_5985,N_5971);
or U6005 (N_6005,N_5597,N_4110);
nor U6006 (N_6006,N_4844,N_5948);
or U6007 (N_6007,N_4962,N_5350);
and U6008 (N_6008,N_4738,N_5303);
or U6009 (N_6009,N_5966,N_4579);
or U6010 (N_6010,N_5392,N_5915);
nand U6011 (N_6011,N_5252,N_5064);
or U6012 (N_6012,N_5004,N_4248);
nand U6013 (N_6013,N_5118,N_5895);
nand U6014 (N_6014,N_4420,N_4651);
nand U6015 (N_6015,N_5804,N_5911);
and U6016 (N_6016,N_5464,N_4907);
and U6017 (N_6017,N_5291,N_5242);
or U6018 (N_6018,N_4170,N_5914);
nor U6019 (N_6019,N_4697,N_5921);
nor U6020 (N_6020,N_5781,N_5529);
and U6021 (N_6021,N_4730,N_5035);
or U6022 (N_6022,N_4943,N_5926);
or U6023 (N_6023,N_4192,N_4635);
or U6024 (N_6024,N_4389,N_5053);
nor U6025 (N_6025,N_4617,N_5862);
nor U6026 (N_6026,N_5705,N_5470);
nor U6027 (N_6027,N_4854,N_5324);
nor U6028 (N_6028,N_4634,N_5606);
and U6029 (N_6029,N_4725,N_4339);
and U6030 (N_6030,N_5651,N_5800);
nand U6031 (N_6031,N_4202,N_5702);
xor U6032 (N_6032,N_5476,N_5851);
or U6033 (N_6033,N_5214,N_5984);
nand U6034 (N_6034,N_4642,N_4869);
nor U6035 (N_6035,N_5263,N_4242);
nor U6036 (N_6036,N_4614,N_5627);
xnor U6037 (N_6037,N_4035,N_4082);
or U6038 (N_6038,N_5473,N_5728);
and U6039 (N_6039,N_5533,N_4498);
nand U6040 (N_6040,N_5058,N_4454);
and U6041 (N_6041,N_5524,N_4033);
nand U6042 (N_6042,N_4994,N_4270);
or U6043 (N_6043,N_5235,N_5858);
or U6044 (N_6044,N_4575,N_5141);
nand U6045 (N_6045,N_4403,N_4118);
nand U6046 (N_6046,N_4536,N_5949);
nand U6047 (N_6047,N_4731,N_5625);
nand U6048 (N_6048,N_4164,N_5538);
and U6049 (N_6049,N_5694,N_5936);
nor U6050 (N_6050,N_5962,N_5247);
or U6051 (N_6051,N_5126,N_5482);
and U6052 (N_6052,N_5873,N_5759);
or U6053 (N_6053,N_5304,N_5772);
xnor U6054 (N_6054,N_4001,N_5789);
and U6055 (N_6055,N_5131,N_4719);
and U6056 (N_6056,N_4762,N_5158);
nor U6057 (N_6057,N_5296,N_4616);
or U6058 (N_6058,N_4947,N_5016);
or U6059 (N_6059,N_5744,N_4224);
or U6060 (N_6060,N_5951,N_5500);
nand U6061 (N_6061,N_4908,N_5047);
xor U6062 (N_6062,N_5506,N_4541);
nand U6063 (N_6063,N_4215,N_4084);
or U6064 (N_6064,N_5777,N_5275);
or U6065 (N_6065,N_4544,N_5821);
or U6066 (N_6066,N_4022,N_4402);
or U6067 (N_6067,N_4254,N_5485);
or U6068 (N_6068,N_4811,N_5318);
nor U6069 (N_6069,N_4729,N_4691);
xor U6070 (N_6070,N_4142,N_4206);
and U6071 (N_6071,N_5959,N_4929);
nand U6072 (N_6072,N_4961,N_4829);
xor U6073 (N_6073,N_5238,N_5188);
and U6074 (N_6074,N_5472,N_4937);
and U6075 (N_6075,N_5471,N_4763);
or U6076 (N_6076,N_4471,N_5913);
or U6077 (N_6077,N_5690,N_5580);
nand U6078 (N_6078,N_4573,N_4465);
nor U6079 (N_6079,N_4081,N_4894);
nand U6080 (N_6080,N_4439,N_4656);
nand U6081 (N_6081,N_5363,N_5273);
or U6082 (N_6082,N_4238,N_5293);
and U6083 (N_6083,N_4292,N_4417);
and U6084 (N_6084,N_5650,N_5590);
xor U6085 (N_6085,N_4695,N_5993);
nand U6086 (N_6086,N_4078,N_4480);
nand U6087 (N_6087,N_4088,N_4783);
nand U6088 (N_6088,N_4329,N_4793);
or U6089 (N_6089,N_4800,N_4542);
nor U6090 (N_6090,N_4151,N_5175);
nor U6091 (N_6091,N_4838,N_5305);
nand U6092 (N_6092,N_5081,N_5498);
nor U6093 (N_6093,N_5049,N_4779);
and U6094 (N_6094,N_4127,N_4421);
and U6095 (N_6095,N_4755,N_4901);
xnor U6096 (N_6096,N_5624,N_4363);
xnor U6097 (N_6097,N_5622,N_4904);
nor U6098 (N_6098,N_4490,N_5411);
or U6099 (N_6099,N_5738,N_5306);
and U6100 (N_6100,N_5784,N_4745);
xor U6101 (N_6101,N_4638,N_4772);
nand U6102 (N_6102,N_4167,N_5267);
nand U6103 (N_6103,N_4419,N_5121);
or U6104 (N_6104,N_5332,N_5331);
nand U6105 (N_6105,N_5319,N_5251);
and U6106 (N_6106,N_5481,N_5423);
and U6107 (N_6107,N_4602,N_5240);
nor U6108 (N_6108,N_5115,N_5073);
nor U6109 (N_6109,N_4426,N_4979);
and U6110 (N_6110,N_4877,N_5725);
and U6111 (N_6111,N_4503,N_5193);
or U6112 (N_6112,N_4592,N_4968);
or U6113 (N_6113,N_4776,N_4765);
or U6114 (N_6114,N_4394,N_5613);
or U6115 (N_6115,N_4186,N_5735);
nand U6116 (N_6116,N_4137,N_5184);
or U6117 (N_6117,N_4611,N_5845);
and U6118 (N_6118,N_5050,N_4505);
nand U6119 (N_6119,N_5107,N_5374);
or U6120 (N_6120,N_5753,N_5120);
or U6121 (N_6121,N_4191,N_5659);
nor U6122 (N_6122,N_4281,N_4585);
and U6123 (N_6123,N_4583,N_4133);
and U6124 (N_6124,N_4196,N_4624);
xor U6125 (N_6125,N_5195,N_4337);
or U6126 (N_6126,N_4474,N_4444);
or U6127 (N_6127,N_5022,N_4134);
nand U6128 (N_6128,N_5142,N_4563);
nand U6129 (N_6129,N_5736,N_5431);
nand U6130 (N_6130,N_5454,N_5674);
and U6131 (N_6131,N_5874,N_4061);
nor U6132 (N_6132,N_5312,N_5274);
xor U6133 (N_6133,N_5731,N_5207);
nor U6134 (N_6134,N_4808,N_4742);
nor U6135 (N_6135,N_4756,N_5180);
or U6136 (N_6136,N_4360,N_5382);
nor U6137 (N_6137,N_5075,N_5764);
nand U6138 (N_6138,N_5525,N_4274);
and U6139 (N_6139,N_5130,N_4068);
nand U6140 (N_6140,N_4213,N_5395);
nand U6141 (N_6141,N_5194,N_5811);
nor U6142 (N_6142,N_4272,N_5892);
nor U6143 (N_6143,N_5512,N_5390);
and U6144 (N_6144,N_5572,N_4491);
or U6145 (N_6145,N_5766,N_4932);
and U6146 (N_6146,N_5366,N_5203);
or U6147 (N_6147,N_5796,N_4569);
or U6148 (N_6148,N_4663,N_4365);
and U6149 (N_6149,N_4458,N_5277);
nor U6150 (N_6150,N_4048,N_4247);
and U6151 (N_6151,N_5593,N_4631);
and U6152 (N_6152,N_5148,N_5614);
nor U6153 (N_6153,N_4633,N_4315);
and U6154 (N_6154,N_5661,N_5909);
xor U6155 (N_6155,N_5540,N_4831);
or U6156 (N_6156,N_4218,N_4059);
nor U6157 (N_6157,N_4194,N_5967);
nand U6158 (N_6158,N_4547,N_5220);
xor U6159 (N_6159,N_4071,N_4423);
nor U6160 (N_6160,N_4355,N_4903);
nor U6161 (N_6161,N_4915,N_5978);
or U6162 (N_6162,N_5860,N_4034);
and U6163 (N_6163,N_4076,N_4146);
nor U6164 (N_6164,N_4311,N_5213);
and U6165 (N_6165,N_5765,N_4307);
or U6166 (N_6166,N_4286,N_5990);
and U6167 (N_6167,N_5850,N_4507);
nor U6168 (N_6168,N_4615,N_4815);
nand U6169 (N_6169,N_5693,N_4550);
nor U6170 (N_6170,N_4845,N_5846);
or U6171 (N_6171,N_4041,N_5187);
or U6172 (N_6172,N_4472,N_5854);
and U6173 (N_6173,N_4030,N_4993);
nor U6174 (N_6174,N_5174,N_4607);
nand U6175 (N_6175,N_4053,N_5885);
nand U6176 (N_6176,N_4873,N_4208);
and U6177 (N_6177,N_5907,N_4367);
nor U6178 (N_6178,N_4231,N_5582);
nor U6179 (N_6179,N_5356,N_4325);
and U6180 (N_6180,N_5636,N_5477);
nand U6181 (N_6181,N_4820,N_5479);
or U6182 (N_6182,N_5550,N_5623);
or U6183 (N_6183,N_4347,N_5603);
and U6184 (N_6184,N_4574,N_5831);
nand U6185 (N_6185,N_4070,N_5268);
or U6186 (N_6186,N_5151,N_5547);
nor U6187 (N_6187,N_4914,N_5147);
or U6188 (N_6188,N_5078,N_5942);
or U6189 (N_6189,N_5445,N_5893);
or U6190 (N_6190,N_5070,N_5552);
nand U6191 (N_6191,N_4063,N_5867);
or U6192 (N_6192,N_5896,N_4711);
and U6193 (N_6193,N_4299,N_5798);
or U6194 (N_6194,N_4488,N_5323);
nor U6195 (N_6195,N_4842,N_5929);
nor U6196 (N_6196,N_5337,N_5373);
and U6197 (N_6197,N_4004,N_4250);
or U6198 (N_6198,N_5934,N_5616);
nand U6199 (N_6199,N_5292,N_5484);
nor U6200 (N_6200,N_4243,N_5008);
or U6201 (N_6201,N_4767,N_5325);
nor U6202 (N_6202,N_5576,N_5317);
nor U6203 (N_6203,N_5103,N_5646);
nor U6204 (N_6204,N_4552,N_5299);
nor U6205 (N_6205,N_4184,N_5450);
or U6206 (N_6206,N_4766,N_4764);
nor U6207 (N_6207,N_4952,N_5090);
nor U6208 (N_6208,N_5780,N_5898);
or U6209 (N_6209,N_4593,N_5475);
or U6210 (N_6210,N_4665,N_5302);
xor U6211 (N_6211,N_5975,N_4159);
nand U6212 (N_6212,N_4219,N_4951);
nand U6213 (N_6213,N_5917,N_5381);
nor U6214 (N_6214,N_4132,N_4954);
or U6215 (N_6215,N_5657,N_5639);
and U6216 (N_6216,N_4020,N_5724);
nor U6217 (N_6217,N_5973,N_4155);
or U6218 (N_6218,N_4580,N_5767);
nand U6219 (N_6219,N_5093,N_5117);
or U6220 (N_6220,N_5160,N_5581);
nand U6221 (N_6221,N_5943,N_4555);
and U6222 (N_6222,N_4324,N_5096);
or U6223 (N_6223,N_4775,N_5236);
nand U6224 (N_6224,N_5432,N_5037);
and U6225 (N_6225,N_5960,N_5726);
nand U6226 (N_6226,N_5976,N_5610);
nor U6227 (N_6227,N_5859,N_5956);
nor U6228 (N_6228,N_4618,N_4761);
and U6229 (N_6229,N_5480,N_4049);
and U6230 (N_6230,N_4760,N_5168);
or U6231 (N_6231,N_4318,N_4753);
or U6232 (N_6232,N_5944,N_5511);
nand U6233 (N_6233,N_4493,N_5461);
xor U6234 (N_6234,N_4099,N_4162);
xor U6235 (N_6235,N_5641,N_5700);
nor U6236 (N_6236,N_4641,N_4898);
nor U6237 (N_6237,N_5589,N_5531);
and U6238 (N_6238,N_5379,N_4628);
nor U6239 (N_6239,N_4917,N_4515);
or U6240 (N_6240,N_4647,N_5742);
nand U6241 (N_6241,N_4933,N_4989);
nand U6242 (N_6242,N_4759,N_5079);
nor U6243 (N_6243,N_4416,N_4888);
or U6244 (N_6244,N_4791,N_4535);
and U6245 (N_6245,N_4996,N_4558);
nor U6246 (N_6246,N_5416,N_5912);
or U6247 (N_6247,N_5905,N_4177);
and U6248 (N_6248,N_5186,N_5199);
nand U6249 (N_6249,N_5666,N_4644);
nor U6250 (N_6250,N_4557,N_4283);
nand U6251 (N_6251,N_4025,N_5278);
or U6252 (N_6252,N_4594,N_4216);
or U6253 (N_6253,N_5536,N_5996);
or U6254 (N_6254,N_4298,N_4335);
nor U6255 (N_6255,N_4668,N_5137);
and U6256 (N_6256,N_5732,N_4096);
nor U6257 (N_6257,N_4862,N_5670);
and U6258 (N_6258,N_4524,N_4824);
or U6259 (N_6259,N_5521,N_5105);
nand U6260 (N_6260,N_4027,N_5169);
and U6261 (N_6261,N_5161,N_5294);
or U6262 (N_6262,N_4523,N_5565);
and U6263 (N_6263,N_4770,N_5361);
and U6264 (N_6264,N_5145,N_5313);
xor U6265 (N_6265,N_4846,N_5649);
and U6266 (N_6266,N_4886,N_4152);
nand U6267 (N_6267,N_5435,N_5428);
and U6268 (N_6268,N_4010,N_4780);
or U6269 (N_6269,N_5882,N_4789);
and U6270 (N_6270,N_5065,N_4391);
nand U6271 (N_6271,N_5842,N_4002);
nor U6272 (N_6272,N_5112,N_4657);
and U6273 (N_6273,N_4896,N_4551);
or U6274 (N_6274,N_4525,N_5908);
nor U6275 (N_6275,N_4237,N_4689);
or U6276 (N_6276,N_4326,N_5528);
and U6277 (N_6277,N_5937,N_5034);
or U6278 (N_6278,N_4136,N_4011);
and U6279 (N_6279,N_4168,N_5030);
nand U6280 (N_6280,N_5847,N_4214);
nand U6281 (N_6281,N_5730,N_4865);
and U6282 (N_6282,N_4424,N_4475);
nor U6283 (N_6283,N_5210,N_4659);
nand U6284 (N_6284,N_5228,N_5046);
or U6285 (N_6285,N_5957,N_5684);
and U6286 (N_6286,N_4290,N_4074);
or U6287 (N_6287,N_5003,N_5823);
nand U6288 (N_6288,N_5110,N_5607);
nor U6289 (N_6289,N_4995,N_4336);
nand U6290 (N_6290,N_5488,N_4539);
nand U6291 (N_6291,N_5612,N_4026);
nand U6292 (N_6292,N_5717,N_4925);
or U6293 (N_6293,N_4926,N_5843);
nand U6294 (N_6294,N_5085,N_4187);
and U6295 (N_6295,N_5011,N_5809);
or U6296 (N_6296,N_5950,N_5033);
nand U6297 (N_6297,N_4222,N_5712);
nor U6298 (N_6298,N_5441,N_4024);
nor U6299 (N_6299,N_5341,N_4372);
or U6300 (N_6300,N_5522,N_5486);
nor U6301 (N_6301,N_5370,N_4875);
xor U6302 (N_6302,N_4807,N_4418);
and U6303 (N_6303,N_5863,N_4453);
or U6304 (N_6304,N_4857,N_4441);
or U6305 (N_6305,N_4157,N_4771);
nand U6306 (N_6306,N_4436,N_5652);
nor U6307 (N_6307,N_5290,N_5328);
nand U6308 (N_6308,N_4964,N_5026);
xnor U6309 (N_6309,N_5491,N_4413);
or U6310 (N_6310,N_4802,N_4090);
xor U6311 (N_6311,N_5760,N_5157);
nor U6312 (N_6312,N_5791,N_4448);
nand U6313 (N_6313,N_5264,N_5579);
nor U6314 (N_6314,N_5038,N_5042);
xor U6315 (N_6315,N_4982,N_4828);
nand U6316 (N_6316,N_4987,N_5094);
nor U6317 (N_6317,N_4473,N_4833);
nand U6318 (N_6318,N_5806,N_4975);
nor U6319 (N_6319,N_4319,N_4064);
nor U6320 (N_6320,N_5710,N_5436);
nand U6321 (N_6321,N_5509,N_4113);
nand U6322 (N_6322,N_4357,N_5647);
or U6323 (N_6323,N_5680,N_4293);
and U6324 (N_6324,N_4210,N_5421);
and U6325 (N_6325,N_4609,N_5626);
nor U6326 (N_6326,N_4652,N_5167);
or U6327 (N_6327,N_5116,N_5301);
or U6328 (N_6328,N_4245,N_5709);
nor U6329 (N_6329,N_4220,N_5387);
or U6330 (N_6330,N_5360,N_4232);
nor U6331 (N_6331,N_4287,N_5629);
nand U6332 (N_6332,N_5752,N_4138);
or U6333 (N_6333,N_5663,N_5244);
nand U6334 (N_6334,N_4970,N_5757);
nand U6335 (N_6335,N_5418,N_4393);
and U6336 (N_6336,N_5216,N_5149);
nor U6337 (N_6337,N_4513,N_4911);
or U6338 (N_6338,N_4456,N_4052);
xor U6339 (N_6339,N_4577,N_4023);
nor U6340 (N_6340,N_4442,N_4385);
or U6341 (N_6341,N_5520,N_4427);
or U6342 (N_6342,N_4769,N_4412);
nand U6343 (N_6343,N_4782,N_4785);
nor U6344 (N_6344,N_4899,N_5134);
and U6345 (N_6345,N_4902,N_4673);
xnor U6346 (N_6346,N_5279,N_4273);
or U6347 (N_6347,N_4042,N_4768);
and U6348 (N_6348,N_5343,N_5808);
or U6349 (N_6349,N_4704,N_5737);
nor U6350 (N_6350,N_4504,N_5190);
xnor U6351 (N_6351,N_4291,N_4835);
and U6352 (N_6352,N_5460,N_4741);
nor U6353 (N_6353,N_4150,N_5836);
and U6354 (N_6354,N_4484,N_5783);
and U6355 (N_6355,N_4489,N_4221);
nand U6356 (N_6356,N_5001,N_4511);
xor U6357 (N_6357,N_5101,N_4249);
nand U6358 (N_6358,N_4226,N_5977);
or U6359 (N_6359,N_5225,N_4255);
or U6360 (N_6360,N_4562,N_4714);
nor U6361 (N_6361,N_5039,N_5879);
and U6362 (N_6362,N_5592,N_4455);
or U6363 (N_6363,N_4227,N_4468);
nor U6364 (N_6364,N_4639,N_4296);
nand U6365 (N_6365,N_5490,N_4397);
nor U6366 (N_6366,N_4406,N_5176);
nand U6367 (N_6367,N_5987,N_4786);
nand U6368 (N_6368,N_5083,N_4487);
nor U6369 (N_6369,N_4540,N_5945);
nand U6370 (N_6370,N_4564,N_5349);
and U6371 (N_6371,N_4459,N_5734);
or U6372 (N_6372,N_4545,N_5514);
or U6373 (N_6373,N_4977,N_5906);
nor U6374 (N_6374,N_5719,N_5316);
or U6375 (N_6375,N_4120,N_5163);
and U6376 (N_6376,N_4410,N_5132);
nor U6377 (N_6377,N_4300,N_4392);
nand U6378 (N_6378,N_5162,N_4799);
xnor U6379 (N_6379,N_4893,N_5812);
nor U6380 (N_6380,N_4649,N_4452);
and U6381 (N_6381,N_5886,N_5594);
nand U6382 (N_6382,N_5793,N_5961);
nand U6383 (N_6383,N_5870,N_5848);
and U6384 (N_6384,N_4105,N_4839);
nor U6385 (N_6385,N_4856,N_4500);
and U6386 (N_6386,N_4913,N_5617);
nor U6387 (N_6387,N_4941,N_4095);
nand U6388 (N_6388,N_5000,N_4876);
xor U6389 (N_6389,N_4726,N_4262);
xnor U6390 (N_6390,N_5333,N_5166);
nand U6391 (N_6391,N_5668,N_4743);
or U6392 (N_6392,N_5814,N_4997);
nand U6393 (N_6393,N_5246,N_5458);
or U6394 (N_6394,N_5825,N_4625);
nor U6395 (N_6395,N_5329,N_5276);
nor U6396 (N_6396,N_4323,N_4384);
nand U6397 (N_6397,N_5234,N_5880);
or U6398 (N_6398,N_4382,N_4864);
nor U6399 (N_6399,N_5855,N_4868);
nand U6400 (N_6400,N_4662,N_5608);
xor U6401 (N_6401,N_5868,N_5822);
or U6402 (N_6402,N_5964,N_5191);
and U6403 (N_6403,N_4566,N_4591);
nand U6404 (N_6404,N_4446,N_5740);
nand U6405 (N_6405,N_5544,N_4294);
nor U6406 (N_6406,N_4748,N_4124);
or U6407 (N_6407,N_5601,N_5013);
and U6408 (N_6408,N_4897,N_5655);
nor U6409 (N_6409,N_5995,N_4295);
nor U6410 (N_6410,N_4945,N_5172);
xor U6411 (N_6411,N_5233,N_4007);
xnor U6412 (N_6412,N_5527,N_4694);
xnor U6413 (N_6413,N_4936,N_5718);
xor U6414 (N_6414,N_4777,N_4740);
and U6415 (N_6415,N_5578,N_4821);
or U6416 (N_6416,N_5872,N_4377);
nand U6417 (N_6417,N_5061,N_5992);
nand U6418 (N_6418,N_5352,N_5136);
nor U6419 (N_6419,N_5982,N_5307);
and U6420 (N_6420,N_5656,N_4934);
and U6421 (N_6421,N_4681,N_4309);
or U6422 (N_6422,N_5334,N_4205);
and U6423 (N_6423,N_4251,N_5840);
and U6424 (N_6424,N_4843,N_4314);
nand U6425 (N_6425,N_5871,N_5628);
nand U6426 (N_6426,N_4924,N_4627);
and U6427 (N_6427,N_4608,N_4112);
and U6428 (N_6428,N_4737,N_5150);
and U6429 (N_6429,N_5749,N_5027);
and U6430 (N_6430,N_5255,N_5795);
or U6431 (N_6431,N_5746,N_5059);
or U6432 (N_6432,N_4344,N_5181);
and U6433 (N_6433,N_4946,N_5989);
and U6434 (N_6434,N_4128,N_4827);
and U6435 (N_6435,N_4310,N_4664);
and U6436 (N_6436,N_5114,N_4565);
and U6437 (N_6437,N_5404,N_4266);
nor U6438 (N_6438,N_5269,N_4094);
nand U6439 (N_6439,N_4450,N_5043);
xnor U6440 (N_6440,N_5023,N_5383);
nor U6441 (N_6441,N_4599,N_4328);
and U6442 (N_6442,N_5819,N_5051);
or U6443 (N_6443,N_4596,N_4141);
nor U6444 (N_6444,N_5029,N_4225);
or U6445 (N_6445,N_5555,N_5173);
nand U6446 (N_6446,N_4193,N_5143);
nand U6447 (N_6447,N_4600,N_5988);
and U6448 (N_6448,N_4905,N_4486);
or U6449 (N_6449,N_5678,N_4431);
nor U6450 (N_6450,N_4878,N_5584);
nand U6451 (N_6451,N_5935,N_5658);
and U6452 (N_6452,N_5447,N_4204);
and U6453 (N_6453,N_5088,N_5683);
and U6454 (N_6454,N_4021,N_5835);
xnor U6455 (N_6455,N_4258,N_4923);
nor U6456 (N_6456,N_5598,N_4342);
or U6457 (N_6457,N_4891,N_4409);
nor U6458 (N_6458,N_4407,N_5197);
and U6459 (N_6459,N_5505,N_4512);
and U6460 (N_6460,N_5219,N_5346);
nand U6461 (N_6461,N_4605,N_4404);
nor U6462 (N_6462,N_5017,N_4739);
nor U6463 (N_6463,N_4510,N_5534);
xnor U6464 (N_6464,N_4077,N_4803);
and U6465 (N_6465,N_4171,N_4718);
nor U6466 (N_6466,N_5315,N_5692);
nand U6467 (N_6467,N_4733,N_4702);
nor U6468 (N_6468,N_4338,N_4978);
and U6469 (N_6469,N_5380,N_4354);
nor U6470 (N_6470,N_5208,N_4746);
and U6471 (N_6471,N_4173,N_4198);
nand U6472 (N_6472,N_4847,N_4620);
nor U6473 (N_6473,N_4122,N_5986);
or U6474 (N_6474,N_5839,N_5832);
nor U6475 (N_6475,N_4429,N_4056);
nor U6476 (N_6476,N_5941,N_5621);
xor U6477 (N_6477,N_5596,N_5701);
nand U6478 (N_6478,N_4796,N_5408);
or U6479 (N_6479,N_4685,N_5257);
or U6480 (N_6480,N_5138,N_4003);
xnor U6481 (N_6481,N_4795,N_5362);
nor U6482 (N_6482,N_5239,N_4313);
and U6483 (N_6483,N_4570,N_5774);
nor U6484 (N_6484,N_4568,N_4390);
xnor U6485 (N_6485,N_4261,N_5551);
nand U6486 (N_6486,N_5440,N_5947);
and U6487 (N_6487,N_4422,N_4462);
nor U6488 (N_6488,N_5559,N_5715);
nand U6489 (N_6489,N_5797,N_4832);
or U6490 (N_6490,N_4981,N_4457);
and U6491 (N_6491,N_4235,N_4008);
or U6492 (N_6492,N_5063,N_4282);
nand U6493 (N_6493,N_5266,N_4587);
or U6494 (N_6494,N_5054,N_5340);
and U6495 (N_6495,N_4597,N_4584);
and U6496 (N_6496,N_5066,N_4721);
nor U6497 (N_6497,N_5171,N_5919);
or U6498 (N_6498,N_4069,N_5571);
or U6499 (N_6499,N_4364,N_5573);
nor U6500 (N_6500,N_4317,N_5097);
or U6501 (N_6501,N_5748,N_5713);
nor U6502 (N_6502,N_4006,N_4851);
xor U6503 (N_6503,N_4713,N_4398);
or U6504 (N_6504,N_4648,N_4306);
nor U6505 (N_6505,N_4810,N_4825);
nor U6506 (N_6506,N_5545,N_5439);
and U6507 (N_6507,N_4973,N_4548);
nor U6508 (N_6508,N_4188,N_5456);
and U6509 (N_6509,N_5703,N_5068);
or U6510 (N_6510,N_5086,N_5569);
and U6511 (N_6511,N_5465,N_4308);
nor U6512 (N_6512,N_4172,N_5014);
nor U6513 (N_6513,N_4710,N_5089);
nand U6514 (N_6514,N_4276,N_5348);
and U6515 (N_6515,N_5419,N_5501);
nand U6516 (N_6516,N_5564,N_5923);
and U6517 (N_6517,N_5104,N_5438);
nand U6518 (N_6518,N_4890,N_4244);
and U6519 (N_6519,N_5015,N_5686);
nor U6520 (N_6520,N_5402,N_4037);
and U6521 (N_6521,N_5635,N_4816);
nand U6522 (N_6522,N_4481,N_5558);
nand U6523 (N_6523,N_4083,N_5644);
nand U6524 (N_6524,N_5351,N_5720);
nand U6525 (N_6525,N_4682,N_5618);
xnor U6526 (N_6526,N_5671,N_5707);
nor U6527 (N_6527,N_5775,N_4352);
nor U6528 (N_6528,N_5600,N_5676);
nand U6529 (N_6529,N_5468,N_5100);
xor U6530 (N_6530,N_5497,N_4841);
nand U6531 (N_6531,N_5587,N_5745);
and U6532 (N_6532,N_5062,N_5747);
nor U6533 (N_6533,N_5270,N_4316);
and U6534 (N_6534,N_5516,N_4667);
nor U6535 (N_6535,N_5224,N_5813);
or U6536 (N_6536,N_4874,N_5357);
or U6537 (N_6537,N_4380,N_4960);
and U6538 (N_6538,N_5124,N_5261);
nand U6539 (N_6539,N_4537,N_4967);
or U6540 (N_6540,N_4999,N_5675);
xnor U6541 (N_6541,N_5810,N_5541);
nor U6542 (N_6542,N_5230,N_5588);
or U6543 (N_6543,N_5452,N_5129);
and U6544 (N_6544,N_4858,N_5769);
or U6545 (N_6545,N_5309,N_5492);
nor U6546 (N_6546,N_5209,N_4533);
nor U6547 (N_6547,N_5820,N_4976);
nand U6548 (N_6548,N_4097,N_4744);
and U6549 (N_6549,N_4400,N_5469);
nor U6550 (N_6550,N_4303,N_4153);
nor U6551 (N_6551,N_4984,N_4396);
and U6552 (N_6552,N_5119,N_5099);
and U6553 (N_6553,N_5076,N_4341);
or U6554 (N_6554,N_5899,N_4289);
or U6555 (N_6555,N_4722,N_5495);
or U6556 (N_6556,N_5425,N_5474);
nor U6557 (N_6557,N_5697,N_5133);
and U6558 (N_6558,N_4054,N_4330);
nor U6559 (N_6559,N_4957,N_4051);
nand U6560 (N_6560,N_5159,N_5901);
nor U6561 (N_6561,N_4499,N_5830);
and U6562 (N_6562,N_5140,N_5095);
and U6563 (N_6563,N_5785,N_4371);
nand U6564 (N_6564,N_4358,N_4492);
or U6565 (N_6565,N_4701,N_4974);
and U6566 (N_6566,N_4102,N_4655);
nand U6567 (N_6567,N_5642,N_4872);
or U6568 (N_6568,N_5721,N_5077);
and U6569 (N_6569,N_4556,N_4388);
nand U6570 (N_6570,N_4228,N_4189);
and U6571 (N_6571,N_4826,N_4958);
or U6572 (N_6572,N_5605,N_4467);
xor U6573 (N_6573,N_4445,N_4603);
nor U6574 (N_6574,N_5444,N_4200);
and U6575 (N_6575,N_4906,N_4180);
and U6576 (N_6576,N_5773,N_5633);
xor U6577 (N_6577,N_5933,N_5448);
and U6578 (N_6578,N_5002,N_5792);
xnor U6579 (N_6579,N_5499,N_5838);
or U6580 (N_6580,N_5770,N_4927);
nand U6581 (N_6581,N_5695,N_4199);
nand U6582 (N_6582,N_4016,N_5198);
and U6583 (N_6583,N_5741,N_4495);
nor U6584 (N_6584,N_4469,N_4209);
or U6585 (N_6585,N_4531,N_4103);
or U6586 (N_6586,N_4207,N_4671);
and U6587 (N_6587,N_5857,N_4246);
and U6588 (N_6588,N_4813,N_4047);
nand U6589 (N_6589,N_4443,N_5189);
nand U6590 (N_6590,N_4060,N_5689);
and U6591 (N_6591,N_5518,N_4114);
or U6592 (N_6592,N_5865,N_5048);
or U6593 (N_6593,N_4279,N_5782);
and U6594 (N_6594,N_4332,N_4794);
nor U6595 (N_6595,N_5417,N_4145);
nor U6596 (N_6596,N_5508,N_4654);
nor U6597 (N_6597,N_4119,N_5164);
xnor U6598 (N_6598,N_4723,N_4229);
or U6599 (N_6599,N_4479,N_4179);
xor U6600 (N_6600,N_4892,N_5217);
xnor U6601 (N_6601,N_4549,N_4860);
nor U6602 (N_6602,N_4571,N_5611);
or U6603 (N_6603,N_4322,N_5052);
nand U6604 (N_6604,N_4709,N_5691);
nand U6605 (N_6605,N_4386,N_5256);
nor U6606 (N_6606,N_4375,N_5801);
and U6607 (N_6607,N_4019,N_5972);
and U6608 (N_6608,N_5231,N_5123);
nand U6609 (N_6609,N_5271,N_5953);
xnor U6610 (N_6610,N_4882,N_4301);
nand U6611 (N_6611,N_4143,N_4201);
nor U6612 (N_6612,N_5212,N_4449);
nor U6613 (N_6613,N_5563,N_5939);
nand U6614 (N_6614,N_4823,N_4058);
and U6615 (N_6615,N_4275,N_5568);
nor U6616 (N_6616,N_5602,N_4433);
nor U6617 (N_6617,N_5245,N_4414);
nor U6618 (N_6618,N_4169,N_4212);
nand U6619 (N_6619,N_4971,N_4900);
nor U6620 (N_6620,N_4528,N_5827);
nor U6621 (N_6621,N_5991,N_4527);
and U6622 (N_6622,N_5409,N_5515);
nor U6623 (N_6623,N_5687,N_4065);
or U6624 (N_6624,N_4728,N_5272);
nor U6625 (N_6625,N_5071,N_5640);
nand U6626 (N_6626,N_5204,N_4239);
xor U6627 (N_6627,N_5637,N_5314);
nor U6628 (N_6628,N_5751,N_5574);
or U6629 (N_6629,N_5669,N_5604);
nor U6630 (N_6630,N_5422,N_4836);
nand U6631 (N_6631,N_4526,N_4861);
nand U6632 (N_6632,N_4277,N_5954);
or U6633 (N_6633,N_5881,N_4362);
and U6634 (N_6634,N_4175,N_4203);
and U6635 (N_6635,N_5615,N_4072);
xor U6636 (N_6636,N_5200,N_4038);
nor U6637 (N_6637,N_5875,N_4948);
nor U6638 (N_6638,N_4885,N_5542);
nor U6639 (N_6639,N_4855,N_4938);
and U6640 (N_6640,N_4751,N_5487);
xor U6641 (N_6641,N_5342,N_5384);
and U6642 (N_6642,N_5952,N_5453);
and U6643 (N_6643,N_5994,N_5903);
nor U6644 (N_6644,N_5248,N_4674);
nor U6645 (N_6645,N_5135,N_4331);
nand U6646 (N_6646,N_4757,N_4581);
nand U6647 (N_6647,N_5786,N_5430);
xnor U6648 (N_6648,N_5834,N_5177);
xnor U6649 (N_6649,N_5560,N_5673);
xor U6650 (N_6650,N_5758,N_5688);
or U6651 (N_6651,N_5768,N_4720);
nand U6652 (N_6652,N_4040,N_4774);
xnor U6653 (N_6653,N_4359,N_5358);
nor U6654 (N_6654,N_4267,N_4518);
and U6655 (N_6655,N_4101,N_5546);
nor U6656 (N_6656,N_4302,N_5462);
nor U6657 (N_6657,N_4956,N_5344);
nor U6658 (N_6658,N_5359,N_5260);
nor U6659 (N_6659,N_5403,N_5523);
nor U6660 (N_6660,N_5005,N_4983);
nand U6661 (N_6661,N_5371,N_4148);
nor U6662 (N_6662,N_5887,N_4285);
and U6663 (N_6663,N_4182,N_5283);
and U6664 (N_6664,N_5146,N_4534);
xor U6665 (N_6665,N_5056,N_5496);
nand U6666 (N_6666,N_5221,N_5653);
nor U6667 (N_6667,N_5376,N_4622);
nor U6668 (N_6668,N_5931,N_4470);
nand U6669 (N_6669,N_5399,N_5837);
or U6670 (N_6670,N_4520,N_5455);
nor U6671 (N_6671,N_5537,N_4884);
or U6672 (N_6672,N_4284,N_5012);
or U6673 (N_6673,N_5466,N_4107);
nand U6674 (N_6674,N_5968,N_4401);
nand U6675 (N_6675,N_5427,N_5020);
or U6676 (N_6676,N_5861,N_4848);
nand U6677 (N_6677,N_4000,N_5413);
and U6678 (N_6678,N_4032,N_5554);
and U6679 (N_6679,N_4532,N_5282);
nor U6680 (N_6680,N_4256,N_4619);
and U6681 (N_6681,N_4126,N_4154);
nand U6682 (N_6682,N_5297,N_5028);
nor U6683 (N_6683,N_4015,N_5510);
and U6684 (N_6684,N_5170,N_5925);
or U6685 (N_6685,N_4098,N_5335);
or U6686 (N_6686,N_5756,N_4115);
nor U6687 (N_6687,N_5761,N_4376);
and U6688 (N_6688,N_4106,N_4787);
and U6689 (N_6689,N_5326,N_4014);
or U6690 (N_6690,N_4699,N_4304);
xnor U6691 (N_6691,N_5983,N_5415);
nand U6692 (N_6692,N_4399,N_4703);
nand U6693 (N_6693,N_5963,N_4483);
or U6694 (N_6694,N_5619,N_5727);
and U6695 (N_6695,N_4140,N_5478);
or U6696 (N_6696,N_4233,N_4125);
and U6697 (N_6697,N_5310,N_5532);
nor U6698 (N_6698,N_4280,N_4606);
nand U6699 (N_6699,N_4612,N_5424);
nand U6700 (N_6700,N_4881,N_4880);
and U6701 (N_6701,N_4696,N_4837);
xor U6702 (N_6702,N_5876,N_5098);
or U6703 (N_6703,N_5347,N_5922);
and U6704 (N_6704,N_4408,N_4129);
nand U6705 (N_6705,N_5467,N_5620);
and U6706 (N_6706,N_4506,N_5833);
and U6707 (N_6707,N_5890,N_4553);
and U6708 (N_6708,N_5549,N_5446);
nor U6709 (N_6709,N_4940,N_5165);
and U6710 (N_6710,N_4676,N_5762);
nand U6711 (N_6711,N_4959,N_5869);
nor U6712 (N_6712,N_4817,N_5122);
nand U6713 (N_6713,N_4830,N_5320);
nand U6714 (N_6714,N_4437,N_4986);
and U6715 (N_6715,N_4411,N_5841);
or U6716 (N_6716,N_4972,N_4012);
or U6717 (N_6717,N_4093,N_5280);
nor U6718 (N_6718,N_4252,N_4075);
or U6719 (N_6719,N_5648,N_4646);
and U6720 (N_6720,N_5575,N_4149);
or U6721 (N_6721,N_5667,N_5414);
and U6722 (N_6722,N_4345,N_4669);
nand U6723 (N_6723,N_4942,N_5045);
and U6724 (N_6724,N_4724,N_4521);
nand U6725 (N_6725,N_4707,N_4305);
nor U6726 (N_6726,N_5364,N_4626);
nand U6727 (N_6727,N_5196,N_4840);
or U6728 (N_6728,N_4130,N_4018);
nor U6729 (N_6729,N_5397,N_5802);
and U6730 (N_6730,N_4108,N_4327);
and U6731 (N_6731,N_5237,N_4749);
nand U6732 (N_6732,N_4109,N_4920);
or U6733 (N_6733,N_5733,N_5463);
nor U6734 (N_6734,N_4379,N_4005);
or U6735 (N_6735,N_5803,N_5677);
and U6736 (N_6736,N_5586,N_4683);
or U6737 (N_6737,N_5599,N_4554);
and U6738 (N_6738,N_4086,N_5375);
or U6739 (N_6739,N_5938,N_5155);
nor U6740 (N_6740,N_5074,N_5009);
nand U6741 (N_6741,N_4440,N_5969);
nor U6742 (N_6742,N_4036,N_4658);
or U6743 (N_6743,N_5932,N_4073);
xnor U6744 (N_6744,N_4477,N_4031);
or U6745 (N_6745,N_4572,N_5970);
and U6746 (N_6746,N_4117,N_4190);
nand U6747 (N_6747,N_5091,N_5327);
and U6748 (N_6748,N_5451,N_4988);
or U6749 (N_6749,N_5739,N_4717);
or U6750 (N_6750,N_4366,N_4271);
nand U6751 (N_6751,N_5698,N_4265);
xnor U6752 (N_6752,N_5087,N_4425);
and U6753 (N_6753,N_4677,N_4043);
or U6754 (N_6754,N_5828,N_4104);
xnor U6755 (N_6755,N_4747,N_5407);
nand U6756 (N_6756,N_4297,N_5562);
nor U6757 (N_6757,N_4089,N_4312);
or U6758 (N_6758,N_4217,N_4451);
and U6759 (N_6759,N_4502,N_4264);
nor U6760 (N_6760,N_5338,N_5853);
or U6761 (N_6761,N_5330,N_4916);
nand U6762 (N_6762,N_4333,N_5681);
nand U6763 (N_6763,N_4223,N_4589);
nand U6764 (N_6764,N_4814,N_5378);
xor U6765 (N_6765,N_5113,N_4812);
or U6766 (N_6766,N_4369,N_4949);
and U6767 (N_6767,N_4139,N_5723);
or U6768 (N_6768,N_4463,N_5750);
xnor U6769 (N_6769,N_4661,N_5910);
and U6770 (N_6770,N_4079,N_4992);
nand U6771 (N_6771,N_4680,N_4930);
nand U6772 (N_6772,N_5946,N_4700);
nand U6773 (N_6773,N_5032,N_5595);
and U6774 (N_6774,N_4066,N_5300);
nor U6775 (N_6775,N_4822,N_5153);
or U6776 (N_6776,N_4863,N_5125);
or U6777 (N_6777,N_4185,N_4123);
or U6778 (N_6778,N_5577,N_5021);
nor U6779 (N_6779,N_5958,N_5722);
nand U6780 (N_6780,N_4181,N_4464);
nor U6781 (N_6781,N_4482,N_5398);
and U6782 (N_6782,N_5716,N_4567);
nand U6783 (N_6783,N_5553,N_5685);
nor U6784 (N_6784,N_5561,N_5824);
nor U6785 (N_6785,N_5281,N_5102);
and U6786 (N_6786,N_4698,N_5706);
nor U6787 (N_6787,N_5965,N_5998);
nor U6788 (N_6788,N_5144,N_4561);
nor U6789 (N_6789,N_5385,N_5111);
nor U6790 (N_6790,N_4260,N_5704);
or U6791 (N_6791,N_5539,N_5036);
xnor U6792 (N_6792,N_5192,N_5106);
or U6793 (N_6793,N_5109,N_4712);
nand U6794 (N_6794,N_5336,N_4735);
nor U6795 (N_6795,N_4395,N_4257);
or U6796 (N_6796,N_4121,N_5243);
or U6797 (N_6797,N_4158,N_4922);
xor U6798 (N_6798,N_5818,N_4754);
nand U6799 (N_6799,N_4356,N_5900);
xor U6800 (N_6800,N_4686,N_5249);
nor U6801 (N_6801,N_5779,N_5503);
and U6802 (N_6802,N_5254,N_5645);
nand U6803 (N_6803,N_5082,N_4909);
nor U6804 (N_6804,N_5585,N_4666);
xnor U6805 (N_6805,N_5816,N_4678);
nor U6806 (N_6806,N_5388,N_5583);
nand U6807 (N_6807,N_5250,N_4590);
nand U6808 (N_6808,N_4918,N_4514);
or U6809 (N_6809,N_4950,N_4643);
nor U6810 (N_6810,N_5924,N_4062);
nand U6811 (N_6811,N_5776,N_5729);
nand U6812 (N_6812,N_5980,N_4080);
or U6813 (N_6813,N_4797,N_4879);
and U6814 (N_6814,N_4867,N_4640);
or U6815 (N_6815,N_4374,N_5412);
nand U6816 (N_6816,N_4497,N_5127);
nand U6817 (N_6817,N_4734,N_5654);
nor U6818 (N_6818,N_5434,N_5287);
nand U6819 (N_6819,N_4809,N_5807);
and U6820 (N_6820,N_5185,N_5799);
xnor U6821 (N_6821,N_5955,N_5672);
or U6822 (N_6822,N_4736,N_5927);
xor U6823 (N_6823,N_5154,N_4428);
and U6824 (N_6824,N_4361,N_4935);
or U6825 (N_6825,N_5682,N_5178);
nand U6826 (N_6826,N_4057,N_4144);
and U6827 (N_6827,N_5080,N_5215);
or U6828 (N_6828,N_4804,N_5567);
nor U6829 (N_6829,N_5401,N_4028);
nand U6830 (N_6830,N_4610,N_5787);
or U6831 (N_6831,N_4165,N_5060);
xor U6832 (N_6832,N_5894,N_5856);
or U6833 (N_6833,N_5889,N_5543);
or U6834 (N_6834,N_5372,N_5891);
nor U6835 (N_6835,N_4919,N_4116);
nor U6836 (N_6836,N_5006,N_4853);
nand U6837 (N_6837,N_4727,N_5632);
nand U6838 (N_6838,N_4517,N_5205);
nand U6839 (N_6839,N_4508,N_5031);
nand U6840 (N_6840,N_4543,N_4156);
nor U6841 (N_6841,N_4708,N_5449);
nor U6842 (N_6842,N_4373,N_4100);
nand U6843 (N_6843,N_4519,N_4350);
or U6844 (N_6844,N_4805,N_4530);
and U6845 (N_6845,N_5389,N_5844);
and U6846 (N_6846,N_4432,N_4050);
nand U6847 (N_6847,N_4653,N_5699);
nand U6848 (N_6848,N_5322,N_5974);
nand U6849 (N_6849,N_4849,N_4955);
and U6850 (N_6850,N_5152,N_5788);
or U6851 (N_6851,N_5285,N_5526);
and U6852 (N_6852,N_5530,N_5778);
or U6853 (N_6853,N_5369,N_4434);
nor U6854 (N_6854,N_5815,N_4781);
or U6855 (N_6855,N_5794,N_4604);
nor U6856 (N_6856,N_4560,N_4017);
or U6857 (N_6857,N_5391,N_5981);
nand U6858 (N_6858,N_5406,N_5367);
nor U6859 (N_6859,N_5679,N_4135);
nor U6860 (N_6860,N_5433,N_4969);
nand U6861 (N_6861,N_4546,N_5298);
nor U6862 (N_6862,N_4636,N_4750);
nand U6863 (N_6863,N_5179,N_5609);
nor U6864 (N_6864,N_4240,N_5437);
nand U6865 (N_6865,N_4819,N_5918);
and U6866 (N_6866,N_4963,N_4921);
xnor U6867 (N_6867,N_5826,N_5459);
and U6868 (N_6868,N_4383,N_5940);
nand U6869 (N_6869,N_4269,N_4912);
or U6870 (N_6870,N_5355,N_5660);
and U6871 (N_6871,N_5904,N_4690);
nand U6872 (N_6872,N_4111,N_5286);
nor U6873 (N_6873,N_4991,N_4321);
nand U6874 (N_6874,N_5007,N_4670);
or U6875 (N_6875,N_4092,N_4939);
nor U6876 (N_6876,N_5930,N_4758);
nand U6877 (N_6877,N_4131,N_5920);
or U6878 (N_6878,N_5548,N_4910);
nand U6879 (N_6879,N_4178,N_4263);
nand U6880 (N_6880,N_4928,N_5696);
nand U6881 (N_6881,N_5222,N_4834);
nor U6882 (N_6882,N_4516,N_4259);
nand U6883 (N_6883,N_5429,N_4621);
and U6884 (N_6884,N_4460,N_5504);
nor U6885 (N_6885,N_4351,N_5289);
or U6886 (N_6886,N_5634,N_4166);
and U6887 (N_6887,N_5393,N_5377);
and U6888 (N_6888,N_5999,N_4931);
xnor U6889 (N_6889,N_5311,N_5258);
nor U6890 (N_6890,N_5232,N_4091);
or U6891 (N_6891,N_5519,N_5502);
nand U6892 (N_6892,N_5024,N_4044);
nor U6893 (N_6893,N_4288,N_4346);
xor U6894 (N_6894,N_5884,N_5849);
xnor U6895 (N_6895,N_5711,N_4966);
xor U6896 (N_6896,N_4405,N_5714);
nand U6897 (N_6897,N_4706,N_5354);
nor U6898 (N_6898,N_4183,N_5057);
and U6899 (N_6899,N_4953,N_5566);
or U6900 (N_6900,N_5763,N_5259);
nand U6901 (N_6901,N_4852,N_4381);
and U6902 (N_6902,N_5108,N_4784);
and U6903 (N_6903,N_4798,N_5755);
or U6904 (N_6904,N_5227,N_5643);
or U6905 (N_6905,N_5483,N_5507);
or U6906 (N_6906,N_4705,N_4496);
nor U6907 (N_6907,N_5010,N_4009);
xnor U6908 (N_6908,N_5664,N_4582);
nand U6909 (N_6909,N_4509,N_4629);
nor U6910 (N_6910,N_5494,N_5443);
and U6911 (N_6911,N_4623,N_4368);
nand U6912 (N_6912,N_5040,N_4588);
and U6913 (N_6913,N_5829,N_4778);
nand U6914 (N_6914,N_4773,N_4538);
nor U6915 (N_6915,N_4716,N_5979);
and U6916 (N_6916,N_4522,N_5556);
nor U6917 (N_6917,N_4067,N_4013);
and U6918 (N_6918,N_4595,N_5708);
or U6919 (N_6919,N_5997,N_4965);
or U6920 (N_6920,N_5019,N_4732);
and U6921 (N_6921,N_5183,N_5883);
or U6922 (N_6922,N_4630,N_4320);
nand U6923 (N_6923,N_4871,N_5771);
nor U6924 (N_6924,N_5665,N_4160);
nand U6925 (N_6925,N_5182,N_5817);
nand U6926 (N_6926,N_5345,N_5790);
nand U6927 (N_6927,N_5630,N_4632);
or U6928 (N_6928,N_4348,N_4887);
nor U6929 (N_6929,N_4529,N_5288);
nand U6930 (N_6930,N_4461,N_4378);
and U6931 (N_6931,N_4370,N_4494);
or U6932 (N_6932,N_4688,N_4790);
and U6933 (N_6933,N_4236,N_5265);
and U6934 (N_6934,N_4085,N_4387);
or U6935 (N_6935,N_5229,N_4687);
nand U6936 (N_6936,N_4415,N_4601);
and U6937 (N_6937,N_5591,N_5211);
or U6938 (N_6938,N_5426,N_4586);
nand U6939 (N_6939,N_4174,N_4430);
or U6940 (N_6940,N_5743,N_4679);
and U6941 (N_6941,N_4866,N_5055);
or U6942 (N_6942,N_4055,N_5754);
or U6943 (N_6943,N_5897,N_4715);
or U6944 (N_6944,N_5902,N_4046);
nand U6945 (N_6945,N_4613,N_5223);
nand U6946 (N_6946,N_4889,N_5535);
and U6947 (N_6947,N_4792,N_5631);
nand U6948 (N_6948,N_4253,N_4476);
xor U6949 (N_6949,N_5888,N_5557);
xnor U6950 (N_6950,N_5513,N_4195);
and U6951 (N_6951,N_5517,N_5368);
nand U6952 (N_6952,N_4197,N_4559);
or U6953 (N_6953,N_5339,N_4343);
and U6954 (N_6954,N_4693,N_5852);
nor U6955 (N_6955,N_4578,N_5202);
nor U6956 (N_6956,N_4435,N_4234);
and U6957 (N_6957,N_5805,N_5025);
nand U6958 (N_6958,N_4147,N_5295);
nand U6959 (N_6959,N_4895,N_5410);
xor U6960 (N_6960,N_5069,N_4850);
nor U6961 (N_6961,N_4268,N_4230);
and U6962 (N_6962,N_5878,N_5570);
or U6963 (N_6963,N_5864,N_5638);
xor U6964 (N_6964,N_5156,N_5041);
nand U6965 (N_6965,N_4598,N_4161);
and U6966 (N_6966,N_5218,N_4466);
nand U6967 (N_6967,N_4087,N_4806);
nand U6968 (N_6968,N_4349,N_4818);
and U6969 (N_6969,N_5241,N_4438);
nand U6970 (N_6970,N_4752,N_4340);
xor U6971 (N_6971,N_5018,N_4990);
and U6972 (N_6972,N_4980,N_4211);
or U6973 (N_6973,N_5420,N_4883);
and U6974 (N_6974,N_4944,N_5253);
nor U6975 (N_6975,N_4684,N_5128);
or U6976 (N_6976,N_5084,N_4672);
and U6977 (N_6977,N_5067,N_4692);
or U6978 (N_6978,N_5442,N_5262);
nand U6979 (N_6979,N_5866,N_5489);
and U6980 (N_6980,N_5139,N_4801);
nand U6981 (N_6981,N_4576,N_4241);
nand U6982 (N_6982,N_4353,N_4278);
nand U6983 (N_6983,N_5457,N_5400);
and U6984 (N_6984,N_5386,N_4650);
or U6985 (N_6985,N_4645,N_4176);
and U6986 (N_6986,N_5916,N_4998);
nor U6987 (N_6987,N_5396,N_5353);
xnor U6988 (N_6988,N_5321,N_5877);
nor U6989 (N_6989,N_4788,N_5206);
and U6990 (N_6990,N_5201,N_4478);
and U6991 (N_6991,N_5662,N_5365);
or U6992 (N_6992,N_5226,N_5394);
or U6993 (N_6993,N_5044,N_4501);
nand U6994 (N_6994,N_5072,N_5092);
or U6995 (N_6995,N_4485,N_4660);
and U6996 (N_6996,N_5405,N_4029);
xor U6997 (N_6997,N_4870,N_4447);
nor U6998 (N_6998,N_4637,N_5308);
and U6999 (N_6999,N_4859,N_4675);
or U7000 (N_7000,N_5066,N_5602);
xnor U7001 (N_7001,N_4940,N_5700);
nor U7002 (N_7002,N_4466,N_4880);
or U7003 (N_7003,N_5628,N_5192);
or U7004 (N_7004,N_4640,N_5156);
and U7005 (N_7005,N_4240,N_5143);
nor U7006 (N_7006,N_5449,N_4789);
and U7007 (N_7007,N_4592,N_5262);
or U7008 (N_7008,N_5781,N_4957);
and U7009 (N_7009,N_4778,N_5528);
or U7010 (N_7010,N_5269,N_5628);
nand U7011 (N_7011,N_4110,N_4968);
or U7012 (N_7012,N_4886,N_4304);
or U7013 (N_7013,N_5356,N_5854);
xnor U7014 (N_7014,N_4153,N_5896);
or U7015 (N_7015,N_5884,N_4059);
or U7016 (N_7016,N_4186,N_4367);
xor U7017 (N_7017,N_4566,N_4607);
and U7018 (N_7018,N_4720,N_4555);
nand U7019 (N_7019,N_5768,N_5177);
and U7020 (N_7020,N_4473,N_5548);
nand U7021 (N_7021,N_4065,N_4797);
nor U7022 (N_7022,N_4268,N_5031);
and U7023 (N_7023,N_4092,N_5462);
nor U7024 (N_7024,N_4084,N_5916);
and U7025 (N_7025,N_4213,N_4342);
and U7026 (N_7026,N_5396,N_4716);
and U7027 (N_7027,N_5359,N_5646);
nor U7028 (N_7028,N_5517,N_4642);
nor U7029 (N_7029,N_4276,N_5617);
nand U7030 (N_7030,N_4533,N_4431);
or U7031 (N_7031,N_4451,N_4395);
or U7032 (N_7032,N_5020,N_5505);
nand U7033 (N_7033,N_4888,N_4047);
nand U7034 (N_7034,N_4605,N_4277);
nor U7035 (N_7035,N_4718,N_5405);
and U7036 (N_7036,N_5562,N_4506);
nor U7037 (N_7037,N_5821,N_5979);
nor U7038 (N_7038,N_5965,N_5533);
or U7039 (N_7039,N_5637,N_4955);
nand U7040 (N_7040,N_5190,N_4306);
nand U7041 (N_7041,N_5879,N_5805);
xor U7042 (N_7042,N_4861,N_5452);
xnor U7043 (N_7043,N_5580,N_5710);
and U7044 (N_7044,N_4389,N_5949);
and U7045 (N_7045,N_4227,N_5864);
xnor U7046 (N_7046,N_4719,N_5006);
nor U7047 (N_7047,N_4736,N_4682);
or U7048 (N_7048,N_4599,N_5156);
nand U7049 (N_7049,N_5538,N_5406);
nand U7050 (N_7050,N_4857,N_4602);
and U7051 (N_7051,N_5556,N_4492);
or U7052 (N_7052,N_5213,N_5169);
nor U7053 (N_7053,N_4702,N_5961);
nand U7054 (N_7054,N_5521,N_5110);
nor U7055 (N_7055,N_4061,N_4560);
and U7056 (N_7056,N_4569,N_4644);
or U7057 (N_7057,N_4261,N_4957);
and U7058 (N_7058,N_5405,N_4285);
nand U7059 (N_7059,N_5374,N_4396);
or U7060 (N_7060,N_4280,N_4294);
or U7061 (N_7061,N_4418,N_4424);
nor U7062 (N_7062,N_4557,N_5839);
and U7063 (N_7063,N_5940,N_5158);
nand U7064 (N_7064,N_4084,N_4293);
and U7065 (N_7065,N_4850,N_4224);
or U7066 (N_7066,N_5527,N_4584);
xor U7067 (N_7067,N_5213,N_5328);
and U7068 (N_7068,N_4789,N_5557);
or U7069 (N_7069,N_4495,N_5108);
or U7070 (N_7070,N_5397,N_5320);
and U7071 (N_7071,N_4702,N_4146);
xor U7072 (N_7072,N_5741,N_4468);
or U7073 (N_7073,N_5625,N_4472);
and U7074 (N_7074,N_4310,N_4189);
or U7075 (N_7075,N_5405,N_4533);
or U7076 (N_7076,N_4570,N_5086);
or U7077 (N_7077,N_4120,N_4237);
nor U7078 (N_7078,N_4568,N_5151);
or U7079 (N_7079,N_5653,N_5624);
and U7080 (N_7080,N_5752,N_4624);
or U7081 (N_7081,N_5379,N_4001);
and U7082 (N_7082,N_4007,N_5369);
or U7083 (N_7083,N_5364,N_4798);
and U7084 (N_7084,N_4273,N_5802);
or U7085 (N_7085,N_4999,N_5730);
and U7086 (N_7086,N_5429,N_4172);
or U7087 (N_7087,N_4450,N_4838);
or U7088 (N_7088,N_5614,N_4635);
nand U7089 (N_7089,N_5899,N_4191);
xnor U7090 (N_7090,N_5867,N_5218);
nand U7091 (N_7091,N_4643,N_4067);
nor U7092 (N_7092,N_5638,N_4282);
nor U7093 (N_7093,N_5372,N_4829);
xnor U7094 (N_7094,N_5071,N_5148);
nand U7095 (N_7095,N_5808,N_4601);
and U7096 (N_7096,N_5719,N_4952);
nor U7097 (N_7097,N_5651,N_5707);
nor U7098 (N_7098,N_5018,N_5086);
xnor U7099 (N_7099,N_4158,N_5104);
nor U7100 (N_7100,N_5826,N_4478);
nor U7101 (N_7101,N_5575,N_4919);
or U7102 (N_7102,N_5435,N_4157);
nor U7103 (N_7103,N_4666,N_4271);
and U7104 (N_7104,N_4840,N_5922);
nand U7105 (N_7105,N_4210,N_5603);
or U7106 (N_7106,N_5447,N_5054);
nand U7107 (N_7107,N_4330,N_5765);
nor U7108 (N_7108,N_4265,N_4309);
nand U7109 (N_7109,N_5023,N_5807);
xnor U7110 (N_7110,N_5396,N_5606);
or U7111 (N_7111,N_5371,N_5907);
and U7112 (N_7112,N_5557,N_4965);
or U7113 (N_7113,N_4372,N_4789);
nand U7114 (N_7114,N_5128,N_4654);
nand U7115 (N_7115,N_4655,N_5162);
nor U7116 (N_7116,N_4728,N_5655);
nand U7117 (N_7117,N_5739,N_5443);
or U7118 (N_7118,N_4723,N_5892);
and U7119 (N_7119,N_4408,N_5346);
or U7120 (N_7120,N_4269,N_5608);
nand U7121 (N_7121,N_4347,N_4756);
nand U7122 (N_7122,N_5100,N_5323);
xor U7123 (N_7123,N_5226,N_5591);
nand U7124 (N_7124,N_4073,N_5667);
or U7125 (N_7125,N_5824,N_4708);
and U7126 (N_7126,N_5504,N_5097);
or U7127 (N_7127,N_5408,N_5388);
and U7128 (N_7128,N_5127,N_4979);
nor U7129 (N_7129,N_4800,N_5417);
or U7130 (N_7130,N_4613,N_5611);
nand U7131 (N_7131,N_5649,N_5473);
or U7132 (N_7132,N_5208,N_4314);
nand U7133 (N_7133,N_4403,N_5919);
nand U7134 (N_7134,N_5102,N_4580);
and U7135 (N_7135,N_5523,N_4632);
xnor U7136 (N_7136,N_5235,N_5031);
and U7137 (N_7137,N_4798,N_5764);
nand U7138 (N_7138,N_4501,N_4769);
and U7139 (N_7139,N_5096,N_4548);
and U7140 (N_7140,N_4554,N_5006);
and U7141 (N_7141,N_4684,N_5225);
and U7142 (N_7142,N_5004,N_4887);
nand U7143 (N_7143,N_4361,N_5027);
nor U7144 (N_7144,N_4486,N_5393);
nand U7145 (N_7145,N_5308,N_4500);
or U7146 (N_7146,N_5843,N_4119);
or U7147 (N_7147,N_4635,N_5498);
or U7148 (N_7148,N_4192,N_4454);
and U7149 (N_7149,N_4762,N_5234);
nand U7150 (N_7150,N_5111,N_4820);
nand U7151 (N_7151,N_4143,N_5575);
or U7152 (N_7152,N_4416,N_4788);
nand U7153 (N_7153,N_5535,N_5990);
nand U7154 (N_7154,N_4623,N_4912);
xor U7155 (N_7155,N_5371,N_5660);
or U7156 (N_7156,N_5251,N_4681);
nor U7157 (N_7157,N_4207,N_4009);
nor U7158 (N_7158,N_4429,N_4736);
or U7159 (N_7159,N_5824,N_5241);
nor U7160 (N_7160,N_5221,N_4301);
nor U7161 (N_7161,N_5826,N_4113);
or U7162 (N_7162,N_5975,N_5199);
nor U7163 (N_7163,N_5279,N_5739);
and U7164 (N_7164,N_4742,N_5349);
and U7165 (N_7165,N_5792,N_5591);
nand U7166 (N_7166,N_5100,N_4415);
or U7167 (N_7167,N_5769,N_5800);
xnor U7168 (N_7168,N_5509,N_4170);
or U7169 (N_7169,N_4950,N_5961);
nand U7170 (N_7170,N_4932,N_5777);
nor U7171 (N_7171,N_5494,N_5000);
and U7172 (N_7172,N_5714,N_4321);
nor U7173 (N_7173,N_4673,N_5677);
or U7174 (N_7174,N_5733,N_5253);
nand U7175 (N_7175,N_4466,N_5385);
nand U7176 (N_7176,N_5663,N_5429);
xor U7177 (N_7177,N_4257,N_4704);
or U7178 (N_7178,N_5746,N_5684);
nand U7179 (N_7179,N_5711,N_5157);
nor U7180 (N_7180,N_5423,N_5480);
nor U7181 (N_7181,N_4079,N_5871);
nand U7182 (N_7182,N_5190,N_5080);
nand U7183 (N_7183,N_5871,N_5506);
or U7184 (N_7184,N_4383,N_4842);
or U7185 (N_7185,N_4254,N_5913);
and U7186 (N_7186,N_4369,N_5033);
and U7187 (N_7187,N_4770,N_5679);
or U7188 (N_7188,N_5045,N_5154);
nand U7189 (N_7189,N_4646,N_4407);
nand U7190 (N_7190,N_5656,N_4322);
and U7191 (N_7191,N_4577,N_5029);
nand U7192 (N_7192,N_4055,N_5779);
xor U7193 (N_7193,N_4913,N_5251);
nand U7194 (N_7194,N_4754,N_4618);
and U7195 (N_7195,N_5810,N_5122);
or U7196 (N_7196,N_4234,N_4656);
nand U7197 (N_7197,N_5520,N_4204);
nor U7198 (N_7198,N_4169,N_4886);
nand U7199 (N_7199,N_5608,N_4655);
and U7200 (N_7200,N_5474,N_5914);
or U7201 (N_7201,N_5092,N_5835);
or U7202 (N_7202,N_5773,N_5218);
nand U7203 (N_7203,N_5037,N_4165);
or U7204 (N_7204,N_5140,N_5991);
or U7205 (N_7205,N_5312,N_4523);
nor U7206 (N_7206,N_5859,N_4684);
nand U7207 (N_7207,N_5472,N_5660);
nor U7208 (N_7208,N_5033,N_5534);
or U7209 (N_7209,N_4299,N_5707);
nand U7210 (N_7210,N_4516,N_4407);
and U7211 (N_7211,N_4266,N_4235);
nand U7212 (N_7212,N_5748,N_5164);
nor U7213 (N_7213,N_5267,N_5558);
nand U7214 (N_7214,N_5615,N_5460);
or U7215 (N_7215,N_4696,N_4398);
nor U7216 (N_7216,N_5027,N_5203);
and U7217 (N_7217,N_4043,N_5128);
or U7218 (N_7218,N_4621,N_5174);
nor U7219 (N_7219,N_5766,N_4665);
or U7220 (N_7220,N_4437,N_4348);
and U7221 (N_7221,N_5692,N_5111);
nor U7222 (N_7222,N_5659,N_4631);
and U7223 (N_7223,N_4173,N_5530);
xor U7224 (N_7224,N_4921,N_5977);
nor U7225 (N_7225,N_5959,N_4601);
or U7226 (N_7226,N_5185,N_4117);
nand U7227 (N_7227,N_5452,N_4591);
and U7228 (N_7228,N_4320,N_5580);
or U7229 (N_7229,N_5666,N_4228);
and U7230 (N_7230,N_4072,N_5449);
nand U7231 (N_7231,N_4396,N_5919);
nor U7232 (N_7232,N_5611,N_5028);
nand U7233 (N_7233,N_4426,N_4323);
and U7234 (N_7234,N_4465,N_5127);
xor U7235 (N_7235,N_5671,N_5467);
nor U7236 (N_7236,N_5531,N_5229);
xnor U7237 (N_7237,N_4378,N_5457);
xor U7238 (N_7238,N_5669,N_4635);
or U7239 (N_7239,N_5197,N_5578);
xnor U7240 (N_7240,N_5471,N_4165);
nand U7241 (N_7241,N_4318,N_5531);
and U7242 (N_7242,N_4542,N_5988);
nand U7243 (N_7243,N_4579,N_5192);
and U7244 (N_7244,N_4099,N_4454);
and U7245 (N_7245,N_5563,N_4009);
and U7246 (N_7246,N_5843,N_5085);
and U7247 (N_7247,N_4552,N_5903);
nor U7248 (N_7248,N_5593,N_4248);
nor U7249 (N_7249,N_5807,N_5052);
nor U7250 (N_7250,N_4264,N_5495);
or U7251 (N_7251,N_5778,N_4478);
or U7252 (N_7252,N_4904,N_5204);
and U7253 (N_7253,N_5917,N_5214);
or U7254 (N_7254,N_5713,N_5014);
nand U7255 (N_7255,N_5102,N_5410);
and U7256 (N_7256,N_4661,N_4436);
nand U7257 (N_7257,N_4751,N_4011);
nand U7258 (N_7258,N_5986,N_5941);
xnor U7259 (N_7259,N_5233,N_4740);
nand U7260 (N_7260,N_4109,N_4196);
or U7261 (N_7261,N_4041,N_5865);
xor U7262 (N_7262,N_5821,N_5191);
and U7263 (N_7263,N_5069,N_5125);
and U7264 (N_7264,N_5976,N_5266);
nand U7265 (N_7265,N_5718,N_4399);
and U7266 (N_7266,N_4915,N_5592);
xnor U7267 (N_7267,N_5607,N_5099);
and U7268 (N_7268,N_5910,N_5147);
nor U7269 (N_7269,N_4636,N_4528);
and U7270 (N_7270,N_5100,N_4311);
or U7271 (N_7271,N_4995,N_5246);
and U7272 (N_7272,N_4954,N_4731);
or U7273 (N_7273,N_5365,N_4812);
and U7274 (N_7274,N_5022,N_4162);
nand U7275 (N_7275,N_4649,N_5150);
nor U7276 (N_7276,N_4534,N_5345);
or U7277 (N_7277,N_5258,N_4921);
or U7278 (N_7278,N_5344,N_5302);
nor U7279 (N_7279,N_4745,N_5218);
or U7280 (N_7280,N_5466,N_4161);
and U7281 (N_7281,N_5534,N_4159);
nand U7282 (N_7282,N_5503,N_5284);
nor U7283 (N_7283,N_4678,N_4728);
or U7284 (N_7284,N_4274,N_4754);
or U7285 (N_7285,N_5460,N_5774);
or U7286 (N_7286,N_4214,N_4796);
nand U7287 (N_7287,N_4207,N_4597);
and U7288 (N_7288,N_5599,N_4874);
nand U7289 (N_7289,N_4103,N_4500);
nand U7290 (N_7290,N_5526,N_4460);
xor U7291 (N_7291,N_5020,N_4952);
or U7292 (N_7292,N_5552,N_4406);
nor U7293 (N_7293,N_5751,N_5601);
nand U7294 (N_7294,N_4707,N_4991);
and U7295 (N_7295,N_4777,N_4488);
or U7296 (N_7296,N_5008,N_4333);
or U7297 (N_7297,N_4598,N_5501);
xnor U7298 (N_7298,N_5717,N_5584);
nor U7299 (N_7299,N_5762,N_5901);
nor U7300 (N_7300,N_4255,N_5203);
nor U7301 (N_7301,N_4166,N_5416);
nor U7302 (N_7302,N_4672,N_5772);
or U7303 (N_7303,N_5339,N_4499);
xnor U7304 (N_7304,N_4010,N_4752);
and U7305 (N_7305,N_5484,N_5752);
xor U7306 (N_7306,N_4801,N_4095);
xor U7307 (N_7307,N_4367,N_4024);
nand U7308 (N_7308,N_5189,N_5544);
or U7309 (N_7309,N_5943,N_4844);
nand U7310 (N_7310,N_5414,N_4565);
and U7311 (N_7311,N_5671,N_5951);
nor U7312 (N_7312,N_4478,N_4008);
nand U7313 (N_7313,N_4742,N_5324);
nor U7314 (N_7314,N_5110,N_5745);
or U7315 (N_7315,N_5666,N_5021);
nand U7316 (N_7316,N_4725,N_5011);
and U7317 (N_7317,N_4614,N_4700);
nor U7318 (N_7318,N_5022,N_5583);
or U7319 (N_7319,N_4343,N_5765);
nand U7320 (N_7320,N_4379,N_4779);
and U7321 (N_7321,N_4642,N_4308);
and U7322 (N_7322,N_5152,N_5525);
or U7323 (N_7323,N_5723,N_4176);
nor U7324 (N_7324,N_4573,N_5899);
or U7325 (N_7325,N_5511,N_5520);
nand U7326 (N_7326,N_4619,N_5402);
xnor U7327 (N_7327,N_4079,N_5097);
nor U7328 (N_7328,N_4446,N_4803);
or U7329 (N_7329,N_5916,N_5727);
nor U7330 (N_7330,N_4850,N_4775);
and U7331 (N_7331,N_4199,N_4328);
and U7332 (N_7332,N_4448,N_4051);
nand U7333 (N_7333,N_5758,N_5289);
or U7334 (N_7334,N_4108,N_5136);
nand U7335 (N_7335,N_5107,N_5101);
and U7336 (N_7336,N_5375,N_4067);
xor U7337 (N_7337,N_5407,N_5762);
nand U7338 (N_7338,N_4571,N_4535);
or U7339 (N_7339,N_5286,N_4481);
or U7340 (N_7340,N_5004,N_4538);
nor U7341 (N_7341,N_4420,N_4542);
or U7342 (N_7342,N_4468,N_5363);
nor U7343 (N_7343,N_5566,N_4240);
xnor U7344 (N_7344,N_4898,N_4968);
nand U7345 (N_7345,N_5650,N_5960);
nand U7346 (N_7346,N_5684,N_5927);
or U7347 (N_7347,N_4237,N_5708);
nand U7348 (N_7348,N_5048,N_4077);
nor U7349 (N_7349,N_4484,N_4705);
nor U7350 (N_7350,N_5927,N_4790);
or U7351 (N_7351,N_5033,N_4933);
and U7352 (N_7352,N_4197,N_5234);
xnor U7353 (N_7353,N_4177,N_5531);
nor U7354 (N_7354,N_4578,N_4503);
xor U7355 (N_7355,N_5248,N_4389);
and U7356 (N_7356,N_5469,N_5986);
or U7357 (N_7357,N_5041,N_5964);
nor U7358 (N_7358,N_5273,N_4134);
nand U7359 (N_7359,N_4125,N_5675);
and U7360 (N_7360,N_5857,N_5932);
and U7361 (N_7361,N_5375,N_5158);
or U7362 (N_7362,N_5034,N_5040);
xnor U7363 (N_7363,N_4501,N_4222);
xnor U7364 (N_7364,N_5334,N_5859);
nand U7365 (N_7365,N_5910,N_5921);
nor U7366 (N_7366,N_5795,N_4478);
nor U7367 (N_7367,N_4652,N_5265);
nor U7368 (N_7368,N_5798,N_4930);
or U7369 (N_7369,N_5512,N_4253);
xnor U7370 (N_7370,N_4665,N_4768);
and U7371 (N_7371,N_4128,N_5977);
and U7372 (N_7372,N_4401,N_5106);
nand U7373 (N_7373,N_5352,N_4692);
nand U7374 (N_7374,N_5889,N_5459);
xor U7375 (N_7375,N_4818,N_5105);
or U7376 (N_7376,N_4082,N_5282);
and U7377 (N_7377,N_5684,N_4163);
nor U7378 (N_7378,N_5946,N_4945);
and U7379 (N_7379,N_4706,N_5823);
nand U7380 (N_7380,N_4628,N_5731);
nor U7381 (N_7381,N_5355,N_4151);
nand U7382 (N_7382,N_4986,N_4387);
and U7383 (N_7383,N_5221,N_5000);
xnor U7384 (N_7384,N_4565,N_4595);
or U7385 (N_7385,N_5407,N_4823);
nor U7386 (N_7386,N_4544,N_4630);
nor U7387 (N_7387,N_5673,N_5525);
nor U7388 (N_7388,N_4421,N_5833);
nand U7389 (N_7389,N_4725,N_4649);
nor U7390 (N_7390,N_5450,N_5217);
nand U7391 (N_7391,N_4977,N_4114);
nand U7392 (N_7392,N_4319,N_4059);
or U7393 (N_7393,N_4286,N_5287);
or U7394 (N_7394,N_4180,N_4333);
or U7395 (N_7395,N_5174,N_5676);
or U7396 (N_7396,N_4576,N_4526);
nor U7397 (N_7397,N_5313,N_4202);
and U7398 (N_7398,N_4132,N_5690);
or U7399 (N_7399,N_5189,N_5416);
nand U7400 (N_7400,N_4669,N_5326);
or U7401 (N_7401,N_5223,N_4804);
nor U7402 (N_7402,N_4696,N_5311);
nor U7403 (N_7403,N_4489,N_4966);
nor U7404 (N_7404,N_5630,N_4275);
nor U7405 (N_7405,N_5529,N_5440);
xnor U7406 (N_7406,N_5077,N_5645);
or U7407 (N_7407,N_5279,N_4517);
nand U7408 (N_7408,N_4576,N_5024);
and U7409 (N_7409,N_5717,N_4272);
or U7410 (N_7410,N_5137,N_4327);
or U7411 (N_7411,N_4906,N_5736);
nand U7412 (N_7412,N_5023,N_5329);
or U7413 (N_7413,N_4488,N_4512);
and U7414 (N_7414,N_4768,N_5769);
nand U7415 (N_7415,N_5649,N_4076);
nor U7416 (N_7416,N_4093,N_5999);
and U7417 (N_7417,N_5962,N_4566);
and U7418 (N_7418,N_5262,N_4608);
nor U7419 (N_7419,N_5043,N_5985);
and U7420 (N_7420,N_5081,N_5538);
or U7421 (N_7421,N_5162,N_4369);
or U7422 (N_7422,N_5746,N_4596);
or U7423 (N_7423,N_4300,N_5620);
or U7424 (N_7424,N_5525,N_5106);
nor U7425 (N_7425,N_4682,N_4088);
or U7426 (N_7426,N_5718,N_5529);
nor U7427 (N_7427,N_4994,N_5387);
nand U7428 (N_7428,N_5297,N_4526);
or U7429 (N_7429,N_4417,N_4341);
nand U7430 (N_7430,N_5348,N_5792);
nand U7431 (N_7431,N_4670,N_4877);
nand U7432 (N_7432,N_4156,N_4409);
and U7433 (N_7433,N_5527,N_5068);
or U7434 (N_7434,N_4812,N_4136);
and U7435 (N_7435,N_4377,N_4171);
or U7436 (N_7436,N_5935,N_4791);
nor U7437 (N_7437,N_5417,N_5908);
nand U7438 (N_7438,N_5512,N_4477);
or U7439 (N_7439,N_5892,N_5833);
or U7440 (N_7440,N_5625,N_5560);
nand U7441 (N_7441,N_5873,N_5680);
nor U7442 (N_7442,N_4657,N_4649);
and U7443 (N_7443,N_4614,N_4895);
nand U7444 (N_7444,N_5127,N_5386);
xor U7445 (N_7445,N_4030,N_5375);
and U7446 (N_7446,N_4002,N_4096);
nand U7447 (N_7447,N_5773,N_4798);
nor U7448 (N_7448,N_4628,N_5113);
nor U7449 (N_7449,N_5434,N_4759);
nand U7450 (N_7450,N_4213,N_5093);
or U7451 (N_7451,N_5898,N_5250);
or U7452 (N_7452,N_5382,N_5018);
nor U7453 (N_7453,N_5261,N_4771);
nand U7454 (N_7454,N_5775,N_4398);
nand U7455 (N_7455,N_5410,N_5161);
xnor U7456 (N_7456,N_4151,N_4528);
nand U7457 (N_7457,N_5060,N_4091);
nand U7458 (N_7458,N_4819,N_4173);
nor U7459 (N_7459,N_4520,N_5238);
nand U7460 (N_7460,N_5170,N_4433);
nand U7461 (N_7461,N_4102,N_5950);
nand U7462 (N_7462,N_5303,N_5653);
and U7463 (N_7463,N_5922,N_4972);
and U7464 (N_7464,N_5944,N_4520);
nand U7465 (N_7465,N_4830,N_5322);
nand U7466 (N_7466,N_4767,N_5499);
nand U7467 (N_7467,N_4641,N_5276);
nor U7468 (N_7468,N_5475,N_4105);
xnor U7469 (N_7469,N_4413,N_5251);
xnor U7470 (N_7470,N_4024,N_5724);
nand U7471 (N_7471,N_4747,N_5082);
nor U7472 (N_7472,N_5457,N_5109);
nand U7473 (N_7473,N_5467,N_4228);
and U7474 (N_7474,N_4681,N_5521);
or U7475 (N_7475,N_5379,N_5595);
and U7476 (N_7476,N_5127,N_4831);
and U7477 (N_7477,N_5461,N_4246);
nand U7478 (N_7478,N_4423,N_4543);
nor U7479 (N_7479,N_4092,N_5825);
and U7480 (N_7480,N_4583,N_5584);
or U7481 (N_7481,N_5558,N_5062);
and U7482 (N_7482,N_5779,N_5827);
nor U7483 (N_7483,N_4401,N_4820);
nand U7484 (N_7484,N_5617,N_5598);
and U7485 (N_7485,N_5794,N_5631);
nor U7486 (N_7486,N_5432,N_4896);
nor U7487 (N_7487,N_4553,N_5913);
and U7488 (N_7488,N_5911,N_4427);
nor U7489 (N_7489,N_5032,N_4605);
and U7490 (N_7490,N_4706,N_4433);
nand U7491 (N_7491,N_4641,N_5525);
nand U7492 (N_7492,N_5998,N_4451);
nand U7493 (N_7493,N_4720,N_4743);
and U7494 (N_7494,N_5960,N_5643);
and U7495 (N_7495,N_5094,N_5007);
and U7496 (N_7496,N_4030,N_4199);
nand U7497 (N_7497,N_5802,N_4018);
nor U7498 (N_7498,N_5082,N_5891);
xor U7499 (N_7499,N_5963,N_5125);
nand U7500 (N_7500,N_4718,N_4881);
or U7501 (N_7501,N_4755,N_5334);
nand U7502 (N_7502,N_5196,N_5135);
or U7503 (N_7503,N_5486,N_5042);
or U7504 (N_7504,N_4723,N_4748);
nand U7505 (N_7505,N_4100,N_4097);
xnor U7506 (N_7506,N_4654,N_5208);
nand U7507 (N_7507,N_5089,N_5530);
or U7508 (N_7508,N_4595,N_5900);
or U7509 (N_7509,N_4124,N_4495);
and U7510 (N_7510,N_5498,N_4065);
nand U7511 (N_7511,N_5279,N_4727);
nor U7512 (N_7512,N_4300,N_5920);
nand U7513 (N_7513,N_5279,N_5020);
or U7514 (N_7514,N_4328,N_5945);
nor U7515 (N_7515,N_4615,N_4918);
and U7516 (N_7516,N_5173,N_5883);
nor U7517 (N_7517,N_5690,N_4011);
nand U7518 (N_7518,N_4256,N_4220);
and U7519 (N_7519,N_4684,N_5436);
nand U7520 (N_7520,N_5848,N_4275);
and U7521 (N_7521,N_5293,N_4211);
or U7522 (N_7522,N_4583,N_4661);
nor U7523 (N_7523,N_5388,N_4035);
or U7524 (N_7524,N_5023,N_4957);
or U7525 (N_7525,N_4032,N_4590);
or U7526 (N_7526,N_4508,N_5495);
and U7527 (N_7527,N_4320,N_4799);
and U7528 (N_7528,N_4059,N_4428);
nand U7529 (N_7529,N_5204,N_4418);
nand U7530 (N_7530,N_5703,N_4625);
nor U7531 (N_7531,N_5412,N_4382);
nand U7532 (N_7532,N_4042,N_4215);
and U7533 (N_7533,N_4507,N_4125);
or U7534 (N_7534,N_5403,N_5839);
nand U7535 (N_7535,N_4408,N_4702);
nand U7536 (N_7536,N_4597,N_5087);
nand U7537 (N_7537,N_5812,N_4572);
nand U7538 (N_7538,N_4058,N_5646);
nor U7539 (N_7539,N_5639,N_5091);
or U7540 (N_7540,N_4547,N_4240);
nand U7541 (N_7541,N_5967,N_5739);
or U7542 (N_7542,N_5309,N_4181);
and U7543 (N_7543,N_4951,N_5120);
nand U7544 (N_7544,N_4037,N_4032);
and U7545 (N_7545,N_4464,N_4991);
nor U7546 (N_7546,N_4779,N_4429);
nand U7547 (N_7547,N_5318,N_5716);
or U7548 (N_7548,N_5170,N_5043);
nor U7549 (N_7549,N_4540,N_5211);
or U7550 (N_7550,N_4642,N_4294);
or U7551 (N_7551,N_4416,N_4537);
nand U7552 (N_7552,N_5756,N_5409);
and U7553 (N_7553,N_5255,N_5159);
nor U7554 (N_7554,N_4543,N_5559);
or U7555 (N_7555,N_4919,N_5804);
and U7556 (N_7556,N_5519,N_5164);
and U7557 (N_7557,N_4639,N_5484);
or U7558 (N_7558,N_5399,N_4652);
and U7559 (N_7559,N_4285,N_5127);
xnor U7560 (N_7560,N_4551,N_4805);
or U7561 (N_7561,N_4730,N_4262);
and U7562 (N_7562,N_4012,N_4912);
or U7563 (N_7563,N_4877,N_5453);
nand U7564 (N_7564,N_4325,N_5948);
nand U7565 (N_7565,N_4515,N_4117);
or U7566 (N_7566,N_5059,N_4336);
nand U7567 (N_7567,N_5643,N_5161);
nor U7568 (N_7568,N_4650,N_4422);
xnor U7569 (N_7569,N_5836,N_4405);
and U7570 (N_7570,N_5416,N_4487);
or U7571 (N_7571,N_4806,N_5317);
and U7572 (N_7572,N_4536,N_5950);
nor U7573 (N_7573,N_5419,N_5757);
nand U7574 (N_7574,N_4533,N_4297);
and U7575 (N_7575,N_4457,N_5712);
nand U7576 (N_7576,N_4521,N_5150);
and U7577 (N_7577,N_4345,N_4135);
or U7578 (N_7578,N_4826,N_4449);
nor U7579 (N_7579,N_4157,N_5583);
or U7580 (N_7580,N_4176,N_5593);
nor U7581 (N_7581,N_4755,N_5201);
nor U7582 (N_7582,N_5557,N_4110);
nor U7583 (N_7583,N_4222,N_5100);
or U7584 (N_7584,N_4734,N_4963);
nor U7585 (N_7585,N_4331,N_4376);
or U7586 (N_7586,N_4189,N_4165);
and U7587 (N_7587,N_4852,N_4555);
nand U7588 (N_7588,N_4995,N_4194);
xor U7589 (N_7589,N_5073,N_5041);
nand U7590 (N_7590,N_4770,N_5671);
or U7591 (N_7591,N_5199,N_5777);
or U7592 (N_7592,N_4101,N_5194);
and U7593 (N_7593,N_5910,N_5349);
xor U7594 (N_7594,N_5503,N_4536);
and U7595 (N_7595,N_5771,N_5291);
nor U7596 (N_7596,N_4053,N_4067);
and U7597 (N_7597,N_5867,N_5588);
nor U7598 (N_7598,N_4550,N_5748);
or U7599 (N_7599,N_4496,N_4629);
or U7600 (N_7600,N_4024,N_5590);
xnor U7601 (N_7601,N_4533,N_5968);
nor U7602 (N_7602,N_4556,N_5839);
and U7603 (N_7603,N_4548,N_4792);
or U7604 (N_7604,N_5577,N_5181);
nor U7605 (N_7605,N_5509,N_4212);
nor U7606 (N_7606,N_4892,N_4484);
nor U7607 (N_7607,N_5211,N_5552);
and U7608 (N_7608,N_5785,N_4918);
nand U7609 (N_7609,N_4482,N_4146);
and U7610 (N_7610,N_4518,N_4838);
nand U7611 (N_7611,N_5575,N_4891);
or U7612 (N_7612,N_4000,N_5287);
or U7613 (N_7613,N_5334,N_4300);
or U7614 (N_7614,N_4233,N_4185);
and U7615 (N_7615,N_4750,N_4496);
or U7616 (N_7616,N_4696,N_4536);
or U7617 (N_7617,N_5514,N_4049);
nand U7618 (N_7618,N_4460,N_5626);
nor U7619 (N_7619,N_5178,N_5867);
nand U7620 (N_7620,N_4035,N_5975);
xnor U7621 (N_7621,N_4224,N_4570);
or U7622 (N_7622,N_5366,N_5009);
nand U7623 (N_7623,N_4420,N_4604);
nand U7624 (N_7624,N_5085,N_4536);
nor U7625 (N_7625,N_5713,N_4976);
xor U7626 (N_7626,N_5265,N_5657);
and U7627 (N_7627,N_4328,N_5733);
and U7628 (N_7628,N_5606,N_5540);
or U7629 (N_7629,N_5122,N_4813);
nand U7630 (N_7630,N_5267,N_5906);
or U7631 (N_7631,N_5633,N_5995);
and U7632 (N_7632,N_5967,N_4926);
xor U7633 (N_7633,N_4536,N_4551);
or U7634 (N_7634,N_5265,N_4536);
nor U7635 (N_7635,N_4503,N_4900);
and U7636 (N_7636,N_5000,N_5736);
and U7637 (N_7637,N_4300,N_5748);
or U7638 (N_7638,N_5755,N_4857);
nor U7639 (N_7639,N_4018,N_4603);
nand U7640 (N_7640,N_4365,N_5287);
or U7641 (N_7641,N_5754,N_5995);
and U7642 (N_7642,N_5280,N_5078);
xnor U7643 (N_7643,N_4590,N_4889);
nand U7644 (N_7644,N_4278,N_5347);
nand U7645 (N_7645,N_5420,N_4652);
and U7646 (N_7646,N_5718,N_4377);
nor U7647 (N_7647,N_5274,N_4680);
nor U7648 (N_7648,N_5000,N_5567);
xor U7649 (N_7649,N_4175,N_5698);
or U7650 (N_7650,N_5811,N_5510);
and U7651 (N_7651,N_4491,N_5216);
xnor U7652 (N_7652,N_4309,N_4331);
or U7653 (N_7653,N_4580,N_4722);
or U7654 (N_7654,N_4275,N_5112);
and U7655 (N_7655,N_5176,N_4052);
and U7656 (N_7656,N_4411,N_4299);
nand U7657 (N_7657,N_5100,N_4220);
xor U7658 (N_7658,N_5343,N_4170);
nand U7659 (N_7659,N_5025,N_4669);
xnor U7660 (N_7660,N_4399,N_4002);
nor U7661 (N_7661,N_4915,N_5023);
nand U7662 (N_7662,N_5970,N_5340);
nor U7663 (N_7663,N_5225,N_5570);
nand U7664 (N_7664,N_4833,N_4187);
xnor U7665 (N_7665,N_5486,N_5098);
nand U7666 (N_7666,N_4178,N_4559);
and U7667 (N_7667,N_4540,N_5270);
and U7668 (N_7668,N_4636,N_4327);
nand U7669 (N_7669,N_5298,N_4922);
or U7670 (N_7670,N_5929,N_5139);
or U7671 (N_7671,N_4502,N_4253);
nor U7672 (N_7672,N_4430,N_5904);
and U7673 (N_7673,N_5166,N_5044);
xnor U7674 (N_7674,N_4620,N_4016);
and U7675 (N_7675,N_5581,N_5038);
nor U7676 (N_7676,N_5461,N_5538);
nor U7677 (N_7677,N_4304,N_4649);
and U7678 (N_7678,N_4545,N_5551);
and U7679 (N_7679,N_4425,N_4490);
nand U7680 (N_7680,N_5590,N_4306);
nand U7681 (N_7681,N_4970,N_4260);
and U7682 (N_7682,N_4248,N_5505);
and U7683 (N_7683,N_5034,N_4529);
or U7684 (N_7684,N_5177,N_4239);
xor U7685 (N_7685,N_4464,N_5117);
nand U7686 (N_7686,N_4238,N_5830);
or U7687 (N_7687,N_4468,N_4741);
and U7688 (N_7688,N_5249,N_5281);
or U7689 (N_7689,N_5331,N_4240);
and U7690 (N_7690,N_5391,N_5798);
nor U7691 (N_7691,N_4053,N_5054);
nor U7692 (N_7692,N_5043,N_4080);
or U7693 (N_7693,N_4523,N_5226);
nand U7694 (N_7694,N_5650,N_5285);
xor U7695 (N_7695,N_5325,N_5647);
and U7696 (N_7696,N_5203,N_5063);
nand U7697 (N_7697,N_5505,N_5067);
and U7698 (N_7698,N_4129,N_5979);
nor U7699 (N_7699,N_5958,N_5707);
or U7700 (N_7700,N_4387,N_4350);
nand U7701 (N_7701,N_4398,N_5040);
and U7702 (N_7702,N_5750,N_5711);
and U7703 (N_7703,N_4813,N_5743);
or U7704 (N_7704,N_4337,N_4076);
and U7705 (N_7705,N_4785,N_5226);
or U7706 (N_7706,N_4748,N_5347);
and U7707 (N_7707,N_5084,N_5134);
and U7708 (N_7708,N_5991,N_5635);
nor U7709 (N_7709,N_5792,N_5168);
nand U7710 (N_7710,N_4659,N_5249);
or U7711 (N_7711,N_5352,N_5409);
or U7712 (N_7712,N_5160,N_4051);
or U7713 (N_7713,N_4313,N_4951);
or U7714 (N_7714,N_4536,N_4394);
nand U7715 (N_7715,N_4780,N_5000);
nor U7716 (N_7716,N_5312,N_4567);
or U7717 (N_7717,N_4190,N_4309);
nand U7718 (N_7718,N_4101,N_4206);
nor U7719 (N_7719,N_5424,N_4511);
and U7720 (N_7720,N_5150,N_4545);
nor U7721 (N_7721,N_5887,N_5924);
nand U7722 (N_7722,N_4946,N_5807);
and U7723 (N_7723,N_4731,N_5752);
or U7724 (N_7724,N_5761,N_4235);
nand U7725 (N_7725,N_5452,N_5538);
and U7726 (N_7726,N_5870,N_4387);
or U7727 (N_7727,N_5608,N_5418);
nand U7728 (N_7728,N_5424,N_5606);
nand U7729 (N_7729,N_4663,N_4650);
and U7730 (N_7730,N_4308,N_4298);
nand U7731 (N_7731,N_5041,N_5914);
nand U7732 (N_7732,N_5551,N_4307);
nand U7733 (N_7733,N_5328,N_5033);
and U7734 (N_7734,N_4805,N_5161);
nor U7735 (N_7735,N_4931,N_5436);
nand U7736 (N_7736,N_5569,N_4123);
nand U7737 (N_7737,N_4833,N_5012);
nand U7738 (N_7738,N_4197,N_4333);
nor U7739 (N_7739,N_5654,N_4032);
nand U7740 (N_7740,N_4793,N_4603);
and U7741 (N_7741,N_4296,N_5994);
nand U7742 (N_7742,N_4722,N_5084);
nor U7743 (N_7743,N_4892,N_4316);
nand U7744 (N_7744,N_5552,N_5496);
xor U7745 (N_7745,N_5007,N_4143);
or U7746 (N_7746,N_5075,N_5783);
or U7747 (N_7747,N_4907,N_5466);
and U7748 (N_7748,N_5299,N_4687);
nor U7749 (N_7749,N_5675,N_5096);
nand U7750 (N_7750,N_5778,N_4450);
nand U7751 (N_7751,N_4120,N_5120);
nor U7752 (N_7752,N_4471,N_4738);
nor U7753 (N_7753,N_5790,N_4719);
nand U7754 (N_7754,N_4595,N_5609);
nand U7755 (N_7755,N_5862,N_5621);
nand U7756 (N_7756,N_4297,N_4811);
nor U7757 (N_7757,N_4902,N_4831);
nor U7758 (N_7758,N_4196,N_4374);
nand U7759 (N_7759,N_4857,N_5190);
nor U7760 (N_7760,N_5375,N_4998);
and U7761 (N_7761,N_4634,N_5927);
nor U7762 (N_7762,N_4467,N_5884);
nand U7763 (N_7763,N_5398,N_4510);
nand U7764 (N_7764,N_4385,N_5770);
xnor U7765 (N_7765,N_4041,N_4631);
and U7766 (N_7766,N_4833,N_5561);
and U7767 (N_7767,N_4435,N_5264);
nor U7768 (N_7768,N_5952,N_5395);
and U7769 (N_7769,N_4713,N_5163);
nand U7770 (N_7770,N_5097,N_5733);
nor U7771 (N_7771,N_5134,N_5055);
nor U7772 (N_7772,N_5724,N_5998);
nand U7773 (N_7773,N_4112,N_5525);
nor U7774 (N_7774,N_4990,N_5256);
and U7775 (N_7775,N_5341,N_5422);
nor U7776 (N_7776,N_5947,N_5398);
or U7777 (N_7777,N_5900,N_4624);
nand U7778 (N_7778,N_5739,N_4945);
nor U7779 (N_7779,N_5742,N_5275);
or U7780 (N_7780,N_4537,N_5248);
nand U7781 (N_7781,N_4680,N_4212);
xor U7782 (N_7782,N_5901,N_4501);
nand U7783 (N_7783,N_4998,N_5886);
or U7784 (N_7784,N_4974,N_5835);
and U7785 (N_7785,N_4231,N_4068);
and U7786 (N_7786,N_4511,N_4056);
and U7787 (N_7787,N_4180,N_5891);
nand U7788 (N_7788,N_4912,N_5227);
nor U7789 (N_7789,N_5577,N_4550);
xor U7790 (N_7790,N_4890,N_5584);
nand U7791 (N_7791,N_4768,N_4010);
or U7792 (N_7792,N_4875,N_5720);
nor U7793 (N_7793,N_5059,N_4034);
nor U7794 (N_7794,N_4102,N_4868);
nor U7795 (N_7795,N_5203,N_5410);
and U7796 (N_7796,N_5452,N_5355);
nand U7797 (N_7797,N_5193,N_4206);
nand U7798 (N_7798,N_5001,N_5909);
xnor U7799 (N_7799,N_5914,N_5621);
nand U7800 (N_7800,N_5641,N_4451);
nor U7801 (N_7801,N_4671,N_4092);
nor U7802 (N_7802,N_5581,N_5419);
or U7803 (N_7803,N_4453,N_4874);
nand U7804 (N_7804,N_4855,N_5665);
and U7805 (N_7805,N_5622,N_4572);
xnor U7806 (N_7806,N_4218,N_4964);
nand U7807 (N_7807,N_5131,N_4427);
nor U7808 (N_7808,N_4732,N_5666);
nor U7809 (N_7809,N_5772,N_5348);
nor U7810 (N_7810,N_4262,N_4501);
or U7811 (N_7811,N_5820,N_5569);
nand U7812 (N_7812,N_5883,N_4826);
or U7813 (N_7813,N_4907,N_4347);
xor U7814 (N_7814,N_5868,N_5354);
nor U7815 (N_7815,N_4601,N_5709);
nand U7816 (N_7816,N_5715,N_5750);
nor U7817 (N_7817,N_5650,N_5924);
and U7818 (N_7818,N_4655,N_5400);
nor U7819 (N_7819,N_4539,N_4829);
and U7820 (N_7820,N_4722,N_4317);
nor U7821 (N_7821,N_5927,N_4173);
nand U7822 (N_7822,N_5713,N_5872);
and U7823 (N_7823,N_4632,N_4729);
and U7824 (N_7824,N_4066,N_5454);
and U7825 (N_7825,N_5808,N_5674);
or U7826 (N_7826,N_5584,N_4736);
nor U7827 (N_7827,N_4549,N_5304);
or U7828 (N_7828,N_5286,N_5559);
xnor U7829 (N_7829,N_4205,N_4928);
and U7830 (N_7830,N_4939,N_4984);
nand U7831 (N_7831,N_5857,N_4227);
or U7832 (N_7832,N_4862,N_5406);
nor U7833 (N_7833,N_5669,N_5535);
nor U7834 (N_7834,N_4202,N_4267);
xor U7835 (N_7835,N_5372,N_4090);
xor U7836 (N_7836,N_5035,N_4257);
or U7837 (N_7837,N_4035,N_5773);
nor U7838 (N_7838,N_4804,N_4320);
and U7839 (N_7839,N_4240,N_4991);
or U7840 (N_7840,N_4781,N_5228);
or U7841 (N_7841,N_4287,N_5397);
nor U7842 (N_7842,N_4794,N_5843);
xor U7843 (N_7843,N_5427,N_4520);
nand U7844 (N_7844,N_5989,N_4398);
xor U7845 (N_7845,N_5109,N_5026);
and U7846 (N_7846,N_5065,N_5187);
or U7847 (N_7847,N_4996,N_5524);
nand U7848 (N_7848,N_5202,N_5571);
nor U7849 (N_7849,N_4278,N_5023);
and U7850 (N_7850,N_5899,N_5540);
nand U7851 (N_7851,N_4063,N_4396);
nor U7852 (N_7852,N_4775,N_5689);
or U7853 (N_7853,N_4498,N_4234);
nor U7854 (N_7854,N_4558,N_4533);
nand U7855 (N_7855,N_5509,N_5728);
nor U7856 (N_7856,N_5053,N_5755);
nor U7857 (N_7857,N_5232,N_4762);
and U7858 (N_7858,N_4780,N_4031);
xnor U7859 (N_7859,N_4418,N_4781);
or U7860 (N_7860,N_5436,N_4319);
and U7861 (N_7861,N_4986,N_5287);
and U7862 (N_7862,N_4600,N_5764);
xnor U7863 (N_7863,N_4520,N_4030);
and U7864 (N_7864,N_5391,N_4890);
or U7865 (N_7865,N_5965,N_5957);
nor U7866 (N_7866,N_5138,N_5510);
xor U7867 (N_7867,N_4890,N_5719);
nor U7868 (N_7868,N_4555,N_4547);
nand U7869 (N_7869,N_5579,N_4065);
or U7870 (N_7870,N_5877,N_5573);
or U7871 (N_7871,N_4801,N_5473);
and U7872 (N_7872,N_4985,N_5846);
or U7873 (N_7873,N_5379,N_5895);
or U7874 (N_7874,N_4061,N_4774);
nand U7875 (N_7875,N_5522,N_4274);
nand U7876 (N_7876,N_5778,N_4752);
or U7877 (N_7877,N_5807,N_5741);
or U7878 (N_7878,N_5970,N_5180);
nor U7879 (N_7879,N_4286,N_5667);
or U7880 (N_7880,N_5540,N_5570);
xnor U7881 (N_7881,N_5523,N_5439);
and U7882 (N_7882,N_5615,N_5736);
and U7883 (N_7883,N_5307,N_4560);
or U7884 (N_7884,N_5725,N_5429);
and U7885 (N_7885,N_4032,N_5517);
or U7886 (N_7886,N_4814,N_5950);
and U7887 (N_7887,N_4181,N_4161);
nor U7888 (N_7888,N_5343,N_4424);
nand U7889 (N_7889,N_5128,N_5336);
nand U7890 (N_7890,N_5296,N_4599);
nor U7891 (N_7891,N_4177,N_4083);
and U7892 (N_7892,N_5645,N_4424);
nand U7893 (N_7893,N_4026,N_4703);
xor U7894 (N_7894,N_5486,N_4841);
and U7895 (N_7895,N_5477,N_5217);
nand U7896 (N_7896,N_4330,N_5534);
and U7897 (N_7897,N_4458,N_4756);
xor U7898 (N_7898,N_4308,N_5518);
nand U7899 (N_7899,N_4980,N_5798);
and U7900 (N_7900,N_5213,N_5349);
and U7901 (N_7901,N_4021,N_5307);
nor U7902 (N_7902,N_5990,N_5882);
nor U7903 (N_7903,N_5860,N_5645);
xor U7904 (N_7904,N_4498,N_4451);
nand U7905 (N_7905,N_4134,N_5935);
nand U7906 (N_7906,N_4689,N_4322);
and U7907 (N_7907,N_5762,N_5951);
or U7908 (N_7908,N_4989,N_5968);
nor U7909 (N_7909,N_5336,N_5287);
xnor U7910 (N_7910,N_4685,N_5123);
nor U7911 (N_7911,N_5794,N_4921);
and U7912 (N_7912,N_4754,N_5705);
or U7913 (N_7913,N_4745,N_5285);
and U7914 (N_7914,N_4621,N_4409);
or U7915 (N_7915,N_5115,N_4141);
and U7916 (N_7916,N_5317,N_4738);
or U7917 (N_7917,N_4200,N_5725);
and U7918 (N_7918,N_4294,N_5771);
nand U7919 (N_7919,N_5027,N_4699);
nor U7920 (N_7920,N_4759,N_4409);
nor U7921 (N_7921,N_4161,N_5735);
nor U7922 (N_7922,N_5011,N_4922);
nand U7923 (N_7923,N_5514,N_4609);
or U7924 (N_7924,N_5903,N_4021);
xor U7925 (N_7925,N_5756,N_5654);
or U7926 (N_7926,N_5509,N_5098);
nand U7927 (N_7927,N_4800,N_4165);
nand U7928 (N_7928,N_5270,N_4520);
or U7929 (N_7929,N_5574,N_5735);
or U7930 (N_7930,N_5359,N_4672);
and U7931 (N_7931,N_5708,N_5604);
and U7932 (N_7932,N_4548,N_5350);
or U7933 (N_7933,N_5460,N_5897);
or U7934 (N_7934,N_5216,N_4367);
and U7935 (N_7935,N_4009,N_5076);
nand U7936 (N_7936,N_5238,N_4050);
nor U7937 (N_7937,N_5949,N_4108);
nand U7938 (N_7938,N_4278,N_5796);
nor U7939 (N_7939,N_5312,N_4023);
xor U7940 (N_7940,N_5154,N_5805);
nor U7941 (N_7941,N_4588,N_4032);
nand U7942 (N_7942,N_4534,N_4759);
nand U7943 (N_7943,N_4798,N_5644);
nor U7944 (N_7944,N_5144,N_4252);
nand U7945 (N_7945,N_5236,N_4816);
or U7946 (N_7946,N_5459,N_4456);
nand U7947 (N_7947,N_5664,N_4695);
and U7948 (N_7948,N_5672,N_5645);
nor U7949 (N_7949,N_5318,N_5447);
xor U7950 (N_7950,N_5132,N_4158);
or U7951 (N_7951,N_5459,N_5969);
and U7952 (N_7952,N_5711,N_5200);
and U7953 (N_7953,N_4995,N_5090);
nor U7954 (N_7954,N_5498,N_4904);
nand U7955 (N_7955,N_5194,N_5464);
nand U7956 (N_7956,N_4993,N_4188);
or U7957 (N_7957,N_4431,N_5824);
nand U7958 (N_7958,N_4932,N_5288);
xnor U7959 (N_7959,N_5846,N_4028);
or U7960 (N_7960,N_4669,N_4592);
nand U7961 (N_7961,N_5778,N_4072);
nor U7962 (N_7962,N_4464,N_5066);
nand U7963 (N_7963,N_5111,N_5650);
or U7964 (N_7964,N_5343,N_5185);
or U7965 (N_7965,N_4850,N_5248);
nor U7966 (N_7966,N_4687,N_5793);
nor U7967 (N_7967,N_5138,N_4733);
nand U7968 (N_7968,N_5906,N_5472);
xnor U7969 (N_7969,N_4618,N_4741);
xor U7970 (N_7970,N_4441,N_5245);
and U7971 (N_7971,N_5164,N_5900);
nor U7972 (N_7972,N_4640,N_5419);
xnor U7973 (N_7973,N_5506,N_5444);
xnor U7974 (N_7974,N_4165,N_4616);
and U7975 (N_7975,N_5849,N_5732);
xor U7976 (N_7976,N_5572,N_4078);
nor U7977 (N_7977,N_4362,N_5581);
and U7978 (N_7978,N_4952,N_5832);
nor U7979 (N_7979,N_4959,N_4821);
nor U7980 (N_7980,N_5129,N_5480);
and U7981 (N_7981,N_5194,N_4081);
and U7982 (N_7982,N_4718,N_5234);
or U7983 (N_7983,N_5643,N_5004);
or U7984 (N_7984,N_5400,N_4751);
or U7985 (N_7985,N_5748,N_5278);
or U7986 (N_7986,N_5507,N_5157);
nand U7987 (N_7987,N_4517,N_5658);
or U7988 (N_7988,N_4373,N_4142);
nand U7989 (N_7989,N_5947,N_5003);
nand U7990 (N_7990,N_5989,N_4607);
and U7991 (N_7991,N_4829,N_4329);
nor U7992 (N_7992,N_5573,N_4390);
nor U7993 (N_7993,N_5607,N_5485);
nand U7994 (N_7994,N_4429,N_5476);
and U7995 (N_7995,N_5838,N_4108);
xnor U7996 (N_7996,N_5389,N_5561);
xor U7997 (N_7997,N_5649,N_4993);
nand U7998 (N_7998,N_5440,N_5732);
nor U7999 (N_7999,N_5235,N_5585);
nand U8000 (N_8000,N_6270,N_6854);
nor U8001 (N_8001,N_7387,N_7162);
xnor U8002 (N_8002,N_6560,N_7248);
and U8003 (N_8003,N_6311,N_6885);
nand U8004 (N_8004,N_6895,N_7568);
nor U8005 (N_8005,N_6918,N_7433);
nand U8006 (N_8006,N_6035,N_6622);
nand U8007 (N_8007,N_6745,N_6778);
nand U8008 (N_8008,N_6104,N_6971);
nand U8009 (N_8009,N_6478,N_7855);
nand U8010 (N_8010,N_6612,N_7756);
and U8011 (N_8011,N_6604,N_6632);
nor U8012 (N_8012,N_7658,N_7915);
xor U8013 (N_8013,N_6715,N_6366);
or U8014 (N_8014,N_7993,N_6923);
and U8015 (N_8015,N_6459,N_7205);
or U8016 (N_8016,N_7633,N_6829);
xnor U8017 (N_8017,N_7075,N_7795);
and U8018 (N_8018,N_6121,N_6406);
or U8019 (N_8019,N_7005,N_6039);
or U8020 (N_8020,N_7213,N_7317);
xor U8021 (N_8021,N_7586,N_7345);
nand U8022 (N_8022,N_6405,N_6484);
and U8023 (N_8023,N_6103,N_6101);
xor U8024 (N_8024,N_7422,N_6008);
and U8025 (N_8025,N_7891,N_7599);
xnor U8026 (N_8026,N_7881,N_7833);
or U8027 (N_8027,N_6142,N_7070);
and U8028 (N_8028,N_6936,N_6900);
nor U8029 (N_8029,N_7437,N_6011);
and U8030 (N_8030,N_7718,N_7973);
or U8031 (N_8031,N_7147,N_6609);
or U8032 (N_8032,N_7747,N_7931);
nor U8033 (N_8033,N_6434,N_7808);
nor U8034 (N_8034,N_7954,N_7304);
nor U8035 (N_8035,N_7136,N_7564);
and U8036 (N_8036,N_7990,N_7853);
and U8037 (N_8037,N_6864,N_6117);
or U8038 (N_8038,N_7521,N_6001);
xor U8039 (N_8039,N_7549,N_6815);
and U8040 (N_8040,N_6664,N_6762);
and U8041 (N_8041,N_6042,N_7047);
nand U8042 (N_8042,N_7082,N_7169);
and U8043 (N_8043,N_7883,N_6631);
nor U8044 (N_8044,N_6274,N_7241);
and U8045 (N_8045,N_6056,N_7464);
xor U8046 (N_8046,N_6666,N_6531);
nand U8047 (N_8047,N_6913,N_6265);
and U8048 (N_8048,N_7286,N_6827);
nor U8049 (N_8049,N_7856,N_7036);
xnor U8050 (N_8050,N_6146,N_6383);
and U8051 (N_8051,N_6528,N_6037);
or U8052 (N_8052,N_6369,N_6650);
nor U8053 (N_8053,N_6718,N_7815);
nor U8054 (N_8054,N_7144,N_6706);
and U8055 (N_8055,N_6315,N_6929);
or U8056 (N_8056,N_6048,N_7593);
nand U8057 (N_8057,N_6947,N_6985);
nand U8058 (N_8058,N_6523,N_7771);
and U8059 (N_8059,N_7763,N_6471);
or U8060 (N_8060,N_7654,N_6520);
nand U8061 (N_8061,N_6770,N_7431);
xor U8062 (N_8062,N_6637,N_7445);
nand U8063 (N_8063,N_6244,N_7092);
nand U8064 (N_8064,N_7327,N_6940);
or U8065 (N_8065,N_7976,N_6671);
nor U8066 (N_8066,N_6570,N_6225);
nor U8067 (N_8067,N_7116,N_7494);
nor U8068 (N_8068,N_6897,N_7006);
or U8069 (N_8069,N_7963,N_6978);
nor U8070 (N_8070,N_7350,N_6557);
or U8071 (N_8071,N_6633,N_7846);
or U8072 (N_8072,N_6380,N_6413);
nor U8073 (N_8073,N_6242,N_7440);
and U8074 (N_8074,N_6803,N_6026);
nand U8075 (N_8075,N_7887,N_6443);
and U8076 (N_8076,N_6521,N_7409);
and U8077 (N_8077,N_7164,N_7752);
and U8078 (N_8078,N_6680,N_7251);
nor U8079 (N_8079,N_7042,N_7481);
nor U8080 (N_8080,N_7310,N_6297);
nor U8081 (N_8081,N_7779,N_7479);
xor U8082 (N_8082,N_6626,N_6399);
xnor U8083 (N_8083,N_6343,N_6354);
nor U8084 (N_8084,N_6140,N_6651);
nor U8085 (N_8085,N_7877,N_7238);
nor U8086 (N_8086,N_6994,N_6364);
and U8087 (N_8087,N_7091,N_6424);
or U8088 (N_8088,N_7154,N_6182);
nor U8089 (N_8089,N_6348,N_6704);
and U8090 (N_8090,N_7017,N_6569);
nor U8091 (N_8091,N_7842,N_6722);
or U8092 (N_8092,N_7418,N_7056);
nor U8093 (N_8093,N_6700,N_6282);
and U8094 (N_8094,N_6120,N_6780);
nor U8095 (N_8095,N_6332,N_6096);
and U8096 (N_8096,N_6307,N_6188);
and U8097 (N_8097,N_7123,N_6813);
or U8098 (N_8098,N_7442,N_6937);
nor U8099 (N_8099,N_6107,N_7622);
and U8100 (N_8100,N_6269,N_6152);
or U8101 (N_8101,N_6759,N_7268);
xor U8102 (N_8102,N_7219,N_7114);
xor U8103 (N_8103,N_6731,N_7383);
or U8104 (N_8104,N_6997,N_6428);
nand U8105 (N_8105,N_6387,N_7516);
and U8106 (N_8106,N_7328,N_7928);
or U8107 (N_8107,N_7605,N_7053);
nand U8108 (N_8108,N_7259,N_7411);
nand U8109 (N_8109,N_7577,N_7696);
nand U8110 (N_8110,N_6655,N_6113);
nor U8111 (N_8111,N_6581,N_6344);
and U8112 (N_8112,N_7027,N_6742);
xor U8113 (N_8113,N_7246,N_7486);
and U8114 (N_8114,N_6059,N_6596);
nor U8115 (N_8115,N_6931,N_7830);
or U8116 (N_8116,N_6993,N_6685);
and U8117 (N_8117,N_6426,N_7712);
or U8118 (N_8118,N_6796,N_7283);
nor U8119 (N_8119,N_7868,N_6533);
nor U8120 (N_8120,N_6972,N_6239);
or U8121 (N_8121,N_7065,N_6732);
or U8122 (N_8122,N_6494,N_7412);
xnor U8123 (N_8123,N_7584,N_6483);
or U8124 (N_8124,N_6810,N_6564);
nor U8125 (N_8125,N_6053,N_7733);
nand U8126 (N_8126,N_7639,N_7828);
nor U8127 (N_8127,N_7836,N_7299);
and U8128 (N_8128,N_7721,N_6719);
xor U8129 (N_8129,N_6360,N_7880);
nand U8130 (N_8130,N_6544,N_7446);
nor U8131 (N_8131,N_6353,N_7052);
nand U8132 (N_8132,N_7555,N_7532);
and U8133 (N_8133,N_6213,N_6433);
or U8134 (N_8134,N_6295,N_6460);
and U8135 (N_8135,N_6587,N_7753);
and U8136 (N_8136,N_6248,N_7168);
nor U8137 (N_8137,N_7189,N_7166);
or U8138 (N_8138,N_6419,N_6743);
or U8139 (N_8139,N_7140,N_7432);
nand U8140 (N_8140,N_7298,N_7414);
xnor U8141 (N_8141,N_7610,N_7757);
nand U8142 (N_8142,N_7982,N_7392);
xor U8143 (N_8143,N_6966,N_6708);
or U8144 (N_8144,N_6259,N_6139);
or U8145 (N_8145,N_7699,N_7273);
xor U8146 (N_8146,N_7352,N_7600);
nand U8147 (N_8147,N_7044,N_7804);
and U8148 (N_8148,N_6748,N_7252);
nor U8149 (N_8149,N_7221,N_7934);
and U8150 (N_8150,N_6954,N_6168);
xnor U8151 (N_8151,N_6691,N_6746);
nand U8152 (N_8152,N_6470,N_7751);
or U8153 (N_8153,N_6862,N_6293);
or U8154 (N_8154,N_7242,N_6497);
or U8155 (N_8155,N_7230,N_6205);
and U8156 (N_8156,N_7155,N_6414);
and U8157 (N_8157,N_6150,N_7417);
and U8158 (N_8158,N_7914,N_6490);
nor U8159 (N_8159,N_7708,N_7714);
or U8160 (N_8160,N_6198,N_7793);
nor U8161 (N_8161,N_7704,N_7745);
nor U8162 (N_8162,N_6616,N_7032);
and U8163 (N_8163,N_7014,N_7308);
nand U8164 (N_8164,N_6502,N_7572);
nor U8165 (N_8165,N_6454,N_6382);
nand U8166 (N_8166,N_6763,N_7986);
nand U8167 (N_8167,N_7774,N_7787);
nor U8168 (N_8168,N_7382,N_7944);
and U8169 (N_8169,N_7790,N_6889);
nand U8170 (N_8170,N_7262,N_7300);
nor U8171 (N_8171,N_7018,N_6850);
and U8172 (N_8172,N_7472,N_6550);
and U8173 (N_8173,N_6701,N_6488);
or U8174 (N_8174,N_7093,N_6105);
nand U8175 (N_8175,N_6373,N_7102);
or U8176 (N_8176,N_6933,N_7571);
or U8177 (N_8177,N_6076,N_6289);
nand U8178 (N_8178,N_6589,N_6014);
nand U8179 (N_8179,N_6572,N_6579);
nor U8180 (N_8180,N_6617,N_7989);
nor U8181 (N_8181,N_7946,N_7827);
and U8182 (N_8182,N_7675,N_7956);
nor U8183 (N_8183,N_7362,N_7457);
nor U8184 (N_8184,N_6368,N_7240);
and U8185 (N_8185,N_6099,N_6316);
nand U8186 (N_8186,N_7870,N_6851);
xor U8187 (N_8187,N_7058,N_7773);
or U8188 (N_8188,N_7509,N_7165);
and U8189 (N_8189,N_7498,N_6092);
nand U8190 (N_8190,N_6679,N_6951);
nor U8191 (N_8191,N_6582,N_7949);
nand U8192 (N_8192,N_6306,N_7907);
and U8193 (N_8193,N_7800,N_6545);
nand U8194 (N_8194,N_7538,N_7111);
or U8195 (N_8195,N_7474,N_6436);
nor U8196 (N_8196,N_7770,N_6216);
nand U8197 (N_8197,N_6075,N_7672);
nand U8198 (N_8198,N_7104,N_7133);
or U8199 (N_8199,N_6578,N_6125);
nor U8200 (N_8200,N_6093,N_7132);
nand U8201 (N_8201,N_6486,N_7844);
or U8202 (N_8202,N_7979,N_7234);
or U8203 (N_8203,N_7084,N_6525);
nand U8204 (N_8204,N_7970,N_6791);
and U8205 (N_8205,N_6530,N_6262);
nor U8206 (N_8206,N_7193,N_7702);
xor U8207 (N_8207,N_6510,N_6822);
and U8208 (N_8208,N_6635,N_7715);
and U8209 (N_8209,N_6884,N_6263);
or U8210 (N_8210,N_6308,N_7443);
nand U8211 (N_8211,N_7608,N_6398);
nand U8212 (N_8212,N_7135,N_7031);
or U8213 (N_8213,N_7066,N_6600);
xor U8214 (N_8214,N_7527,N_6890);
nand U8215 (N_8215,N_7468,N_7279);
nand U8216 (N_8216,N_6017,N_7182);
nand U8217 (N_8217,N_6737,N_7918);
and U8218 (N_8218,N_6773,N_6444);
nand U8219 (N_8219,N_7628,N_7746);
nor U8220 (N_8220,N_6894,N_7235);
nand U8221 (N_8221,N_7875,N_6605);
xor U8222 (N_8222,N_6736,N_6031);
xnor U8223 (N_8223,N_6590,N_6181);
and U8224 (N_8224,N_7947,N_6839);
nor U8225 (N_8225,N_6466,N_6721);
and U8226 (N_8226,N_6267,N_7062);
and U8227 (N_8227,N_6148,N_7627);
or U8228 (N_8228,N_6568,N_7174);
nor U8229 (N_8229,N_7079,N_7203);
nor U8230 (N_8230,N_7818,N_7434);
xnor U8231 (N_8231,N_7488,N_7583);
xor U8232 (N_8232,N_7528,N_7260);
or U8233 (N_8233,N_7685,N_6089);
nor U8234 (N_8234,N_6684,N_7054);
nor U8235 (N_8235,N_7687,N_7517);
and U8236 (N_8236,N_7531,N_6760);
xor U8237 (N_8237,N_7372,N_6656);
and U8238 (N_8238,N_7603,N_6534);
nor U8239 (N_8239,N_6944,N_7161);
or U8240 (N_8240,N_7236,N_6955);
nand U8241 (N_8241,N_7636,N_7886);
nor U8242 (N_8242,N_7288,N_7638);
and U8243 (N_8243,N_7634,N_6509);
nand U8244 (N_8244,N_6823,N_7832);
nand U8245 (N_8245,N_6811,N_6640);
and U8246 (N_8246,N_7739,N_7644);
nand U8247 (N_8247,N_6789,N_6403);
nand U8248 (N_8248,N_6597,N_6326);
or U8249 (N_8249,N_7280,N_7899);
nor U8250 (N_8250,N_7237,N_7146);
nor U8251 (N_8251,N_6379,N_6143);
nor U8252 (N_8252,N_7816,N_6032);
nor U8253 (N_8253,N_7512,N_7063);
or U8254 (N_8254,N_7840,N_6887);
nand U8255 (N_8255,N_6625,N_6879);
and U8256 (N_8256,N_7177,N_7332);
and U8257 (N_8257,N_7037,N_6601);
nand U8258 (N_8258,N_7788,N_6527);
nor U8259 (N_8259,N_6677,N_6892);
nor U8260 (N_8260,N_6709,N_7218);
and U8261 (N_8261,N_7676,N_6402);
nor U8262 (N_8262,N_7256,N_7223);
nand U8263 (N_8263,N_7912,N_7305);
nor U8264 (N_8264,N_6234,N_6291);
nor U8265 (N_8265,N_6891,N_7502);
and U8266 (N_8266,N_6040,N_6197);
or U8267 (N_8267,N_7285,N_7271);
nand U8268 (N_8268,N_6898,N_7157);
nor U8269 (N_8269,N_7284,N_7178);
nor U8270 (N_8270,N_6855,N_7101);
and U8271 (N_8271,N_7023,N_6986);
or U8272 (N_8272,N_6464,N_6300);
and U8273 (N_8273,N_7019,N_6324);
nor U8274 (N_8274,N_7348,N_6939);
xor U8275 (N_8275,N_6847,N_6602);
and U8276 (N_8276,N_7728,N_6452);
and U8277 (N_8277,N_7179,N_7334);
or U8278 (N_8278,N_7476,N_7785);
nand U8279 (N_8279,N_6273,N_6689);
nor U8280 (N_8280,N_7072,N_6196);
or U8281 (N_8281,N_6835,N_6946);
and U8282 (N_8282,N_7959,N_7071);
or U8283 (N_8283,N_7962,N_7688);
nand U8284 (N_8284,N_6930,N_6208);
xnor U8285 (N_8285,N_6726,N_6271);
or U8286 (N_8286,N_7192,N_7496);
nor U8287 (N_8287,N_7185,N_7001);
and U8288 (N_8288,N_6134,N_6781);
nand U8289 (N_8289,N_7439,N_6904);
nand U8290 (N_8290,N_6586,N_6318);
nand U8291 (N_8291,N_7247,N_6171);
nor U8292 (N_8292,N_6613,N_6438);
nand U8293 (N_8293,N_6462,N_6286);
xor U8294 (N_8294,N_6337,N_6673);
xor U8295 (N_8295,N_6974,N_7690);
and U8296 (N_8296,N_6162,N_6174);
nor U8297 (N_8297,N_7402,N_6005);
or U8298 (N_8298,N_7731,N_7449);
nand U8299 (N_8299,N_7210,N_7831);
nand U8300 (N_8300,N_7519,N_6756);
or U8301 (N_8301,N_6606,N_7086);
nor U8302 (N_8302,N_6979,N_6764);
nor U8303 (N_8303,N_7789,N_7493);
and U8304 (N_8304,N_6166,N_7408);
xnor U8305 (N_8305,N_6953,N_7380);
and U8306 (N_8306,N_6410,N_7729);
or U8307 (N_8307,N_6358,N_7999);
nand U8308 (N_8308,N_6575,N_6943);
nand U8309 (N_8309,N_7024,N_7768);
nand U8310 (N_8310,N_7222,N_6404);
nor U8311 (N_8311,N_7239,N_6629);
or U8312 (N_8312,N_7119,N_7138);
nor U8313 (N_8313,N_6830,N_7370);
nor U8314 (N_8314,N_7822,N_7755);
or U8315 (N_8315,N_7204,N_7319);
nor U8316 (N_8316,N_7792,N_7543);
and U8317 (N_8317,N_6312,N_7821);
and U8318 (N_8318,N_6435,N_6838);
and U8319 (N_8319,N_6508,N_6309);
and U8320 (N_8320,N_6591,N_7043);
and U8321 (N_8321,N_6775,N_7720);
or U8322 (N_8322,N_6202,N_7615);
or U8323 (N_8323,N_6285,N_6340);
nand U8324 (N_8324,N_7171,N_7341);
or U8325 (N_8325,N_7264,N_6055);
or U8326 (N_8326,N_6962,N_7371);
and U8327 (N_8327,N_6257,N_7000);
nor U8328 (N_8328,N_7373,N_6804);
nand U8329 (N_8329,N_7368,N_7865);
or U8330 (N_8330,N_7682,N_6919);
and U8331 (N_8331,N_7553,N_6421);
xnor U8332 (N_8332,N_7150,N_6821);
nand U8333 (N_8333,N_6389,N_7401);
xor U8334 (N_8334,N_6160,N_6193);
nand U8335 (N_8335,N_6959,N_7513);
nor U8336 (N_8336,N_6214,N_7261);
xnor U8337 (N_8337,N_7888,N_7911);
nor U8338 (N_8338,N_7301,N_7767);
and U8339 (N_8339,N_6697,N_7094);
nand U8340 (N_8340,N_7389,N_7130);
nor U8341 (N_8341,N_6194,N_7647);
and U8342 (N_8342,N_6319,N_7009);
nand U8343 (N_8343,N_6958,N_6730);
nor U8344 (N_8344,N_6047,N_6173);
and U8345 (N_8345,N_6294,N_7563);
nor U8346 (N_8346,N_7670,N_7625);
nand U8347 (N_8347,N_6290,N_6422);
nand U8348 (N_8348,N_6548,N_7399);
nor U8349 (N_8349,N_7561,N_6571);
or U8350 (N_8350,N_7632,N_6694);
nor U8351 (N_8351,N_6411,N_7245);
nor U8352 (N_8352,N_6739,N_6950);
nor U8353 (N_8353,N_7450,N_6006);
or U8354 (N_8354,N_6952,N_6541);
nand U8355 (N_8355,N_7738,N_7620);
nor U8356 (N_8356,N_6472,N_6754);
and U8357 (N_8357,N_7742,N_7274);
or U8358 (N_8358,N_7852,N_6425);
or U8359 (N_8359,N_6317,N_6546);
nand U8360 (N_8360,N_7611,N_7397);
nor U8361 (N_8361,N_6672,N_7758);
and U8362 (N_8362,N_7678,N_7289);
and U8363 (N_8363,N_7621,N_7405);
nor U8364 (N_8364,N_7961,N_7197);
nand U8365 (N_8365,N_7339,N_7810);
and U8366 (N_8366,N_7320,N_6755);
or U8367 (N_8367,N_6836,N_7691);
nand U8368 (N_8368,N_6250,N_6068);
xor U8369 (N_8369,N_7736,N_7909);
and U8370 (N_8370,N_6322,N_6566);
or U8371 (N_8371,N_6705,N_7172);
nor U8372 (N_8372,N_7484,N_7085);
nand U8373 (N_8373,N_7734,N_6751);
or U8374 (N_8374,N_7303,N_6185);
and U8375 (N_8375,N_7506,N_7186);
nor U8376 (N_8376,N_6787,N_7713);
and U8377 (N_8377,N_6473,N_6223);
or U8378 (N_8378,N_6206,N_6608);
and U8379 (N_8379,N_6499,N_7074);
or U8380 (N_8380,N_6574,N_6676);
and U8381 (N_8381,N_6072,N_6416);
nand U8382 (N_8382,N_6503,N_7048);
and U8383 (N_8383,N_6716,N_6457);
and U8384 (N_8384,N_6859,N_7932);
or U8385 (N_8385,N_7866,N_7551);
or U8386 (N_8386,N_6681,N_7904);
nor U8387 (N_8387,N_7663,N_7988);
or U8388 (N_8388,N_6837,N_7525);
and U8389 (N_8389,N_6915,N_7287);
and U8390 (N_8390,N_6938,N_6386);
nor U8391 (N_8391,N_6302,N_7478);
xnor U8392 (N_8392,N_6853,N_6828);
and U8393 (N_8393,N_6507,N_7709);
nor U8394 (N_8394,N_6108,N_7906);
nand U8395 (N_8395,N_7175,N_6178);
and U8396 (N_8396,N_6310,N_7134);
xor U8397 (N_8397,N_7152,N_7689);
and U8398 (N_8398,N_7338,N_7022);
nand U8399 (N_8399,N_7180,N_7522);
nand U8400 (N_8400,N_7083,N_7969);
and U8401 (N_8401,N_6935,N_7460);
and U8402 (N_8402,N_6711,N_7129);
nand U8403 (N_8403,N_7325,N_7253);
nor U8404 (N_8404,N_6809,N_7249);
nor U8405 (N_8405,N_7657,N_6987);
or U8406 (N_8406,N_6374,N_7985);
and U8407 (N_8407,N_6982,N_6747);
nand U8408 (N_8408,N_7859,N_7200);
or U8409 (N_8409,N_7606,N_6272);
or U8410 (N_8410,N_7537,N_6529);
or U8411 (N_8411,N_6603,N_7597);
and U8412 (N_8412,N_7604,N_6649);
xnor U8413 (N_8413,N_7356,N_6896);
and U8414 (N_8414,N_7013,N_7873);
or U8415 (N_8415,N_6834,N_6080);
or U8416 (N_8416,N_7126,N_7344);
and U8417 (N_8417,N_6800,N_7475);
or U8418 (N_8418,N_7269,N_6329);
and U8419 (N_8419,N_6999,N_7290);
nand U8420 (N_8420,N_7601,N_7347);
xnor U8421 (N_8421,N_6449,N_6130);
or U8422 (N_8422,N_6903,N_6767);
xnor U8423 (N_8423,N_6236,N_7375);
nor U8424 (N_8424,N_6448,N_7557);
nand U8425 (N_8425,N_7293,N_7049);
and U8426 (N_8426,N_7737,N_6235);
nor U8427 (N_8427,N_6067,N_7849);
nor U8428 (N_8428,N_6255,N_7575);
or U8429 (N_8429,N_6774,N_6824);
or U8430 (N_8430,N_6034,N_7735);
and U8431 (N_8431,N_7666,N_6292);
and U8432 (N_8432,N_6361,N_7576);
or U8433 (N_8433,N_7232,N_7231);
nor U8434 (N_8434,N_6973,N_7754);
xnor U8435 (N_8435,N_6907,N_6367);
nand U8436 (N_8436,N_6945,N_7125);
nor U8437 (N_8437,N_7003,N_6514);
or U8438 (N_8438,N_6585,N_6519);
or U8439 (N_8439,N_6376,N_6356);
nand U8440 (N_8440,N_6210,N_6749);
or U8441 (N_8441,N_6074,N_7515);
nor U8442 (N_8442,N_6082,N_7744);
nor U8443 (N_8443,N_7750,N_6819);
nand U8444 (N_8444,N_7614,N_6647);
or U8445 (N_8445,N_6222,N_7794);
nand U8446 (N_8446,N_6325,N_7225);
nor U8447 (N_8447,N_7447,N_6917);
and U8448 (N_8448,N_7088,N_6816);
xor U8449 (N_8449,N_7170,N_6049);
and U8450 (N_8450,N_7984,N_7069);
and U8451 (N_8451,N_7163,N_6840);
or U8452 (N_8452,N_7797,N_7010);
nor U8453 (N_8453,N_7216,N_6515);
nand U8454 (N_8454,N_7080,N_7889);
and U8455 (N_8455,N_6842,N_6893);
nand U8456 (N_8456,N_6752,N_6639);
nand U8457 (N_8457,N_7087,N_6558);
xnor U8458 (N_8458,N_6431,N_6069);
nand U8459 (N_8459,N_6183,N_7465);
or U8460 (N_8460,N_6036,N_6381);
xnor U8461 (N_8461,N_6518,N_7034);
nand U8462 (N_8462,N_7103,N_6702);
nor U8463 (N_8463,N_6619,N_6857);
or U8464 (N_8464,N_7206,N_6692);
or U8465 (N_8465,N_7364,N_6264);
xnor U8466 (N_8466,N_7643,N_7960);
nand U8467 (N_8467,N_7648,N_7395);
or U8468 (N_8468,N_7366,N_6203);
nor U8469 (N_8469,N_6061,N_6351);
nor U8470 (N_8470,N_6963,N_6170);
and U8471 (N_8471,N_6693,N_7558);
or U8472 (N_8472,N_7410,N_7851);
xnor U8473 (N_8473,N_6427,N_6253);
or U8474 (N_8474,N_7631,N_7127);
or U8475 (N_8475,N_7867,N_6167);
xnor U8476 (N_8476,N_6733,N_6323);
and U8477 (N_8477,N_6977,N_7196);
and U8478 (N_8478,N_7772,N_7587);
nand U8479 (N_8479,N_7882,N_7424);
and U8480 (N_8480,N_7967,N_6618);
nor U8481 (N_8481,N_7722,N_6338);
or U8482 (N_8482,N_7578,N_6741);
xor U8483 (N_8483,N_7214,N_7095);
nor U8484 (N_8484,N_7927,N_6397);
xor U8485 (N_8485,N_7524,N_7765);
xor U8486 (N_8486,N_6504,N_7428);
and U8487 (N_8487,N_7766,N_7671);
nor U8488 (N_8488,N_6018,N_7384);
or U8489 (N_8489,N_7548,N_6846);
and U8490 (N_8490,N_7326,N_6138);
nor U8491 (N_8491,N_6339,N_6636);
or U8492 (N_8492,N_7573,N_7761);
or U8493 (N_8493,N_7910,N_7707);
and U8494 (N_8494,N_7938,N_6990);
or U8495 (N_8495,N_7674,N_7589);
or U8496 (N_8496,N_6407,N_6690);
and U8497 (N_8497,N_6260,N_7340);
nor U8498 (N_8498,N_6882,N_6016);
or U8499 (N_8499,N_7514,N_7115);
nand U8500 (N_8500,N_6653,N_6345);
nor U8501 (N_8501,N_7937,N_6880);
and U8502 (N_8502,N_6420,N_7198);
nor U8503 (N_8503,N_7646,N_6535);
nor U8504 (N_8504,N_7933,N_6698);
and U8505 (N_8505,N_6129,N_6565);
or U8506 (N_8506,N_6965,N_7462);
xor U8507 (N_8507,N_7958,N_7511);
and U8508 (N_8508,N_7660,N_6371);
and U8509 (N_8509,N_6975,N_6740);
xor U8510 (N_8510,N_7324,N_6686);
and U8511 (N_8511,N_6275,N_7624);
nor U8512 (N_8512,N_7441,N_7505);
and U8513 (N_8513,N_6221,N_7567);
nand U8514 (N_8514,N_7361,N_6628);
or U8515 (N_8515,N_6451,N_6794);
nor U8516 (N_8516,N_6243,N_6921);
or U8517 (N_8517,N_6594,N_7267);
and U8518 (N_8518,N_7233,N_6218);
nand U8519 (N_8519,N_6097,N_7004);
nor U8520 (N_8520,N_7664,N_7980);
and U8521 (N_8521,N_7276,N_6577);
or U8522 (N_8522,N_6245,N_6865);
nor U8523 (N_8523,N_6644,N_7917);
nand U8524 (N_8524,N_6131,N_6869);
or U8525 (N_8525,N_6482,N_6735);
nand U8526 (N_8526,N_7151,N_6720);
nor U8527 (N_8527,N_6765,N_7526);
xor U8528 (N_8528,N_7534,N_6330);
nand U8529 (N_8529,N_7322,N_7697);
nand U8530 (N_8530,N_6401,N_7379);
nor U8531 (N_8531,N_7991,N_7459);
and U8532 (N_8532,N_7435,N_6512);
xor U8533 (N_8533,N_6948,N_6696);
xor U8534 (N_8534,N_7748,N_7902);
or U8535 (N_8535,N_7570,N_6229);
nand U8536 (N_8536,N_6538,N_7542);
xnor U8537 (N_8537,N_7108,N_6077);
or U8538 (N_8538,N_6333,N_6230);
nor U8539 (N_8539,N_7330,N_6788);
nand U8540 (N_8540,N_7596,N_6710);
xnor U8541 (N_8541,N_7266,N_7706);
nor U8542 (N_8542,N_7510,N_6874);
nand U8543 (N_8543,N_6807,N_6848);
or U8544 (N_8544,N_7518,N_7975);
xnor U8545 (N_8545,N_6003,N_6662);
or U8546 (N_8546,N_7124,N_7580);
and U8547 (N_8547,N_6045,N_7318);
or U8548 (N_8548,N_6607,N_6109);
nor U8549 (N_8549,N_6916,N_7798);
nor U8550 (N_8550,N_7935,N_7861);
nor U8551 (N_8551,N_7694,N_6876);
and U8552 (N_8552,N_7495,N_7461);
nand U8553 (N_8553,N_7025,N_6623);
nand U8554 (N_8554,N_7469,N_6136);
nor U8555 (N_8555,N_7916,N_7695);
xnor U8556 (N_8556,N_7942,N_7097);
nand U8557 (N_8557,N_7547,N_7905);
nand U8558 (N_8558,N_6724,N_6934);
nand U8559 (N_8559,N_7780,N_7471);
nor U8560 (N_8560,N_6249,N_6233);
and U8561 (N_8561,N_6878,N_7209);
and U8562 (N_8562,N_6327,N_7781);
nor U8563 (N_8563,N_6062,N_6501);
nand U8564 (N_8564,N_6220,N_6199);
and U8565 (N_8565,N_6246,N_7595);
or U8566 (N_8566,N_7292,N_6070);
and U8567 (N_8567,N_7426,N_6638);
or U8568 (N_8568,N_7466,N_6856);
and U8569 (N_8569,N_7921,N_7559);
and U8570 (N_8570,N_7501,N_6284);
xnor U8571 (N_8571,N_7540,N_7943);
nand U8572 (N_8572,N_6172,N_7677);
nor U8573 (N_8573,N_6667,N_7307);
and U8574 (N_8574,N_6010,N_7981);
nand U8575 (N_8575,N_7363,N_6362);
nand U8576 (N_8576,N_6725,N_6630);
nor U8577 (N_8577,N_7971,N_6555);
and U8578 (N_8578,N_7679,N_7030);
and U8579 (N_8579,N_7805,N_6019);
nor U8580 (N_8580,N_6727,N_7535);
nor U8581 (N_8581,N_7617,N_6744);
nor U8582 (N_8582,N_7227,N_7807);
nor U8583 (N_8583,N_7591,N_7413);
or U8584 (N_8584,N_7281,N_6675);
nor U8585 (N_8585,N_7467,N_6212);
or U8586 (N_8586,N_7801,N_6429);
or U8587 (N_8587,N_7533,N_7974);
and U8588 (N_8588,N_7073,N_6118);
and U8589 (N_8589,N_7343,N_7473);
nand U8590 (N_8590,N_6189,N_7396);
nand U8591 (N_8591,N_7427,N_6522);
nor U8592 (N_8592,N_6867,N_7602);
or U8593 (N_8593,N_6224,N_7862);
or U8594 (N_8594,N_6905,N_6396);
and U8595 (N_8595,N_6779,N_7385);
nand U8596 (N_8596,N_7497,N_7953);
or U8597 (N_8597,N_7270,N_7845);
or U8598 (N_8598,N_6025,N_7920);
nor U8599 (N_8599,N_7500,N_7309);
nand U8600 (N_8600,N_6157,N_7354);
nor U8601 (N_8601,N_6347,N_7499);
xnor U8602 (N_8602,N_7419,N_6098);
or U8603 (N_8603,N_6191,N_6217);
xnor U8604 (N_8604,N_6161,N_6088);
xor U8605 (N_8605,N_6084,N_7415);
nor U8606 (N_8606,N_7541,N_6079);
or U8607 (N_8607,N_6911,N_6044);
nand U8608 (N_8608,N_7448,N_6439);
or U8609 (N_8609,N_7275,N_6831);
or U8610 (N_8610,N_7665,N_6247);
nand U8611 (N_8611,N_6927,N_7160);
or U8612 (N_8612,N_7477,N_7444);
nor U8613 (N_8613,N_7153,N_6872);
and U8614 (N_8614,N_7529,N_7841);
xnor U8615 (N_8615,N_6661,N_7964);
nand U8616 (N_8616,N_6346,N_7936);
or U8617 (N_8617,N_7416,N_7545);
nand U8618 (N_8618,N_7775,N_6992);
and U8619 (N_8619,N_7297,N_7640);
or U8620 (N_8620,N_7719,N_6562);
and U8621 (N_8621,N_7107,N_6852);
nor U8622 (N_8622,N_7507,N_7900);
and U8623 (N_8623,N_6446,N_6799);
nand U8624 (N_8624,N_7202,N_6186);
and U8625 (N_8625,N_7381,N_6798);
or U8626 (N_8626,N_6516,N_6474);
nor U8627 (N_8627,N_6391,N_6766);
nand U8628 (N_8628,N_6350,N_7220);
and U8629 (N_8629,N_6119,N_7924);
or U8630 (N_8630,N_6707,N_7423);
or U8631 (N_8631,N_6776,N_6888);
or U8632 (N_8632,N_6485,N_6832);
and U8633 (N_8633,N_6481,N_7100);
xnor U8634 (N_8634,N_6180,N_6437);
nor U8635 (N_8635,N_7968,N_7145);
and U8636 (N_8636,N_6144,N_7406);
xnor U8637 (N_8637,N_6232,N_7741);
nor U8638 (N_8638,N_6231,N_6258);
nand U8639 (N_8639,N_7045,N_6703);
nor U8640 (N_8640,N_7007,N_6768);
xor U8641 (N_8641,N_7612,N_7732);
nand U8642 (N_8642,N_6976,N_6941);
or U8643 (N_8643,N_6761,N_7076);
or U8644 (N_8644,N_7579,N_7952);
or U8645 (N_8645,N_6729,N_6517);
or U8646 (N_8646,N_6052,N_7858);
or U8647 (N_8647,N_7311,N_6674);
nor U8648 (N_8648,N_7759,N_6447);
nand U8649 (N_8649,N_6355,N_6091);
xnor U8650 (N_8650,N_6505,N_7141);
or U8651 (N_8651,N_6914,N_7046);
nand U8652 (N_8652,N_6015,N_6256);
nand U8653 (N_8653,N_6995,N_7892);
or U8654 (N_8654,N_7106,N_7609);
or U8655 (N_8655,N_7265,N_6137);
xnor U8656 (N_8656,N_7847,N_6802);
nor U8657 (N_8657,N_6469,N_7487);
nand U8658 (N_8658,N_7769,N_7425);
xnor U8659 (N_8659,N_6207,N_7812);
or U8660 (N_8660,N_7229,N_6784);
or U8661 (N_8661,N_7913,N_7725);
nand U8662 (N_8662,N_6542,N_6094);
and U8663 (N_8663,N_6688,N_7099);
and U8664 (N_8664,N_7552,N_6849);
or U8665 (N_8665,N_7874,N_6000);
and U8666 (N_8666,N_7588,N_6728);
nand U8667 (N_8667,N_6417,N_7201);
nor U8668 (N_8668,N_6479,N_6352);
or U8669 (N_8669,N_6314,N_7705);
or U8670 (N_8670,N_7365,N_7893);
nand U8671 (N_8671,N_6331,N_7349);
nand U8672 (N_8672,N_6620,N_7263);
or U8673 (N_8673,N_6734,N_6187);
nand U8674 (N_8674,N_7799,N_7616);
or U8675 (N_8675,N_7112,N_7582);
or U8676 (N_8676,N_7456,N_6349);
and U8677 (N_8677,N_6165,N_6909);
and U8678 (N_8678,N_6021,N_6683);
nand U8679 (N_8679,N_7908,N_6370);
or U8680 (N_8680,N_7398,N_6204);
nor U8681 (N_8681,N_7860,N_7925);
nand U8682 (N_8682,N_6753,N_6359);
and U8683 (N_8683,N_7139,N_7554);
or U8684 (N_8684,N_6400,N_6432);
or U8685 (N_8685,N_6030,N_6114);
and U8686 (N_8686,N_6717,N_6611);
nand U8687 (N_8687,N_7336,N_6305);
or U8688 (N_8688,N_6467,N_6554);
nand U8689 (N_8689,N_7825,N_7565);
xor U8690 (N_8690,N_7776,N_7823);
and U8691 (N_8691,N_6669,N_7008);
nand U8692 (N_8692,N_6964,N_6493);
nand U8693 (N_8693,N_7955,N_7028);
or U8694 (N_8694,N_6363,N_6342);
nand U8695 (N_8695,N_6970,N_6877);
nand U8696 (N_8696,N_6211,N_7067);
or U8697 (N_8697,N_6806,N_7998);
nor U8698 (N_8698,N_7081,N_7623);
and U8699 (N_8699,N_7651,N_7983);
xor U8700 (N_8700,N_6190,N_6111);
nand U8701 (N_8701,N_6227,N_7783);
and U8702 (N_8702,N_7346,N_6536);
nor U8703 (N_8703,N_6820,N_7388);
or U8704 (N_8704,N_6135,N_7492);
or U8705 (N_8705,N_7957,N_7296);
or U8706 (N_8706,N_7782,N_6991);
nand U8707 (N_8707,N_7167,N_6024);
nor U8708 (N_8708,N_6610,N_6908);
nand U8709 (N_8709,N_6296,N_6106);
nor U8710 (N_8710,N_6648,N_6298);
nor U8711 (N_8711,N_7977,N_6785);
nand U8712 (N_8712,N_7390,N_7762);
and U8713 (N_8713,N_6041,N_6643);
or U8714 (N_8714,N_7277,N_6226);
nor U8715 (N_8715,N_6812,N_7560);
or U8716 (N_8716,N_7011,N_7820);
nor U8717 (N_8717,N_6949,N_7661);
or U8718 (N_8718,N_6461,N_6122);
and U8719 (N_8719,N_6537,N_7826);
or U8720 (N_8720,N_7040,N_7039);
or U8721 (N_8721,N_6007,N_6524);
nor U8722 (N_8722,N_7701,N_7760);
nand U8723 (N_8723,N_7098,N_6268);
nor U8724 (N_8724,N_7791,N_7613);
nor U8725 (N_8725,N_7316,N_7857);
nor U8726 (N_8726,N_6159,N_7191);
nor U8727 (N_8727,N_6925,N_6660);
nor U8728 (N_8728,N_6228,N_7885);
and U8729 (N_8729,N_6988,N_7333);
and U8730 (N_8730,N_6465,N_6238);
nand U8731 (N_8731,N_7814,N_6883);
and U8732 (N_8732,N_7562,N_7041);
nor U8733 (N_8733,N_6552,N_6409);
or U8734 (N_8734,N_7539,N_7619);
nand U8735 (N_8735,N_6654,N_6155);
nand U8736 (N_8736,N_7897,N_7211);
nand U8737 (N_8737,N_7149,N_6147);
or U8738 (N_8738,N_7653,N_6158);
nand U8739 (N_8739,N_7420,N_7941);
or U8740 (N_8740,N_7159,N_6455);
nand U8741 (N_8741,N_6124,N_7254);
nand U8742 (N_8742,N_7951,N_7294);
nor U8743 (N_8743,N_6164,N_7142);
nand U8744 (N_8744,N_7727,N_6492);
xor U8745 (N_8745,N_6110,N_6539);
nor U8746 (N_8746,N_6145,N_7403);
or U8747 (N_8747,N_7581,N_6573);
nor U8748 (N_8748,N_6588,N_6912);
nand U8749 (N_8749,N_7394,N_7454);
nand U8750 (N_8750,N_7207,N_6928);
xnor U8751 (N_8751,N_7480,N_6659);
nand U8752 (N_8752,N_7652,N_6981);
nor U8753 (N_8753,N_6614,N_7838);
nand U8754 (N_8754,N_6090,N_6445);
and U8755 (N_8755,N_6156,N_6141);
and U8756 (N_8756,N_6450,N_6054);
and U8757 (N_8757,N_7829,N_7212);
nor U8758 (N_8758,N_6814,N_7896);
nor U8759 (N_8759,N_7105,N_7374);
nor U8760 (N_8760,N_7817,N_6060);
and U8761 (N_8761,N_7351,N_7618);
or U8762 (N_8762,N_6151,N_6866);
nand U8763 (N_8763,N_6390,N_7077);
nand U8764 (N_8764,N_7367,N_6980);
nand U8765 (N_8765,N_6027,N_7376);
or U8766 (N_8766,N_7594,N_6920);
nand U8767 (N_8767,N_6453,N_6480);
and U8768 (N_8768,N_6321,N_6580);
and U8769 (N_8769,N_6634,N_6682);
and U8770 (N_8770,N_7020,N_7360);
or U8771 (N_8771,N_7109,N_6299);
xnor U8772 (N_8772,N_7508,N_7217);
nand U8773 (N_8773,N_7656,N_6910);
and U8774 (N_8774,N_7692,N_6169);
nor U8775 (N_8775,N_7055,N_6020);
nand U8776 (N_8776,N_6886,N_6279);
xor U8777 (N_8777,N_6219,N_7978);
or U8778 (N_8778,N_6004,N_6750);
or U8779 (N_8779,N_7700,N_7504);
or U8780 (N_8780,N_7683,N_7485);
or U8781 (N_8781,N_7470,N_6468);
and U8782 (N_8782,N_7786,N_7536);
nand U8783 (N_8783,N_7452,N_6547);
nand U8784 (N_8784,N_6561,N_7015);
nand U8785 (N_8785,N_7386,N_6393);
or U8786 (N_8786,N_7796,N_6116);
and U8787 (N_8787,N_7994,N_6050);
nor U8788 (N_8788,N_6254,N_6078);
and U8789 (N_8789,N_6576,N_7113);
nand U8790 (N_8790,N_6808,N_7190);
or U8791 (N_8791,N_6983,N_7717);
nand U8792 (N_8792,N_7002,N_6624);
or U8793 (N_8793,N_6128,N_6738);
nand U8794 (N_8794,N_7667,N_7090);
and U8795 (N_8795,N_7272,N_6932);
and U8796 (N_8796,N_7393,N_7342);
nand U8797 (N_8797,N_6957,N_6984);
or U8798 (N_8798,N_7035,N_6844);
or U8799 (N_8799,N_7926,N_6063);
and U8800 (N_8800,N_7057,N_7684);
and U8801 (N_8801,N_7668,N_6477);
or U8802 (N_8802,N_6495,N_6177);
xor U8803 (N_8803,N_7337,N_6365);
or U8804 (N_8804,N_6786,N_7183);
xor U8805 (N_8805,N_6463,N_6320);
and U8806 (N_8806,N_6906,N_6002);
xor U8807 (N_8807,N_7740,N_6304);
or U8808 (N_8808,N_6066,N_6153);
xnor U8809 (N_8809,N_6665,N_7291);
nor U8810 (N_8810,N_7295,N_6127);
or U8811 (N_8811,N_7876,N_6073);
xor U8812 (N_8812,N_6922,N_7187);
nand U8813 (N_8813,N_6372,N_6593);
or U8814 (N_8814,N_7458,N_6085);
and U8815 (N_8815,N_7255,N_7026);
or U8816 (N_8816,N_6237,N_7060);
or U8817 (N_8817,N_7181,N_6029);
nand U8818 (N_8818,N_7598,N_7258);
nand U8819 (N_8819,N_6009,N_6871);
xor U8820 (N_8820,N_6215,N_7730);
or U8821 (N_8821,N_7879,N_7655);
xnor U8822 (N_8822,N_6845,N_6678);
nor U8823 (N_8823,N_6377,N_7369);
and U8824 (N_8824,N_7863,N_7490);
nand U8825 (N_8825,N_6777,N_6713);
nand U8826 (N_8826,N_6095,N_6652);
xor U8827 (N_8827,N_7839,N_6065);
xnor U8828 (N_8828,N_6489,N_7637);
xor U8829 (N_8829,N_6642,N_6801);
nand U8830 (N_8830,N_6087,N_7669);
nor U8831 (N_8831,N_7726,N_7778);
xor U8832 (N_8832,N_7038,N_6598);
or U8833 (N_8833,N_6663,N_7224);
or U8834 (N_8834,N_7118,N_7686);
xor U8835 (N_8835,N_6968,N_6818);
nor U8836 (N_8836,N_7021,N_6057);
nor U8837 (N_8837,N_6658,N_6496);
or U8838 (N_8838,N_7199,N_7939);
nand U8839 (N_8839,N_7819,N_7585);
and U8840 (N_8840,N_7429,N_7607);
and U8841 (N_8841,N_6209,N_6442);
xnor U8842 (N_8842,N_7650,N_6415);
or U8843 (N_8843,N_7358,N_6792);
or U8844 (N_8844,N_7890,N_7997);
nand U8845 (N_8845,N_6378,N_7226);
nor U8846 (N_8846,N_7710,N_7698);
and U8847 (N_8847,N_6526,N_7029);
or U8848 (N_8848,N_6328,N_6797);
nand U8849 (N_8849,N_6790,N_6102);
or U8850 (N_8850,N_7803,N_7315);
nor U8851 (N_8851,N_7033,N_7703);
and U8852 (N_8852,N_6712,N_6592);
nor U8853 (N_8853,N_7121,N_7483);
nor U8854 (N_8854,N_6303,N_7743);
or U8855 (N_8855,N_7966,N_6418);
and U8856 (N_8856,N_6942,N_6192);
xor U8857 (N_8857,N_6758,N_6394);
xor U8858 (N_8858,N_7764,N_7569);
nand U8859 (N_8859,N_7421,N_6334);
nor U8860 (N_8860,N_6154,N_7156);
nand U8861 (N_8861,N_6868,N_7430);
and U8862 (N_8862,N_7110,N_7929);
nand U8863 (N_8863,N_7811,N_7089);
nor U8864 (N_8864,N_7919,N_7641);
nand U8865 (N_8865,N_6699,N_7250);
xnor U8866 (N_8866,N_6873,N_7930);
or U8867 (N_8867,N_6956,N_7050);
or U8868 (N_8868,N_6176,N_6771);
nor U8869 (N_8869,N_7482,N_7550);
nor U8870 (N_8870,N_6861,N_7802);
nor U8871 (N_8871,N_6195,N_6083);
nand U8872 (N_8872,N_6392,N_6870);
nor U8873 (N_8873,N_7965,N_7945);
nand U8874 (N_8874,N_7523,N_7813);
or U8875 (N_8875,N_7451,N_6441);
or U8876 (N_8876,N_6567,N_6998);
and U8877 (N_8877,N_7463,N_6513);
nand U8878 (N_8878,N_7131,N_6043);
or U8879 (N_8879,N_6385,N_6200);
nand U8880 (N_8880,N_7282,N_7546);
nand U8881 (N_8881,N_6487,N_7681);
and U8882 (N_8882,N_7629,N_7923);
nor U8883 (N_8883,N_6126,N_6551);
nand U8884 (N_8884,N_7806,N_6769);
and U8885 (N_8885,N_6714,N_7950);
nand U8886 (N_8886,N_6563,N_6583);
and U8887 (N_8887,N_6549,N_7455);
nor U8888 (N_8888,N_6201,N_6500);
nor U8889 (N_8889,N_7096,N_7148);
nand U8890 (N_8890,N_6081,N_7188);
and U8891 (N_8891,N_6252,N_7884);
nand U8892 (N_8892,N_7068,N_7940);
nand U8893 (N_8893,N_7137,N_6841);
or U8894 (N_8894,N_6833,N_7662);
or U8895 (N_8895,N_7894,N_6599);
xnor U8896 (N_8896,N_7302,N_6408);
nand U8897 (N_8897,N_6695,N_6266);
and U8898 (N_8898,N_6071,N_7331);
nand U8899 (N_8899,N_7673,N_6283);
xor U8900 (N_8900,N_7243,N_6278);
nand U8901 (N_8901,N_7834,N_6645);
nand U8902 (N_8902,N_6023,N_6423);
nand U8903 (N_8903,N_7854,N_6013);
and U8904 (N_8904,N_7898,N_7407);
nor U8905 (N_8905,N_7173,N_7078);
and U8906 (N_8906,N_6038,N_7228);
nor U8907 (N_8907,N_7257,N_6795);
and U8908 (N_8908,N_7872,N_6313);
nor U8909 (N_8909,N_7059,N_7848);
nor U8910 (N_8910,N_6532,N_7995);
nor U8911 (N_8911,N_6280,N_6335);
and U8912 (N_8912,N_7278,N_6989);
nand U8913 (N_8913,N_6240,N_6858);
xor U8914 (N_8914,N_6123,N_7948);
or U8915 (N_8915,N_6863,N_7404);
nor U8916 (N_8916,N_6012,N_7061);
and U8917 (N_8917,N_6901,N_7128);
nand U8918 (N_8918,N_6556,N_7377);
nand U8919 (N_8919,N_6179,N_6668);
nor U8920 (N_8920,N_6670,N_7724);
nand U8921 (N_8921,N_7436,N_7064);
nor U8922 (N_8922,N_6277,N_6133);
nand U8923 (N_8923,N_6860,N_6276);
nor U8924 (N_8924,N_6621,N_7544);
nor U8925 (N_8925,N_7306,N_7143);
xnor U8926 (N_8926,N_6288,N_6341);
or U8927 (N_8927,N_6772,N_7649);
nand U8928 (N_8928,N_6657,N_7996);
and U8929 (N_8929,N_7215,N_6584);
nand U8930 (N_8930,N_7711,N_7903);
or U8931 (N_8931,N_6595,N_7400);
nor U8932 (N_8932,N_6641,N_7922);
and U8933 (N_8933,N_6086,N_6028);
nand U8934 (N_8934,N_6033,N_7244);
nor U8935 (N_8935,N_7357,N_7329);
nor U8936 (N_8936,N_7837,N_7194);
xnor U8937 (N_8937,N_7530,N_7592);
or U8938 (N_8938,N_6506,N_7359);
nor U8939 (N_8939,N_6961,N_6559);
and U8940 (N_8940,N_6440,N_7453);
nor U8941 (N_8941,N_7645,N_6996);
nor U8942 (N_8942,N_7784,N_7693);
nand U8943 (N_8943,N_6491,N_7120);
and U8944 (N_8944,N_7824,N_6783);
and U8945 (N_8945,N_6540,N_7176);
xnor U8946 (N_8946,N_6498,N_7635);
nor U8947 (N_8947,N_7590,N_6926);
and U8948 (N_8948,N_7987,N_6757);
or U8949 (N_8949,N_6967,N_6022);
nand U8950 (N_8950,N_7438,N_6825);
and U8951 (N_8951,N_7871,N_7659);
nand U8952 (N_8952,N_7184,N_7195);
nor U8953 (N_8953,N_6969,N_6384);
and U8954 (N_8954,N_7850,N_7489);
and U8955 (N_8955,N_6476,N_6100);
or U8956 (N_8956,N_6163,N_6553);
and U8957 (N_8957,N_6782,N_6458);
nor U8958 (N_8958,N_6817,N_7680);
and U8959 (N_8959,N_6646,N_7313);
or U8960 (N_8960,N_7323,N_7777);
or U8961 (N_8961,N_6843,N_7051);
or U8962 (N_8962,N_6902,N_7901);
nand U8963 (N_8963,N_6430,N_6388);
nand U8964 (N_8964,N_7491,N_7972);
nand U8965 (N_8965,N_6875,N_7208);
and U8966 (N_8966,N_6241,N_7749);
and U8967 (N_8967,N_7122,N_6184);
and U8968 (N_8968,N_6115,N_6175);
or U8969 (N_8969,N_6046,N_6627);
and U8970 (N_8970,N_6723,N_7992);
or U8971 (N_8971,N_6336,N_6112);
nor U8972 (N_8972,N_6357,N_7723);
and U8973 (N_8973,N_7878,N_7321);
and U8974 (N_8974,N_7012,N_6251);
nand U8975 (N_8975,N_7520,N_6899);
or U8976 (N_8976,N_6793,N_6543);
or U8977 (N_8977,N_7016,N_7566);
or U8978 (N_8978,N_7314,N_7556);
nor U8979 (N_8979,N_7378,N_6395);
or U8980 (N_8980,N_6149,N_6881);
or U8981 (N_8981,N_7117,N_7895);
xnor U8982 (N_8982,N_6051,N_6615);
or U8983 (N_8983,N_6375,N_7391);
nand U8984 (N_8984,N_7312,N_6826);
nand U8985 (N_8985,N_6058,N_7503);
nor U8986 (N_8986,N_7158,N_7630);
and U8987 (N_8987,N_7869,N_6924);
or U8988 (N_8988,N_6456,N_6281);
and U8989 (N_8989,N_6511,N_6412);
nand U8990 (N_8990,N_7843,N_7642);
and U8991 (N_8991,N_7809,N_7716);
or U8992 (N_8992,N_7353,N_6132);
nor U8993 (N_8993,N_6475,N_6960);
or U8994 (N_8994,N_7355,N_6064);
or U8995 (N_8995,N_6687,N_7626);
and U8996 (N_8996,N_6287,N_7835);
nor U8997 (N_8997,N_6301,N_7864);
nor U8998 (N_8998,N_6261,N_7335);
and U8999 (N_8999,N_6805,N_7574);
or U9000 (N_9000,N_7100,N_7969);
xor U9001 (N_9001,N_7473,N_6323);
nand U9002 (N_9002,N_7487,N_6924);
nand U9003 (N_9003,N_6006,N_6343);
nand U9004 (N_9004,N_7312,N_6109);
or U9005 (N_9005,N_6288,N_6909);
nand U9006 (N_9006,N_7373,N_6646);
nor U9007 (N_9007,N_7388,N_6387);
or U9008 (N_9008,N_6730,N_6315);
and U9009 (N_9009,N_7473,N_6488);
nor U9010 (N_9010,N_6390,N_7845);
and U9011 (N_9011,N_7007,N_6590);
or U9012 (N_9012,N_7101,N_7156);
nand U9013 (N_9013,N_7892,N_6521);
nor U9014 (N_9014,N_7812,N_7900);
and U9015 (N_9015,N_6109,N_7805);
or U9016 (N_9016,N_6250,N_6761);
nand U9017 (N_9017,N_7867,N_7155);
nand U9018 (N_9018,N_6125,N_7348);
and U9019 (N_9019,N_6038,N_6324);
nor U9020 (N_9020,N_6970,N_6901);
xnor U9021 (N_9021,N_6697,N_7285);
nor U9022 (N_9022,N_6814,N_7715);
nor U9023 (N_9023,N_6537,N_6085);
or U9024 (N_9024,N_6263,N_7823);
nand U9025 (N_9025,N_6646,N_6812);
xnor U9026 (N_9026,N_7873,N_7826);
xnor U9027 (N_9027,N_7115,N_6290);
and U9028 (N_9028,N_7061,N_6771);
nor U9029 (N_9029,N_6725,N_7157);
or U9030 (N_9030,N_6554,N_7358);
nor U9031 (N_9031,N_7535,N_6554);
xnor U9032 (N_9032,N_7331,N_7656);
and U9033 (N_9033,N_6256,N_6768);
nand U9034 (N_9034,N_7517,N_7748);
and U9035 (N_9035,N_6978,N_6093);
nand U9036 (N_9036,N_6899,N_6639);
nor U9037 (N_9037,N_7802,N_6306);
or U9038 (N_9038,N_7699,N_6201);
nand U9039 (N_9039,N_6098,N_6167);
or U9040 (N_9040,N_7436,N_6527);
nand U9041 (N_9041,N_7121,N_6751);
nand U9042 (N_9042,N_7136,N_7114);
nand U9043 (N_9043,N_7034,N_6566);
nor U9044 (N_9044,N_6908,N_6755);
or U9045 (N_9045,N_7553,N_6508);
or U9046 (N_9046,N_6797,N_7543);
xnor U9047 (N_9047,N_7079,N_7170);
or U9048 (N_9048,N_6172,N_6552);
nand U9049 (N_9049,N_7875,N_6205);
nor U9050 (N_9050,N_6745,N_7321);
xor U9051 (N_9051,N_7997,N_7867);
or U9052 (N_9052,N_6357,N_6483);
and U9053 (N_9053,N_6133,N_7436);
and U9054 (N_9054,N_6014,N_7539);
or U9055 (N_9055,N_7341,N_6379);
and U9056 (N_9056,N_7430,N_6093);
and U9057 (N_9057,N_6816,N_7336);
nand U9058 (N_9058,N_7850,N_7710);
nand U9059 (N_9059,N_6746,N_7915);
nor U9060 (N_9060,N_7042,N_7992);
or U9061 (N_9061,N_7451,N_7746);
nand U9062 (N_9062,N_6500,N_6301);
xor U9063 (N_9063,N_7580,N_6140);
nand U9064 (N_9064,N_7639,N_6687);
nand U9065 (N_9065,N_7478,N_6642);
and U9066 (N_9066,N_6940,N_6702);
nand U9067 (N_9067,N_6820,N_6962);
and U9068 (N_9068,N_7066,N_7787);
nand U9069 (N_9069,N_7981,N_7539);
nor U9070 (N_9070,N_7646,N_7206);
or U9071 (N_9071,N_6376,N_6137);
nor U9072 (N_9072,N_6249,N_7664);
xor U9073 (N_9073,N_6390,N_6569);
nor U9074 (N_9074,N_6564,N_6777);
nor U9075 (N_9075,N_7590,N_6945);
nor U9076 (N_9076,N_7415,N_6004);
and U9077 (N_9077,N_7850,N_6879);
or U9078 (N_9078,N_7301,N_7610);
or U9079 (N_9079,N_7929,N_7375);
or U9080 (N_9080,N_6663,N_6480);
or U9081 (N_9081,N_6525,N_6467);
nand U9082 (N_9082,N_6927,N_6865);
nor U9083 (N_9083,N_7894,N_6571);
nand U9084 (N_9084,N_6926,N_7616);
or U9085 (N_9085,N_6459,N_6898);
xnor U9086 (N_9086,N_7288,N_6186);
nand U9087 (N_9087,N_7348,N_6514);
or U9088 (N_9088,N_6163,N_7270);
xor U9089 (N_9089,N_6240,N_7058);
and U9090 (N_9090,N_6364,N_7502);
nor U9091 (N_9091,N_7913,N_6925);
nand U9092 (N_9092,N_6233,N_7695);
nand U9093 (N_9093,N_6801,N_6603);
or U9094 (N_9094,N_6589,N_7424);
or U9095 (N_9095,N_7798,N_7300);
nor U9096 (N_9096,N_7437,N_7601);
nand U9097 (N_9097,N_7013,N_6870);
nor U9098 (N_9098,N_6385,N_6857);
nor U9099 (N_9099,N_6594,N_7906);
and U9100 (N_9100,N_7097,N_6186);
nor U9101 (N_9101,N_6255,N_7658);
nand U9102 (N_9102,N_6803,N_6784);
and U9103 (N_9103,N_7897,N_6790);
and U9104 (N_9104,N_7505,N_6745);
nor U9105 (N_9105,N_6289,N_6625);
or U9106 (N_9106,N_7829,N_7495);
and U9107 (N_9107,N_7215,N_6221);
nor U9108 (N_9108,N_7032,N_6763);
or U9109 (N_9109,N_6795,N_7650);
or U9110 (N_9110,N_6012,N_7198);
nand U9111 (N_9111,N_7964,N_7632);
nand U9112 (N_9112,N_6460,N_7278);
or U9113 (N_9113,N_6675,N_7502);
xnor U9114 (N_9114,N_6516,N_6977);
and U9115 (N_9115,N_6747,N_6831);
and U9116 (N_9116,N_6669,N_7624);
nand U9117 (N_9117,N_6330,N_6671);
and U9118 (N_9118,N_7094,N_6496);
or U9119 (N_9119,N_7109,N_6139);
nand U9120 (N_9120,N_7295,N_7052);
and U9121 (N_9121,N_6322,N_6064);
nor U9122 (N_9122,N_6156,N_6572);
and U9123 (N_9123,N_6795,N_6125);
and U9124 (N_9124,N_6708,N_7887);
nand U9125 (N_9125,N_6825,N_7718);
or U9126 (N_9126,N_6241,N_6733);
or U9127 (N_9127,N_7290,N_7491);
or U9128 (N_9128,N_7297,N_7505);
nor U9129 (N_9129,N_7859,N_6325);
or U9130 (N_9130,N_6800,N_7518);
nand U9131 (N_9131,N_6636,N_7409);
nand U9132 (N_9132,N_6467,N_6873);
nor U9133 (N_9133,N_7298,N_7611);
or U9134 (N_9134,N_7517,N_7121);
or U9135 (N_9135,N_6630,N_7452);
or U9136 (N_9136,N_6470,N_7721);
and U9137 (N_9137,N_7955,N_6119);
and U9138 (N_9138,N_6404,N_6960);
and U9139 (N_9139,N_6193,N_6293);
or U9140 (N_9140,N_6284,N_6871);
and U9141 (N_9141,N_7379,N_7825);
nand U9142 (N_9142,N_7982,N_6004);
xor U9143 (N_9143,N_7902,N_6363);
or U9144 (N_9144,N_6761,N_7307);
and U9145 (N_9145,N_7463,N_7677);
or U9146 (N_9146,N_6253,N_6873);
xnor U9147 (N_9147,N_7801,N_7031);
and U9148 (N_9148,N_7313,N_7505);
or U9149 (N_9149,N_7556,N_6942);
and U9150 (N_9150,N_7798,N_6729);
nor U9151 (N_9151,N_6879,N_6267);
nor U9152 (N_9152,N_7577,N_6315);
nand U9153 (N_9153,N_7982,N_7044);
nor U9154 (N_9154,N_6317,N_6119);
xnor U9155 (N_9155,N_6580,N_7193);
and U9156 (N_9156,N_6848,N_6309);
and U9157 (N_9157,N_7196,N_7531);
nand U9158 (N_9158,N_6802,N_6408);
nor U9159 (N_9159,N_6479,N_7156);
and U9160 (N_9160,N_7215,N_6211);
nor U9161 (N_9161,N_7707,N_6864);
nor U9162 (N_9162,N_7144,N_7054);
nor U9163 (N_9163,N_7598,N_6872);
nor U9164 (N_9164,N_7061,N_6088);
and U9165 (N_9165,N_6828,N_7169);
nor U9166 (N_9166,N_7471,N_6699);
or U9167 (N_9167,N_6987,N_6448);
nand U9168 (N_9168,N_7392,N_6628);
nor U9169 (N_9169,N_6105,N_7497);
nand U9170 (N_9170,N_6597,N_7715);
or U9171 (N_9171,N_7221,N_7927);
nor U9172 (N_9172,N_7451,N_6687);
xnor U9173 (N_9173,N_6454,N_7442);
nor U9174 (N_9174,N_6293,N_6255);
and U9175 (N_9175,N_6509,N_7966);
and U9176 (N_9176,N_6673,N_6630);
or U9177 (N_9177,N_6118,N_7115);
nor U9178 (N_9178,N_7199,N_7448);
xnor U9179 (N_9179,N_6613,N_7858);
nor U9180 (N_9180,N_6420,N_7671);
and U9181 (N_9181,N_7166,N_7968);
or U9182 (N_9182,N_7994,N_6860);
xnor U9183 (N_9183,N_7278,N_7177);
nand U9184 (N_9184,N_6557,N_6462);
nor U9185 (N_9185,N_6941,N_7738);
or U9186 (N_9186,N_7119,N_7631);
and U9187 (N_9187,N_6171,N_6351);
and U9188 (N_9188,N_7238,N_6780);
or U9189 (N_9189,N_7180,N_7875);
nor U9190 (N_9190,N_7721,N_7648);
nor U9191 (N_9191,N_6647,N_6403);
xnor U9192 (N_9192,N_7917,N_6868);
nand U9193 (N_9193,N_6376,N_6428);
nor U9194 (N_9194,N_6232,N_6968);
or U9195 (N_9195,N_6037,N_7398);
nor U9196 (N_9196,N_7116,N_6019);
or U9197 (N_9197,N_6637,N_6115);
nor U9198 (N_9198,N_6931,N_7502);
or U9199 (N_9199,N_7027,N_6433);
xor U9200 (N_9200,N_6050,N_6731);
nor U9201 (N_9201,N_7267,N_6396);
nor U9202 (N_9202,N_7948,N_6110);
xnor U9203 (N_9203,N_7415,N_7276);
nor U9204 (N_9204,N_7552,N_7982);
or U9205 (N_9205,N_7814,N_6959);
nand U9206 (N_9206,N_7073,N_6697);
or U9207 (N_9207,N_6452,N_6753);
nand U9208 (N_9208,N_7215,N_6043);
or U9209 (N_9209,N_6609,N_6651);
and U9210 (N_9210,N_6700,N_7956);
or U9211 (N_9211,N_6367,N_7938);
xnor U9212 (N_9212,N_7958,N_7260);
nor U9213 (N_9213,N_6423,N_7313);
xor U9214 (N_9214,N_7377,N_7196);
nand U9215 (N_9215,N_7654,N_6584);
xnor U9216 (N_9216,N_6714,N_7144);
nand U9217 (N_9217,N_6093,N_7046);
xnor U9218 (N_9218,N_7265,N_6436);
nor U9219 (N_9219,N_6298,N_7567);
and U9220 (N_9220,N_7879,N_7430);
nand U9221 (N_9221,N_7885,N_7145);
nand U9222 (N_9222,N_6179,N_7658);
and U9223 (N_9223,N_6342,N_7072);
nand U9224 (N_9224,N_7329,N_6940);
and U9225 (N_9225,N_7718,N_7017);
nand U9226 (N_9226,N_6256,N_6677);
and U9227 (N_9227,N_6491,N_7394);
or U9228 (N_9228,N_7664,N_7908);
and U9229 (N_9229,N_6195,N_7643);
or U9230 (N_9230,N_6131,N_7067);
nor U9231 (N_9231,N_6529,N_7986);
nor U9232 (N_9232,N_7849,N_7816);
and U9233 (N_9233,N_7529,N_6920);
and U9234 (N_9234,N_6016,N_7689);
and U9235 (N_9235,N_6779,N_7291);
and U9236 (N_9236,N_6609,N_7944);
and U9237 (N_9237,N_7399,N_6895);
xor U9238 (N_9238,N_6140,N_7221);
or U9239 (N_9239,N_7098,N_7545);
nor U9240 (N_9240,N_7376,N_7743);
and U9241 (N_9241,N_7940,N_6731);
and U9242 (N_9242,N_7964,N_6204);
or U9243 (N_9243,N_6063,N_6006);
nand U9244 (N_9244,N_6500,N_6534);
and U9245 (N_9245,N_7468,N_7743);
or U9246 (N_9246,N_6318,N_7823);
nor U9247 (N_9247,N_6965,N_7559);
xnor U9248 (N_9248,N_7111,N_6190);
and U9249 (N_9249,N_7821,N_7365);
nor U9250 (N_9250,N_7051,N_6270);
and U9251 (N_9251,N_6648,N_7210);
xnor U9252 (N_9252,N_7058,N_6083);
nand U9253 (N_9253,N_7593,N_7761);
nor U9254 (N_9254,N_7231,N_6145);
and U9255 (N_9255,N_6475,N_7283);
xnor U9256 (N_9256,N_7760,N_6481);
and U9257 (N_9257,N_7399,N_6335);
and U9258 (N_9258,N_7801,N_6001);
nor U9259 (N_9259,N_7389,N_6009);
nand U9260 (N_9260,N_7999,N_7248);
or U9261 (N_9261,N_6346,N_6986);
and U9262 (N_9262,N_6394,N_6145);
nor U9263 (N_9263,N_6911,N_6514);
nand U9264 (N_9264,N_6376,N_6697);
or U9265 (N_9265,N_7089,N_7389);
nor U9266 (N_9266,N_6104,N_7430);
nand U9267 (N_9267,N_6622,N_7384);
and U9268 (N_9268,N_6165,N_6287);
xnor U9269 (N_9269,N_7655,N_7408);
or U9270 (N_9270,N_7836,N_7420);
nand U9271 (N_9271,N_7273,N_6894);
nor U9272 (N_9272,N_6604,N_6996);
or U9273 (N_9273,N_6704,N_7395);
or U9274 (N_9274,N_7264,N_6631);
or U9275 (N_9275,N_6115,N_6957);
and U9276 (N_9276,N_6082,N_6583);
nand U9277 (N_9277,N_6764,N_6227);
and U9278 (N_9278,N_7337,N_7845);
nor U9279 (N_9279,N_6841,N_6750);
and U9280 (N_9280,N_7053,N_7464);
or U9281 (N_9281,N_7115,N_7852);
nand U9282 (N_9282,N_6378,N_6133);
nor U9283 (N_9283,N_7006,N_6148);
and U9284 (N_9284,N_7657,N_7409);
nor U9285 (N_9285,N_7999,N_6816);
nand U9286 (N_9286,N_7576,N_7215);
or U9287 (N_9287,N_7633,N_6673);
nor U9288 (N_9288,N_6517,N_6927);
nor U9289 (N_9289,N_7102,N_6949);
nor U9290 (N_9290,N_6273,N_7781);
xor U9291 (N_9291,N_6066,N_7498);
nor U9292 (N_9292,N_7738,N_6549);
and U9293 (N_9293,N_7365,N_7145);
or U9294 (N_9294,N_7966,N_6468);
nand U9295 (N_9295,N_6334,N_6350);
or U9296 (N_9296,N_7352,N_7130);
xnor U9297 (N_9297,N_7524,N_7514);
and U9298 (N_9298,N_7597,N_6660);
and U9299 (N_9299,N_6151,N_7431);
or U9300 (N_9300,N_6637,N_6682);
or U9301 (N_9301,N_7062,N_6490);
and U9302 (N_9302,N_7767,N_7187);
or U9303 (N_9303,N_6591,N_6287);
nand U9304 (N_9304,N_7880,N_7431);
nand U9305 (N_9305,N_6168,N_6017);
or U9306 (N_9306,N_6001,N_6157);
or U9307 (N_9307,N_6366,N_7833);
and U9308 (N_9308,N_7460,N_6685);
nor U9309 (N_9309,N_6150,N_6402);
or U9310 (N_9310,N_6649,N_7459);
and U9311 (N_9311,N_6009,N_6395);
or U9312 (N_9312,N_6561,N_7661);
nand U9313 (N_9313,N_7120,N_6605);
nand U9314 (N_9314,N_6437,N_7735);
nand U9315 (N_9315,N_7098,N_6310);
nand U9316 (N_9316,N_7593,N_7139);
or U9317 (N_9317,N_7918,N_6448);
nor U9318 (N_9318,N_7299,N_7344);
nand U9319 (N_9319,N_7323,N_7200);
nor U9320 (N_9320,N_6325,N_6854);
nand U9321 (N_9321,N_7951,N_6438);
or U9322 (N_9322,N_7755,N_7650);
xnor U9323 (N_9323,N_7501,N_7734);
xor U9324 (N_9324,N_6121,N_6548);
or U9325 (N_9325,N_7814,N_6621);
or U9326 (N_9326,N_7255,N_6881);
nor U9327 (N_9327,N_6516,N_7629);
xnor U9328 (N_9328,N_7437,N_7626);
nor U9329 (N_9329,N_6542,N_7524);
nor U9330 (N_9330,N_7825,N_7817);
or U9331 (N_9331,N_7549,N_7327);
nor U9332 (N_9332,N_7968,N_7641);
nand U9333 (N_9333,N_6980,N_7712);
or U9334 (N_9334,N_7846,N_7697);
nand U9335 (N_9335,N_6634,N_7386);
xor U9336 (N_9336,N_6242,N_6801);
or U9337 (N_9337,N_7222,N_7585);
or U9338 (N_9338,N_6012,N_6711);
nor U9339 (N_9339,N_7320,N_6076);
xor U9340 (N_9340,N_6960,N_6030);
or U9341 (N_9341,N_7046,N_6299);
nor U9342 (N_9342,N_7227,N_6823);
xnor U9343 (N_9343,N_6394,N_7507);
nor U9344 (N_9344,N_6556,N_6594);
or U9345 (N_9345,N_6770,N_7289);
nand U9346 (N_9346,N_6137,N_7298);
or U9347 (N_9347,N_6349,N_6317);
or U9348 (N_9348,N_7041,N_6969);
nor U9349 (N_9349,N_7245,N_6519);
nor U9350 (N_9350,N_7896,N_7358);
or U9351 (N_9351,N_7020,N_6823);
and U9352 (N_9352,N_6592,N_7726);
and U9353 (N_9353,N_6703,N_6002);
or U9354 (N_9354,N_6252,N_6460);
and U9355 (N_9355,N_7750,N_6240);
xnor U9356 (N_9356,N_7822,N_6679);
nand U9357 (N_9357,N_6318,N_6390);
nor U9358 (N_9358,N_7546,N_6882);
and U9359 (N_9359,N_6299,N_7202);
nor U9360 (N_9360,N_6065,N_7511);
or U9361 (N_9361,N_7957,N_6955);
and U9362 (N_9362,N_6208,N_6246);
nand U9363 (N_9363,N_7541,N_6774);
or U9364 (N_9364,N_6145,N_6892);
or U9365 (N_9365,N_6372,N_7737);
nand U9366 (N_9366,N_6887,N_7778);
and U9367 (N_9367,N_7645,N_6231);
nand U9368 (N_9368,N_7314,N_7951);
nand U9369 (N_9369,N_6669,N_7184);
or U9370 (N_9370,N_7651,N_6748);
and U9371 (N_9371,N_6061,N_6985);
and U9372 (N_9372,N_6538,N_6748);
and U9373 (N_9373,N_6731,N_6227);
xnor U9374 (N_9374,N_7821,N_6567);
or U9375 (N_9375,N_7626,N_6608);
nand U9376 (N_9376,N_7960,N_7479);
nand U9377 (N_9377,N_7780,N_6111);
and U9378 (N_9378,N_7469,N_6801);
and U9379 (N_9379,N_7168,N_7312);
or U9380 (N_9380,N_6145,N_7824);
or U9381 (N_9381,N_7245,N_7612);
nor U9382 (N_9382,N_6422,N_7512);
or U9383 (N_9383,N_7629,N_6229);
or U9384 (N_9384,N_7466,N_6820);
nand U9385 (N_9385,N_6116,N_6776);
nor U9386 (N_9386,N_7672,N_7067);
nor U9387 (N_9387,N_7360,N_6385);
or U9388 (N_9388,N_6873,N_6995);
nor U9389 (N_9389,N_6325,N_7568);
or U9390 (N_9390,N_7071,N_7310);
nand U9391 (N_9391,N_7473,N_7714);
xnor U9392 (N_9392,N_7006,N_6964);
nor U9393 (N_9393,N_6148,N_6030);
or U9394 (N_9394,N_6354,N_6631);
or U9395 (N_9395,N_6923,N_6253);
and U9396 (N_9396,N_6846,N_6185);
xnor U9397 (N_9397,N_6322,N_6168);
nor U9398 (N_9398,N_6635,N_7776);
and U9399 (N_9399,N_6144,N_6914);
or U9400 (N_9400,N_6084,N_6351);
nor U9401 (N_9401,N_7890,N_7868);
xnor U9402 (N_9402,N_6032,N_6832);
or U9403 (N_9403,N_7964,N_7772);
nor U9404 (N_9404,N_7669,N_7556);
nor U9405 (N_9405,N_7804,N_6948);
nand U9406 (N_9406,N_7348,N_7893);
or U9407 (N_9407,N_6793,N_7713);
and U9408 (N_9408,N_6268,N_6273);
nor U9409 (N_9409,N_6222,N_6607);
xor U9410 (N_9410,N_7319,N_7624);
or U9411 (N_9411,N_7847,N_7232);
nand U9412 (N_9412,N_6283,N_6772);
nand U9413 (N_9413,N_6250,N_7104);
nor U9414 (N_9414,N_7058,N_6364);
nor U9415 (N_9415,N_7919,N_6023);
nand U9416 (N_9416,N_6975,N_7133);
nand U9417 (N_9417,N_7838,N_7160);
or U9418 (N_9418,N_6378,N_7152);
nand U9419 (N_9419,N_6683,N_7069);
nand U9420 (N_9420,N_7346,N_7345);
xor U9421 (N_9421,N_7129,N_7948);
nor U9422 (N_9422,N_6661,N_7431);
nor U9423 (N_9423,N_6249,N_7096);
or U9424 (N_9424,N_7349,N_6469);
or U9425 (N_9425,N_6154,N_6290);
nand U9426 (N_9426,N_6179,N_7593);
nor U9427 (N_9427,N_6347,N_7086);
and U9428 (N_9428,N_7088,N_7515);
and U9429 (N_9429,N_6175,N_7658);
nand U9430 (N_9430,N_7538,N_7607);
and U9431 (N_9431,N_6504,N_6721);
and U9432 (N_9432,N_7387,N_6787);
nor U9433 (N_9433,N_7213,N_7063);
or U9434 (N_9434,N_6553,N_7612);
and U9435 (N_9435,N_6879,N_7659);
and U9436 (N_9436,N_6441,N_6579);
nand U9437 (N_9437,N_6827,N_6924);
and U9438 (N_9438,N_7576,N_6378);
or U9439 (N_9439,N_6211,N_6151);
and U9440 (N_9440,N_7991,N_7463);
nor U9441 (N_9441,N_7716,N_7213);
or U9442 (N_9442,N_7715,N_6577);
nand U9443 (N_9443,N_7189,N_6682);
nand U9444 (N_9444,N_7156,N_7889);
xnor U9445 (N_9445,N_6560,N_6066);
nand U9446 (N_9446,N_6145,N_7658);
or U9447 (N_9447,N_6279,N_7701);
xnor U9448 (N_9448,N_7734,N_7503);
and U9449 (N_9449,N_6732,N_6830);
or U9450 (N_9450,N_6861,N_6678);
nand U9451 (N_9451,N_7708,N_6139);
or U9452 (N_9452,N_7240,N_7393);
and U9453 (N_9453,N_7325,N_7127);
nand U9454 (N_9454,N_7658,N_6779);
nand U9455 (N_9455,N_7424,N_6446);
xor U9456 (N_9456,N_6278,N_6683);
or U9457 (N_9457,N_6510,N_6131);
nor U9458 (N_9458,N_6591,N_7260);
nand U9459 (N_9459,N_7919,N_7441);
or U9460 (N_9460,N_6700,N_7192);
nand U9461 (N_9461,N_7764,N_7621);
nand U9462 (N_9462,N_6335,N_7208);
or U9463 (N_9463,N_7382,N_6886);
nand U9464 (N_9464,N_7321,N_7686);
and U9465 (N_9465,N_6490,N_7257);
nor U9466 (N_9466,N_7576,N_6623);
and U9467 (N_9467,N_7797,N_6492);
or U9468 (N_9468,N_7016,N_6395);
xor U9469 (N_9469,N_6816,N_7639);
nor U9470 (N_9470,N_7614,N_6954);
or U9471 (N_9471,N_7368,N_7118);
nor U9472 (N_9472,N_7650,N_7252);
and U9473 (N_9473,N_7303,N_7926);
xor U9474 (N_9474,N_7995,N_6090);
nand U9475 (N_9475,N_7982,N_7920);
xnor U9476 (N_9476,N_6066,N_7772);
nand U9477 (N_9477,N_7025,N_7006);
nand U9478 (N_9478,N_6238,N_6290);
xor U9479 (N_9479,N_6881,N_7442);
nor U9480 (N_9480,N_6375,N_7956);
or U9481 (N_9481,N_7771,N_6516);
or U9482 (N_9482,N_7066,N_7877);
and U9483 (N_9483,N_6114,N_6777);
and U9484 (N_9484,N_6524,N_6795);
nand U9485 (N_9485,N_7304,N_7329);
nand U9486 (N_9486,N_6308,N_6469);
nand U9487 (N_9487,N_7816,N_6220);
and U9488 (N_9488,N_7727,N_7053);
nor U9489 (N_9489,N_6660,N_6115);
nor U9490 (N_9490,N_7167,N_7246);
nor U9491 (N_9491,N_6900,N_7125);
nand U9492 (N_9492,N_6832,N_7226);
or U9493 (N_9493,N_7729,N_6430);
nor U9494 (N_9494,N_6768,N_6605);
or U9495 (N_9495,N_7275,N_7397);
nor U9496 (N_9496,N_6315,N_7685);
and U9497 (N_9497,N_7976,N_6501);
nor U9498 (N_9498,N_6008,N_7035);
and U9499 (N_9499,N_7488,N_6508);
or U9500 (N_9500,N_6192,N_6198);
or U9501 (N_9501,N_7494,N_7595);
nand U9502 (N_9502,N_6125,N_6449);
xnor U9503 (N_9503,N_6779,N_6365);
xor U9504 (N_9504,N_7942,N_6274);
and U9505 (N_9505,N_7489,N_7039);
nor U9506 (N_9506,N_7537,N_7867);
xor U9507 (N_9507,N_7742,N_6209);
nor U9508 (N_9508,N_7250,N_7330);
or U9509 (N_9509,N_6487,N_7810);
nor U9510 (N_9510,N_6787,N_6100);
nor U9511 (N_9511,N_6409,N_7010);
and U9512 (N_9512,N_7221,N_6726);
and U9513 (N_9513,N_7463,N_6767);
nand U9514 (N_9514,N_6847,N_7859);
nand U9515 (N_9515,N_6010,N_6486);
nor U9516 (N_9516,N_6070,N_6833);
nand U9517 (N_9517,N_7259,N_6656);
and U9518 (N_9518,N_7148,N_7624);
nor U9519 (N_9519,N_6918,N_7144);
and U9520 (N_9520,N_7042,N_7162);
nor U9521 (N_9521,N_6814,N_6133);
nor U9522 (N_9522,N_6163,N_7789);
nand U9523 (N_9523,N_6628,N_6137);
xnor U9524 (N_9524,N_7210,N_7343);
nand U9525 (N_9525,N_7017,N_6061);
and U9526 (N_9526,N_6127,N_6051);
nand U9527 (N_9527,N_6496,N_7382);
nor U9528 (N_9528,N_7132,N_6255);
nand U9529 (N_9529,N_7242,N_6647);
or U9530 (N_9530,N_6967,N_7932);
and U9531 (N_9531,N_6334,N_7606);
and U9532 (N_9532,N_6037,N_6205);
and U9533 (N_9533,N_7904,N_7724);
or U9534 (N_9534,N_7106,N_6841);
nand U9535 (N_9535,N_7613,N_6614);
nand U9536 (N_9536,N_6571,N_6209);
or U9537 (N_9537,N_6184,N_7912);
nor U9538 (N_9538,N_6881,N_6916);
nor U9539 (N_9539,N_6265,N_6735);
or U9540 (N_9540,N_7965,N_7614);
nor U9541 (N_9541,N_7760,N_7821);
nor U9542 (N_9542,N_6170,N_6614);
nor U9543 (N_9543,N_7171,N_7323);
and U9544 (N_9544,N_7231,N_6280);
xnor U9545 (N_9545,N_6280,N_6311);
or U9546 (N_9546,N_6725,N_7042);
xor U9547 (N_9547,N_6761,N_7128);
and U9548 (N_9548,N_7682,N_7715);
nand U9549 (N_9549,N_7588,N_7000);
or U9550 (N_9550,N_7779,N_6433);
xor U9551 (N_9551,N_7912,N_7771);
nand U9552 (N_9552,N_7207,N_7542);
and U9553 (N_9553,N_7101,N_6426);
or U9554 (N_9554,N_7137,N_7139);
nand U9555 (N_9555,N_7482,N_7779);
nor U9556 (N_9556,N_7590,N_6536);
nor U9557 (N_9557,N_6193,N_7782);
xnor U9558 (N_9558,N_6302,N_6932);
nand U9559 (N_9559,N_6025,N_7004);
nor U9560 (N_9560,N_7287,N_7543);
nor U9561 (N_9561,N_6110,N_6100);
nor U9562 (N_9562,N_7885,N_6358);
and U9563 (N_9563,N_6991,N_7749);
nor U9564 (N_9564,N_7107,N_7336);
nor U9565 (N_9565,N_6397,N_7353);
xor U9566 (N_9566,N_6466,N_7768);
nand U9567 (N_9567,N_6886,N_6994);
or U9568 (N_9568,N_7900,N_6017);
and U9569 (N_9569,N_6939,N_6718);
nand U9570 (N_9570,N_7806,N_7769);
and U9571 (N_9571,N_7009,N_7191);
or U9572 (N_9572,N_7551,N_7558);
or U9573 (N_9573,N_7939,N_6343);
nand U9574 (N_9574,N_7242,N_6815);
or U9575 (N_9575,N_7306,N_6604);
or U9576 (N_9576,N_6418,N_6694);
nor U9577 (N_9577,N_6067,N_7172);
nor U9578 (N_9578,N_7467,N_6215);
and U9579 (N_9579,N_6210,N_7185);
and U9580 (N_9580,N_7386,N_6278);
and U9581 (N_9581,N_6110,N_7037);
and U9582 (N_9582,N_6321,N_7615);
and U9583 (N_9583,N_6643,N_7824);
xnor U9584 (N_9584,N_6577,N_6623);
nand U9585 (N_9585,N_7894,N_6050);
and U9586 (N_9586,N_6002,N_7774);
or U9587 (N_9587,N_6192,N_7109);
or U9588 (N_9588,N_6780,N_7165);
nand U9589 (N_9589,N_7667,N_6806);
nor U9590 (N_9590,N_6393,N_6423);
or U9591 (N_9591,N_7581,N_7854);
nor U9592 (N_9592,N_7183,N_7432);
xor U9593 (N_9593,N_6547,N_7145);
nand U9594 (N_9594,N_6509,N_6162);
or U9595 (N_9595,N_6589,N_7902);
xor U9596 (N_9596,N_7577,N_7913);
nor U9597 (N_9597,N_7478,N_6027);
and U9598 (N_9598,N_6538,N_6461);
or U9599 (N_9599,N_7795,N_6823);
or U9600 (N_9600,N_7781,N_7896);
nor U9601 (N_9601,N_6318,N_7773);
nand U9602 (N_9602,N_6208,N_6146);
and U9603 (N_9603,N_7094,N_6564);
and U9604 (N_9604,N_6223,N_6258);
nor U9605 (N_9605,N_6138,N_6849);
nand U9606 (N_9606,N_6871,N_6976);
and U9607 (N_9607,N_6694,N_7452);
and U9608 (N_9608,N_7023,N_7929);
nand U9609 (N_9609,N_7883,N_7585);
or U9610 (N_9610,N_6031,N_6398);
or U9611 (N_9611,N_7405,N_6448);
nor U9612 (N_9612,N_6998,N_7776);
and U9613 (N_9613,N_6697,N_7228);
nor U9614 (N_9614,N_6210,N_6510);
nor U9615 (N_9615,N_7595,N_6854);
xnor U9616 (N_9616,N_7047,N_6769);
and U9617 (N_9617,N_7311,N_6510);
and U9618 (N_9618,N_7308,N_6519);
and U9619 (N_9619,N_6035,N_6697);
nand U9620 (N_9620,N_7821,N_7751);
and U9621 (N_9621,N_7842,N_6817);
and U9622 (N_9622,N_7231,N_7407);
or U9623 (N_9623,N_7297,N_7040);
and U9624 (N_9624,N_7870,N_6308);
nand U9625 (N_9625,N_7601,N_7523);
nor U9626 (N_9626,N_7522,N_6321);
or U9627 (N_9627,N_7202,N_7006);
or U9628 (N_9628,N_6412,N_7884);
xnor U9629 (N_9629,N_7290,N_7001);
and U9630 (N_9630,N_6964,N_6366);
nand U9631 (N_9631,N_7503,N_6174);
xnor U9632 (N_9632,N_7567,N_7356);
xor U9633 (N_9633,N_7381,N_6582);
and U9634 (N_9634,N_7723,N_6073);
nand U9635 (N_9635,N_7287,N_7895);
xnor U9636 (N_9636,N_7161,N_7589);
nand U9637 (N_9637,N_6598,N_7525);
nor U9638 (N_9638,N_6918,N_7661);
and U9639 (N_9639,N_6561,N_6048);
or U9640 (N_9640,N_7750,N_6528);
or U9641 (N_9641,N_7243,N_6117);
and U9642 (N_9642,N_6055,N_7930);
or U9643 (N_9643,N_7084,N_7070);
and U9644 (N_9644,N_7494,N_6942);
nor U9645 (N_9645,N_6151,N_6132);
nand U9646 (N_9646,N_6550,N_6718);
and U9647 (N_9647,N_6776,N_6353);
or U9648 (N_9648,N_6299,N_6619);
and U9649 (N_9649,N_6538,N_7178);
nor U9650 (N_9650,N_6932,N_6687);
xnor U9651 (N_9651,N_6081,N_6143);
or U9652 (N_9652,N_6823,N_6469);
nand U9653 (N_9653,N_7890,N_6917);
nor U9654 (N_9654,N_6350,N_6272);
xnor U9655 (N_9655,N_7642,N_6836);
xor U9656 (N_9656,N_7276,N_7857);
nor U9657 (N_9657,N_6956,N_6892);
and U9658 (N_9658,N_7340,N_6913);
nand U9659 (N_9659,N_6664,N_6949);
nor U9660 (N_9660,N_7827,N_6581);
and U9661 (N_9661,N_6106,N_7675);
nor U9662 (N_9662,N_7145,N_7919);
nand U9663 (N_9663,N_7475,N_7260);
xnor U9664 (N_9664,N_6767,N_7648);
nand U9665 (N_9665,N_7400,N_6245);
or U9666 (N_9666,N_7425,N_6702);
or U9667 (N_9667,N_6627,N_6049);
nand U9668 (N_9668,N_6309,N_7811);
and U9669 (N_9669,N_6605,N_7908);
or U9670 (N_9670,N_7136,N_7032);
or U9671 (N_9671,N_6863,N_6825);
or U9672 (N_9672,N_6403,N_7681);
nor U9673 (N_9673,N_7119,N_6869);
and U9674 (N_9674,N_6847,N_7680);
nor U9675 (N_9675,N_7790,N_6107);
or U9676 (N_9676,N_6773,N_7221);
and U9677 (N_9677,N_6351,N_6620);
nand U9678 (N_9678,N_7488,N_6782);
xor U9679 (N_9679,N_6594,N_6602);
nand U9680 (N_9680,N_7628,N_6384);
and U9681 (N_9681,N_6638,N_7451);
xnor U9682 (N_9682,N_7937,N_6134);
nor U9683 (N_9683,N_6810,N_6296);
nand U9684 (N_9684,N_6919,N_6222);
and U9685 (N_9685,N_6854,N_6133);
xnor U9686 (N_9686,N_6856,N_7070);
and U9687 (N_9687,N_7385,N_7175);
nand U9688 (N_9688,N_7813,N_7118);
nand U9689 (N_9689,N_7113,N_7506);
and U9690 (N_9690,N_7448,N_6655);
nor U9691 (N_9691,N_7929,N_7984);
or U9692 (N_9692,N_7002,N_6252);
or U9693 (N_9693,N_6377,N_6125);
or U9694 (N_9694,N_6029,N_7432);
and U9695 (N_9695,N_7781,N_7876);
nand U9696 (N_9696,N_7949,N_7058);
or U9697 (N_9697,N_6054,N_6502);
and U9698 (N_9698,N_6558,N_6077);
or U9699 (N_9699,N_6308,N_7742);
and U9700 (N_9700,N_6741,N_6040);
xnor U9701 (N_9701,N_7702,N_6524);
or U9702 (N_9702,N_6405,N_7231);
and U9703 (N_9703,N_7628,N_7448);
nand U9704 (N_9704,N_7136,N_7663);
nor U9705 (N_9705,N_6908,N_6451);
nor U9706 (N_9706,N_6543,N_7901);
nor U9707 (N_9707,N_6199,N_6848);
nand U9708 (N_9708,N_6582,N_6603);
nor U9709 (N_9709,N_7702,N_6752);
nand U9710 (N_9710,N_6716,N_7655);
nor U9711 (N_9711,N_7010,N_6953);
xor U9712 (N_9712,N_6522,N_7206);
nor U9713 (N_9713,N_7464,N_6418);
and U9714 (N_9714,N_7089,N_6150);
or U9715 (N_9715,N_6933,N_7531);
nand U9716 (N_9716,N_7178,N_7026);
xnor U9717 (N_9717,N_6522,N_6121);
nand U9718 (N_9718,N_6507,N_6709);
and U9719 (N_9719,N_7181,N_7489);
nand U9720 (N_9720,N_7758,N_6719);
nand U9721 (N_9721,N_7893,N_6921);
or U9722 (N_9722,N_7183,N_6252);
nand U9723 (N_9723,N_7369,N_6073);
nor U9724 (N_9724,N_7892,N_7451);
or U9725 (N_9725,N_6885,N_6399);
or U9726 (N_9726,N_7358,N_7969);
nand U9727 (N_9727,N_7095,N_6463);
nor U9728 (N_9728,N_6951,N_7726);
nor U9729 (N_9729,N_7822,N_6342);
or U9730 (N_9730,N_7251,N_6179);
nand U9731 (N_9731,N_6382,N_6716);
xnor U9732 (N_9732,N_6083,N_6414);
or U9733 (N_9733,N_6031,N_6197);
and U9734 (N_9734,N_6749,N_6493);
or U9735 (N_9735,N_6206,N_6536);
or U9736 (N_9736,N_7935,N_7650);
and U9737 (N_9737,N_6692,N_7351);
xor U9738 (N_9738,N_7990,N_6778);
or U9739 (N_9739,N_7120,N_7538);
nor U9740 (N_9740,N_7259,N_7911);
nor U9741 (N_9741,N_6295,N_7844);
or U9742 (N_9742,N_6796,N_6024);
nand U9743 (N_9743,N_7243,N_6272);
or U9744 (N_9744,N_6759,N_6643);
and U9745 (N_9745,N_7222,N_7114);
or U9746 (N_9746,N_6315,N_7764);
nor U9747 (N_9747,N_6975,N_7494);
or U9748 (N_9748,N_6181,N_7587);
and U9749 (N_9749,N_6327,N_6130);
nor U9750 (N_9750,N_7440,N_7537);
nand U9751 (N_9751,N_6218,N_6820);
or U9752 (N_9752,N_7056,N_7011);
nand U9753 (N_9753,N_7080,N_6930);
nand U9754 (N_9754,N_7944,N_7488);
or U9755 (N_9755,N_7844,N_7305);
nand U9756 (N_9756,N_7097,N_6273);
nor U9757 (N_9757,N_7566,N_7785);
nand U9758 (N_9758,N_6216,N_7999);
nand U9759 (N_9759,N_7995,N_6173);
xnor U9760 (N_9760,N_7685,N_7190);
and U9761 (N_9761,N_7898,N_7079);
xnor U9762 (N_9762,N_6346,N_7623);
nand U9763 (N_9763,N_7502,N_6015);
and U9764 (N_9764,N_7021,N_6758);
or U9765 (N_9765,N_6421,N_6255);
and U9766 (N_9766,N_6619,N_6727);
and U9767 (N_9767,N_7134,N_7627);
nand U9768 (N_9768,N_7683,N_6749);
and U9769 (N_9769,N_6322,N_7445);
and U9770 (N_9770,N_7040,N_7198);
or U9771 (N_9771,N_6152,N_6532);
and U9772 (N_9772,N_7007,N_6580);
or U9773 (N_9773,N_7568,N_6108);
or U9774 (N_9774,N_6468,N_7048);
or U9775 (N_9775,N_7604,N_7459);
and U9776 (N_9776,N_6863,N_7195);
or U9777 (N_9777,N_6761,N_7125);
xnor U9778 (N_9778,N_7049,N_7318);
or U9779 (N_9779,N_7915,N_7534);
or U9780 (N_9780,N_7780,N_7969);
nand U9781 (N_9781,N_7042,N_6537);
nor U9782 (N_9782,N_7412,N_6672);
xnor U9783 (N_9783,N_6803,N_6650);
nand U9784 (N_9784,N_6604,N_7627);
or U9785 (N_9785,N_7005,N_7022);
or U9786 (N_9786,N_6372,N_7257);
or U9787 (N_9787,N_6704,N_7128);
or U9788 (N_9788,N_6595,N_7519);
and U9789 (N_9789,N_7311,N_7860);
and U9790 (N_9790,N_6556,N_7359);
nand U9791 (N_9791,N_6867,N_6010);
and U9792 (N_9792,N_7070,N_7921);
nor U9793 (N_9793,N_6785,N_7391);
and U9794 (N_9794,N_7438,N_7372);
nand U9795 (N_9795,N_7836,N_7531);
xor U9796 (N_9796,N_6701,N_7123);
or U9797 (N_9797,N_6278,N_6203);
nand U9798 (N_9798,N_6138,N_7690);
or U9799 (N_9799,N_6331,N_7777);
nand U9800 (N_9800,N_7856,N_6239);
nor U9801 (N_9801,N_6662,N_7515);
and U9802 (N_9802,N_7000,N_7665);
or U9803 (N_9803,N_7237,N_7148);
nor U9804 (N_9804,N_7735,N_7320);
and U9805 (N_9805,N_7276,N_6456);
nand U9806 (N_9806,N_6328,N_6534);
or U9807 (N_9807,N_7191,N_6100);
or U9808 (N_9808,N_6777,N_6606);
nor U9809 (N_9809,N_6161,N_6182);
and U9810 (N_9810,N_7768,N_6021);
and U9811 (N_9811,N_7282,N_7345);
and U9812 (N_9812,N_7207,N_6240);
nor U9813 (N_9813,N_6613,N_6953);
nand U9814 (N_9814,N_6128,N_6146);
or U9815 (N_9815,N_6765,N_7505);
or U9816 (N_9816,N_7368,N_7162);
nand U9817 (N_9817,N_7732,N_6883);
nand U9818 (N_9818,N_7565,N_7540);
nand U9819 (N_9819,N_7637,N_7449);
or U9820 (N_9820,N_6967,N_7012);
nor U9821 (N_9821,N_7707,N_7163);
nor U9822 (N_9822,N_7729,N_7259);
and U9823 (N_9823,N_7261,N_7080);
nand U9824 (N_9824,N_7174,N_6443);
nand U9825 (N_9825,N_6970,N_7242);
xor U9826 (N_9826,N_6593,N_7227);
and U9827 (N_9827,N_7576,N_7219);
and U9828 (N_9828,N_7150,N_7280);
nand U9829 (N_9829,N_7491,N_7988);
or U9830 (N_9830,N_6829,N_7708);
and U9831 (N_9831,N_6254,N_6559);
nand U9832 (N_9832,N_7921,N_7808);
or U9833 (N_9833,N_7266,N_6151);
nor U9834 (N_9834,N_7003,N_6455);
nor U9835 (N_9835,N_6374,N_7971);
and U9836 (N_9836,N_6102,N_7939);
or U9837 (N_9837,N_6990,N_7634);
nand U9838 (N_9838,N_7972,N_7189);
or U9839 (N_9839,N_7146,N_7268);
nor U9840 (N_9840,N_6368,N_7456);
or U9841 (N_9841,N_6192,N_7870);
nand U9842 (N_9842,N_6094,N_6826);
nand U9843 (N_9843,N_6617,N_6407);
and U9844 (N_9844,N_7570,N_6032);
xnor U9845 (N_9845,N_6322,N_6795);
nor U9846 (N_9846,N_6904,N_6372);
and U9847 (N_9847,N_6288,N_7220);
or U9848 (N_9848,N_6296,N_7586);
or U9849 (N_9849,N_6586,N_7809);
nand U9850 (N_9850,N_7071,N_6562);
nand U9851 (N_9851,N_7716,N_6542);
nand U9852 (N_9852,N_6918,N_6426);
nand U9853 (N_9853,N_7003,N_6265);
and U9854 (N_9854,N_7893,N_6753);
and U9855 (N_9855,N_7466,N_6570);
and U9856 (N_9856,N_6483,N_6698);
nand U9857 (N_9857,N_7241,N_6530);
and U9858 (N_9858,N_6535,N_7018);
nand U9859 (N_9859,N_6733,N_6237);
nand U9860 (N_9860,N_6546,N_6245);
nand U9861 (N_9861,N_7208,N_7933);
nor U9862 (N_9862,N_6916,N_7548);
xor U9863 (N_9863,N_7505,N_6223);
or U9864 (N_9864,N_7000,N_6236);
or U9865 (N_9865,N_7751,N_6131);
nor U9866 (N_9866,N_6697,N_6780);
and U9867 (N_9867,N_6815,N_7125);
nor U9868 (N_9868,N_7822,N_7187);
or U9869 (N_9869,N_7501,N_7084);
xor U9870 (N_9870,N_7375,N_7609);
or U9871 (N_9871,N_6198,N_6159);
nand U9872 (N_9872,N_6423,N_7090);
nand U9873 (N_9873,N_6929,N_7368);
nor U9874 (N_9874,N_6663,N_6840);
nor U9875 (N_9875,N_6167,N_7411);
nor U9876 (N_9876,N_6266,N_7825);
and U9877 (N_9877,N_7048,N_7738);
nand U9878 (N_9878,N_6378,N_6577);
and U9879 (N_9879,N_7481,N_6802);
or U9880 (N_9880,N_7755,N_6035);
nand U9881 (N_9881,N_7458,N_7342);
or U9882 (N_9882,N_6376,N_6124);
or U9883 (N_9883,N_6018,N_7946);
and U9884 (N_9884,N_7576,N_6484);
xor U9885 (N_9885,N_6691,N_7539);
xor U9886 (N_9886,N_7597,N_7446);
or U9887 (N_9887,N_6296,N_6593);
nor U9888 (N_9888,N_7292,N_6249);
xor U9889 (N_9889,N_7201,N_7570);
nand U9890 (N_9890,N_6437,N_6738);
nand U9891 (N_9891,N_7921,N_7018);
nand U9892 (N_9892,N_7791,N_6881);
nor U9893 (N_9893,N_6978,N_7435);
nor U9894 (N_9894,N_7138,N_6939);
or U9895 (N_9895,N_6708,N_7571);
or U9896 (N_9896,N_6665,N_7536);
nand U9897 (N_9897,N_7910,N_6817);
xnor U9898 (N_9898,N_7885,N_7336);
and U9899 (N_9899,N_6759,N_7719);
nor U9900 (N_9900,N_6517,N_6568);
nand U9901 (N_9901,N_6446,N_6140);
or U9902 (N_9902,N_7692,N_7355);
xnor U9903 (N_9903,N_7487,N_6448);
nor U9904 (N_9904,N_6849,N_6180);
nor U9905 (N_9905,N_6308,N_6243);
and U9906 (N_9906,N_6625,N_7775);
or U9907 (N_9907,N_6580,N_6563);
nand U9908 (N_9908,N_6245,N_7965);
nand U9909 (N_9909,N_6244,N_7418);
and U9910 (N_9910,N_7268,N_6864);
or U9911 (N_9911,N_6363,N_7899);
nand U9912 (N_9912,N_6688,N_7986);
nor U9913 (N_9913,N_6766,N_7979);
and U9914 (N_9914,N_6629,N_6901);
nor U9915 (N_9915,N_6176,N_6115);
nand U9916 (N_9916,N_7832,N_7651);
nand U9917 (N_9917,N_6741,N_7950);
nor U9918 (N_9918,N_6307,N_6187);
nor U9919 (N_9919,N_7554,N_7050);
nor U9920 (N_9920,N_6796,N_7526);
and U9921 (N_9921,N_7244,N_6222);
xnor U9922 (N_9922,N_7734,N_7952);
nand U9923 (N_9923,N_7465,N_7170);
nor U9924 (N_9924,N_7739,N_6522);
and U9925 (N_9925,N_6252,N_6844);
and U9926 (N_9926,N_6832,N_7723);
or U9927 (N_9927,N_6548,N_7866);
and U9928 (N_9928,N_6696,N_6191);
xor U9929 (N_9929,N_7776,N_7866);
nor U9930 (N_9930,N_7762,N_7113);
nand U9931 (N_9931,N_7439,N_7126);
nand U9932 (N_9932,N_6218,N_7117);
xor U9933 (N_9933,N_7983,N_6951);
or U9934 (N_9934,N_6509,N_6809);
and U9935 (N_9935,N_7134,N_7978);
and U9936 (N_9936,N_6571,N_6396);
and U9937 (N_9937,N_6521,N_7407);
or U9938 (N_9938,N_6197,N_7127);
or U9939 (N_9939,N_6139,N_6182);
and U9940 (N_9940,N_6777,N_6089);
nand U9941 (N_9941,N_7748,N_7962);
or U9942 (N_9942,N_6405,N_7926);
or U9943 (N_9943,N_7520,N_7154);
and U9944 (N_9944,N_7450,N_6513);
and U9945 (N_9945,N_6281,N_6831);
or U9946 (N_9946,N_7423,N_7483);
or U9947 (N_9947,N_7978,N_7890);
nand U9948 (N_9948,N_6224,N_6500);
nand U9949 (N_9949,N_6150,N_6182);
nor U9950 (N_9950,N_6123,N_6528);
nand U9951 (N_9951,N_7209,N_7779);
or U9952 (N_9952,N_7366,N_6123);
or U9953 (N_9953,N_6944,N_7522);
nand U9954 (N_9954,N_6965,N_6796);
nand U9955 (N_9955,N_7049,N_6000);
or U9956 (N_9956,N_6582,N_6976);
xor U9957 (N_9957,N_7122,N_7155);
and U9958 (N_9958,N_7239,N_6104);
and U9959 (N_9959,N_6505,N_7652);
nor U9960 (N_9960,N_6501,N_7996);
xor U9961 (N_9961,N_7353,N_7375);
nor U9962 (N_9962,N_7116,N_6868);
xor U9963 (N_9963,N_6325,N_7726);
nor U9964 (N_9964,N_7230,N_7142);
nand U9965 (N_9965,N_6179,N_7933);
nor U9966 (N_9966,N_7974,N_6745);
and U9967 (N_9967,N_7426,N_7501);
and U9968 (N_9968,N_6137,N_7574);
nor U9969 (N_9969,N_6252,N_7498);
and U9970 (N_9970,N_7962,N_7671);
and U9971 (N_9971,N_7893,N_7232);
nand U9972 (N_9972,N_6693,N_7275);
or U9973 (N_9973,N_6834,N_7261);
xor U9974 (N_9974,N_7253,N_7191);
and U9975 (N_9975,N_7017,N_6244);
or U9976 (N_9976,N_7176,N_7754);
nand U9977 (N_9977,N_7953,N_6580);
nor U9978 (N_9978,N_7064,N_6961);
or U9979 (N_9979,N_6885,N_7331);
or U9980 (N_9980,N_6143,N_7298);
and U9981 (N_9981,N_7320,N_7930);
nand U9982 (N_9982,N_7469,N_7619);
and U9983 (N_9983,N_7542,N_7260);
nor U9984 (N_9984,N_7741,N_6988);
nor U9985 (N_9985,N_7611,N_7383);
nand U9986 (N_9986,N_6063,N_7397);
or U9987 (N_9987,N_7469,N_6611);
xnor U9988 (N_9988,N_7297,N_7906);
nor U9989 (N_9989,N_6926,N_7646);
nand U9990 (N_9990,N_6691,N_7347);
and U9991 (N_9991,N_7212,N_6345);
nand U9992 (N_9992,N_7216,N_7854);
or U9993 (N_9993,N_7419,N_6676);
and U9994 (N_9994,N_7983,N_6383);
and U9995 (N_9995,N_6166,N_7746);
nor U9996 (N_9996,N_6575,N_7714);
xor U9997 (N_9997,N_7268,N_7584);
nor U9998 (N_9998,N_6792,N_6368);
or U9999 (N_9999,N_7310,N_6404);
nand UO_0 (O_0,N_8107,N_8420);
and UO_1 (O_1,N_9716,N_8919);
or UO_2 (O_2,N_9555,N_8678);
or UO_3 (O_3,N_8576,N_8566);
nand UO_4 (O_4,N_8248,N_8859);
and UO_5 (O_5,N_9668,N_8251);
nand UO_6 (O_6,N_9418,N_9886);
nand UO_7 (O_7,N_8591,N_8256);
and UO_8 (O_8,N_9752,N_8060);
and UO_9 (O_9,N_8224,N_8374);
nand UO_10 (O_10,N_9049,N_8476);
and UO_11 (O_11,N_9657,N_8550);
nand UO_12 (O_12,N_9805,N_9816);
or UO_13 (O_13,N_8607,N_8118);
nand UO_14 (O_14,N_9496,N_8604);
nor UO_15 (O_15,N_8483,N_8429);
or UO_16 (O_16,N_8026,N_8069);
xor UO_17 (O_17,N_8117,N_8729);
nor UO_18 (O_18,N_8524,N_9952);
nor UO_19 (O_19,N_9377,N_9803);
xor UO_20 (O_20,N_8596,N_8095);
or UO_21 (O_21,N_8774,N_8580);
and UO_22 (O_22,N_9387,N_8275);
or UO_23 (O_23,N_8058,N_9264);
nor UO_24 (O_24,N_9055,N_9028);
and UO_25 (O_25,N_9380,N_8521);
nand UO_26 (O_26,N_9004,N_9990);
nand UO_27 (O_27,N_9212,N_9619);
nand UO_28 (O_28,N_9611,N_8219);
nand UO_29 (O_29,N_8985,N_8245);
nand UO_30 (O_30,N_9840,N_8048);
and UO_31 (O_31,N_9726,N_8862);
xnor UO_32 (O_32,N_9615,N_8939);
nor UO_33 (O_33,N_8489,N_9930);
and UO_34 (O_34,N_8254,N_9665);
nor UO_35 (O_35,N_8873,N_8883);
xor UO_36 (O_36,N_9591,N_8769);
nand UO_37 (O_37,N_8694,N_9642);
and UO_38 (O_38,N_9164,N_9355);
and UO_39 (O_39,N_8396,N_9104);
nor UO_40 (O_40,N_8974,N_9799);
xnor UO_41 (O_41,N_9117,N_8920);
or UO_42 (O_42,N_8361,N_8298);
xnor UO_43 (O_43,N_8595,N_9776);
or UO_44 (O_44,N_8104,N_8629);
xor UO_45 (O_45,N_9465,N_8031);
xor UO_46 (O_46,N_8153,N_9648);
nor UO_47 (O_47,N_9133,N_9181);
xnor UO_48 (O_48,N_8589,N_8053);
nor UO_49 (O_49,N_9997,N_8549);
xnor UO_50 (O_50,N_8913,N_8150);
nor UO_51 (O_51,N_8714,N_8705);
nor UO_52 (O_52,N_9834,N_8370);
or UO_53 (O_53,N_9519,N_8240);
and UO_54 (O_54,N_8141,N_9570);
or UO_55 (O_55,N_8309,N_8706);
and UO_56 (O_56,N_8916,N_9596);
and UO_57 (O_57,N_9787,N_8843);
xor UO_58 (O_58,N_8393,N_9281);
and UO_59 (O_59,N_9132,N_9372);
nor UO_60 (O_60,N_9206,N_8543);
nor UO_61 (O_61,N_8713,N_9824);
and UO_62 (O_62,N_8941,N_9622);
nor UO_63 (O_63,N_8501,N_9883);
or UO_64 (O_64,N_9548,N_9340);
nor UO_65 (O_65,N_8132,N_9289);
xnor UO_66 (O_66,N_8562,N_8269);
and UO_67 (O_67,N_9934,N_9987);
nand UO_68 (O_68,N_9124,N_8848);
and UO_69 (O_69,N_8431,N_9394);
and UO_70 (O_70,N_8316,N_9159);
nand UO_71 (O_71,N_9180,N_8575);
and UO_72 (O_72,N_9488,N_9178);
and UO_73 (O_73,N_8888,N_8894);
or UO_74 (O_74,N_9962,N_8295);
or UO_75 (O_75,N_8324,N_9533);
or UO_76 (O_76,N_9674,N_8367);
or UO_77 (O_77,N_8574,N_8340);
nor UO_78 (O_78,N_9551,N_8113);
or UO_79 (O_79,N_8745,N_9325);
nand UO_80 (O_80,N_8379,N_9298);
and UO_81 (O_81,N_9501,N_9107);
nand UO_82 (O_82,N_8433,N_8285);
or UO_83 (O_83,N_8034,N_9953);
nand UO_84 (O_84,N_9142,N_8636);
or UO_85 (O_85,N_9365,N_9587);
and UO_86 (O_86,N_8539,N_8164);
nor UO_87 (O_87,N_8086,N_8276);
and UO_88 (O_88,N_8992,N_8389);
nand UO_89 (O_89,N_8671,N_9924);
nand UO_90 (O_90,N_8481,N_9835);
and UO_91 (O_91,N_8668,N_8516);
xnor UO_92 (O_92,N_8001,N_9639);
and UO_93 (O_93,N_9530,N_9774);
xor UO_94 (O_94,N_8517,N_8651);
and UO_95 (O_95,N_9445,N_9867);
or UO_96 (O_96,N_8934,N_9228);
nor UO_97 (O_97,N_9306,N_9819);
and UO_98 (O_98,N_8151,N_9802);
or UO_99 (O_99,N_8626,N_9894);
and UO_100 (O_100,N_9236,N_8376);
nor UO_101 (O_101,N_9388,N_8014);
or UO_102 (O_102,N_9096,N_8447);
xnor UO_103 (O_103,N_8402,N_8868);
nor UO_104 (O_104,N_8812,N_8226);
nor UO_105 (O_105,N_9420,N_8124);
nand UO_106 (O_106,N_9994,N_9652);
or UO_107 (O_107,N_9021,N_9778);
nor UO_108 (O_108,N_8189,N_8453);
xnor UO_109 (O_109,N_9419,N_9862);
and UO_110 (O_110,N_8231,N_9019);
nand UO_111 (O_111,N_8710,N_9705);
or UO_112 (O_112,N_8695,N_9916);
nor UO_113 (O_113,N_8750,N_9368);
and UO_114 (O_114,N_8752,N_8892);
nor UO_115 (O_115,N_8753,N_9827);
nor UO_116 (O_116,N_9832,N_8593);
or UO_117 (O_117,N_9956,N_8464);
or UO_118 (O_118,N_8649,N_9771);
nor UO_119 (O_119,N_8147,N_9856);
and UO_120 (O_120,N_8454,N_9099);
and UO_121 (O_121,N_8565,N_9552);
nand UO_122 (O_122,N_9196,N_8239);
nand UO_123 (O_123,N_8907,N_8392);
and UO_124 (O_124,N_9669,N_8762);
nand UO_125 (O_125,N_9711,N_8040);
nor UO_126 (O_126,N_8866,N_9540);
nor UO_127 (O_127,N_8290,N_9877);
nand UO_128 (O_128,N_8732,N_8138);
or UO_129 (O_129,N_9579,N_8789);
and UO_130 (O_130,N_9853,N_9031);
nor UO_131 (O_131,N_9059,N_9979);
xnor UO_132 (O_132,N_9972,N_8469);
nor UO_133 (O_133,N_8146,N_9982);
or UO_134 (O_134,N_8620,N_8378);
nor UO_135 (O_135,N_9315,N_8200);
and UO_136 (O_136,N_8300,N_8704);
nand UO_137 (O_137,N_9123,N_9731);
and UO_138 (O_138,N_9506,N_8485);
nand UO_139 (O_139,N_8938,N_9135);
nor UO_140 (O_140,N_9350,N_8904);
xor UO_141 (O_141,N_9014,N_9201);
nor UO_142 (O_142,N_8455,N_8929);
nand UO_143 (O_143,N_8423,N_9082);
and UO_144 (O_144,N_9728,N_8188);
nand UO_145 (O_145,N_8299,N_9502);
nand UO_146 (O_146,N_9455,N_9753);
nor UO_147 (O_147,N_8764,N_8969);
nor UO_148 (O_148,N_9042,N_8749);
and UO_149 (O_149,N_8784,N_8080);
nor UO_150 (O_150,N_9527,N_8327);
and UO_151 (O_151,N_9662,N_9061);
nand UO_152 (O_152,N_9334,N_8103);
nand UO_153 (O_153,N_8864,N_9308);
nor UO_154 (O_154,N_8137,N_8247);
or UO_155 (O_155,N_9850,N_9079);
nor UO_156 (O_156,N_9250,N_9905);
nand UO_157 (O_157,N_8820,N_8957);
nor UO_158 (O_158,N_9663,N_9713);
or UO_159 (O_159,N_8070,N_8858);
or UO_160 (O_160,N_9227,N_8682);
nor UO_161 (O_161,N_8215,N_9745);
nor UO_162 (O_162,N_8057,N_9213);
xnor UO_163 (O_163,N_9874,N_8643);
xnor UO_164 (O_164,N_9473,N_9275);
nor UO_165 (O_165,N_9670,N_9483);
nor UO_166 (O_166,N_8946,N_8442);
nand UO_167 (O_167,N_9115,N_8191);
nand UO_168 (O_168,N_9471,N_9432);
nand UO_169 (O_169,N_9878,N_8409);
nand UO_170 (O_170,N_9442,N_9561);
nor UO_171 (O_171,N_9153,N_9041);
nand UO_172 (O_172,N_8965,N_9882);
or UO_173 (O_173,N_8403,N_9928);
nand UO_174 (O_174,N_8612,N_9628);
nand UO_175 (O_175,N_9450,N_8768);
nor UO_176 (O_176,N_8701,N_9288);
nor UO_177 (O_177,N_8551,N_8826);
or UO_178 (O_178,N_9682,N_9136);
xor UO_179 (O_179,N_9703,N_8488);
and UO_180 (O_180,N_9125,N_9024);
nor UO_181 (O_181,N_9661,N_9709);
or UO_182 (O_182,N_9433,N_8531);
xnor UO_183 (O_183,N_8507,N_9242);
and UO_184 (O_184,N_8723,N_9106);
nand UO_185 (O_185,N_8301,N_9400);
nor UO_186 (O_186,N_9382,N_9456);
and UO_187 (O_187,N_9459,N_8518);
nand UO_188 (O_188,N_8783,N_9801);
and UO_189 (O_189,N_9446,N_8220);
nand UO_190 (O_190,N_9790,N_8538);
and UO_191 (O_191,N_8600,N_8616);
nor UO_192 (O_192,N_8405,N_8047);
nand UO_193 (O_193,N_9904,N_9659);
nor UO_194 (O_194,N_9186,N_9892);
and UO_195 (O_195,N_9087,N_9841);
nand UO_196 (O_196,N_9574,N_8925);
nor UO_197 (O_197,N_8667,N_9147);
and UO_198 (O_198,N_9785,N_8956);
nand UO_199 (O_199,N_9371,N_8711);
nor UO_200 (O_200,N_8372,N_9461);
xnor UO_201 (O_201,N_8754,N_8746);
and UO_202 (O_202,N_8152,N_9158);
and UO_203 (O_203,N_8079,N_9183);
or UO_204 (O_204,N_8180,N_8953);
and UO_205 (O_205,N_9640,N_9435);
or UO_206 (O_206,N_9534,N_9163);
nor UO_207 (O_207,N_8025,N_9454);
nand UO_208 (O_208,N_9337,N_9470);
or UO_209 (O_209,N_8045,N_8097);
and UO_210 (O_210,N_8815,N_9976);
nor UO_211 (O_211,N_9706,N_8805);
and UO_212 (O_212,N_9958,N_8614);
nand UO_213 (O_213,N_9205,N_8296);
nand UO_214 (O_214,N_8470,N_8202);
nor UO_215 (O_215,N_8197,N_8498);
nand UO_216 (O_216,N_8294,N_8187);
and UO_217 (O_217,N_9815,N_9073);
nor UO_218 (O_218,N_8062,N_9397);
nand UO_219 (O_219,N_8257,N_8326);
or UO_220 (O_220,N_8093,N_8131);
nor UO_221 (O_221,N_8716,N_9961);
xnor UO_222 (O_222,N_8005,N_9252);
nor UO_223 (O_223,N_9266,N_8874);
nor UO_224 (O_224,N_8082,N_8194);
or UO_225 (O_225,N_9244,N_8412);
or UO_226 (O_226,N_8356,N_8793);
nand UO_227 (O_227,N_8303,N_8051);
nand UO_228 (O_228,N_9557,N_8617);
or UO_229 (O_229,N_8166,N_8828);
nand UO_230 (O_230,N_8661,N_9597);
xnor UO_231 (O_231,N_9809,N_9416);
or UO_232 (O_232,N_8725,N_8149);
and UO_233 (O_233,N_8777,N_9908);
nor UO_234 (O_234,N_9093,N_9008);
xnor UO_235 (O_235,N_8807,N_8120);
xor UO_236 (O_236,N_8609,N_9872);
nor UO_237 (O_237,N_9373,N_8624);
nor UO_238 (O_238,N_8487,N_9320);
nand UO_239 (O_239,N_8757,N_8717);
nor UO_240 (O_240,N_9311,N_8391);
nor UO_241 (O_241,N_9495,N_8613);
or UO_242 (O_242,N_8832,N_8185);
and UO_243 (O_243,N_9406,N_9245);
nor UO_244 (O_244,N_9520,N_9563);
and UO_245 (O_245,N_8398,N_9974);
nor UO_246 (O_246,N_8932,N_8597);
or UO_247 (O_247,N_9396,N_8760);
or UO_248 (O_248,N_8362,N_8145);
xnor UO_249 (O_249,N_8666,N_9179);
nand UO_250 (O_250,N_8473,N_9078);
nand UO_251 (O_251,N_9410,N_8533);
nor UO_252 (O_252,N_9441,N_8625);
and UO_253 (O_253,N_8756,N_9068);
nor UO_254 (O_254,N_8462,N_9270);
nor UO_255 (O_255,N_8313,N_9550);
nor UO_256 (O_256,N_9421,N_9666);
xnor UO_257 (O_257,N_9062,N_8927);
or UO_258 (O_258,N_9437,N_8193);
nor UO_259 (O_259,N_8335,N_9685);
nand UO_260 (O_260,N_9297,N_9900);
nand UO_261 (O_261,N_8640,N_8134);
nor UO_262 (O_262,N_9255,N_8981);
xnor UO_263 (O_263,N_8451,N_9750);
nand UO_264 (O_264,N_9238,N_9282);
or UO_265 (O_265,N_8743,N_8204);
and UO_266 (O_266,N_9876,N_9192);
nand UO_267 (O_267,N_8621,N_8853);
nor UO_268 (O_268,N_9813,N_8144);
or UO_269 (O_269,N_9317,N_8216);
xor UO_270 (O_270,N_8515,N_9671);
and UO_271 (O_271,N_9312,N_9415);
and UO_272 (O_272,N_8496,N_9542);
and UO_273 (O_273,N_8664,N_8881);
or UO_274 (O_274,N_8681,N_8333);
nor UO_275 (O_275,N_9343,N_9528);
xnor UO_276 (O_276,N_8639,N_8017);
nand UO_277 (O_277,N_8237,N_9097);
nand UO_278 (O_278,N_9048,N_8253);
nand UO_279 (O_279,N_9174,N_9873);
or UO_280 (O_280,N_8836,N_9467);
nand UO_281 (O_281,N_8731,N_8262);
nand UO_282 (O_282,N_9765,N_9616);
or UO_283 (O_283,N_9708,N_9044);
xnor UO_284 (O_284,N_8980,N_9268);
or UO_285 (O_285,N_8686,N_9865);
and UO_286 (O_286,N_8312,N_9921);
nand UO_287 (O_287,N_9170,N_9942);
nand UO_288 (O_288,N_8910,N_8792);
nor UO_289 (O_289,N_8320,N_8441);
or UO_290 (O_290,N_8148,N_9656);
and UO_291 (O_291,N_8810,N_8905);
or UO_292 (O_292,N_9702,N_9169);
nor UO_293 (O_293,N_8424,N_8252);
and UO_294 (O_294,N_8457,N_8735);
nand UO_295 (O_295,N_9469,N_9885);
nor UO_296 (O_296,N_9945,N_9769);
xnor UO_297 (O_297,N_8229,N_8886);
and UO_298 (O_298,N_8942,N_9653);
and UO_299 (O_299,N_9128,N_8278);
or UO_300 (O_300,N_8937,N_9814);
or UO_301 (O_301,N_9220,N_8426);
and UO_302 (O_302,N_8797,N_9022);
or UO_303 (O_303,N_9464,N_8122);
and UO_304 (O_304,N_9697,N_9920);
or UO_305 (O_305,N_8924,N_9973);
xnor UO_306 (O_306,N_8066,N_9764);
or UO_307 (O_307,N_9584,N_8976);
and UO_308 (O_308,N_9485,N_9229);
or UO_309 (O_309,N_8344,N_8406);
nor UO_310 (O_310,N_9338,N_9571);
nor UO_311 (O_311,N_8978,N_8734);
or UO_312 (O_312,N_8542,N_8090);
or UO_313 (O_313,N_9207,N_8841);
xor UO_314 (O_314,N_9466,N_8394);
xor UO_315 (O_315,N_9804,N_8986);
or UO_316 (O_316,N_8126,N_9260);
nand UO_317 (O_317,N_9763,N_9276);
or UO_318 (O_318,N_8887,N_9434);
or UO_319 (O_319,N_9447,N_8650);
or UO_320 (O_320,N_9361,N_8203);
nor UO_321 (O_321,N_8400,N_8647);
xor UO_322 (O_322,N_8570,N_9052);
or UO_323 (O_323,N_8174,N_9515);
nand UO_324 (O_324,N_9003,N_8342);
nand UO_325 (O_325,N_9422,N_8584);
or UO_326 (O_326,N_9738,N_8438);
nor UO_327 (O_327,N_9202,N_9793);
nor UO_328 (O_328,N_9523,N_9614);
nand UO_329 (O_329,N_9629,N_9772);
or UO_330 (O_330,N_8077,N_8446);
and UO_331 (O_331,N_9510,N_8380);
and UO_332 (O_332,N_8315,N_9767);
and UO_333 (O_333,N_9166,N_9016);
and UO_334 (O_334,N_8013,N_9940);
and UO_335 (O_335,N_9937,N_8763);
and UO_336 (O_336,N_9025,N_9633);
nor UO_337 (O_337,N_8813,N_8791);
or UO_338 (O_338,N_9808,N_8540);
or UO_339 (O_339,N_8125,N_9296);
or UO_340 (O_340,N_9468,N_9864);
nor UO_341 (O_341,N_8519,N_8293);
and UO_342 (O_342,N_9429,N_8523);
nand UO_343 (O_343,N_8261,N_8255);
nand UO_344 (O_344,N_9509,N_8889);
nor UO_345 (O_345,N_9092,N_8954);
nor UO_346 (O_346,N_9589,N_9909);
nand UO_347 (O_347,N_8444,N_9758);
nand UO_348 (O_348,N_9303,N_8355);
and UO_349 (O_349,N_9655,N_8195);
nand UO_350 (O_350,N_8545,N_8747);
and UO_351 (O_351,N_9914,N_8670);
nand UO_352 (O_352,N_8790,N_9727);
nand UO_353 (O_353,N_8363,N_8139);
nor UO_354 (O_354,N_9230,N_8837);
and UO_355 (O_355,N_9830,N_9345);
xnor UO_356 (O_356,N_9687,N_9218);
or UO_357 (O_357,N_8437,N_8004);
or UO_358 (O_358,N_8977,N_9988);
nor UO_359 (O_359,N_9011,N_9013);
nor UO_360 (O_360,N_8201,N_9754);
and UO_361 (O_361,N_8885,N_9782);
xnor UO_362 (O_362,N_8708,N_8067);
xor UO_363 (O_363,N_8578,N_9595);
nor UO_364 (O_364,N_8842,N_9072);
nand UO_365 (O_365,N_9634,N_9849);
nor UO_366 (O_366,N_9146,N_8780);
and UO_367 (O_367,N_9526,N_9980);
nand UO_368 (O_368,N_9152,N_8684);
or UO_369 (O_369,N_8029,N_9103);
nand UO_370 (O_370,N_9037,N_9902);
or UO_371 (O_371,N_9243,N_9842);
or UO_372 (O_372,N_8020,N_8430);
and UO_373 (O_373,N_9583,N_9462);
nor UO_374 (O_374,N_9081,N_8078);
xor UO_375 (O_375,N_8765,N_9593);
and UO_376 (O_376,N_9448,N_8648);
nand UO_377 (O_377,N_8435,N_9300);
and UO_378 (O_378,N_9392,N_8988);
xor UO_379 (O_379,N_8787,N_8581);
and UO_380 (O_380,N_9675,N_9910);
and UO_381 (O_381,N_8991,N_8821);
and UO_382 (O_382,N_9710,N_8785);
nand UO_383 (O_383,N_9991,N_8720);
nand UO_384 (O_384,N_8136,N_9741);
nand UO_385 (O_385,N_8258,N_8806);
nor UO_386 (O_386,N_8655,N_8690);
or UO_387 (O_387,N_9636,N_9119);
and UO_388 (O_388,N_8967,N_9066);
and UO_389 (O_389,N_9613,N_9010);
and UO_390 (O_390,N_9829,N_8970);
or UO_391 (O_391,N_8738,N_9247);
nand UO_392 (O_392,N_8582,N_8235);
nand UO_393 (O_393,N_9603,N_9277);
nand UO_394 (O_394,N_8458,N_9221);
nand UO_395 (O_395,N_8349,N_8627);
nor UO_396 (O_396,N_8931,N_9836);
or UO_397 (O_397,N_9002,N_8641);
nor UO_398 (O_398,N_9293,N_9766);
or UO_399 (O_399,N_9319,N_9036);
nand UO_400 (O_400,N_9113,N_8009);
and UO_401 (O_401,N_9390,N_9947);
xnor UO_402 (O_402,N_8896,N_9984);
and UO_403 (O_403,N_9363,N_9009);
or UO_404 (O_404,N_9643,N_9981);
or UO_405 (O_405,N_8751,N_8675);
nor UO_406 (O_406,N_8884,N_9582);
or UO_407 (O_407,N_8829,N_9807);
and UO_408 (O_408,N_8377,N_8915);
nand UO_409 (O_409,N_9929,N_9474);
nand UO_410 (O_410,N_9328,N_8950);
and UO_411 (O_411,N_9919,N_9518);
or UO_412 (O_412,N_9493,N_9553);
nor UO_413 (O_413,N_9572,N_9694);
nand UO_414 (O_414,N_8715,N_9038);
or UO_415 (O_415,N_8703,N_8744);
nor UO_416 (O_416,N_9695,N_9262);
or UO_417 (O_417,N_9332,N_8602);
xor UO_418 (O_418,N_9499,N_9975);
or UO_419 (O_419,N_9719,N_8339);
nand UO_420 (O_420,N_8211,N_9630);
nor UO_421 (O_421,N_8951,N_9118);
nor UO_422 (O_422,N_9100,N_9736);
xnor UO_423 (O_423,N_8346,N_9686);
nor UO_424 (O_424,N_8632,N_9992);
and UO_425 (O_425,N_8850,N_8983);
and UO_426 (O_426,N_8733,N_9822);
or UO_427 (O_427,N_9575,N_9393);
and UO_428 (O_428,N_8758,N_9209);
or UO_429 (O_429,N_8012,N_9532);
and UO_430 (O_430,N_9232,N_8691);
or UO_431 (O_431,N_8281,N_9272);
and UO_432 (O_432,N_8042,N_9931);
nand UO_433 (O_433,N_8506,N_8857);
and UO_434 (O_434,N_8949,N_8359);
xor UO_435 (O_435,N_9417,N_9223);
and UO_436 (O_436,N_8657,N_8952);
nand UO_437 (O_437,N_9789,N_8646);
or UO_438 (O_438,N_8637,N_8039);
and UO_439 (O_439,N_8234,N_8906);
xnor UO_440 (O_440,N_9884,N_8116);
and UO_441 (O_441,N_9524,N_8917);
nand UO_442 (O_442,N_9098,N_9517);
and UO_443 (O_443,N_9412,N_9131);
nor UO_444 (O_444,N_8129,N_8172);
xnor UO_445 (O_445,N_9443,N_9781);
xor UO_446 (O_446,N_9033,N_8169);
nor UO_447 (O_447,N_8851,N_9998);
xnor UO_448 (O_448,N_8555,N_9875);
or UO_449 (O_449,N_8021,N_8016);
or UO_450 (O_450,N_8825,N_9529);
or UO_451 (O_451,N_9254,N_8317);
xnor UO_452 (O_452,N_8503,N_8814);
nor UO_453 (O_453,N_9609,N_8286);
nor UO_454 (O_454,N_9821,N_9215);
nor UO_455 (O_455,N_9211,N_9116);
nand UO_456 (O_456,N_9681,N_8572);
or UO_457 (O_457,N_9546,N_8727);
or UO_458 (O_458,N_9080,N_9954);
xor UO_459 (O_459,N_9959,N_9811);
and UO_460 (O_460,N_9698,N_9556);
nand UO_461 (O_461,N_9143,N_9134);
xor UO_462 (O_462,N_9649,N_9346);
or UO_463 (O_463,N_9941,N_9354);
nand UO_464 (O_464,N_8244,N_9182);
and UO_465 (O_465,N_8534,N_8500);
and UO_466 (O_466,N_9627,N_9012);
nor UO_467 (O_467,N_8808,N_9017);
or UO_468 (O_468,N_8795,N_8073);
nand UO_469 (O_469,N_9839,N_8241);
nand UO_470 (O_470,N_8522,N_8492);
and UO_471 (O_471,N_8486,N_9915);
or UO_472 (O_472,N_8770,N_8121);
nor UO_473 (O_473,N_9301,N_9599);
nor UO_474 (O_474,N_8182,N_8155);
and UO_475 (O_475,N_9562,N_9374);
nor UO_476 (O_476,N_8341,N_9472);
nor UO_477 (O_477,N_9779,N_9065);
nor UO_478 (O_478,N_8399,N_8961);
nand UO_479 (O_479,N_9057,N_8083);
or UO_480 (O_480,N_9898,N_9349);
and UO_481 (O_481,N_9278,N_9197);
nor UO_482 (O_482,N_8638,N_9331);
nor UO_483 (O_483,N_8375,N_9043);
nor UO_484 (O_484,N_8217,N_9544);
and UO_485 (O_485,N_8334,N_9187);
nor UO_486 (O_486,N_9399,N_9326);
nor UO_487 (O_487,N_8844,N_9105);
nor UO_488 (O_488,N_9148,N_8386);
or UO_489 (O_489,N_9309,N_8722);
nand UO_490 (O_490,N_8432,N_8497);
and UO_491 (O_491,N_9253,N_9249);
nor UO_492 (O_492,N_9171,N_8822);
or UO_493 (O_493,N_8106,N_9537);
or UO_494 (O_494,N_9487,N_9034);
and UO_495 (O_495,N_8461,N_9985);
and UO_496 (O_496,N_9737,N_8900);
and UO_497 (O_497,N_8502,N_9889);
or UO_498 (O_498,N_9318,N_9175);
xor UO_499 (O_499,N_9859,N_9127);
or UO_500 (O_500,N_8631,N_9364);
nor UO_501 (O_501,N_8065,N_8074);
or UO_502 (O_502,N_9101,N_8418);
xnor UO_503 (O_503,N_8702,N_9500);
and UO_504 (O_504,N_8767,N_9069);
or UO_505 (O_505,N_8130,N_8623);
and UO_506 (O_506,N_9715,N_9219);
nor UO_507 (O_507,N_9095,N_8345);
or UO_508 (O_508,N_8782,N_9660);
nand UO_509 (O_509,N_8383,N_9070);
xnor UO_510 (O_510,N_9513,N_9457);
and UO_511 (O_511,N_8353,N_9925);
nand UO_512 (O_512,N_8871,N_8802);
nor UO_513 (O_513,N_9746,N_9088);
xnor UO_514 (O_514,N_9225,N_9440);
and UO_515 (O_515,N_8178,N_8673);
nand UO_516 (O_516,N_8413,N_8328);
nand UO_517 (O_517,N_9323,N_9775);
nor UO_518 (O_518,N_8171,N_8943);
and UO_519 (O_519,N_9258,N_9880);
and UO_520 (O_520,N_9203,N_8494);
xor UO_521 (O_521,N_9837,N_9360);
nor UO_522 (O_522,N_8371,N_9887);
or UO_523 (O_523,N_9729,N_9983);
xnor UO_524 (O_524,N_9525,N_9054);
or UO_525 (O_525,N_8043,N_8050);
nand UO_526 (O_526,N_8436,N_8033);
or UO_527 (O_527,N_8603,N_9451);
nor UO_528 (O_528,N_8823,N_9679);
and UO_529 (O_529,N_9505,N_9749);
and UO_530 (O_530,N_8800,N_8221);
nand UO_531 (O_531,N_8525,N_8416);
nor UO_532 (O_532,N_8947,N_9967);
or UO_533 (O_533,N_9516,N_9993);
or UO_534 (O_534,N_8509,N_8979);
nor UO_535 (O_535,N_8036,N_8443);
nand UO_536 (O_536,N_9351,N_9423);
and UO_537 (O_537,N_9732,N_9046);
or UO_538 (O_538,N_9251,N_8307);
nand UO_539 (O_539,N_8484,N_9559);
or UO_540 (O_540,N_9672,N_8585);
nand UO_541 (O_541,N_8699,N_9806);
and UO_542 (O_542,N_8912,N_8781);
or UO_543 (O_543,N_9723,N_9112);
nand UO_544 (O_544,N_9384,N_9751);
and UO_545 (O_545,N_9549,N_9431);
or UO_546 (O_546,N_8480,N_9151);
or UO_547 (O_547,N_8179,N_8973);
and UO_548 (O_548,N_9743,N_9333);
and UO_549 (O_549,N_9307,N_8337);
nor UO_550 (O_550,N_8645,N_9623);
and UO_551 (O_551,N_9932,N_8831);
xnor UO_552 (O_552,N_8590,N_8971);
xor UO_553 (O_553,N_8030,N_8490);
nand UO_554 (O_554,N_9658,N_8998);
nand UO_555 (O_555,N_9291,N_9798);
or UO_556 (O_556,N_9140,N_8692);
nor UO_557 (O_557,N_8366,N_9463);
and UO_558 (O_558,N_8833,N_8605);
nand UO_559 (O_559,N_9699,N_9403);
nand UO_560 (O_560,N_8809,N_8181);
nor UO_561 (O_561,N_8914,N_9507);
nor UO_562 (O_562,N_8959,N_8456);
xor UO_563 (O_563,N_8936,N_8055);
or UO_564 (O_564,N_8306,N_8154);
nor UO_565 (O_565,N_9600,N_9491);
and UO_566 (O_566,N_8803,N_9408);
nand UO_567 (O_567,N_8495,N_8279);
or UO_568 (O_568,N_8076,N_8654);
xnor UO_569 (O_569,N_9160,N_9367);
and UO_570 (O_570,N_9114,N_8213);
or UO_571 (O_571,N_8945,N_9000);
xor UO_572 (O_572,N_9005,N_9404);
nand UO_573 (O_573,N_8840,N_8742);
xnor UO_574 (O_574,N_9176,N_8011);
nand UO_575 (O_575,N_8331,N_8041);
or UO_576 (O_576,N_9504,N_9001);
xor UO_577 (O_577,N_9773,N_9358);
xor UO_578 (O_578,N_8984,N_9233);
nand UO_579 (O_579,N_8520,N_8679);
or UO_580 (O_580,N_9045,N_9302);
nor UO_581 (O_581,N_8242,N_8899);
nor UO_582 (O_582,N_9381,N_9680);
nor UO_583 (O_583,N_9757,N_9436);
nor UO_584 (O_584,N_8297,N_8465);
nor UO_585 (O_585,N_9482,N_8855);
nand UO_586 (O_586,N_8388,N_9718);
or UO_587 (O_587,N_9511,N_9383);
nor UO_588 (O_588,N_8876,N_9292);
or UO_589 (O_589,N_8475,N_8861);
nand UO_590 (O_590,N_9585,N_9963);
and UO_591 (O_591,N_8587,N_9362);
or UO_592 (O_592,N_9522,N_9149);
nor UO_593 (O_593,N_8608,N_8618);
or UO_594 (O_594,N_8287,N_8165);
nor UO_595 (O_595,N_9939,N_9797);
and UO_596 (O_596,N_8948,N_9786);
nor UO_597 (O_597,N_9359,N_9015);
nor UO_598 (O_598,N_9673,N_8845);
nor UO_599 (O_599,N_8351,N_9376);
or UO_600 (O_600,N_8422,N_9978);
or UO_601 (O_601,N_8192,N_9352);
or UO_602 (O_602,N_9762,N_8583);
or UO_603 (O_603,N_8878,N_9895);
and UO_604 (O_604,N_9812,N_9479);
nand UO_605 (O_605,N_9449,N_8175);
nor UO_606 (O_606,N_8730,N_9968);
nor UO_607 (O_607,N_8292,N_8264);
xor UO_608 (O_608,N_9185,N_9794);
or UO_609 (O_609,N_8478,N_8209);
or UO_610 (O_610,N_8926,N_9427);
nor UO_611 (O_611,N_9800,N_9299);
and UO_612 (O_612,N_9050,N_9535);
nor UO_613 (O_613,N_8816,N_9780);
and UO_614 (O_614,N_8846,N_9208);
and UO_615 (O_615,N_9691,N_9026);
nor UO_616 (O_616,N_8196,N_9734);
xor UO_617 (O_617,N_9989,N_9826);
nand UO_618 (O_618,N_8830,N_9594);
nor UO_619 (O_619,N_9335,N_9508);
nor UO_620 (O_620,N_9888,N_8084);
and UO_621 (O_621,N_8662,N_9224);
nand UO_622 (O_622,N_9906,N_8736);
nand UO_623 (O_623,N_8964,N_8536);
and UO_624 (O_624,N_9141,N_8003);
xor UO_625 (O_625,N_9545,N_8163);
nand UO_626 (O_626,N_9426,N_8064);
nand UO_627 (O_627,N_8689,N_8962);
nor UO_628 (O_628,N_8071,N_8923);
nand UO_629 (O_629,N_8529,N_9999);
or UO_630 (O_630,N_9110,N_8291);
nand UO_631 (O_631,N_9168,N_8267);
nor UO_632 (O_632,N_8505,N_9489);
or UO_633 (O_633,N_8839,N_9911);
and UO_634 (O_634,N_9861,N_9475);
nor UO_635 (O_635,N_8417,N_8236);
xor UO_636 (O_636,N_9739,N_8477);
nor UO_637 (O_637,N_9111,N_8198);
nand UO_638 (O_638,N_9091,N_9855);
nor UO_639 (O_639,N_9217,N_8232);
nor UO_640 (O_640,N_9927,N_9858);
nor UO_641 (O_641,N_9503,N_9344);
nor UO_642 (O_642,N_8308,N_9645);
nor UO_643 (O_643,N_9130,N_8601);
nand UO_644 (O_644,N_9700,N_8019);
and UO_645 (O_645,N_9692,N_9188);
or UO_646 (O_646,N_9690,N_9950);
or UO_647 (O_647,N_9618,N_9122);
or UO_648 (O_648,N_9701,N_8397);
and UO_649 (O_649,N_8230,N_8527);
and UO_650 (O_650,N_8922,N_8918);
and UO_651 (O_651,N_9027,N_9683);
or UO_652 (O_652,N_9901,N_9411);
nor UO_653 (O_653,N_9818,N_8284);
xnor UO_654 (O_654,N_9608,N_9313);
or UO_655 (O_655,N_8425,N_8369);
nor UO_656 (O_656,N_8683,N_8002);
nor UO_657 (O_657,N_8577,N_9460);
nor UO_658 (O_658,N_8061,N_8271);
nor UO_659 (O_659,N_8778,N_9341);
nand UO_660 (O_660,N_8622,N_8908);
and UO_661 (O_661,N_9414,N_9305);
and UO_662 (O_662,N_8225,N_8250);
or UO_663 (O_663,N_8467,N_8700);
nand UO_664 (O_664,N_9768,N_9401);
or UO_665 (O_665,N_8737,N_9759);
and UO_666 (O_666,N_9071,N_9214);
and UO_667 (O_667,N_8559,N_9286);
xnor UO_668 (O_668,N_8963,N_9210);
xor UO_669 (O_669,N_9316,N_9156);
or UO_670 (O_670,N_9369,N_9560);
and UO_671 (O_671,N_8579,N_8314);
nand UO_672 (O_672,N_8571,N_9257);
xnor UO_673 (O_673,N_8092,N_9329);
nand UO_674 (O_674,N_9285,N_8504);
or UO_675 (O_675,N_9018,N_9407);
nor UO_676 (O_676,N_8108,N_8512);
and UO_677 (O_677,N_8199,N_9607);
nand UO_678 (O_678,N_8996,N_8799);
and UO_679 (O_679,N_8008,N_8594);
or UO_680 (O_680,N_9347,N_9650);
or UO_681 (O_681,N_9481,N_8428);
nor UO_682 (O_682,N_9857,N_8088);
nor UO_683 (O_683,N_9792,N_8096);
or UO_684 (O_684,N_8159,N_8056);
or UO_685 (O_685,N_9558,N_8847);
xnor UO_686 (O_686,N_9379,N_8280);
nand UO_687 (O_687,N_8445,N_8212);
and UO_688 (O_688,N_9053,N_9274);
nand UO_689 (O_689,N_9918,N_8176);
xnor UO_690 (O_690,N_9290,N_8755);
nor UO_691 (O_691,N_9295,N_8270);
nor UO_692 (O_692,N_9755,N_8897);
and UO_693 (O_693,N_9960,N_9051);
nor UO_694 (O_694,N_8989,N_9644);
and UO_695 (O_695,N_9631,N_8227);
nand UO_696 (O_696,N_8909,N_8027);
or UO_697 (O_697,N_9588,N_8669);
or UO_698 (O_698,N_8414,N_8696);
nor UO_699 (O_699,N_8698,N_8592);
xor UO_700 (O_700,N_9949,N_8548);
nand UO_701 (O_701,N_8160,N_8119);
xnor UO_702 (O_702,N_8158,N_9926);
nand UO_703 (O_703,N_8310,N_9944);
nand UO_704 (O_704,N_9621,N_9881);
nand UO_705 (O_705,N_8091,N_9547);
nor UO_706 (O_706,N_9735,N_8870);
xor UO_707 (O_707,N_8530,N_9199);
or UO_708 (O_708,N_9833,N_8382);
nand UO_709 (O_709,N_9102,N_9035);
or UO_710 (O_710,N_9592,N_9756);
xor UO_711 (O_711,N_9531,N_9637);
nor UO_712 (O_712,N_8087,N_9267);
nand UO_713 (O_713,N_8046,N_8387);
or UO_714 (O_714,N_8343,N_8135);
and UO_715 (O_715,N_9725,N_9848);
nor UO_716 (O_716,N_9246,N_8891);
nor UO_717 (O_717,N_9395,N_9724);
and UO_718 (O_718,N_9714,N_9846);
or UO_719 (O_719,N_9074,N_9173);
xor UO_720 (O_720,N_9704,N_9612);
nand UO_721 (O_721,N_9678,N_9490);
nor UO_722 (O_722,N_9324,N_8000);
and UO_723 (O_723,N_8373,N_9554);
nand UO_724 (O_724,N_8993,N_8898);
nor UO_725 (O_725,N_8032,N_8995);
and UO_726 (O_726,N_8776,N_9321);
or UO_727 (O_727,N_9327,N_8233);
nor UO_728 (O_728,N_8660,N_9817);
xnor UO_729 (O_729,N_9707,N_9896);
and UO_730 (O_730,N_8526,N_8123);
and UO_731 (O_731,N_8218,N_8852);
and UO_732 (O_732,N_8289,N_9971);
and UO_733 (O_733,N_8381,N_8038);
nor UO_734 (O_734,N_8395,N_9386);
and UO_735 (O_735,N_8493,N_9538);
xor UO_736 (O_736,N_8177,N_9453);
nand UO_737 (O_737,N_9086,N_8085);
and UO_738 (O_738,N_8068,N_8466);
nand UO_739 (O_739,N_9964,N_8390);
or UO_740 (O_740,N_9795,N_8586);
or UO_741 (O_741,N_9890,N_8268);
xnor UO_742 (O_742,N_9933,N_9239);
and UO_743 (O_743,N_8911,N_9943);
nor UO_744 (O_744,N_8246,N_8676);
xor UO_745 (O_745,N_9860,N_8471);
or UO_746 (O_746,N_8059,N_9165);
nand UO_747 (O_747,N_9497,N_8882);
or UO_748 (O_748,N_9409,N_9831);
xor UO_749 (O_749,N_8697,N_9040);
or UO_750 (O_750,N_9995,N_8552);
and UO_751 (O_751,N_8434,N_9606);
nor UO_752 (O_752,N_9586,N_8332);
nand UO_753 (O_753,N_8207,N_8111);
or UO_754 (O_754,N_8665,N_8472);
nand UO_755 (O_755,N_8266,N_8880);
or UO_756 (O_756,N_9788,N_8094);
nand UO_757 (O_757,N_8546,N_8274);
nand UO_758 (O_758,N_9241,N_8558);
or UO_759 (O_759,N_9083,N_9039);
xor UO_760 (O_760,N_8537,N_8024);
nand UO_761 (O_761,N_8459,N_9913);
nand UO_762 (O_762,N_9090,N_9056);
or UO_763 (O_763,N_8685,N_8168);
or UO_764 (O_764,N_8958,N_8719);
or UO_765 (O_765,N_9654,N_9075);
and UO_766 (O_766,N_9263,N_8449);
or UO_767 (O_767,N_8161,N_8081);
or UO_768 (O_768,N_8611,N_9868);
or UO_769 (O_769,N_8350,N_8157);
or UO_770 (O_770,N_9620,N_9076);
and UO_771 (O_771,N_9957,N_9256);
nor UO_772 (O_772,N_8321,N_8933);
nor UO_773 (O_773,N_9145,N_8766);
or UO_774 (O_774,N_8170,N_8771);
or UO_775 (O_775,N_9273,N_8619);
nand UO_776 (O_776,N_8072,N_9689);
and UO_777 (O_777,N_8824,N_9624);
xnor UO_778 (O_778,N_8112,N_9539);
nand UO_779 (O_779,N_9067,N_9512);
or UO_780 (O_780,N_8569,N_9094);
nor UO_781 (O_781,N_9058,N_9577);
nand UO_782 (O_782,N_8634,N_9425);
xor UO_783 (O_783,N_8863,N_8348);
or UO_784 (O_784,N_9129,N_8474);
nand UO_785 (O_785,N_9342,N_8183);
nor UO_786 (O_786,N_9120,N_8368);
xor UO_787 (O_787,N_8867,N_8672);
nand UO_788 (O_788,N_8879,N_8100);
nor UO_789 (O_789,N_8133,N_8628);
xnor UO_790 (O_790,N_8838,N_8656);
and UO_791 (O_791,N_9851,N_9677);
nor UO_792 (O_792,N_8687,N_9951);
or UO_793 (O_793,N_8098,N_8759);
nor UO_794 (O_794,N_8052,N_8156);
nor UO_795 (O_795,N_9742,N_8184);
nand UO_796 (O_796,N_9541,N_9986);
and UO_797 (O_797,N_9138,N_9157);
or UO_798 (O_798,N_9085,N_9280);
nand UO_799 (O_799,N_8968,N_8427);
nor UO_800 (O_800,N_8779,N_8726);
and UO_801 (O_801,N_9744,N_8089);
nor UO_802 (O_802,N_9720,N_8547);
and UO_803 (O_803,N_8712,N_8302);
nand UO_804 (O_804,N_8568,N_9063);
xor UO_805 (O_805,N_9651,N_9647);
or UO_806 (O_806,N_9733,N_8688);
nor UO_807 (O_807,N_9271,N_8352);
or UO_808 (O_808,N_9965,N_8798);
nand UO_809 (O_809,N_8944,N_9696);
nand UO_810 (O_810,N_8653,N_8190);
nand UO_811 (O_811,N_9398,N_9375);
nor UO_812 (O_812,N_9235,N_8819);
nand UO_813 (O_813,N_8940,N_9646);
nor UO_814 (O_814,N_8557,N_9190);
nand UO_815 (O_815,N_9310,N_9844);
nand UO_816 (O_816,N_9602,N_8054);
or UO_817 (O_817,N_8304,N_9477);
xnor UO_818 (O_818,N_9155,N_8901);
or UO_819 (O_819,N_8018,N_8354);
nand UO_820 (O_820,N_9478,N_8564);
nand UO_821 (O_821,N_8128,N_9154);
nand UO_822 (O_822,N_8263,N_8560);
and UO_823 (O_823,N_9632,N_8273);
or UO_824 (O_824,N_8511,N_9167);
or UO_825 (O_825,N_9838,N_8869);
nor UO_826 (O_826,N_8544,N_9378);
xor UO_827 (O_827,N_8338,N_8063);
and UO_828 (O_828,N_8265,N_9139);
and UO_829 (O_829,N_8243,N_9617);
nand UO_830 (O_830,N_8006,N_8748);
nor UO_831 (O_831,N_9339,N_9237);
and UO_832 (O_832,N_8856,N_9370);
or UO_833 (O_833,N_8610,N_9294);
nor UO_834 (O_834,N_8510,N_8210);
or UO_835 (O_835,N_8114,N_9194);
nand UO_836 (O_836,N_9567,N_8563);
or UO_837 (O_837,N_8410,N_8930);
nand UO_838 (O_838,N_9907,N_8357);
and UO_839 (O_839,N_8630,N_9077);
or UO_840 (O_840,N_9476,N_8288);
or UO_841 (O_841,N_9330,N_8282);
or UO_842 (O_842,N_9688,N_8028);
nand UO_843 (O_843,N_8238,N_9879);
xor UO_844 (O_844,N_8801,N_8554);
nor UO_845 (O_845,N_8615,N_9216);
nor UO_846 (O_846,N_9828,N_9162);
nand UO_847 (O_847,N_9684,N_8606);
and UO_848 (O_848,N_8347,N_8482);
nor UO_849 (O_849,N_9521,N_8804);
nor UO_850 (O_850,N_8044,N_8322);
xnor UO_851 (O_851,N_8674,N_9604);
and UO_852 (O_852,N_9893,N_8460);
and UO_853 (O_853,N_8818,N_8407);
xor UO_854 (O_854,N_8972,N_8663);
or UO_855 (O_855,N_9566,N_8567);
and UO_856 (O_856,N_9903,N_9641);
nor UO_857 (O_857,N_9590,N_8994);
or UO_858 (O_858,N_8479,N_8109);
and UO_859 (O_859,N_9428,N_8633);
or UO_860 (O_860,N_9322,N_9193);
nor UO_861 (O_861,N_9047,N_9498);
nand UO_862 (O_862,N_8902,N_9287);
and UO_863 (O_863,N_8277,N_9693);
and UO_864 (O_864,N_8775,N_8223);
or UO_865 (O_865,N_9265,N_9946);
or UO_866 (O_866,N_9626,N_9740);
nand UO_867 (O_867,N_8167,N_8075);
and UO_868 (O_868,N_9543,N_8872);
nand UO_869 (O_869,N_9269,N_8834);
and UO_870 (O_870,N_8854,N_8794);
xnor UO_871 (O_871,N_8411,N_9717);
or UO_872 (O_872,N_8508,N_9969);
and UO_873 (O_873,N_8960,N_8817);
and UO_874 (O_874,N_9897,N_8718);
nor UO_875 (O_875,N_8249,N_9777);
nand UO_876 (O_876,N_8419,N_8272);
and UO_877 (O_877,N_9664,N_9356);
or UO_878 (O_878,N_8921,N_9006);
nand UO_879 (O_879,N_9748,N_9108);
nand UO_880 (O_880,N_8023,N_9064);
xnor UO_881 (O_881,N_8811,N_9177);
nand UO_882 (O_882,N_9576,N_9722);
nor UO_883 (O_883,N_9007,N_9430);
nand UO_884 (O_884,N_9825,N_8827);
nor UO_885 (O_885,N_8598,N_8877);
xor UO_886 (O_886,N_8788,N_9810);
and UO_887 (O_887,N_9770,N_8761);
and UO_888 (O_888,N_8588,N_8127);
and UO_889 (O_889,N_8214,N_8305);
nand UO_890 (O_890,N_9783,N_9938);
nor UO_891 (O_891,N_8740,N_8865);
or UO_892 (O_892,N_9970,N_8860);
or UO_893 (O_893,N_8642,N_8528);
nor UO_894 (O_894,N_9912,N_8228);
or UO_895 (O_895,N_9480,N_8658);
nand UO_896 (O_896,N_8385,N_8890);
nand UO_897 (O_897,N_9023,N_9385);
and UO_898 (O_898,N_9084,N_8997);
nor UO_899 (O_899,N_8336,N_8022);
nor UO_900 (O_900,N_9854,N_8115);
nand UO_901 (O_901,N_9996,N_9843);
and UO_902 (O_902,N_8448,N_8401);
nor UO_903 (O_903,N_9845,N_9283);
nor UO_904 (O_904,N_8928,N_8463);
and UO_905 (O_905,N_8439,N_9796);
or UO_906 (O_906,N_9240,N_8535);
nor UO_907 (O_907,N_8404,N_8599);
and UO_908 (O_908,N_9284,N_8739);
and UO_909 (O_909,N_8895,N_9150);
or UO_910 (O_910,N_8010,N_9869);
nand UO_911 (O_911,N_8384,N_8573);
or UO_912 (O_912,N_9638,N_8499);
and UO_913 (O_913,N_9747,N_9366);
xor UO_914 (O_914,N_8955,N_8709);
xor UO_915 (O_915,N_8990,N_9189);
and UO_916 (O_916,N_9581,N_9891);
nor UO_917 (O_917,N_9184,N_8556);
and UO_918 (O_918,N_9452,N_9923);
nand UO_919 (O_919,N_8903,N_9413);
xor UO_920 (O_920,N_8102,N_8105);
and UO_921 (O_921,N_8007,N_9304);
and UO_922 (O_922,N_8875,N_8421);
and UO_923 (O_923,N_9823,N_9899);
xor UO_924 (O_924,N_8205,N_8541);
xor UO_925 (O_925,N_9144,N_8329);
xnor UO_926 (O_926,N_8966,N_8360);
nand UO_927 (O_927,N_8162,N_9172);
nor UO_928 (O_928,N_9761,N_9917);
and UO_929 (O_929,N_9444,N_9402);
or UO_930 (O_930,N_9195,N_9580);
and UO_931 (O_931,N_9578,N_8935);
and UO_932 (O_932,N_9030,N_9784);
nor UO_933 (O_933,N_9635,N_8015);
or UO_934 (O_934,N_8049,N_9676);
nor UO_935 (O_935,N_8849,N_9610);
and UO_936 (O_936,N_8553,N_9492);
and UO_937 (O_937,N_9605,N_9955);
and UO_938 (O_938,N_9222,N_9226);
nand UO_939 (O_939,N_9198,N_9977);
nand UO_940 (O_940,N_8773,N_9514);
and UO_941 (O_941,N_8796,N_8415);
or UO_942 (O_942,N_9863,N_9060);
or UO_943 (O_943,N_9935,N_9424);
nor UO_944 (O_944,N_9852,N_8772);
and UO_945 (O_945,N_9730,N_8532);
nand UO_946 (O_946,N_8440,N_8260);
and UO_947 (O_947,N_8693,N_8222);
nand UO_948 (O_948,N_9721,N_9029);
or UO_949 (O_949,N_8408,N_9439);
and UO_950 (O_950,N_9089,N_8677);
nor UO_951 (O_951,N_8893,N_9922);
nor UO_952 (O_952,N_8035,N_9791);
nor UO_953 (O_953,N_9948,N_9820);
or UO_954 (O_954,N_9389,N_8110);
nand UO_955 (O_955,N_9625,N_8318);
nor UO_956 (O_956,N_8311,N_8259);
nor UO_957 (O_957,N_9204,N_8491);
and UO_958 (O_958,N_8468,N_8143);
xor UO_959 (O_959,N_9391,N_8186);
xor UO_960 (O_960,N_8835,N_9248);
nand UO_961 (O_961,N_9137,N_8208);
or UO_962 (O_962,N_9261,N_9231);
nand UO_963 (O_963,N_9598,N_9191);
nand UO_964 (O_964,N_8561,N_8452);
and UO_965 (O_965,N_8099,N_9126);
nand UO_966 (O_966,N_8513,N_8173);
nor UO_967 (O_967,N_8330,N_8659);
nand UO_968 (O_968,N_8987,N_9234);
and UO_969 (O_969,N_8741,N_9494);
and UO_970 (O_970,N_8975,N_9760);
or UO_971 (O_971,N_9484,N_9568);
nor UO_972 (O_972,N_9866,N_8707);
nor UO_973 (O_973,N_9438,N_8999);
nor UO_974 (O_974,N_9348,N_9336);
nand UO_975 (O_975,N_9279,N_9847);
or UO_976 (O_976,N_9109,N_8652);
xor UO_977 (O_977,N_9573,N_8364);
nor UO_978 (O_978,N_9936,N_9161);
nand UO_979 (O_979,N_9353,N_9870);
nand UO_980 (O_980,N_9712,N_9259);
or UO_981 (O_981,N_9020,N_8142);
or UO_982 (O_982,N_9121,N_9871);
and UO_983 (O_983,N_9405,N_9032);
nand UO_984 (O_984,N_8786,N_8101);
and UO_985 (O_985,N_8323,N_8644);
and UO_986 (O_986,N_9536,N_9357);
nor UO_987 (O_987,N_9564,N_8982);
nand UO_988 (O_988,N_9966,N_8358);
and UO_989 (O_989,N_9569,N_8037);
nand UO_990 (O_990,N_9667,N_9565);
xnor UO_991 (O_991,N_9458,N_9601);
and UO_992 (O_992,N_8319,N_9486);
nor UO_993 (O_993,N_8514,N_8680);
and UO_994 (O_994,N_8283,N_9314);
or UO_995 (O_995,N_9200,N_8635);
nor UO_996 (O_996,N_8206,N_8721);
nand UO_997 (O_997,N_8140,N_8724);
or UO_998 (O_998,N_8728,N_8450);
nand UO_999 (O_999,N_8325,N_8365);
and UO_1000 (O_1000,N_9592,N_9229);
nor UO_1001 (O_1001,N_8024,N_8094);
nor UO_1002 (O_1002,N_8417,N_9878);
and UO_1003 (O_1003,N_9683,N_8438);
and UO_1004 (O_1004,N_9661,N_8163);
and UO_1005 (O_1005,N_9667,N_9750);
and UO_1006 (O_1006,N_8893,N_9171);
or UO_1007 (O_1007,N_9080,N_8666);
xor UO_1008 (O_1008,N_9320,N_9350);
nor UO_1009 (O_1009,N_8912,N_9926);
or UO_1010 (O_1010,N_9143,N_9251);
nor UO_1011 (O_1011,N_9021,N_8605);
nand UO_1012 (O_1012,N_8471,N_8723);
nor UO_1013 (O_1013,N_8310,N_9445);
or UO_1014 (O_1014,N_9411,N_9571);
nor UO_1015 (O_1015,N_9331,N_8208);
nor UO_1016 (O_1016,N_9055,N_9059);
xor UO_1017 (O_1017,N_8750,N_9722);
or UO_1018 (O_1018,N_8225,N_8465);
nor UO_1019 (O_1019,N_8928,N_8408);
nor UO_1020 (O_1020,N_8952,N_9769);
and UO_1021 (O_1021,N_8924,N_8109);
nand UO_1022 (O_1022,N_9832,N_9821);
or UO_1023 (O_1023,N_8286,N_8566);
or UO_1024 (O_1024,N_8531,N_9103);
and UO_1025 (O_1025,N_9648,N_9085);
nor UO_1026 (O_1026,N_8794,N_8004);
nor UO_1027 (O_1027,N_9494,N_8481);
nand UO_1028 (O_1028,N_9706,N_9392);
xor UO_1029 (O_1029,N_8563,N_8828);
or UO_1030 (O_1030,N_8237,N_9796);
nand UO_1031 (O_1031,N_9777,N_9252);
or UO_1032 (O_1032,N_9617,N_8975);
or UO_1033 (O_1033,N_8938,N_9528);
or UO_1034 (O_1034,N_9701,N_8813);
nor UO_1035 (O_1035,N_8991,N_9900);
or UO_1036 (O_1036,N_8988,N_8804);
and UO_1037 (O_1037,N_9946,N_9851);
nand UO_1038 (O_1038,N_8135,N_8472);
and UO_1039 (O_1039,N_8788,N_9746);
and UO_1040 (O_1040,N_8099,N_9905);
and UO_1041 (O_1041,N_8313,N_8380);
xor UO_1042 (O_1042,N_8944,N_8218);
nor UO_1043 (O_1043,N_9208,N_9509);
and UO_1044 (O_1044,N_8469,N_8368);
nand UO_1045 (O_1045,N_9987,N_9617);
or UO_1046 (O_1046,N_9756,N_9034);
nand UO_1047 (O_1047,N_8791,N_8606);
xnor UO_1048 (O_1048,N_9209,N_8587);
or UO_1049 (O_1049,N_8165,N_8289);
and UO_1050 (O_1050,N_9649,N_8907);
xor UO_1051 (O_1051,N_9078,N_8331);
and UO_1052 (O_1052,N_9405,N_8950);
xnor UO_1053 (O_1053,N_9700,N_9984);
nand UO_1054 (O_1054,N_9302,N_8622);
or UO_1055 (O_1055,N_8643,N_9970);
or UO_1056 (O_1056,N_8885,N_8172);
or UO_1057 (O_1057,N_8795,N_8703);
or UO_1058 (O_1058,N_8541,N_9437);
and UO_1059 (O_1059,N_9601,N_9432);
or UO_1060 (O_1060,N_9142,N_8339);
or UO_1061 (O_1061,N_8408,N_8125);
nor UO_1062 (O_1062,N_8592,N_9533);
and UO_1063 (O_1063,N_9911,N_8239);
nand UO_1064 (O_1064,N_8379,N_8475);
or UO_1065 (O_1065,N_8082,N_8746);
and UO_1066 (O_1066,N_8989,N_8069);
nand UO_1067 (O_1067,N_9519,N_8566);
nor UO_1068 (O_1068,N_9956,N_8433);
or UO_1069 (O_1069,N_8653,N_9802);
or UO_1070 (O_1070,N_9078,N_8113);
and UO_1071 (O_1071,N_8484,N_8768);
or UO_1072 (O_1072,N_9106,N_8067);
nand UO_1073 (O_1073,N_9005,N_8564);
xor UO_1074 (O_1074,N_8549,N_9025);
nor UO_1075 (O_1075,N_8078,N_9264);
and UO_1076 (O_1076,N_8436,N_8395);
nor UO_1077 (O_1077,N_8319,N_8059);
or UO_1078 (O_1078,N_8719,N_9928);
xnor UO_1079 (O_1079,N_9233,N_8228);
nor UO_1080 (O_1080,N_8969,N_9163);
and UO_1081 (O_1081,N_9514,N_9395);
and UO_1082 (O_1082,N_9506,N_8445);
and UO_1083 (O_1083,N_9337,N_8816);
nor UO_1084 (O_1084,N_9747,N_9274);
and UO_1085 (O_1085,N_9605,N_9544);
and UO_1086 (O_1086,N_8771,N_9921);
and UO_1087 (O_1087,N_9503,N_8342);
and UO_1088 (O_1088,N_8244,N_9735);
nand UO_1089 (O_1089,N_8928,N_9887);
or UO_1090 (O_1090,N_8712,N_8306);
or UO_1091 (O_1091,N_9597,N_8696);
nor UO_1092 (O_1092,N_9906,N_9125);
or UO_1093 (O_1093,N_8165,N_9654);
xnor UO_1094 (O_1094,N_9519,N_8548);
nor UO_1095 (O_1095,N_8562,N_8398);
or UO_1096 (O_1096,N_8169,N_9638);
xnor UO_1097 (O_1097,N_9420,N_8809);
nor UO_1098 (O_1098,N_8183,N_9542);
nand UO_1099 (O_1099,N_8806,N_8891);
or UO_1100 (O_1100,N_9175,N_9495);
or UO_1101 (O_1101,N_8249,N_9824);
or UO_1102 (O_1102,N_8382,N_9048);
nand UO_1103 (O_1103,N_9255,N_8562);
nand UO_1104 (O_1104,N_8237,N_9516);
nor UO_1105 (O_1105,N_9368,N_9235);
xor UO_1106 (O_1106,N_8199,N_8295);
nor UO_1107 (O_1107,N_8699,N_8236);
or UO_1108 (O_1108,N_9859,N_8642);
or UO_1109 (O_1109,N_9600,N_9610);
xnor UO_1110 (O_1110,N_8009,N_9433);
or UO_1111 (O_1111,N_8435,N_9341);
nand UO_1112 (O_1112,N_9186,N_9332);
xnor UO_1113 (O_1113,N_9110,N_9187);
nand UO_1114 (O_1114,N_9645,N_9077);
and UO_1115 (O_1115,N_8323,N_9224);
nor UO_1116 (O_1116,N_8193,N_8943);
or UO_1117 (O_1117,N_9571,N_9114);
nand UO_1118 (O_1118,N_8512,N_9863);
and UO_1119 (O_1119,N_8976,N_9787);
or UO_1120 (O_1120,N_8012,N_8997);
xnor UO_1121 (O_1121,N_9595,N_9075);
and UO_1122 (O_1122,N_8300,N_9185);
and UO_1123 (O_1123,N_8431,N_8045);
or UO_1124 (O_1124,N_9026,N_8437);
nor UO_1125 (O_1125,N_9521,N_8217);
or UO_1126 (O_1126,N_8263,N_9693);
nand UO_1127 (O_1127,N_9624,N_9866);
and UO_1128 (O_1128,N_8099,N_9145);
or UO_1129 (O_1129,N_9738,N_9375);
nand UO_1130 (O_1130,N_9616,N_8984);
nor UO_1131 (O_1131,N_9090,N_8515);
nor UO_1132 (O_1132,N_9730,N_8931);
nand UO_1133 (O_1133,N_8565,N_9198);
xor UO_1134 (O_1134,N_9582,N_8165);
nor UO_1135 (O_1135,N_8856,N_9031);
nor UO_1136 (O_1136,N_8495,N_9111);
nand UO_1137 (O_1137,N_9073,N_9645);
nor UO_1138 (O_1138,N_8324,N_9121);
nand UO_1139 (O_1139,N_9940,N_8604);
or UO_1140 (O_1140,N_9297,N_9070);
and UO_1141 (O_1141,N_8669,N_9677);
or UO_1142 (O_1142,N_9191,N_8929);
nand UO_1143 (O_1143,N_9438,N_8148);
nor UO_1144 (O_1144,N_9434,N_9776);
nand UO_1145 (O_1145,N_8366,N_8309);
nor UO_1146 (O_1146,N_9399,N_9709);
or UO_1147 (O_1147,N_9263,N_8892);
nand UO_1148 (O_1148,N_9467,N_8162);
nor UO_1149 (O_1149,N_8313,N_8558);
xnor UO_1150 (O_1150,N_8422,N_8245);
nor UO_1151 (O_1151,N_8058,N_9975);
and UO_1152 (O_1152,N_8841,N_8173);
and UO_1153 (O_1153,N_8550,N_9607);
nand UO_1154 (O_1154,N_8328,N_8356);
nor UO_1155 (O_1155,N_8168,N_8320);
nand UO_1156 (O_1156,N_8299,N_8206);
or UO_1157 (O_1157,N_9591,N_8730);
nand UO_1158 (O_1158,N_9088,N_8629);
and UO_1159 (O_1159,N_8881,N_9487);
or UO_1160 (O_1160,N_9057,N_9110);
nor UO_1161 (O_1161,N_9622,N_8427);
nor UO_1162 (O_1162,N_8538,N_8137);
nand UO_1163 (O_1163,N_8642,N_8737);
or UO_1164 (O_1164,N_9764,N_9949);
nor UO_1165 (O_1165,N_8427,N_9478);
nand UO_1166 (O_1166,N_8330,N_9439);
nand UO_1167 (O_1167,N_8158,N_8397);
or UO_1168 (O_1168,N_8762,N_8738);
nor UO_1169 (O_1169,N_9190,N_9431);
nand UO_1170 (O_1170,N_9329,N_9106);
and UO_1171 (O_1171,N_9858,N_8530);
nor UO_1172 (O_1172,N_8182,N_9009);
or UO_1173 (O_1173,N_9466,N_9497);
or UO_1174 (O_1174,N_8861,N_9078);
nor UO_1175 (O_1175,N_8498,N_9186);
nand UO_1176 (O_1176,N_8401,N_8643);
and UO_1177 (O_1177,N_8513,N_8610);
nand UO_1178 (O_1178,N_8325,N_9923);
or UO_1179 (O_1179,N_9103,N_8460);
or UO_1180 (O_1180,N_9239,N_8170);
nor UO_1181 (O_1181,N_8760,N_8798);
nor UO_1182 (O_1182,N_8572,N_8118);
nand UO_1183 (O_1183,N_8239,N_9593);
nor UO_1184 (O_1184,N_9570,N_9259);
nand UO_1185 (O_1185,N_9190,N_8883);
or UO_1186 (O_1186,N_8620,N_8124);
xor UO_1187 (O_1187,N_8064,N_8220);
and UO_1188 (O_1188,N_9051,N_9251);
nand UO_1189 (O_1189,N_9815,N_8008);
or UO_1190 (O_1190,N_8548,N_8822);
nand UO_1191 (O_1191,N_9140,N_9167);
and UO_1192 (O_1192,N_8225,N_9756);
xor UO_1193 (O_1193,N_8137,N_8325);
xnor UO_1194 (O_1194,N_9895,N_9771);
nor UO_1195 (O_1195,N_8961,N_8835);
and UO_1196 (O_1196,N_9288,N_9508);
and UO_1197 (O_1197,N_9144,N_9790);
nor UO_1198 (O_1198,N_9788,N_9568);
xnor UO_1199 (O_1199,N_9012,N_8338);
or UO_1200 (O_1200,N_9964,N_8991);
or UO_1201 (O_1201,N_8867,N_8268);
nand UO_1202 (O_1202,N_9978,N_9881);
or UO_1203 (O_1203,N_8426,N_9789);
nand UO_1204 (O_1204,N_8044,N_8601);
and UO_1205 (O_1205,N_8231,N_9192);
nor UO_1206 (O_1206,N_8859,N_8514);
nor UO_1207 (O_1207,N_8878,N_9543);
and UO_1208 (O_1208,N_9833,N_9651);
and UO_1209 (O_1209,N_8930,N_9618);
nand UO_1210 (O_1210,N_8214,N_9873);
nand UO_1211 (O_1211,N_8704,N_8933);
nand UO_1212 (O_1212,N_8567,N_9583);
or UO_1213 (O_1213,N_9544,N_8043);
and UO_1214 (O_1214,N_8101,N_8450);
and UO_1215 (O_1215,N_8756,N_8382);
nand UO_1216 (O_1216,N_9316,N_9040);
and UO_1217 (O_1217,N_8631,N_9986);
and UO_1218 (O_1218,N_9467,N_9246);
nand UO_1219 (O_1219,N_8605,N_8603);
and UO_1220 (O_1220,N_8467,N_8560);
and UO_1221 (O_1221,N_8832,N_8288);
nand UO_1222 (O_1222,N_9200,N_8103);
or UO_1223 (O_1223,N_9593,N_8276);
or UO_1224 (O_1224,N_9595,N_9156);
xor UO_1225 (O_1225,N_8805,N_8874);
nor UO_1226 (O_1226,N_9552,N_9248);
xor UO_1227 (O_1227,N_8884,N_9166);
nand UO_1228 (O_1228,N_8534,N_9533);
and UO_1229 (O_1229,N_8020,N_8320);
nand UO_1230 (O_1230,N_8791,N_9973);
nor UO_1231 (O_1231,N_9867,N_9774);
xor UO_1232 (O_1232,N_9508,N_8202);
nor UO_1233 (O_1233,N_8671,N_9954);
and UO_1234 (O_1234,N_8537,N_8603);
or UO_1235 (O_1235,N_8491,N_9691);
or UO_1236 (O_1236,N_9463,N_8981);
nor UO_1237 (O_1237,N_8447,N_8927);
and UO_1238 (O_1238,N_8415,N_9747);
nor UO_1239 (O_1239,N_8377,N_8577);
xor UO_1240 (O_1240,N_8115,N_8615);
nand UO_1241 (O_1241,N_8566,N_9484);
nand UO_1242 (O_1242,N_8367,N_8240);
or UO_1243 (O_1243,N_8311,N_9141);
nand UO_1244 (O_1244,N_9810,N_9317);
nor UO_1245 (O_1245,N_9132,N_8898);
nand UO_1246 (O_1246,N_8129,N_9001);
nand UO_1247 (O_1247,N_9157,N_9120);
nand UO_1248 (O_1248,N_9136,N_8940);
nand UO_1249 (O_1249,N_8578,N_8600);
nand UO_1250 (O_1250,N_8868,N_9637);
nand UO_1251 (O_1251,N_8651,N_9021);
nor UO_1252 (O_1252,N_8455,N_8038);
nand UO_1253 (O_1253,N_9276,N_8261);
or UO_1254 (O_1254,N_8068,N_9060);
nor UO_1255 (O_1255,N_8747,N_9738);
nor UO_1256 (O_1256,N_9900,N_8113);
nand UO_1257 (O_1257,N_9949,N_8872);
nand UO_1258 (O_1258,N_8131,N_9305);
and UO_1259 (O_1259,N_8832,N_8825);
and UO_1260 (O_1260,N_8411,N_9092);
or UO_1261 (O_1261,N_9611,N_9805);
nor UO_1262 (O_1262,N_9943,N_9644);
xnor UO_1263 (O_1263,N_9260,N_9791);
nor UO_1264 (O_1264,N_9585,N_8451);
nor UO_1265 (O_1265,N_9801,N_9248);
nor UO_1266 (O_1266,N_8560,N_9834);
nand UO_1267 (O_1267,N_9174,N_8332);
or UO_1268 (O_1268,N_9519,N_8037);
nor UO_1269 (O_1269,N_8672,N_9610);
nand UO_1270 (O_1270,N_8404,N_8790);
or UO_1271 (O_1271,N_8796,N_8920);
or UO_1272 (O_1272,N_8746,N_8000);
nor UO_1273 (O_1273,N_9575,N_8222);
or UO_1274 (O_1274,N_9984,N_9462);
nor UO_1275 (O_1275,N_8390,N_8191);
nor UO_1276 (O_1276,N_8604,N_9037);
xor UO_1277 (O_1277,N_9383,N_8265);
xor UO_1278 (O_1278,N_8338,N_9520);
and UO_1279 (O_1279,N_9631,N_9916);
nand UO_1280 (O_1280,N_8496,N_8559);
nor UO_1281 (O_1281,N_8330,N_9572);
nor UO_1282 (O_1282,N_9861,N_9652);
and UO_1283 (O_1283,N_8360,N_8820);
nor UO_1284 (O_1284,N_9595,N_8939);
or UO_1285 (O_1285,N_9226,N_9420);
and UO_1286 (O_1286,N_9686,N_9585);
and UO_1287 (O_1287,N_8139,N_9922);
nor UO_1288 (O_1288,N_8511,N_8680);
nor UO_1289 (O_1289,N_8018,N_9194);
and UO_1290 (O_1290,N_8452,N_8335);
xor UO_1291 (O_1291,N_9145,N_8585);
or UO_1292 (O_1292,N_9661,N_9827);
and UO_1293 (O_1293,N_9966,N_9634);
xor UO_1294 (O_1294,N_9573,N_9085);
nor UO_1295 (O_1295,N_9051,N_9062);
and UO_1296 (O_1296,N_9451,N_9792);
and UO_1297 (O_1297,N_8684,N_9236);
or UO_1298 (O_1298,N_8687,N_9761);
nand UO_1299 (O_1299,N_8453,N_8834);
and UO_1300 (O_1300,N_8848,N_9113);
xor UO_1301 (O_1301,N_8937,N_8897);
nor UO_1302 (O_1302,N_9643,N_9864);
nor UO_1303 (O_1303,N_8897,N_9361);
and UO_1304 (O_1304,N_9345,N_8929);
or UO_1305 (O_1305,N_8933,N_9914);
nand UO_1306 (O_1306,N_9229,N_8107);
nand UO_1307 (O_1307,N_8725,N_9969);
or UO_1308 (O_1308,N_9006,N_8737);
and UO_1309 (O_1309,N_9022,N_9967);
xor UO_1310 (O_1310,N_8489,N_8067);
and UO_1311 (O_1311,N_8634,N_8279);
nand UO_1312 (O_1312,N_8391,N_9495);
and UO_1313 (O_1313,N_9705,N_9382);
nand UO_1314 (O_1314,N_9345,N_9793);
and UO_1315 (O_1315,N_9187,N_9014);
nand UO_1316 (O_1316,N_9417,N_9450);
or UO_1317 (O_1317,N_8194,N_9002);
nand UO_1318 (O_1318,N_9107,N_9788);
xnor UO_1319 (O_1319,N_9377,N_9132);
nand UO_1320 (O_1320,N_9264,N_8378);
or UO_1321 (O_1321,N_9314,N_8699);
nand UO_1322 (O_1322,N_8222,N_8186);
or UO_1323 (O_1323,N_8381,N_8506);
nand UO_1324 (O_1324,N_8554,N_9590);
nor UO_1325 (O_1325,N_8960,N_8786);
nor UO_1326 (O_1326,N_9997,N_8877);
and UO_1327 (O_1327,N_8201,N_8849);
nor UO_1328 (O_1328,N_8113,N_8923);
xor UO_1329 (O_1329,N_9590,N_9275);
and UO_1330 (O_1330,N_9750,N_8604);
or UO_1331 (O_1331,N_9848,N_8924);
and UO_1332 (O_1332,N_8212,N_8474);
or UO_1333 (O_1333,N_9224,N_8850);
nand UO_1334 (O_1334,N_9508,N_8122);
nor UO_1335 (O_1335,N_9320,N_9053);
nor UO_1336 (O_1336,N_8916,N_9828);
or UO_1337 (O_1337,N_9456,N_8629);
xnor UO_1338 (O_1338,N_9181,N_9339);
or UO_1339 (O_1339,N_8364,N_8748);
xor UO_1340 (O_1340,N_9013,N_9974);
and UO_1341 (O_1341,N_9168,N_8748);
xor UO_1342 (O_1342,N_8751,N_8779);
nand UO_1343 (O_1343,N_8719,N_9356);
and UO_1344 (O_1344,N_9831,N_9268);
nand UO_1345 (O_1345,N_9317,N_9870);
or UO_1346 (O_1346,N_9925,N_9274);
and UO_1347 (O_1347,N_9089,N_8428);
nor UO_1348 (O_1348,N_8403,N_8743);
or UO_1349 (O_1349,N_9856,N_8318);
nor UO_1350 (O_1350,N_9311,N_8549);
nor UO_1351 (O_1351,N_8652,N_9121);
and UO_1352 (O_1352,N_8317,N_8473);
nand UO_1353 (O_1353,N_9437,N_9440);
nand UO_1354 (O_1354,N_9857,N_8154);
or UO_1355 (O_1355,N_9675,N_9084);
nand UO_1356 (O_1356,N_8378,N_9726);
and UO_1357 (O_1357,N_8321,N_9611);
and UO_1358 (O_1358,N_9620,N_8806);
or UO_1359 (O_1359,N_9833,N_9978);
nor UO_1360 (O_1360,N_8032,N_8036);
or UO_1361 (O_1361,N_8166,N_9190);
nor UO_1362 (O_1362,N_8551,N_9972);
and UO_1363 (O_1363,N_9718,N_9596);
nor UO_1364 (O_1364,N_8405,N_9410);
or UO_1365 (O_1365,N_8189,N_9547);
nand UO_1366 (O_1366,N_8713,N_8786);
or UO_1367 (O_1367,N_8364,N_8916);
nor UO_1368 (O_1368,N_9281,N_8622);
nor UO_1369 (O_1369,N_8590,N_9843);
xnor UO_1370 (O_1370,N_8279,N_8574);
nor UO_1371 (O_1371,N_8882,N_9204);
xnor UO_1372 (O_1372,N_8598,N_9291);
nand UO_1373 (O_1373,N_8655,N_8157);
nand UO_1374 (O_1374,N_9075,N_8731);
nand UO_1375 (O_1375,N_9995,N_9450);
and UO_1376 (O_1376,N_8954,N_8371);
or UO_1377 (O_1377,N_9682,N_9588);
nand UO_1378 (O_1378,N_8588,N_9896);
or UO_1379 (O_1379,N_8978,N_9237);
nor UO_1380 (O_1380,N_9851,N_9090);
xnor UO_1381 (O_1381,N_9552,N_9196);
and UO_1382 (O_1382,N_9446,N_9708);
or UO_1383 (O_1383,N_8642,N_8607);
nand UO_1384 (O_1384,N_8299,N_9333);
nand UO_1385 (O_1385,N_9335,N_8211);
or UO_1386 (O_1386,N_8898,N_9565);
nand UO_1387 (O_1387,N_8019,N_8582);
nand UO_1388 (O_1388,N_8735,N_8061);
nor UO_1389 (O_1389,N_9714,N_8045);
or UO_1390 (O_1390,N_9035,N_8805);
xnor UO_1391 (O_1391,N_8955,N_9759);
nor UO_1392 (O_1392,N_8199,N_9846);
nor UO_1393 (O_1393,N_9432,N_9077);
or UO_1394 (O_1394,N_9618,N_8317);
nand UO_1395 (O_1395,N_8248,N_9995);
and UO_1396 (O_1396,N_8200,N_8000);
xnor UO_1397 (O_1397,N_8727,N_9504);
or UO_1398 (O_1398,N_9415,N_8441);
nor UO_1399 (O_1399,N_9614,N_8570);
xnor UO_1400 (O_1400,N_9177,N_8093);
xor UO_1401 (O_1401,N_9439,N_9344);
or UO_1402 (O_1402,N_8841,N_9117);
nand UO_1403 (O_1403,N_9488,N_8672);
and UO_1404 (O_1404,N_9028,N_9395);
nor UO_1405 (O_1405,N_8106,N_9905);
nand UO_1406 (O_1406,N_8499,N_9599);
or UO_1407 (O_1407,N_9661,N_9159);
or UO_1408 (O_1408,N_9946,N_9167);
nor UO_1409 (O_1409,N_9739,N_9520);
nor UO_1410 (O_1410,N_9812,N_9140);
nor UO_1411 (O_1411,N_8594,N_9054);
xor UO_1412 (O_1412,N_8808,N_8036);
nand UO_1413 (O_1413,N_8451,N_9040);
xor UO_1414 (O_1414,N_8932,N_8023);
nand UO_1415 (O_1415,N_9211,N_8553);
nor UO_1416 (O_1416,N_9466,N_8568);
or UO_1417 (O_1417,N_9406,N_8539);
or UO_1418 (O_1418,N_8139,N_9260);
and UO_1419 (O_1419,N_9999,N_8442);
nor UO_1420 (O_1420,N_8936,N_9971);
xor UO_1421 (O_1421,N_8691,N_9896);
or UO_1422 (O_1422,N_8470,N_8545);
nor UO_1423 (O_1423,N_8086,N_8032);
and UO_1424 (O_1424,N_8659,N_9588);
xor UO_1425 (O_1425,N_9300,N_9088);
or UO_1426 (O_1426,N_8841,N_8906);
xor UO_1427 (O_1427,N_9356,N_8088);
and UO_1428 (O_1428,N_8293,N_9243);
and UO_1429 (O_1429,N_8038,N_8563);
and UO_1430 (O_1430,N_8385,N_8444);
or UO_1431 (O_1431,N_9163,N_9310);
nand UO_1432 (O_1432,N_9709,N_9225);
or UO_1433 (O_1433,N_8200,N_8431);
nor UO_1434 (O_1434,N_8550,N_9876);
and UO_1435 (O_1435,N_9293,N_8783);
nor UO_1436 (O_1436,N_8450,N_8366);
nand UO_1437 (O_1437,N_9112,N_8268);
xnor UO_1438 (O_1438,N_8246,N_9028);
xor UO_1439 (O_1439,N_9644,N_8629);
xnor UO_1440 (O_1440,N_8126,N_9486);
xor UO_1441 (O_1441,N_8856,N_8235);
or UO_1442 (O_1442,N_8254,N_8645);
nor UO_1443 (O_1443,N_8111,N_9864);
and UO_1444 (O_1444,N_9843,N_9364);
nand UO_1445 (O_1445,N_9506,N_8743);
and UO_1446 (O_1446,N_9679,N_8978);
and UO_1447 (O_1447,N_8086,N_8479);
and UO_1448 (O_1448,N_9748,N_9805);
or UO_1449 (O_1449,N_8963,N_9603);
nand UO_1450 (O_1450,N_8674,N_8168);
nor UO_1451 (O_1451,N_9394,N_9278);
or UO_1452 (O_1452,N_9018,N_9295);
and UO_1453 (O_1453,N_8422,N_9750);
nand UO_1454 (O_1454,N_8158,N_9848);
nand UO_1455 (O_1455,N_8362,N_9383);
and UO_1456 (O_1456,N_9625,N_9770);
or UO_1457 (O_1457,N_9404,N_9120);
nor UO_1458 (O_1458,N_9515,N_8579);
nand UO_1459 (O_1459,N_9886,N_8818);
nor UO_1460 (O_1460,N_9241,N_8072);
nor UO_1461 (O_1461,N_8179,N_8917);
or UO_1462 (O_1462,N_9757,N_8573);
or UO_1463 (O_1463,N_8167,N_8444);
or UO_1464 (O_1464,N_9281,N_9517);
nand UO_1465 (O_1465,N_9751,N_9797);
nand UO_1466 (O_1466,N_8910,N_9021);
nand UO_1467 (O_1467,N_8534,N_9305);
and UO_1468 (O_1468,N_9891,N_8610);
and UO_1469 (O_1469,N_9778,N_8188);
nand UO_1470 (O_1470,N_8756,N_8617);
nand UO_1471 (O_1471,N_8318,N_9237);
or UO_1472 (O_1472,N_8979,N_9921);
and UO_1473 (O_1473,N_8841,N_8790);
nor UO_1474 (O_1474,N_9450,N_8542);
nor UO_1475 (O_1475,N_9391,N_9063);
nor UO_1476 (O_1476,N_9723,N_9199);
and UO_1477 (O_1477,N_8196,N_8703);
xnor UO_1478 (O_1478,N_8655,N_9391);
or UO_1479 (O_1479,N_9972,N_9341);
nand UO_1480 (O_1480,N_8166,N_8742);
or UO_1481 (O_1481,N_8621,N_9581);
and UO_1482 (O_1482,N_8457,N_8212);
or UO_1483 (O_1483,N_8910,N_9042);
nand UO_1484 (O_1484,N_8578,N_8774);
or UO_1485 (O_1485,N_9339,N_9176);
xor UO_1486 (O_1486,N_9479,N_9820);
nand UO_1487 (O_1487,N_9640,N_9367);
nor UO_1488 (O_1488,N_8398,N_9737);
nand UO_1489 (O_1489,N_8412,N_8161);
nor UO_1490 (O_1490,N_9300,N_9242);
and UO_1491 (O_1491,N_8998,N_9613);
xnor UO_1492 (O_1492,N_9475,N_8100);
xnor UO_1493 (O_1493,N_9390,N_8186);
nor UO_1494 (O_1494,N_8037,N_8482);
or UO_1495 (O_1495,N_8238,N_8492);
or UO_1496 (O_1496,N_9281,N_9801);
nor UO_1497 (O_1497,N_9061,N_9111);
nor UO_1498 (O_1498,N_9812,N_8764);
xnor UO_1499 (O_1499,N_9421,N_9535);
endmodule