module basic_2000_20000_2500_50_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xnor U0 (N_0,In_1606,In_568);
nor U1 (N_1,In_1704,In_217);
or U2 (N_2,In_500,In_1556);
and U3 (N_3,In_431,In_1714);
nand U4 (N_4,In_716,In_841);
and U5 (N_5,In_222,In_1375);
nor U6 (N_6,In_1695,In_1669);
and U7 (N_7,In_119,In_1931);
xor U8 (N_8,In_1469,In_1200);
and U9 (N_9,In_1333,In_984);
or U10 (N_10,In_871,In_408);
xnor U11 (N_11,In_1531,In_619);
xnor U12 (N_12,In_1829,In_1914);
xnor U13 (N_13,In_1495,In_985);
or U14 (N_14,In_1516,In_822);
nor U15 (N_15,In_1102,In_668);
and U16 (N_16,In_1786,In_116);
nor U17 (N_17,In_1872,In_1146);
nand U18 (N_18,In_70,In_1559);
nor U19 (N_19,In_1944,In_1153);
nor U20 (N_20,In_1139,In_862);
xnor U21 (N_21,In_977,In_1911);
nor U22 (N_22,In_115,In_461);
xor U23 (N_23,In_1848,In_953);
nor U24 (N_24,In_875,In_760);
nor U25 (N_25,In_979,In_368);
nand U26 (N_26,In_1191,In_316);
nor U27 (N_27,In_1756,In_1255);
xor U28 (N_28,In_1710,In_1780);
xnor U29 (N_29,In_1818,In_1446);
and U30 (N_30,In_750,In_1171);
nor U31 (N_31,In_53,In_166);
or U32 (N_32,In_48,In_1048);
nor U33 (N_33,In_663,In_1555);
nor U34 (N_34,In_880,In_1128);
xnor U35 (N_35,In_1750,In_1765);
nand U36 (N_36,In_1697,In_1712);
nand U37 (N_37,In_1003,In_302);
nand U38 (N_38,In_318,In_739);
and U39 (N_39,In_653,In_1465);
xnor U40 (N_40,In_417,In_1511);
nor U41 (N_41,In_343,In_1239);
nand U42 (N_42,In_208,In_1185);
nor U43 (N_43,In_136,In_375);
or U44 (N_44,In_349,In_891);
and U45 (N_45,In_83,In_1973);
nand U46 (N_46,In_28,In_1266);
xor U47 (N_47,In_1376,In_602);
and U48 (N_48,In_697,In_1194);
or U49 (N_49,In_1863,In_873);
nor U50 (N_50,In_978,In_1478);
nand U51 (N_51,In_1644,In_1915);
or U52 (N_52,In_1135,In_1419);
and U53 (N_53,In_1421,In_694);
nand U54 (N_54,In_1213,In_596);
nor U55 (N_55,In_1783,In_341);
nor U56 (N_56,In_1834,In_1594);
nand U57 (N_57,In_1089,In_689);
or U58 (N_58,In_1462,In_1209);
xor U59 (N_59,In_1835,In_1387);
xor U60 (N_60,In_198,In_882);
nor U61 (N_61,In_1691,In_403);
and U62 (N_62,In_1051,In_929);
and U63 (N_63,In_877,In_1867);
or U64 (N_64,In_1988,In_1832);
or U65 (N_65,In_1242,In_1836);
xnor U66 (N_66,In_27,In_1345);
or U67 (N_67,In_453,In_1002);
or U68 (N_68,In_845,In_1087);
nor U69 (N_69,In_1943,In_39);
nor U70 (N_70,In_272,In_1916);
nand U71 (N_71,In_1922,In_1875);
and U72 (N_72,In_502,In_179);
and U73 (N_73,In_129,In_1106);
xnor U74 (N_74,In_1251,In_279);
and U75 (N_75,In_571,In_575);
nand U76 (N_76,In_1974,In_838);
nand U77 (N_77,In_1958,In_815);
nor U78 (N_78,In_1389,In_935);
xor U79 (N_79,In_68,In_1796);
and U80 (N_80,In_128,In_738);
xnor U81 (N_81,In_1014,In_510);
and U82 (N_82,In_1463,In_1535);
nand U83 (N_83,In_1711,In_567);
or U84 (N_84,In_324,In_1521);
and U85 (N_85,In_1476,In_1184);
xnor U86 (N_86,In_1605,In_487);
and U87 (N_87,In_491,In_329);
nor U88 (N_88,In_181,In_586);
xor U89 (N_89,In_856,In_1634);
nor U90 (N_90,In_1212,In_614);
or U91 (N_91,In_1777,In_1530);
or U92 (N_92,In_1949,In_295);
and U93 (N_93,In_226,In_418);
nand U94 (N_94,In_162,In_147);
nand U95 (N_95,In_1891,In_1533);
or U96 (N_96,In_1545,In_1764);
and U97 (N_97,In_1405,In_553);
or U98 (N_98,In_1201,In_958);
or U99 (N_99,In_1055,In_1896);
nand U100 (N_100,In_1932,In_1151);
or U101 (N_101,In_168,In_534);
and U102 (N_102,In_1668,In_737);
or U103 (N_103,In_1580,In_1284);
or U104 (N_104,In_1698,In_827);
xnor U105 (N_105,In_1553,In_1587);
xor U106 (N_106,In_661,In_1012);
nand U107 (N_107,In_92,In_851);
xor U108 (N_108,In_949,In_1134);
nor U109 (N_109,In_1293,In_522);
xnor U110 (N_110,In_1276,In_1913);
and U111 (N_111,In_1772,In_701);
nand U112 (N_112,In_693,In_429);
xor U113 (N_113,In_687,In_1941);
xor U114 (N_114,In_1554,In_1402);
and U115 (N_115,In_1850,In_299);
xnor U116 (N_116,In_347,In_1379);
nand U117 (N_117,In_1749,In_247);
nand U118 (N_118,In_564,In_1787);
or U119 (N_119,In_1100,In_243);
xnor U120 (N_120,In_1391,In_1329);
and U121 (N_121,In_538,In_1203);
and U122 (N_122,In_1022,In_1408);
nand U123 (N_123,In_598,In_1315);
nand U124 (N_124,In_1013,In_1600);
xnor U125 (N_125,In_0,In_1444);
nand U126 (N_126,In_326,In_1456);
xnor U127 (N_127,In_1884,In_1149);
nand U128 (N_128,In_1466,In_894);
or U129 (N_129,In_1997,In_1240);
xor U130 (N_130,In_1803,In_1534);
xnor U131 (N_131,In_266,In_1053);
and U132 (N_132,In_806,In_886);
xor U133 (N_133,In_1497,In_350);
xor U134 (N_134,In_1038,In_1720);
nand U135 (N_135,In_42,In_1674);
nor U136 (N_136,In_997,In_164);
nor U137 (N_137,In_1339,In_37);
and U138 (N_138,In_847,In_145);
nor U139 (N_139,In_358,In_910);
nor U140 (N_140,In_323,In_1437);
nor U141 (N_141,In_764,In_855);
xor U142 (N_142,In_1541,In_629);
or U143 (N_143,In_808,In_36);
xnor U144 (N_144,In_853,In_742);
nand U145 (N_145,In_1570,In_1747);
nor U146 (N_146,In_612,In_646);
nor U147 (N_147,In_1621,In_1813);
nand U148 (N_148,In_1853,In_455);
nand U149 (N_149,In_1581,In_913);
and U150 (N_150,In_816,In_259);
xnor U151 (N_151,In_98,In_1532);
nor U152 (N_152,In_1847,In_576);
nor U153 (N_153,In_526,In_63);
nor U154 (N_154,In_1589,In_700);
xnor U155 (N_155,In_1342,In_938);
and U156 (N_156,In_1340,In_1385);
xnor U157 (N_157,In_157,In_1748);
xnor U158 (N_158,In_321,In_1833);
xnor U159 (N_159,In_19,In_71);
and U160 (N_160,In_15,In_496);
xnor U161 (N_161,In_1152,In_1991);
nor U162 (N_162,In_830,In_1394);
nor U163 (N_163,In_1373,In_1027);
xor U164 (N_164,In_351,In_747);
or U165 (N_165,In_1309,In_1138);
or U166 (N_166,In_398,In_1348);
and U167 (N_167,In_695,In_1977);
nor U168 (N_168,In_1649,In_263);
nor U169 (N_169,In_1507,In_789);
nand U170 (N_170,In_959,In_1679);
nand U171 (N_171,In_1283,In_401);
nand U172 (N_172,In_1295,In_1671);
nor U173 (N_173,In_138,In_1114);
xnor U174 (N_174,In_260,In_99);
xor U175 (N_175,In_1393,In_1418);
and U176 (N_176,In_1980,In_1816);
and U177 (N_177,In_623,In_1214);
nor U178 (N_178,In_1677,In_1351);
nand U179 (N_179,In_1039,In_748);
or U180 (N_180,In_276,In_1252);
nand U181 (N_181,In_190,In_1886);
or U182 (N_182,In_1091,In_963);
nand U183 (N_183,In_369,In_112);
xor U184 (N_184,In_1860,In_647);
nor U185 (N_185,In_21,In_1945);
or U186 (N_186,In_973,In_199);
and U187 (N_187,In_892,In_665);
nor U188 (N_188,In_1312,In_559);
xnor U189 (N_189,In_1180,In_727);
nor U190 (N_190,In_1494,In_471);
and U191 (N_191,In_1007,In_723);
xor U192 (N_192,In_139,In_1036);
nor U193 (N_193,In_627,In_656);
xnor U194 (N_194,In_1707,In_1604);
and U195 (N_195,In_1414,In_1936);
xor U196 (N_196,In_834,In_187);
xor U197 (N_197,In_1830,In_1121);
xnor U198 (N_198,In_1107,In_757);
xor U199 (N_199,In_1360,In_896);
nand U200 (N_200,In_1410,In_223);
or U201 (N_201,In_1186,In_545);
xor U202 (N_202,In_241,In_1726);
or U203 (N_203,In_783,In_1500);
nand U204 (N_204,In_282,In_885);
nor U205 (N_205,In_122,In_1820);
or U206 (N_206,In_183,In_585);
xnor U207 (N_207,In_391,In_1618);
or U208 (N_208,In_460,In_1841);
xor U209 (N_209,In_1609,In_813);
xnor U210 (N_210,In_952,In_483);
nand U211 (N_211,In_1355,In_1996);
nand U212 (N_212,In_409,In_1208);
xor U213 (N_213,In_1520,In_1095);
or U214 (N_214,In_717,In_1064);
xnor U215 (N_215,In_943,In_1565);
nand U216 (N_216,In_5,In_1613);
nand U217 (N_217,In_1804,In_881);
nand U218 (N_218,In_1093,In_1165);
xnor U219 (N_219,In_1739,In_710);
nand U220 (N_220,In_1072,In_1573);
xor U221 (N_221,In_163,In_1705);
xor U222 (N_222,In_599,In_579);
nand U223 (N_223,In_721,In_1727);
and U224 (N_224,In_609,In_1612);
and U225 (N_225,In_1751,In_923);
or U226 (N_226,In_1904,In_308);
or U227 (N_227,In_558,In_1978);
xnor U228 (N_228,In_174,In_640);
and U229 (N_229,In_327,In_1682);
and U230 (N_230,In_580,In_1862);
xnor U231 (N_231,In_1399,In_776);
nand U232 (N_232,In_311,In_50);
or U233 (N_233,In_1985,In_1524);
xor U234 (N_234,In_74,In_758);
xnor U235 (N_235,In_1096,In_44);
nand U236 (N_236,In_879,In_137);
nand U237 (N_237,In_1837,In_1322);
and U238 (N_238,In_1032,In_459);
xnor U239 (N_239,In_1983,In_519);
xor U240 (N_240,In_56,In_901);
or U241 (N_241,In_1610,In_1912);
and U242 (N_242,In_11,In_1386);
or U243 (N_243,In_1549,In_546);
and U244 (N_244,In_535,In_273);
or U245 (N_245,In_1859,In_986);
xnor U246 (N_246,In_1031,In_798);
nand U247 (N_247,In_336,In_1784);
and U248 (N_248,In_1488,In_1718);
nand U249 (N_249,In_792,In_992);
nand U250 (N_250,In_837,In_1041);
nand U251 (N_251,In_312,In_1407);
xor U252 (N_252,In_1449,In_1241);
nor U253 (N_253,In_1332,In_107);
and U254 (N_254,In_968,In_306);
or U255 (N_255,In_540,In_1287);
xnor U256 (N_256,In_672,In_1008);
xnor U257 (N_257,In_172,In_1127);
xor U258 (N_258,In_1046,In_509);
and U259 (N_259,In_607,In_69);
nor U260 (N_260,In_1177,In_1131);
and U261 (N_261,In_1023,In_1908);
nand U262 (N_262,In_682,In_1797);
or U263 (N_263,In_1249,In_994);
nand U264 (N_264,In_1737,In_1626);
or U265 (N_265,In_1229,In_1652);
nand U266 (N_266,In_1642,In_1189);
or U267 (N_267,In_313,In_604);
xnor U268 (N_268,In_1793,In_1415);
nor U269 (N_269,In_1432,In_594);
or U270 (N_270,In_1665,In_1044);
and U271 (N_271,In_307,In_1546);
xor U272 (N_272,In_246,In_1263);
nand U273 (N_273,In_1164,In_1261);
xor U274 (N_274,In_1368,In_876);
nor U275 (N_275,In_280,In_1771);
nand U276 (N_276,In_1403,In_205);
and U277 (N_277,In_231,In_632);
and U278 (N_278,In_52,In_1489);
or U279 (N_279,In_819,In_1715);
xnor U280 (N_280,In_613,In_1721);
xnor U281 (N_281,In_503,In_1412);
and U282 (N_282,In_895,In_230);
nand U283 (N_283,In_1272,In_1431);
or U284 (N_284,In_761,In_652);
nand U285 (N_285,In_1130,In_152);
nand U286 (N_286,In_1075,In_383);
and U287 (N_287,In_1986,In_1150);
xor U288 (N_288,In_1819,In_1708);
nor U289 (N_289,In_1817,In_1956);
and U290 (N_290,In_946,In_1951);
and U291 (N_291,In_1330,In_642);
xor U292 (N_292,In_1125,In_1752);
xor U293 (N_293,In_645,In_447);
xor U294 (N_294,In_1159,In_1390);
nor U295 (N_295,In_531,In_1675);
nand U296 (N_296,In_440,In_1893);
nand U297 (N_297,In_1105,In_622);
xnor U298 (N_298,In_319,In_96);
and U299 (N_299,In_188,In_1248);
nor U300 (N_300,In_592,In_269);
or U301 (N_301,In_775,In_328);
xor U302 (N_302,In_1890,In_1745);
or U303 (N_303,In_10,In_823);
nor U304 (N_304,In_1527,In_1923);
nor U305 (N_305,In_511,In_557);
nand U306 (N_306,In_1047,In_1145);
or U307 (N_307,In_1901,In_651);
or U308 (N_308,In_1948,In_1592);
nand U309 (N_309,In_1919,In_1232);
nand U310 (N_310,In_826,In_920);
xor U311 (N_311,In_330,In_244);
xnor U312 (N_312,In_1499,In_472);
and U313 (N_313,In_1597,In_624);
nor U314 (N_314,In_846,In_1320);
nor U315 (N_315,In_974,In_463);
xor U316 (N_316,In_1078,In_805);
nand U317 (N_317,In_1030,In_61);
nand U318 (N_318,In_1111,In_488);
or U319 (N_319,In_593,In_1660);
or U320 (N_320,In_1323,In_1924);
xor U321 (N_321,In_1289,In_987);
or U322 (N_322,In_1103,In_1987);
and U323 (N_323,In_1979,In_449);
and U324 (N_324,In_1506,In_634);
nor U325 (N_325,In_141,In_692);
and U326 (N_326,In_1801,In_659);
nand U327 (N_327,In_1805,In_1493);
and U328 (N_328,In_1370,In_444);
or U329 (N_329,In_26,In_1243);
or U330 (N_330,In_786,In_79);
nand U331 (N_331,In_671,In_667);
or U332 (N_332,In_1733,In_1955);
nor U333 (N_333,In_1730,In_1004);
and U334 (N_334,In_1616,In_591);
nor U335 (N_335,In_541,In_255);
nor U336 (N_336,In_1678,In_1477);
nand U337 (N_337,In_1062,In_338);
xnor U338 (N_338,In_78,In_1961);
xnor U339 (N_339,In_412,In_1857);
and U340 (N_340,In_184,In_560);
and U341 (N_341,In_466,In_1080);
or U342 (N_342,In_774,In_1161);
xor U343 (N_343,In_490,In_1785);
and U344 (N_344,In_1338,In_1880);
nor U345 (N_345,In_497,In_911);
xor U346 (N_346,In_1350,In_1663);
nand U347 (N_347,In_1868,In_1074);
nand U348 (N_348,In_345,In_600);
nand U349 (N_349,In_960,In_309);
or U350 (N_350,In_1256,In_1356);
or U351 (N_351,In_334,In_698);
nor U352 (N_352,In_1349,In_915);
xor U353 (N_353,In_722,In_8);
or U354 (N_354,In_1754,In_1098);
or U355 (N_355,In_196,In_288);
nand U356 (N_356,In_512,In_1503);
xor U357 (N_357,In_1066,In_1092);
and U358 (N_358,In_353,In_569);
or U359 (N_359,In_228,In_1197);
and U360 (N_360,In_1434,In_1845);
xor U361 (N_361,In_220,In_1811);
and U362 (N_362,In_1906,In_1380);
or U363 (N_363,In_1158,In_339);
xor U364 (N_364,In_1362,In_1395);
nand U365 (N_365,In_1118,In_521);
or U366 (N_366,In_724,In_696);
nand U367 (N_367,In_1167,In_1190);
or U368 (N_368,In_756,In_373);
xor U369 (N_369,In_211,In_1547);
nand U370 (N_370,In_1451,In_1426);
and U371 (N_371,In_1473,In_1578);
xor U372 (N_372,In_1846,In_513);
or U373 (N_373,In_1006,In_31);
and U374 (N_374,In_1404,In_1398);
and U375 (N_375,In_293,In_1552);
xnor U376 (N_376,In_850,In_1);
and U377 (N_377,In_989,In_1328);
nand U378 (N_378,In_1821,In_478);
or U379 (N_379,In_1800,In_411);
and U380 (N_380,In_1228,In_180);
xor U381 (N_381,In_527,In_1439);
xor U382 (N_382,In_1353,In_930);
or U383 (N_383,In_990,In_110);
or U384 (N_384,In_961,In_1441);
nor U385 (N_385,In_1540,In_908);
nor U386 (N_386,In_1265,In_1170);
xnor U387 (N_387,In_1172,In_888);
and U388 (N_388,In_1822,In_485);
nor U389 (N_389,In_1782,In_1060);
and U390 (N_390,In_1575,In_736);
xnor U391 (N_391,In_421,In_104);
and U392 (N_392,In_215,In_1166);
nor U393 (N_393,In_1043,In_45);
nand U394 (N_394,In_1005,In_884);
nor U395 (N_395,In_883,In_1728);
and U396 (N_396,In_1067,In_572);
nor U397 (N_397,In_1672,In_257);
and U398 (N_398,In_1651,In_499);
nor U399 (N_399,In_772,In_1938);
and U400 (N_400,In_1928,In_1684);
nand U401 (N_401,N_176,In_611);
or U402 (N_402,In_237,In_1598);
nand U403 (N_403,In_1779,N_50);
and U404 (N_404,N_20,N_229);
nand U405 (N_405,N_138,In_479);
or U406 (N_406,In_673,N_35);
nor U407 (N_407,In_155,In_1723);
xnor U408 (N_408,In_1761,In_530);
xnor U409 (N_409,In_242,N_362);
or U410 (N_410,In_457,N_368);
xnor U411 (N_411,In_718,In_1318);
or U412 (N_412,In_918,In_554);
and U413 (N_413,In_67,N_204);
nand U414 (N_414,In_1085,In_870);
nor U415 (N_415,In_945,In_1601);
or U416 (N_416,In_1878,In_404);
xor U417 (N_417,In_1020,In_1174);
xor U418 (N_418,In_1069,In_941);
xor U419 (N_419,In_1016,In_590);
and U420 (N_420,In_1560,In_1422);
xnor U421 (N_421,In_1420,In_844);
nor U422 (N_422,In_1413,In_1492);
or U423 (N_423,In_381,In_286);
nor U424 (N_424,In_1781,N_161);
nor U425 (N_425,In_836,N_129);
xor U426 (N_426,In_1812,In_1133);
and U427 (N_427,In_1425,N_391);
and U428 (N_428,N_381,In_317);
xnor U429 (N_429,In_254,In_705);
and U430 (N_430,In_389,In_386);
xnor U431 (N_431,N_183,In_1480);
xnor U432 (N_432,N_133,In_1231);
and U433 (N_433,In_674,N_168);
nand U434 (N_434,In_1537,N_252);
xor U435 (N_435,N_237,In_1686);
nand U436 (N_436,N_360,In_1400);
or U437 (N_437,N_172,In_548);
and U438 (N_438,N_122,In_1490);
and U439 (N_439,In_144,In_1505);
or U440 (N_440,In_420,In_1094);
nand U441 (N_441,In_897,N_38);
nor U442 (N_442,In_523,In_1467);
nand U443 (N_443,In_73,In_1648);
nor U444 (N_444,N_112,N_126);
nand U445 (N_445,N_17,In_1579);
or U446 (N_446,N_103,N_119);
nor U447 (N_447,In_1964,N_349);
or U448 (N_448,In_236,N_353);
and U449 (N_449,In_702,N_175);
or U450 (N_450,In_514,In_426);
nor U451 (N_451,N_181,In_1713);
xnor U452 (N_452,In_456,N_359);
xor U453 (N_453,In_1319,In_66);
nand U454 (N_454,In_926,N_207);
nor U455 (N_455,N_146,In_1258);
xor U456 (N_456,In_1759,In_1461);
and U457 (N_457,In_1742,In_1794);
nor U458 (N_458,N_210,In_785);
nand U459 (N_459,In_265,In_189);
or U460 (N_460,In_1316,N_66);
xnor U461 (N_461,In_1306,In_800);
or U462 (N_462,In_1192,N_162);
xor U463 (N_463,N_385,In_1343);
or U464 (N_464,N_64,In_708);
or U465 (N_465,N_219,In_1934);
nand U466 (N_466,N_124,In_1468);
nand U467 (N_467,In_1104,In_197);
nor U468 (N_468,N_281,In_1282);
xnor U469 (N_469,In_1603,In_762);
or U470 (N_470,In_648,In_270);
nand U471 (N_471,In_1484,In_1169);
and U472 (N_472,N_334,In_1544);
nand U473 (N_473,In_956,In_1654);
or U474 (N_474,N_167,In_161);
nor U475 (N_475,In_1971,In_1851);
or U476 (N_476,In_146,In_108);
nor U477 (N_477,N_72,In_1876);
and U478 (N_478,N_282,In_1994);
nor U479 (N_479,N_163,In_264);
nand U480 (N_480,In_1314,In_900);
or U481 (N_481,In_962,In_12);
nor U482 (N_482,N_141,In_506);
nor U483 (N_483,In_1253,In_749);
nand U484 (N_484,In_356,In_176);
and U485 (N_485,In_473,In_33);
or U486 (N_486,In_1308,In_843);
xnor U487 (N_487,In_1696,N_248);
and U488 (N_488,In_238,In_1061);
xnor U489 (N_489,N_285,In_1302);
or U490 (N_490,N_102,In_1551);
nor U491 (N_491,In_781,N_398);
or U492 (N_492,In_556,In_729);
nand U493 (N_493,In_16,N_177);
nor U494 (N_494,In_928,In_711);
nand U495 (N_495,N_107,In_258);
xnor U496 (N_496,N_4,In_993);
nand U497 (N_497,In_1155,In_799);
nor U498 (N_498,N_260,In_1635);
or U499 (N_499,In_706,In_1457);
nand U500 (N_500,In_1963,In_388);
and U501 (N_501,N_155,In_1296);
nor U502 (N_502,In_520,In_224);
xnor U503 (N_503,In_818,In_1501);
nand U504 (N_504,N_91,In_1147);
or U505 (N_505,In_159,In_638);
nor U506 (N_506,N_256,In_423);
and U507 (N_507,In_34,N_232);
and U508 (N_508,In_1869,In_641);
and U509 (N_509,In_290,In_1357);
nor U510 (N_510,In_1753,In_1854);
nand U511 (N_511,In_763,In_1861);
xor U512 (N_512,In_86,In_1992);
xor U513 (N_513,In_1337,In_1278);
and U514 (N_514,In_858,In_1143);
nand U515 (N_515,In_1870,In_1388);
nand U516 (N_516,In_1548,In_1940);
and U517 (N_517,In_1815,In_1286);
and U518 (N_518,In_1905,In_734);
or U519 (N_519,In_1068,In_123);
nor U520 (N_520,In_1939,In_1221);
or U521 (N_521,In_442,In_1702);
or U522 (N_522,In_1019,In_422);
xnor U523 (N_523,In_1810,In_565);
or U524 (N_524,In_58,In_1257);
nor U525 (N_525,In_796,In_151);
nor U526 (N_526,In_1999,In_720);
nand U527 (N_527,In_903,In_1459);
and U528 (N_528,N_30,N_150);
nand U529 (N_529,In_919,N_173);
nand U530 (N_530,In_1056,In_1195);
nand U531 (N_531,In_1205,In_310);
and U532 (N_532,In_1722,N_99);
or U533 (N_533,N_190,In_606);
nor U534 (N_534,In_1790,In_1717);
and U535 (N_535,N_342,In_1305);
nand U536 (N_536,N_340,In_1364);
or U537 (N_537,In_85,In_156);
nand U538 (N_538,In_1427,In_995);
and U539 (N_539,In_766,In_469);
and U540 (N_540,N_78,N_12);
and U541 (N_541,In_964,In_942);
nor U542 (N_542,In_1897,In_195);
nand U543 (N_543,In_1776,In_51);
nand U544 (N_544,In_1602,In_643);
xnor U545 (N_545,In_1866,N_32);
and U546 (N_546,In_1998,N_193);
or U547 (N_547,In_686,In_778);
xnor U548 (N_548,N_389,In_287);
or U549 (N_549,In_1508,In_869);
nor U550 (N_550,N_36,In_154);
or U551 (N_551,N_139,In_1198);
nor U552 (N_552,In_1975,In_1132);
nor U553 (N_553,In_1766,N_104);
nor U554 (N_554,In_1010,In_400);
and U555 (N_555,In_1168,N_189);
and U556 (N_556,N_128,In_1453);
nor U557 (N_557,In_924,In_1825);
nor U558 (N_558,In_1976,In_1599);
xor U559 (N_559,In_120,In_1294);
nand U560 (N_560,In_1352,In_294);
or U561 (N_561,In_1307,In_382);
xor U562 (N_562,N_15,In_113);
and U563 (N_563,N_98,In_1950);
xor U564 (N_564,N_67,N_214);
or U565 (N_565,In_357,In_493);
nand U566 (N_566,In_1429,In_88);
xor U567 (N_567,In_782,N_286);
xnor U568 (N_568,In_893,In_1619);
xor U569 (N_569,In_1223,N_377);
or U570 (N_570,N_392,N_187);
and U571 (N_571,N_242,N_171);
or U572 (N_572,In_1428,In_182);
or U573 (N_573,In_1244,In_971);
nor U574 (N_574,N_352,In_1157);
nor U575 (N_575,N_387,In_1562);
and U576 (N_576,In_384,In_476);
nor U577 (N_577,In_1755,In_1536);
nor U578 (N_578,In_1090,In_636);
nand U579 (N_579,In_1115,N_196);
nor U580 (N_580,In_7,In_1491);
and U581 (N_581,In_1636,N_238);
and U582 (N_582,N_367,In_127);
xor U583 (N_583,In_424,In_755);
or U584 (N_584,In_1799,In_249);
or U585 (N_585,In_547,In_160);
or U586 (N_586,In_410,In_1063);
or U587 (N_587,In_371,N_23);
and U588 (N_588,In_861,In_544);
or U589 (N_589,In_966,In_1865);
nor U590 (N_590,N_294,N_21);
and U591 (N_591,In_486,In_1281);
nand U592 (N_592,In_1719,In_361);
or U593 (N_593,N_331,In_948);
or U594 (N_594,N_48,In_1625);
nand U595 (N_595,N_116,In_1433);
and U596 (N_596,N_290,In_1081);
xor U597 (N_597,In_124,N_393);
or U598 (N_598,In_1798,In_1732);
or U599 (N_599,N_96,In_1001);
xnor U600 (N_600,In_169,In_1518);
and U601 (N_601,In_1571,In_936);
xor U602 (N_602,N_253,In_1227);
nand U603 (N_603,N_225,N_65);
or U604 (N_604,In_793,In_1317);
and U605 (N_605,In_1887,N_335);
or U606 (N_606,N_93,N_135);
xor U607 (N_607,In_1273,In_454);
or U608 (N_608,In_899,In_379);
nand U609 (N_609,N_369,In_1037);
nand U610 (N_610,In_1181,N_264);
or U611 (N_611,In_840,In_283);
nor U612 (N_612,In_1271,In_178);
nand U613 (N_613,In_707,N_194);
and U614 (N_614,In_1079,In_770);
xor U615 (N_615,In_1633,N_111);
xnor U616 (N_616,In_1042,In_22);
nand U617 (N_617,In_1666,In_1054);
or U618 (N_618,In_524,In_1658);
nand U619 (N_619,In_539,N_106);
nor U620 (N_620,In_103,In_620);
or U621 (N_621,In_203,In_1895);
or U622 (N_622,N_380,In_829);
xor U623 (N_623,N_118,In_1617);
nor U624 (N_624,In_654,In_811);
nor U625 (N_625,In_1445,In_1290);
nor U626 (N_626,N_344,In_1734);
xor U627 (N_627,N_273,N_291);
nand U628 (N_628,N_170,In_1700);
and U629 (N_629,In_430,In_922);
nand U630 (N_630,In_1140,In_887);
and U631 (N_631,In_292,In_810);
nor U632 (N_632,In_1741,In_1823);
xor U633 (N_633,N_57,In_1270);
nor U634 (N_634,N_63,In_14);
xor U635 (N_635,In_29,In_1543);
and U636 (N_636,In_1744,N_227);
nor U637 (N_637,In_1656,N_166);
and U638 (N_638,In_480,N_308);
xnor U639 (N_639,In_904,In_378);
or U640 (N_640,N_18,In_1568);
or U641 (N_641,N_304,In_1372);
or U642 (N_642,In_1539,In_937);
nor U643 (N_643,In_117,N_217);
nor U644 (N_644,In_399,N_87);
or U645 (N_645,In_406,In_1363);
or U646 (N_646,In_165,In_1028);
nor U647 (N_647,In_787,In_1517);
nor U648 (N_648,In_528,In_1358);
nand U649 (N_649,In_344,In_1452);
and U650 (N_650,In_1806,In_828);
xnor U651 (N_651,N_258,N_114);
or U652 (N_652,In_1933,In_325);
nand U653 (N_653,In_1653,N_240);
and U654 (N_654,In_1206,N_49);
nor U655 (N_655,N_14,N_164);
and U656 (N_656,In_1569,In_65);
nor U657 (N_657,N_188,In_43);
and U658 (N_658,In_628,In_704);
xor U659 (N_659,In_542,In_297);
xnor U660 (N_660,In_1129,In_1879);
nand U661 (N_661,In_494,In_562);
nand U662 (N_662,N_366,N_364);
and U663 (N_663,In_1773,N_6);
xnor U664 (N_664,In_1381,In_1298);
nor U665 (N_665,In_1529,N_399);
nand U666 (N_666,In_1585,In_582);
nand U667 (N_667,In_462,N_218);
and U668 (N_668,In_1615,In_233);
nand U669 (N_669,In_109,In_914);
and U670 (N_670,N_73,In_1347);
nor U671 (N_671,In_773,N_350);
and U672 (N_672,In_1331,In_232);
nand U673 (N_673,N_88,In_1855);
nor U674 (N_674,N_143,In_1760);
nand U675 (N_675,In_111,N_84);
nand U676 (N_676,In_866,In_969);
or U677 (N_677,In_1667,In_1324);
nand U678 (N_678,In_1564,In_1464);
nand U679 (N_679,In_1334,In_981);
nor U680 (N_680,In_1768,In_1035);
nand U681 (N_681,In_1424,N_330);
and U682 (N_682,In_1515,In_1071);
nand U683 (N_683,In_285,In_550);
nor U684 (N_684,N_153,In_1965);
nor U685 (N_685,In_1470,N_53);
or U686 (N_686,In_1225,In_731);
nand U687 (N_687,In_1304,N_277);
xnor U688 (N_688,In_1631,In_803);
or U689 (N_689,In_245,In_1970);
nor U690 (N_690,In_1109,N_339);
and U691 (N_691,In_1052,In_954);
xor U692 (N_692,In_1083,N_372);
nor U693 (N_693,N_59,N_371);
xor U694 (N_694,In_1455,In_105);
nor U695 (N_695,In_1238,In_1479);
xor U696 (N_696,In_967,In_1611);
xnor U697 (N_697,In_536,N_68);
xor U698 (N_698,In_1163,In_878);
and U699 (N_699,In_1301,In_191);
and U700 (N_700,In_225,In_1148);
or U701 (N_701,N_191,N_270);
and U702 (N_702,In_1365,In_1957);
and U703 (N_703,In_1925,In_1065);
nor U704 (N_704,N_94,N_251);
nand U705 (N_705,In_996,N_346);
xnor U706 (N_706,In_1900,In_1584);
or U707 (N_707,In_824,In_751);
and U708 (N_708,In_1967,In_759);
nor U709 (N_709,In_1681,In_207);
or U710 (N_710,In_779,N_74);
nand U711 (N_711,In_452,In_1738);
and U712 (N_712,N_206,In_518);
nor U713 (N_713,In_947,N_215);
and U714 (N_714,In_477,N_345);
nor U715 (N_715,N_309,In_1187);
nand U716 (N_716,In_644,In_1011);
and U717 (N_717,In_374,N_382);
nor U718 (N_718,In_387,In_1789);
and U719 (N_719,In_342,In_1736);
nor U720 (N_720,In_82,N_243);
nand U721 (N_721,In_1960,N_305);
or U722 (N_722,In_1984,N_77);
xnor U723 (N_723,N_396,In_1260);
nor U724 (N_724,N_31,N_376);
and U725 (N_725,In_470,In_1367);
or U726 (N_726,In_402,N_70);
nor U727 (N_727,In_999,In_669);
and U728 (N_728,In_40,In_1366);
and U729 (N_729,In_1844,In_666);
nand U730 (N_730,In_1995,In_395);
xnor U731 (N_731,N_259,In_148);
or U732 (N_732,In_1321,In_1250);
nand U733 (N_733,In_305,N_37);
xnor U734 (N_734,In_1645,In_595);
or U735 (N_735,N_58,N_2);
nor U736 (N_736,N_257,In_281);
and U737 (N_737,In_1740,In_566);
nand U738 (N_738,In_1542,N_374);
or U739 (N_739,In_1442,N_101);
or U740 (N_740,In_448,In_714);
nor U741 (N_741,In_1629,N_239);
and U742 (N_742,In_170,In_679);
xor U743 (N_743,In_745,In_465);
or U744 (N_744,In_1852,N_254);
nor U745 (N_745,In_446,N_307);
or U746 (N_746,In_814,In_9);
or U747 (N_747,In_1694,In_235);
nor U748 (N_748,In_1475,In_18);
xnor U749 (N_749,N_255,In_320);
xor U750 (N_750,In_140,In_346);
nand U751 (N_751,In_1397,In_1382);
and U752 (N_752,In_62,In_626);
and U753 (N_753,In_1117,N_39);
xor U754 (N_754,In_1907,N_315);
or U755 (N_755,In_1614,In_1059);
or U756 (N_756,In_1264,In_1778);
nor U757 (N_757,N_85,In_1018);
xnor U758 (N_758,N_25,In_427);
nor U759 (N_759,In_603,In_1471);
nand U760 (N_760,In_1591,In_1522);
or U761 (N_761,In_852,In_394);
and U762 (N_762,In_428,N_263);
nand U763 (N_763,In_1122,In_425);
nor U764 (N_764,N_40,In_376);
or U765 (N_765,In_352,In_414);
xnor U766 (N_766,In_1510,In_1196);
nor U767 (N_767,N_55,In_1406);
and U768 (N_768,In_55,In_746);
nand U769 (N_769,In_218,N_24);
and U770 (N_770,In_1788,In_482);
xnor U771 (N_771,In_1826,In_267);
nand U772 (N_772,N_75,N_265);
nand U773 (N_773,In_587,In_917);
nand U774 (N_774,N_299,In_458);
xor U775 (N_775,In_1024,In_1254);
nor U776 (N_776,In_1483,In_635);
or U777 (N_777,In_551,In_574);
nand U778 (N_778,In_186,In_331);
nand U779 (N_779,In_1460,N_92);
nor U780 (N_780,In_200,In_1015);
xor U781 (N_781,In_32,In_250);
nor U782 (N_782,In_38,N_160);
and U783 (N_783,N_272,In_1246);
nor U784 (N_784,In_940,In_1369);
nor U785 (N_785,In_1341,N_115);
nor U786 (N_786,In_451,N_151);
and U787 (N_787,N_313,In_131);
and U788 (N_788,In_1676,In_1354);
and U789 (N_789,In_1566,In_741);
or U790 (N_790,N_147,In_153);
xor U791 (N_791,In_802,N_250);
or U792 (N_792,N_51,In_1162);
or U793 (N_793,In_91,N_56);
or U794 (N_794,N_336,N_184);
nor U795 (N_795,In_1045,In_601);
xnor U796 (N_796,In_1877,In_239);
xnor U797 (N_797,N_245,N_327);
nor U798 (N_798,N_1,In_754);
xnor U799 (N_799,N_298,In_1447);
nor U800 (N_800,N_622,N_477);
xor U801 (N_801,In_867,N_692);
xor U802 (N_802,N_443,N_739);
and U803 (N_803,N_656,In_54);
nor U804 (N_804,N_541,N_148);
xnor U805 (N_805,In_1017,N_576);
nand U806 (N_806,In_854,In_944);
nor U807 (N_807,In_1673,N_724);
and U808 (N_808,In_508,In_794);
nor U809 (N_809,N_598,N_459);
or U810 (N_810,N_600,In_35);
nand U811 (N_811,N_221,N_784);
nand U812 (N_812,In_1112,In_980);
nand U813 (N_813,In_1454,In_1486);
and U814 (N_814,N_267,N_130);
xnor U815 (N_815,In_683,N_16);
and U816 (N_816,In_84,N_696);
xor U817 (N_817,N_659,N_761);
nand U818 (N_818,N_121,N_492);
nor U819 (N_819,In_1701,In_102);
nand U820 (N_820,In_902,In_171);
nand U821 (N_821,In_1918,N_311);
and U822 (N_822,In_1839,N_535);
and U823 (N_823,N_416,N_198);
nand U824 (N_824,In_517,In_1942);
xor U825 (N_825,N_677,N_131);
and U826 (N_826,N_685,In_630);
xor U827 (N_827,N_404,In_291);
or U828 (N_828,In_1882,In_1930);
nand U829 (N_829,N_543,In_664);
nand U830 (N_830,N_203,In_1077);
nor U831 (N_831,In_1519,In_1116);
or U832 (N_832,In_1359,In_121);
nor U833 (N_833,In_97,N_714);
and U834 (N_834,N_479,N_787);
xnor U835 (N_835,In_49,N_793);
or U836 (N_836,In_1990,N_413);
nand U837 (N_837,In_1514,In_1156);
or U838 (N_838,In_142,In_1383);
nand U839 (N_839,N_633,In_784);
or U840 (N_840,N_288,In_1210);
nor U841 (N_841,In_965,N_347);
nor U842 (N_842,In_676,In_1746);
nand U843 (N_843,In_72,N_510);
or U844 (N_844,In_1892,In_443);
or U845 (N_845,N_213,In_364);
xor U846 (N_846,In_450,In_1838);
and U847 (N_847,N_408,In_1808);
or U848 (N_848,N_743,N_442);
and U849 (N_849,In_1335,In_1222);
and U850 (N_850,N_581,N_792);
xnor U851 (N_851,In_298,N_552);
and U852 (N_852,In_573,In_1966);
xnor U853 (N_853,N_708,N_691);
or U854 (N_854,N_783,In_289);
xnor U855 (N_855,In_1888,In_1699);
xnor U856 (N_856,In_1595,In_563);
nand U857 (N_857,N_681,N_363);
and U858 (N_858,In_726,N_236);
nand U859 (N_859,N_796,In_972);
or U860 (N_860,N_329,In_268);
xnor U861 (N_861,N_631,N_199);
and U862 (N_862,In_617,N_729);
or U863 (N_863,In_1962,N_202);
xnor U864 (N_864,In_1275,In_439);
nor U865 (N_865,N_657,N_611);
nor U866 (N_866,In_498,In_210);
xor U867 (N_867,N_458,N_706);
nand U868 (N_868,N_310,N_292);
nor U869 (N_869,N_476,N_684);
or U870 (N_870,N_223,N_425);
and U871 (N_871,In_1894,In_95);
and U872 (N_872,In_229,In_1482);
or U873 (N_873,N_583,In_874);
or U874 (N_874,In_777,N_481);
xor U875 (N_875,N_537,In_1623);
or U876 (N_876,N_324,N_612);
nor U877 (N_877,In_616,In_1458);
xor U878 (N_878,In_681,N_421);
nand U879 (N_879,N_178,N_637);
and U880 (N_880,N_603,N_627);
nor U881 (N_881,In_1226,N_497);
xnor U882 (N_882,In_1881,N_428);
or U883 (N_883,In_1207,In_921);
and U884 (N_884,In_939,N_47);
or U885 (N_885,In_1858,N_8);
or U886 (N_886,N_544,N_658);
or U887 (N_887,N_332,In_360);
xor U888 (N_888,N_664,N_244);
nor U889 (N_889,In_1378,N_763);
xor U890 (N_890,N_670,In_1346);
or U891 (N_891,N_186,In_890);
nand U892 (N_892,In_1199,In_13);
and U893 (N_893,N_27,In_588);
nand U894 (N_894,In_1280,N_798);
nand U895 (N_895,In_1076,In_752);
or U896 (N_896,In_322,N_361);
xor U897 (N_897,In_1033,N_142);
nor U898 (N_898,In_77,N_516);
nand U899 (N_899,In_1709,N_486);
nor U900 (N_900,In_684,In_1683);
xnor U901 (N_901,In_1989,N_450);
or U902 (N_902,In_365,N_701);
nand U903 (N_903,N_224,N_750);
or U904 (N_904,N_453,N_41);
and U905 (N_905,N_704,In_392);
xnor U906 (N_906,In_216,N_76);
and U907 (N_907,In_436,In_931);
xor U908 (N_908,N_233,In_1550);
xor U909 (N_909,In_1716,In_277);
nor U910 (N_910,In_1182,In_1292);
nand U911 (N_911,N_539,N_781);
xor U912 (N_912,N_429,N_468);
and U913 (N_913,In_370,In_354);
nand U914 (N_914,N_565,In_1952);
xnor U915 (N_915,In_769,In_934);
xor U916 (N_916,In_1596,N_149);
and U917 (N_917,In_413,N_652);
or U918 (N_918,N_69,N_275);
and U919 (N_919,In_1947,In_1202);
nor U920 (N_920,In_1770,N_568);
nor U921 (N_921,In_3,In_1909);
xnor U922 (N_922,N_419,In_134);
and U923 (N_923,In_201,N_727);
nor U924 (N_924,N_745,In_1300);
nor U925 (N_925,In_1247,In_468);
xor U926 (N_926,In_1842,In_605);
xor U927 (N_927,N_636,In_505);
and U928 (N_928,In_584,N_513);
nand U929 (N_929,In_405,N_445);
and U930 (N_930,N_158,In_335);
nand U931 (N_931,N_618,N_318);
or U932 (N_932,N_653,N_0);
or U933 (N_933,N_351,In_1274);
and U934 (N_934,In_1523,N_140);
or U935 (N_935,N_83,N_731);
or U936 (N_936,In_6,N_680);
nand U937 (N_937,N_22,In_177);
and U938 (N_938,N_493,In_1188);
or U939 (N_939,N_337,In_1224);
and U940 (N_940,In_1724,N_591);
nand U941 (N_941,N_9,In_868);
nor U942 (N_942,In_1299,In_1291);
nor U943 (N_943,In_788,In_662);
nor U944 (N_944,In_1123,N_674);
nand U945 (N_945,N_648,N_452);
xor U946 (N_946,N_512,N_378);
nand U947 (N_947,N_296,In_76);
nor U948 (N_948,In_284,N_707);
nor U949 (N_949,In_355,In_543);
xor U950 (N_950,In_1099,N_280);
xor U951 (N_951,In_982,In_1160);
xnor U952 (N_952,In_1136,In_24);
xor U953 (N_953,N_672,In_1443);
nor U954 (N_954,In_57,N_7);
nand U955 (N_955,In_1889,In_1110);
nand U956 (N_956,N_105,N_110);
xor U957 (N_957,N_526,N_89);
nor U958 (N_958,N_60,N_201);
nor U959 (N_959,In_577,N_791);
or U960 (N_960,In_393,N_735);
and U961 (N_961,In_1440,N_303);
nor U962 (N_962,N_588,In_1843);
or U963 (N_963,N_222,In_1899);
or U964 (N_964,In_278,N_575);
or U965 (N_965,In_1026,N_123);
nand U966 (N_966,In_842,N_782);
xor U967 (N_967,N_144,In_1336);
or U968 (N_968,N_538,N_770);
nand U969 (N_969,N_386,N_640);
and U970 (N_970,N_52,N_406);
nor U971 (N_971,In_1245,In_118);
or U972 (N_972,In_1920,In_597);
or U973 (N_973,In_1624,In_975);
or U974 (N_974,In_655,In_1485);
nand U975 (N_975,N_654,In_1154);
xnor U976 (N_976,In_744,In_1968);
xor U977 (N_977,N_441,In_271);
nor U978 (N_978,N_617,N_523);
or U979 (N_979,In_631,In_1448);
or U980 (N_980,N_200,In_340);
nor U981 (N_981,In_976,In_1082);
and U982 (N_982,In_1655,In_1417);
nand U983 (N_983,In_719,In_132);
or U984 (N_984,In_133,N_328);
or U985 (N_985,N_621,In_1436);
or U986 (N_986,N_323,In_525);
or U987 (N_987,N_597,N_461);
or U988 (N_988,N_638,N_578);
xor U989 (N_989,N_675,In_1685);
nor U990 (N_990,In_1620,N_192);
xnor U991 (N_991,In_149,N_650);
xnor U992 (N_992,In_59,In_1049);
nand U993 (N_993,In_933,In_1557);
or U994 (N_994,N_730,In_709);
nand U995 (N_995,N_534,In_839);
or U996 (N_996,In_561,In_1183);
nand U997 (N_997,In_657,In_1910);
xor U998 (N_998,N_678,In_690);
or U999 (N_999,N_62,In_988);
and U1000 (N_1000,N_287,In_1898);
or U1001 (N_1001,In_1525,In_728);
nor U1002 (N_1002,N_137,N_616);
nand U1003 (N_1003,N_712,In_1607);
and U1004 (N_1004,In_1731,N_506);
xnor U1005 (N_1005,N_306,N_709);
or U1006 (N_1006,In_1630,In_25);
nand U1007 (N_1007,In_1775,N_697);
or U1008 (N_1008,N_370,In_4);
xor U1009 (N_1009,In_670,N_574);
nor U1010 (N_1010,In_589,In_1767);
nand U1011 (N_1011,In_1903,In_296);
or U1012 (N_1012,In_1025,In_791);
xor U1013 (N_1013,In_1670,N_495);
and U1014 (N_1014,N_517,N_436);
and U1015 (N_1015,In_955,N_216);
xnor U1016 (N_1016,N_749,In_795);
nor U1017 (N_1017,N_531,N_717);
nand U1018 (N_1018,N_649,N_356);
and U1019 (N_1019,N_779,In_1108);
or U1020 (N_1020,N_590,In_1582);
nand U1021 (N_1021,In_467,In_1220);
nor U1022 (N_1022,In_1972,In_1735);
and U1023 (N_1023,N_390,N_580);
nor U1024 (N_1024,N_566,In_219);
or U1025 (N_1025,N_768,N_533);
nand U1026 (N_1026,N_82,In_1650);
nor U1027 (N_1027,N_619,N_775);
or U1028 (N_1028,In_675,N_325);
xor U1029 (N_1029,N_235,N_728);
nor U1030 (N_1030,In_150,N_427);
or U1031 (N_1031,In_1502,In_925);
nand U1032 (N_1032,N_769,In_864);
and U1033 (N_1033,N_499,In_1230);
nor U1034 (N_1034,N_584,In_1344);
nand U1035 (N_1035,In_1237,N_639);
and U1036 (N_1036,N_197,N_645);
nor U1037 (N_1037,In_1688,In_1641);
nand U1038 (N_1038,N_5,N_579);
or U1039 (N_1039,N_54,In_1590);
xor U1040 (N_1040,In_46,N_610);
and U1041 (N_1041,In_677,In_1288);
and U1042 (N_1042,N_208,N_693);
xnor U1043 (N_1043,N_705,N_134);
nand U1044 (N_1044,In_1814,N_773);
xnor U1045 (N_1045,In_907,N_607);
xor U1046 (N_1046,N_751,N_756);
nor U1047 (N_1047,N_647,N_10);
xnor U1048 (N_1048,N_577,N_460);
nand U1049 (N_1049,N_722,In_849);
nor U1050 (N_1050,In_261,N_758);
or U1051 (N_1051,N_322,N_587);
or U1052 (N_1052,N_759,N_230);
and U1053 (N_1053,In_204,In_1874);
nand U1054 (N_1054,In_1481,N_753);
and U1055 (N_1055,N_589,N_373);
and U1056 (N_1056,In_193,In_555);
nand U1057 (N_1057,N_467,In_1807);
nor U1058 (N_1058,In_481,N_417);
or U1059 (N_1059,N_766,In_1073);
nor U1060 (N_1060,N_508,In_1588);
nand U1061 (N_1061,N_551,In_315);
nand U1062 (N_1062,In_533,N_569);
nand U1063 (N_1063,In_1917,N_503);
nand U1064 (N_1064,N_505,In_625);
and U1065 (N_1065,In_1954,N_549);
nand U1066 (N_1066,In_1792,N_570);
or U1067 (N_1067,N_521,N_439);
or U1068 (N_1068,N_246,In_60);
nor U1069 (N_1069,In_1574,In_1982);
and U1070 (N_1070,N_472,N_757);
or U1071 (N_1071,In_703,In_1144);
nor U1072 (N_1072,N_679,In_363);
xnor U1073 (N_1073,In_1509,In_821);
nand U1074 (N_1074,N_13,In_507);
nand U1075 (N_1075,In_1689,In_1311);
nor U1076 (N_1076,In_1474,In_1703);
nor U1077 (N_1077,In_725,In_415);
nand U1078 (N_1078,N_117,N_293);
nor U1079 (N_1079,In_1774,N_29);
nand U1080 (N_1080,N_624,N_614);
and U1081 (N_1081,In_1937,In_1687);
nand U1082 (N_1082,N_655,In_1757);
nand U1083 (N_1083,N_487,In_1849);
nand U1084 (N_1084,N_231,In_1277);
or U1085 (N_1085,In_691,In_807);
or U1086 (N_1086,In_1743,N_358);
and U1087 (N_1087,In_685,N_407);
or U1088 (N_1088,N_490,In_1504);
or U1089 (N_1089,In_809,N_261);
and U1090 (N_1090,In_1034,N_564);
nand U1091 (N_1091,N_405,N_737);
and U1092 (N_1092,N_426,In_1690);
nor U1093 (N_1093,N_456,In_435);
nor U1094 (N_1094,N_511,In_1929);
nor U1095 (N_1095,N_145,In_1215);
xnor U1096 (N_1096,N_585,In_475);
nor U1097 (N_1097,In_1558,In_889);
or U1098 (N_1098,N_715,N_45);
and U1099 (N_1099,In_234,N_713);
nand U1100 (N_1100,N_409,N_435);
or U1101 (N_1101,In_1572,In_143);
or U1102 (N_1102,In_464,In_441);
xor U1103 (N_1103,N_312,In_957);
nand U1104 (N_1104,N_651,N_341);
nor U1105 (N_1105,In_1583,N_524);
or U1106 (N_1106,N_156,In_492);
nand U1107 (N_1107,In_1137,In_1659);
xor U1108 (N_1108,N_249,N_454);
and U1109 (N_1109,N_752,In_419);
or U1110 (N_1110,N_494,In_484);
or U1111 (N_1111,In_1953,N_542);
and U1112 (N_1112,In_256,In_300);
nand U1113 (N_1113,N_437,In_167);
nor U1114 (N_1114,In_367,In_1430);
nand U1115 (N_1115,N_220,N_343);
and U1116 (N_1116,N_212,N_771);
and U1117 (N_1117,N_491,N_470);
nor U1118 (N_1118,N_397,In_1586);
and U1119 (N_1119,In_114,N_469);
and U1120 (N_1120,In_820,In_1327);
and U1121 (N_1121,N_289,In_94);
and U1122 (N_1122,In_1233,In_303);
xnor U1123 (N_1123,In_474,In_1643);
nand U1124 (N_1124,In_1374,In_768);
nor U1125 (N_1125,N_668,In_790);
xor U1126 (N_1126,N_626,In_1795);
nor U1127 (N_1127,N_496,N_433);
nor U1128 (N_1128,N_179,N_686);
nand U1129 (N_1129,In_304,In_832);
and U1130 (N_1130,N_646,N_643);
and U1131 (N_1131,In_1496,N_726);
or U1132 (N_1132,N_732,N_412);
nand U1133 (N_1133,In_377,In_680);
nand U1134 (N_1134,In_1021,N_394);
and U1135 (N_1135,In_608,In_983);
or U1136 (N_1136,N_557,N_776);
nand U1137 (N_1137,In_135,N_165);
or U1138 (N_1138,In_583,In_825);
nor U1139 (N_1139,N_605,N_234);
nor U1140 (N_1140,N_662,N_447);
or U1141 (N_1141,N_211,In_712);
nand U1142 (N_1142,In_1563,N_466);
nor U1143 (N_1143,In_1680,In_1409);
nor U1144 (N_1144,In_1235,In_214);
or U1145 (N_1145,In_1637,In_780);
nor U1146 (N_1146,In_1173,N_642);
nand U1147 (N_1147,In_1628,In_1935);
xor U1148 (N_1148,N_620,N_698);
nor U1149 (N_1149,In_1411,In_90);
nor U1150 (N_1150,In_390,N_665);
xnor U1151 (N_1151,N_300,N_682);
xnor U1152 (N_1152,In_1809,In_771);
and U1153 (N_1153,In_516,N_725);
and U1154 (N_1154,In_126,In_865);
xnor U1155 (N_1155,In_835,N_113);
xnor U1156 (N_1156,N_473,N_424);
nand U1157 (N_1157,In_1086,N_594);
or U1158 (N_1158,In_87,N_716);
xor U1159 (N_1159,N_582,N_348);
or U1160 (N_1160,In_1029,In_1050);
or U1161 (N_1161,In_1009,In_1377);
nand U1162 (N_1162,In_1762,In_1576);
nor U1163 (N_1163,N_785,In_2);
nand U1164 (N_1164,In_1423,In_1758);
xnor U1165 (N_1165,N_748,N_444);
xnor U1166 (N_1166,N_777,N_689);
xor U1167 (N_1167,N_786,N_43);
xnor U1168 (N_1168,In_1864,In_380);
xnor U1169 (N_1169,In_432,N_451);
xor U1170 (N_1170,In_610,In_1593);
or U1171 (N_1171,In_1392,N_634);
xor U1172 (N_1172,N_635,N_284);
or U1173 (N_1173,In_1946,In_212);
or U1174 (N_1174,In_106,N_448);
or U1175 (N_1175,In_970,N_632);
and U1176 (N_1176,N_241,In_1236);
nor U1177 (N_1177,In_385,In_1661);
xnor U1178 (N_1178,In_372,N_790);
and U1179 (N_1179,In_1126,N_283);
or U1180 (N_1180,N_738,N_667);
nand U1181 (N_1181,In_438,N_507);
nor U1182 (N_1182,N_794,In_812);
and U1183 (N_1183,In_621,N_797);
xor U1184 (N_1184,N_604,In_797);
or U1185 (N_1185,In_1303,N_268);
and U1186 (N_1186,N_630,In_1512);
nand U1187 (N_1187,N_586,N_247);
nand U1188 (N_1188,In_733,N_518);
and U1189 (N_1189,In_1981,N_95);
nor U1190 (N_1190,In_1124,N_548);
nor U1191 (N_1191,In_1840,N_561);
xor U1192 (N_1192,In_905,N_596);
and U1193 (N_1193,N_663,In_699);
nand U1194 (N_1194,In_1538,In_1873);
or U1195 (N_1195,In_1706,In_804);
nor U1196 (N_1196,N_379,N_778);
nor U1197 (N_1197,N_295,N_320);
or U1198 (N_1198,N_61,In_75);
nand U1199 (N_1199,In_1120,In_1371);
and U1200 (N_1200,N_660,N_866);
or U1201 (N_1201,N_1168,In_1269);
nor U1202 (N_1202,N_501,N_936);
nand U1203 (N_1203,N_859,In_1664);
or U1204 (N_1204,N_316,N_550);
and U1205 (N_1205,In_860,N_1188);
or U1206 (N_1206,N_1086,In_1097);
xnor U1207 (N_1207,N_868,N_1043);
nand U1208 (N_1208,N_504,In_765);
and U1209 (N_1209,N_1184,N_1023);
and U1210 (N_1210,N_1112,In_101);
nor U1211 (N_1211,N_834,N_1132);
or U1212 (N_1212,N_520,N_671);
xnor U1213 (N_1213,N_683,N_478);
and U1214 (N_1214,N_1169,N_1196);
and U1215 (N_1215,N_810,N_961);
nand U1216 (N_1216,N_1040,N_1030);
or U1217 (N_1217,In_1234,In_253);
xor U1218 (N_1218,In_274,N_560);
xor U1219 (N_1219,N_109,N_423);
and U1220 (N_1220,N_885,In_730);
and U1221 (N_1221,N_848,N_317);
nor U1222 (N_1222,N_1031,In_618);
and U1223 (N_1223,N_865,In_532);
xor U1224 (N_1224,In_1640,N_801);
and U1225 (N_1225,N_554,N_609);
nor U1226 (N_1226,N_530,N_1095);
nand U1227 (N_1227,In_1326,N_874);
or U1228 (N_1228,In_1361,N_1101);
xnor U1229 (N_1229,N_933,N_1079);
xnor U1230 (N_1230,In_1831,In_817);
nor U1231 (N_1231,N_157,N_1021);
nor U1232 (N_1232,N_529,In_537);
and U1233 (N_1233,N_1042,N_1115);
and U1234 (N_1234,N_120,N_338);
xor U1235 (N_1235,In_173,N_1087);
nand U1236 (N_1236,N_1078,N_1110);
and U1237 (N_1237,In_1802,N_856);
xor U1238 (N_1238,N_319,N_838);
nor U1239 (N_1239,In_1921,N_895);
or U1240 (N_1240,In_831,In_1219);
or U1241 (N_1241,N_365,In_1310);
and U1242 (N_1242,N_953,In_1608);
nand U1243 (N_1243,N_1048,N_772);
and U1244 (N_1244,N_195,N_1126);
nand U1245 (N_1245,In_17,N_498);
nor U1246 (N_1246,N_977,In_912);
nand U1247 (N_1247,N_1038,N_924);
and U1248 (N_1248,N_480,N_1069);
or U1249 (N_1249,N_918,N_887);
and U1250 (N_1250,In_1000,N_297);
and U1251 (N_1251,N_1085,N_1116);
nand U1252 (N_1252,N_734,N_573);
nor U1253 (N_1253,N_799,N_185);
nor U1254 (N_1254,N_1187,N_1122);
nand U1255 (N_1255,N_741,N_440);
and U1256 (N_1256,N_1176,N_964);
or U1257 (N_1257,N_913,N_980);
and U1258 (N_1258,N_525,N_976);
nand U1259 (N_1259,N_1104,N_965);
and U1260 (N_1260,N_1035,N_1134);
or U1261 (N_1261,N_998,N_981);
nor U1262 (N_1262,N_851,In_337);
nor U1263 (N_1263,N_1174,In_89);
nand U1264 (N_1264,N_906,N_1044);
nand U1265 (N_1265,In_125,N_608);
xnor U1266 (N_1266,N_710,N_828);
xor U1267 (N_1267,N_1056,In_833);
and U1268 (N_1268,N_1139,N_962);
or U1269 (N_1269,N_746,In_1435);
nor U1270 (N_1270,N_1046,N_931);
or U1271 (N_1271,In_732,In_1401);
and U1272 (N_1272,In_1561,N_1049);
nor U1273 (N_1273,N_1103,In_1216);
or U1274 (N_1274,N_821,N_1105);
and U1275 (N_1275,N_886,N_438);
xnor U1276 (N_1276,In_1969,N_1155);
xnor U1277 (N_1277,N_1075,N_383);
nor U1278 (N_1278,N_905,In_637);
nor U1279 (N_1279,N_108,N_997);
nand U1280 (N_1280,N_415,N_960);
nor U1281 (N_1281,N_1183,In_93);
nand U1282 (N_1282,N_125,N_788);
nor U1283 (N_1283,N_1162,In_1211);
nor U1284 (N_1284,N_837,N_1163);
or U1285 (N_1285,In_872,N_28);
and U1286 (N_1286,In_688,N_1076);
and U1287 (N_1287,N_971,N_1009);
nor U1288 (N_1288,In_1883,N_606);
or U1289 (N_1289,N_760,N_867);
and U1290 (N_1290,N_1178,N_921);
nor U1291 (N_1291,N_883,N_850);
xor U1292 (N_1292,N_375,N_465);
and U1293 (N_1293,N_817,N_687);
nand U1294 (N_1294,N_959,N_941);
nand U1295 (N_1295,In_1297,N_1028);
and U1296 (N_1296,N_1008,N_1130);
and U1297 (N_1297,N_1053,N_872);
or U1298 (N_1298,N_978,N_1182);
nor U1299 (N_1299,N_950,N_1144);
nor U1300 (N_1300,N_894,In_713);
or U1301 (N_1301,N_702,N_1088);
xnor U1302 (N_1302,N_402,N_744);
and U1303 (N_1303,N_690,N_845);
nor U1304 (N_1304,N_999,N_1161);
and U1305 (N_1305,N_484,N_1054);
or U1306 (N_1306,N_1034,N_276);
xnor U1307 (N_1307,In_715,N_1055);
nor U1308 (N_1308,N_907,N_11);
xor U1309 (N_1309,N_266,N_1141);
and U1310 (N_1310,In_445,N_988);
and U1311 (N_1311,N_1064,In_192);
or U1312 (N_1312,N_431,In_1646);
xnor U1313 (N_1313,N_81,N_26);
or U1314 (N_1314,In_47,In_248);
and U1315 (N_1315,In_1268,N_860);
nor U1316 (N_1316,N_972,In_1262);
and U1317 (N_1317,N_922,In_275);
nor U1318 (N_1318,N_1007,N_871);
or U1319 (N_1319,N_1003,N_1071);
xor U1320 (N_1320,In_1725,In_1993);
or U1321 (N_1321,N_832,N_1073);
nor U1322 (N_1322,In_1084,N_279);
xnor U1323 (N_1323,N_1091,N_1047);
xnor U1324 (N_1324,N_1145,In_81);
nand U1325 (N_1325,In_639,N_559);
xor U1326 (N_1326,N_930,N_774);
nor U1327 (N_1327,In_1176,N_1192);
nor U1328 (N_1328,In_1325,N_540);
and U1329 (N_1329,N_482,In_1828);
and U1330 (N_1330,N_1061,N_742);
and U1331 (N_1331,N_1131,N_900);
or U1332 (N_1332,N_418,In_658);
and U1333 (N_1333,In_41,N_46);
nand U1334 (N_1334,N_762,N_1070);
xnor U1335 (N_1335,N_483,N_820);
and U1336 (N_1336,N_937,N_1066);
and U1337 (N_1337,N_889,N_736);
or U1338 (N_1338,N_488,N_80);
xor U1339 (N_1339,N_430,N_1157);
or U1340 (N_1340,In_100,N_864);
nor U1341 (N_1341,N_944,In_1487);
xnor U1342 (N_1342,N_446,N_829);
nor U1343 (N_1343,N_1142,N_882);
and U1344 (N_1344,In_927,In_397);
and U1345 (N_1345,In_407,N_355);
xor U1346 (N_1346,N_1050,N_528);
nor U1347 (N_1347,In_909,N_100);
nand U1348 (N_1348,N_695,N_1102);
nand U1349 (N_1349,N_1135,In_1175);
xor U1350 (N_1350,N_1032,N_1026);
and U1351 (N_1351,N_946,In_515);
nor U1352 (N_1352,In_552,N_916);
nor U1353 (N_1353,N_878,N_824);
nor U1354 (N_1354,N_395,N_1140);
and U1355 (N_1355,N_789,N_814);
or U1356 (N_1356,In_649,N_849);
nor U1357 (N_1357,N_136,N_226);
nor U1358 (N_1358,N_464,In_1657);
nor U1359 (N_1359,N_615,N_1033);
nand U1360 (N_1360,N_852,N_1195);
nor U1361 (N_1361,N_982,In_1141);
nor U1362 (N_1362,N_842,N_613);
nor U1363 (N_1363,N_822,N_515);
and U1364 (N_1364,In_1179,N_942);
nand U1365 (N_1365,N_485,N_754);
or U1366 (N_1366,N_901,N_987);
nor U1367 (N_1367,N_914,N_1017);
nor U1368 (N_1368,N_1197,In_1927);
xor U1369 (N_1369,N_1194,N_547);
nand U1370 (N_1370,N_967,N_1100);
or U1371 (N_1371,N_1011,N_826);
nand U1372 (N_1372,N_180,In_1729);
nor U1373 (N_1373,N_992,N_1107);
xor U1374 (N_1374,In_314,In_857);
xor U1375 (N_1375,N_805,N_947);
or U1376 (N_1376,N_841,In_633);
or U1377 (N_1377,N_996,N_733);
and U1378 (N_1378,In_753,N_326);
nand U1379 (N_1379,In_1450,In_251);
and U1380 (N_1380,N_1022,N_475);
xor U1381 (N_1381,N_546,N_926);
and U1382 (N_1382,N_809,N_870);
xnor U1383 (N_1383,N_269,In_1416);
nand U1384 (N_1384,In_130,In_863);
xor U1385 (N_1385,N_401,In_30);
nor U1386 (N_1386,N_1128,N_314);
and U1387 (N_1387,N_302,N_1098);
and U1388 (N_1388,In_194,N_765);
nand U1389 (N_1389,N_1059,N_1153);
xnor U1390 (N_1390,N_857,N_847);
nand U1391 (N_1391,In_1926,In_1662);
nand U1392 (N_1392,N_1015,N_811);
or U1393 (N_1393,N_897,In_906);
and U1394 (N_1394,N_920,N_463);
and U1395 (N_1395,In_1259,N_1151);
and U1396 (N_1396,N_862,N_1175);
nor U1397 (N_1397,N_278,N_1012);
nor U1398 (N_1398,N_545,N_949);
nand U1399 (N_1399,N_966,N_703);
and U1400 (N_1400,N_623,N_985);
and U1401 (N_1401,N_1037,N_892);
or U1402 (N_1402,N_911,N_1179);
and U1403 (N_1403,N_1001,N_904);
nand U1404 (N_1404,N_209,N_602);
and U1405 (N_1405,N_673,N_1080);
or U1406 (N_1406,In_801,N_1096);
xor U1407 (N_1407,N_1036,N_1094);
nor U1408 (N_1408,N_1189,In_1526);
or U1409 (N_1409,N_935,N_1005);
nand U1410 (N_1410,In_362,N_909);
xor U1411 (N_1411,N_1010,In_348);
nor U1412 (N_1412,In_64,In_1101);
xor U1413 (N_1413,N_79,N_1120);
xor U1414 (N_1414,N_1186,In_1142);
nor U1415 (N_1415,In_743,N_1159);
and U1416 (N_1416,N_274,N_1006);
and U1417 (N_1417,N_893,In_1119);
and U1418 (N_1418,N_127,N_803);
or U1419 (N_1419,In_950,N_1117);
xor U1420 (N_1420,In_175,N_1138);
or U1421 (N_1421,In_262,N_532);
and U1422 (N_1422,N_384,In_359);
xor U1423 (N_1423,N_1173,N_555);
xor U1424 (N_1424,N_875,N_815);
or U1425 (N_1425,In_366,N_228);
and U1426 (N_1426,N_915,N_843);
xor U1427 (N_1427,N_995,N_71);
nor U1428 (N_1428,N_357,In_1827);
and U1429 (N_1429,In_396,N_880);
or U1430 (N_1430,N_669,N_928);
and U1431 (N_1431,N_823,N_1004);
nor U1432 (N_1432,N_400,N_489);
and U1433 (N_1433,N_927,N_553);
or U1434 (N_1434,N_1039,N_174);
or U1435 (N_1435,In_1113,N_877);
and U1436 (N_1436,N_767,In_1267);
or U1437 (N_1437,In_1693,In_1438);
and U1438 (N_1438,N_846,In_1040);
xnor U1439 (N_1439,In_1528,N_301);
or U1440 (N_1440,In_332,N_1150);
and U1441 (N_1441,In_1769,N_840);
nand U1442 (N_1442,N_951,In_489);
and U1443 (N_1443,In_213,N_19);
and U1444 (N_1444,N_994,N_780);
or U1445 (N_1445,In_202,In_998);
xor U1446 (N_1446,N_571,In_570);
and U1447 (N_1447,N_943,N_1172);
or U1448 (N_1448,N_593,N_721);
xor U1449 (N_1449,N_262,N_1027);
nor U1450 (N_1450,N_979,N_807);
nand U1451 (N_1451,N_1180,In_227);
nor U1452 (N_1452,N_1018,In_1285);
xnor U1453 (N_1453,In_185,N_898);
or U1454 (N_1454,N_969,In_433);
or U1455 (N_1455,In_333,In_416);
nor U1456 (N_1456,N_411,N_388);
and U1457 (N_1457,N_333,N_747);
nor U1458 (N_1458,N_1165,N_929);
nor U1459 (N_1459,N_957,N_958);
nand U1460 (N_1460,N_1072,In_240);
nand U1461 (N_1461,N_984,N_34);
and U1462 (N_1462,N_1058,N_502);
xnor U1463 (N_1463,N_934,N_955);
nor U1464 (N_1464,N_896,N_1109);
nor U1465 (N_1465,N_795,N_804);
and U1466 (N_1466,N_831,In_1791);
nor U1467 (N_1467,N_835,N_833);
xnor U1468 (N_1468,N_1129,N_1118);
xnor U1469 (N_1469,In_1622,N_1148);
or U1470 (N_1470,In_1639,N_970);
xnor U1471 (N_1471,N_1124,N_986);
nand U1472 (N_1472,N_1185,In_898);
and U1473 (N_1473,N_558,N_812);
nand U1474 (N_1474,N_563,N_562);
and U1475 (N_1475,N_271,In_20);
xnor U1476 (N_1476,N_152,In_678);
nor U1477 (N_1477,N_975,N_806);
or U1478 (N_1478,In_1692,N_572);
nor U1479 (N_1479,N_514,In_1384);
xor U1480 (N_1480,N_1114,N_945);
xor U1481 (N_1481,In_767,N_509);
xnor U1482 (N_1482,N_1089,In_735);
and U1483 (N_1483,In_1577,N_1166);
or U1484 (N_1484,N_1065,N_932);
and U1485 (N_1485,In_1513,N_595);
or U1486 (N_1486,In_206,N_939);
nor U1487 (N_1487,In_1218,In_1178);
nand U1488 (N_1488,N_1002,N_556);
or U1489 (N_1489,In_1313,N_462);
and U1490 (N_1490,In_549,N_1081);
or U1491 (N_1491,In_1627,N_159);
or U1492 (N_1492,In_859,N_625);
nor U1493 (N_1493,N_205,In_437);
and U1494 (N_1494,N_1019,In_740);
nand U1495 (N_1495,N_1149,N_873);
or U1496 (N_1496,In_660,N_1000);
and U1497 (N_1497,N_963,N_1025);
nand U1498 (N_1498,N_410,N_1090);
xor U1499 (N_1499,N_989,In_252);
nand U1500 (N_1500,In_1217,N_1198);
nor U1501 (N_1501,In_495,N_414);
or U1502 (N_1502,N_923,N_1014);
nand U1503 (N_1503,N_1190,N_1013);
nand U1504 (N_1504,N_876,In_1638);
and U1505 (N_1505,N_1029,N_827);
or U1506 (N_1506,N_808,N_973);
nand U1507 (N_1507,N_1016,N_455);
nand U1508 (N_1508,N_1154,N_1063);
xnor U1509 (N_1509,In_1058,N_1051);
xnor U1510 (N_1510,N_1167,N_816);
and U1511 (N_1511,N_863,N_474);
or U1512 (N_1512,N_764,N_1146);
nor U1513 (N_1513,N_44,N_1106);
xor U1514 (N_1514,N_991,N_432);
nand U1515 (N_1515,N_1067,N_1068);
or U1516 (N_1516,N_1143,In_529);
nor U1517 (N_1517,N_974,N_154);
nor U1518 (N_1518,N_1164,N_844);
nand U1519 (N_1519,N_599,N_519);
xor U1520 (N_1520,N_471,N_1152);
and U1521 (N_1521,N_917,N_33);
and U1522 (N_1522,N_903,N_855);
nor U1523 (N_1523,N_912,N_899);
xnor U1524 (N_1524,N_1199,N_1125);
nand U1525 (N_1525,In_1204,N_661);
or U1526 (N_1526,In_1763,N_522);
or U1527 (N_1527,N_1156,N_536);
xor U1528 (N_1528,N_567,N_641);
or U1529 (N_1529,N_755,N_861);
or U1530 (N_1530,N_910,N_422);
or U1531 (N_1531,In_158,In_1088);
nand U1532 (N_1532,N_925,N_983);
nand U1533 (N_1533,N_819,N_1077);
xnor U1534 (N_1534,N_592,N_1171);
nand U1535 (N_1535,In_434,In_615);
and U1536 (N_1536,N_825,N_1082);
nand U1537 (N_1537,N_813,N_740);
or U1538 (N_1538,N_818,N_720);
and U1539 (N_1539,In_1567,N_1133);
and U1540 (N_1540,N_1136,N_802);
nor U1541 (N_1541,N_457,N_1158);
nand U1542 (N_1542,N_718,N_836);
nor U1543 (N_1543,In_504,In_209);
nand U1544 (N_1544,N_527,N_666);
nand U1545 (N_1545,N_1119,N_1083);
nand U1546 (N_1546,In_848,N_1127);
and U1547 (N_1547,N_434,N_1137);
xnor U1548 (N_1548,N_1045,N_952);
xnor U1549 (N_1549,In_1279,N_1060);
nand U1550 (N_1550,In_1871,N_940);
nor U1551 (N_1551,N_1191,N_1062);
xor U1552 (N_1552,N_830,N_97);
and U1553 (N_1553,In_991,In_1885);
nor U1554 (N_1554,N_86,N_1093);
or U1555 (N_1555,N_879,N_858);
nor U1556 (N_1556,N_956,In_1902);
xor U1557 (N_1557,N_90,N_919);
or U1558 (N_1558,In_1959,N_1170);
and U1559 (N_1559,N_1160,In_1632);
xnor U1560 (N_1560,N_890,In_932);
and U1561 (N_1561,N_711,In_1647);
xnor U1562 (N_1562,In_916,N_644);
nand U1563 (N_1563,N_853,N_688);
xor U1564 (N_1564,N_854,N_1024);
and U1565 (N_1565,N_869,In_23);
and U1566 (N_1566,In_951,N_1181);
nor U1567 (N_1567,N_676,In_1824);
xnor U1568 (N_1568,N_1193,N_182);
xnor U1569 (N_1569,In_578,N_700);
or U1570 (N_1570,In_1193,N_1074);
nand U1571 (N_1571,N_908,N_169);
or U1572 (N_1572,N_420,N_3);
or U1573 (N_1573,N_1147,N_1097);
or U1574 (N_1574,N_601,In_221);
and U1575 (N_1575,N_403,N_1121);
nand U1576 (N_1576,N_1099,In_1057);
and U1577 (N_1577,In_501,N_891);
nor U1578 (N_1578,N_354,N_1020);
and U1579 (N_1579,N_954,N_800);
and U1580 (N_1580,N_132,In_301);
nor U1581 (N_1581,N_1052,In_581);
or U1582 (N_1582,In_1070,N_694);
or U1583 (N_1583,In_1856,N_1113);
nand U1584 (N_1584,N_993,N_948);
nor U1585 (N_1585,In_1498,N_1123);
nand U1586 (N_1586,N_449,In_80);
xor U1587 (N_1587,N_839,N_719);
and U1588 (N_1588,In_650,N_1092);
nor U1589 (N_1589,N_902,N_321);
nand U1590 (N_1590,N_1057,N_1111);
and U1591 (N_1591,N_629,N_1041);
and U1592 (N_1592,N_888,N_699);
nand U1593 (N_1593,N_968,N_1177);
xor U1594 (N_1594,N_881,N_500);
xnor U1595 (N_1595,N_723,N_938);
nand U1596 (N_1596,N_1108,In_1396);
or U1597 (N_1597,In_1472,N_884);
and U1598 (N_1598,N_990,N_42);
and U1599 (N_1599,N_1084,N_628);
nand U1600 (N_1600,N_1382,N_1304);
nor U1601 (N_1601,N_1437,N_1515);
xor U1602 (N_1602,N_1340,N_1541);
nand U1603 (N_1603,N_1488,N_1267);
nor U1604 (N_1604,N_1457,N_1396);
nor U1605 (N_1605,N_1246,N_1463);
nand U1606 (N_1606,N_1429,N_1263);
nand U1607 (N_1607,N_1313,N_1392);
and U1608 (N_1608,N_1512,N_1308);
nand U1609 (N_1609,N_1534,N_1579);
and U1610 (N_1610,N_1228,N_1368);
nor U1611 (N_1611,N_1493,N_1478);
xnor U1612 (N_1612,N_1558,N_1214);
or U1613 (N_1613,N_1241,N_1530);
xor U1614 (N_1614,N_1443,N_1568);
or U1615 (N_1615,N_1444,N_1551);
nor U1616 (N_1616,N_1365,N_1328);
nand U1617 (N_1617,N_1484,N_1434);
xnor U1618 (N_1618,N_1449,N_1282);
nor U1619 (N_1619,N_1486,N_1581);
nand U1620 (N_1620,N_1315,N_1350);
or U1621 (N_1621,N_1435,N_1317);
and U1622 (N_1622,N_1371,N_1285);
or U1623 (N_1623,N_1465,N_1335);
xnor U1624 (N_1624,N_1270,N_1599);
xnor U1625 (N_1625,N_1527,N_1519);
and U1626 (N_1626,N_1283,N_1320);
nor U1627 (N_1627,N_1569,N_1381);
nor U1628 (N_1628,N_1497,N_1580);
and U1629 (N_1629,N_1255,N_1409);
nand U1630 (N_1630,N_1563,N_1573);
xnor U1631 (N_1631,N_1464,N_1204);
xnor U1632 (N_1632,N_1362,N_1375);
nor U1633 (N_1633,N_1510,N_1404);
or U1634 (N_1634,N_1383,N_1532);
nor U1635 (N_1635,N_1230,N_1298);
or U1636 (N_1636,N_1252,N_1289);
nor U1637 (N_1637,N_1203,N_1379);
nor U1638 (N_1638,N_1215,N_1394);
xor U1639 (N_1639,N_1451,N_1248);
nand U1640 (N_1640,N_1456,N_1454);
nand U1641 (N_1641,N_1250,N_1413);
xnor U1642 (N_1642,N_1301,N_1278);
nor U1643 (N_1643,N_1397,N_1567);
and U1644 (N_1644,N_1591,N_1574);
xor U1645 (N_1645,N_1277,N_1296);
and U1646 (N_1646,N_1374,N_1555);
or U1647 (N_1647,N_1483,N_1564);
nand U1648 (N_1648,N_1407,N_1238);
and U1649 (N_1649,N_1535,N_1207);
nand U1650 (N_1650,N_1405,N_1229);
nor U1651 (N_1651,N_1560,N_1205);
and U1652 (N_1652,N_1377,N_1403);
nor U1653 (N_1653,N_1467,N_1244);
xor U1654 (N_1654,N_1254,N_1466);
nand U1655 (N_1655,N_1516,N_1589);
and U1656 (N_1656,N_1453,N_1299);
or U1657 (N_1657,N_1520,N_1480);
or U1658 (N_1658,N_1327,N_1352);
or U1659 (N_1659,N_1210,N_1505);
xnor U1660 (N_1660,N_1337,N_1208);
nand U1661 (N_1661,N_1524,N_1256);
and U1662 (N_1662,N_1369,N_1471);
and U1663 (N_1663,N_1389,N_1357);
or U1664 (N_1664,N_1408,N_1576);
nor U1665 (N_1665,N_1399,N_1414);
and U1666 (N_1666,N_1595,N_1543);
or U1667 (N_1667,N_1216,N_1312);
nor U1668 (N_1668,N_1322,N_1274);
xor U1669 (N_1669,N_1213,N_1552);
and U1670 (N_1670,N_1331,N_1334);
or U1671 (N_1671,N_1565,N_1354);
or U1672 (N_1672,N_1384,N_1499);
nand U1673 (N_1673,N_1423,N_1587);
nand U1674 (N_1674,N_1319,N_1291);
and U1675 (N_1675,N_1477,N_1487);
nor U1676 (N_1676,N_1273,N_1427);
and U1677 (N_1677,N_1592,N_1430);
nor U1678 (N_1678,N_1415,N_1475);
nand U1679 (N_1679,N_1523,N_1269);
nor U1680 (N_1680,N_1537,N_1402);
nand U1681 (N_1681,N_1432,N_1546);
or U1682 (N_1682,N_1549,N_1330);
nand U1683 (N_1683,N_1355,N_1458);
or U1684 (N_1684,N_1518,N_1293);
and U1685 (N_1685,N_1522,N_1421);
nor U1686 (N_1686,N_1266,N_1496);
nand U1687 (N_1687,N_1542,N_1440);
and U1688 (N_1688,N_1206,N_1276);
and U1689 (N_1689,N_1588,N_1485);
and U1690 (N_1690,N_1309,N_1598);
or U1691 (N_1691,N_1502,N_1287);
or U1692 (N_1692,N_1231,N_1221);
nand U1693 (N_1693,N_1566,N_1200);
nor U1694 (N_1694,N_1366,N_1332);
or U1695 (N_1695,N_1424,N_1311);
nor U1696 (N_1696,N_1233,N_1286);
xnor U1697 (N_1697,N_1412,N_1442);
nor U1698 (N_1698,N_1361,N_1462);
nor U1699 (N_1699,N_1447,N_1257);
or U1700 (N_1700,N_1224,N_1209);
nand U1701 (N_1701,N_1344,N_1279);
xor U1702 (N_1702,N_1507,N_1586);
or U1703 (N_1703,N_1211,N_1585);
xnor U1704 (N_1704,N_1501,N_1358);
and U1705 (N_1705,N_1220,N_1479);
and U1706 (N_1706,N_1219,N_1339);
or U1707 (N_1707,N_1259,N_1540);
and U1708 (N_1708,N_1336,N_1547);
nor U1709 (N_1709,N_1245,N_1324);
and U1710 (N_1710,N_1387,N_1356);
nand U1711 (N_1711,N_1262,N_1450);
nand U1712 (N_1712,N_1461,N_1316);
nor U1713 (N_1713,N_1329,N_1393);
and U1714 (N_1714,N_1295,N_1333);
and U1715 (N_1715,N_1420,N_1468);
nand U1716 (N_1716,N_1584,N_1575);
nor U1717 (N_1717,N_1326,N_1378);
xor U1718 (N_1718,N_1218,N_1416);
xnor U1719 (N_1719,N_1526,N_1400);
xnor U1720 (N_1720,N_1417,N_1239);
xnor U1721 (N_1721,N_1275,N_1441);
or U1722 (N_1722,N_1436,N_1360);
xnor U1723 (N_1723,N_1446,N_1272);
nand U1724 (N_1724,N_1232,N_1554);
or U1725 (N_1725,N_1583,N_1281);
xnor U1726 (N_1726,N_1376,N_1292);
nor U1727 (N_1727,N_1370,N_1433);
xor U1728 (N_1728,N_1338,N_1452);
and U1729 (N_1729,N_1556,N_1445);
and U1730 (N_1730,N_1422,N_1504);
and U1731 (N_1731,N_1348,N_1506);
xor U1732 (N_1732,N_1284,N_1226);
xor U1733 (N_1733,N_1325,N_1438);
nand U1734 (N_1734,N_1533,N_1492);
xor U1735 (N_1735,N_1349,N_1280);
and U1736 (N_1736,N_1528,N_1521);
or U1737 (N_1737,N_1428,N_1470);
nand U1738 (N_1738,N_1388,N_1237);
nand U1739 (N_1739,N_1513,N_1582);
nor U1740 (N_1740,N_1343,N_1517);
xor U1741 (N_1741,N_1559,N_1596);
xnor U1742 (N_1742,N_1491,N_1353);
nor U1743 (N_1743,N_1345,N_1290);
and U1744 (N_1744,N_1225,N_1495);
and U1745 (N_1745,N_1247,N_1472);
xor U1746 (N_1746,N_1390,N_1227);
nand U1747 (N_1747,N_1395,N_1508);
nor U1748 (N_1748,N_1489,N_1538);
and U1749 (N_1749,N_1260,N_1411);
nand U1750 (N_1750,N_1529,N_1323);
and U1751 (N_1751,N_1212,N_1373);
nand U1752 (N_1752,N_1372,N_1271);
nand U1753 (N_1753,N_1439,N_1481);
and U1754 (N_1754,N_1391,N_1494);
or U1755 (N_1755,N_1511,N_1455);
nor U1756 (N_1756,N_1473,N_1570);
or U1757 (N_1757,N_1297,N_1498);
nand U1758 (N_1758,N_1294,N_1305);
or U1759 (N_1759,N_1321,N_1341);
nor U1760 (N_1760,N_1572,N_1268);
nand U1761 (N_1761,N_1469,N_1557);
xor U1762 (N_1762,N_1240,N_1385);
nor U1763 (N_1763,N_1550,N_1406);
or U1764 (N_1764,N_1243,N_1500);
and U1765 (N_1765,N_1590,N_1426);
and U1766 (N_1766,N_1474,N_1578);
nand U1767 (N_1767,N_1431,N_1597);
or U1768 (N_1768,N_1544,N_1562);
nor U1769 (N_1769,N_1380,N_1490);
xnor U1770 (N_1770,N_1223,N_1242);
and U1771 (N_1771,N_1236,N_1201);
and U1772 (N_1772,N_1347,N_1460);
or U1773 (N_1773,N_1425,N_1548);
nor U1774 (N_1774,N_1418,N_1261);
xnor U1775 (N_1775,N_1410,N_1482);
xnor U1776 (N_1776,N_1251,N_1264);
and U1777 (N_1777,N_1419,N_1539);
or U1778 (N_1778,N_1386,N_1545);
or U1779 (N_1779,N_1363,N_1525);
and U1780 (N_1780,N_1594,N_1514);
nor U1781 (N_1781,N_1593,N_1314);
and U1782 (N_1782,N_1359,N_1258);
xnor U1783 (N_1783,N_1398,N_1367);
or U1784 (N_1784,N_1346,N_1265);
nor U1785 (N_1785,N_1342,N_1577);
and U1786 (N_1786,N_1476,N_1459);
nand U1787 (N_1787,N_1503,N_1202);
nand U1788 (N_1788,N_1561,N_1448);
or U1789 (N_1789,N_1300,N_1553);
and U1790 (N_1790,N_1571,N_1303);
nor U1791 (N_1791,N_1234,N_1351);
and U1792 (N_1792,N_1222,N_1249);
and U1793 (N_1793,N_1253,N_1364);
and U1794 (N_1794,N_1536,N_1288);
or U1795 (N_1795,N_1217,N_1318);
nor U1796 (N_1796,N_1310,N_1235);
and U1797 (N_1797,N_1306,N_1302);
nor U1798 (N_1798,N_1307,N_1509);
xor U1799 (N_1799,N_1531,N_1401);
nor U1800 (N_1800,N_1378,N_1232);
or U1801 (N_1801,N_1484,N_1257);
nor U1802 (N_1802,N_1504,N_1341);
nand U1803 (N_1803,N_1201,N_1591);
and U1804 (N_1804,N_1503,N_1322);
nor U1805 (N_1805,N_1535,N_1358);
nand U1806 (N_1806,N_1554,N_1247);
or U1807 (N_1807,N_1243,N_1502);
xnor U1808 (N_1808,N_1541,N_1584);
nor U1809 (N_1809,N_1266,N_1567);
and U1810 (N_1810,N_1404,N_1446);
nor U1811 (N_1811,N_1352,N_1594);
nor U1812 (N_1812,N_1206,N_1220);
and U1813 (N_1813,N_1368,N_1232);
and U1814 (N_1814,N_1274,N_1277);
or U1815 (N_1815,N_1245,N_1479);
and U1816 (N_1816,N_1219,N_1592);
nor U1817 (N_1817,N_1507,N_1344);
nand U1818 (N_1818,N_1352,N_1395);
nor U1819 (N_1819,N_1503,N_1216);
nand U1820 (N_1820,N_1566,N_1217);
or U1821 (N_1821,N_1378,N_1384);
nor U1822 (N_1822,N_1525,N_1341);
and U1823 (N_1823,N_1458,N_1564);
and U1824 (N_1824,N_1596,N_1509);
and U1825 (N_1825,N_1254,N_1366);
xor U1826 (N_1826,N_1270,N_1263);
nand U1827 (N_1827,N_1476,N_1317);
xnor U1828 (N_1828,N_1301,N_1274);
nor U1829 (N_1829,N_1566,N_1564);
nor U1830 (N_1830,N_1272,N_1534);
and U1831 (N_1831,N_1446,N_1385);
xnor U1832 (N_1832,N_1486,N_1476);
and U1833 (N_1833,N_1232,N_1364);
and U1834 (N_1834,N_1295,N_1332);
and U1835 (N_1835,N_1377,N_1517);
or U1836 (N_1836,N_1374,N_1263);
xor U1837 (N_1837,N_1299,N_1451);
and U1838 (N_1838,N_1400,N_1494);
xnor U1839 (N_1839,N_1228,N_1441);
nand U1840 (N_1840,N_1468,N_1257);
nor U1841 (N_1841,N_1367,N_1275);
xnor U1842 (N_1842,N_1469,N_1211);
xnor U1843 (N_1843,N_1311,N_1227);
and U1844 (N_1844,N_1504,N_1206);
or U1845 (N_1845,N_1547,N_1493);
xor U1846 (N_1846,N_1480,N_1321);
xnor U1847 (N_1847,N_1532,N_1500);
and U1848 (N_1848,N_1345,N_1447);
nand U1849 (N_1849,N_1290,N_1373);
nand U1850 (N_1850,N_1251,N_1482);
xnor U1851 (N_1851,N_1546,N_1319);
or U1852 (N_1852,N_1438,N_1592);
nor U1853 (N_1853,N_1262,N_1485);
or U1854 (N_1854,N_1209,N_1489);
nor U1855 (N_1855,N_1272,N_1345);
nand U1856 (N_1856,N_1540,N_1233);
nor U1857 (N_1857,N_1288,N_1256);
or U1858 (N_1858,N_1596,N_1503);
nor U1859 (N_1859,N_1443,N_1338);
xor U1860 (N_1860,N_1531,N_1542);
nand U1861 (N_1861,N_1493,N_1462);
xnor U1862 (N_1862,N_1232,N_1222);
and U1863 (N_1863,N_1336,N_1465);
nor U1864 (N_1864,N_1214,N_1293);
or U1865 (N_1865,N_1231,N_1228);
nand U1866 (N_1866,N_1536,N_1315);
or U1867 (N_1867,N_1211,N_1349);
nor U1868 (N_1868,N_1230,N_1470);
or U1869 (N_1869,N_1376,N_1488);
and U1870 (N_1870,N_1381,N_1209);
xor U1871 (N_1871,N_1511,N_1357);
and U1872 (N_1872,N_1349,N_1208);
xnor U1873 (N_1873,N_1298,N_1530);
nor U1874 (N_1874,N_1597,N_1566);
xor U1875 (N_1875,N_1556,N_1451);
nand U1876 (N_1876,N_1211,N_1450);
or U1877 (N_1877,N_1204,N_1521);
and U1878 (N_1878,N_1469,N_1365);
nand U1879 (N_1879,N_1337,N_1233);
and U1880 (N_1880,N_1582,N_1330);
nor U1881 (N_1881,N_1450,N_1323);
nor U1882 (N_1882,N_1307,N_1470);
xnor U1883 (N_1883,N_1553,N_1547);
xnor U1884 (N_1884,N_1520,N_1218);
nand U1885 (N_1885,N_1212,N_1433);
nor U1886 (N_1886,N_1330,N_1204);
nand U1887 (N_1887,N_1323,N_1366);
nand U1888 (N_1888,N_1375,N_1580);
or U1889 (N_1889,N_1332,N_1244);
nor U1890 (N_1890,N_1477,N_1334);
nor U1891 (N_1891,N_1200,N_1360);
nand U1892 (N_1892,N_1221,N_1535);
or U1893 (N_1893,N_1428,N_1472);
nand U1894 (N_1894,N_1346,N_1403);
nor U1895 (N_1895,N_1587,N_1581);
or U1896 (N_1896,N_1237,N_1292);
nand U1897 (N_1897,N_1245,N_1346);
xnor U1898 (N_1898,N_1336,N_1470);
nand U1899 (N_1899,N_1204,N_1428);
and U1900 (N_1900,N_1383,N_1505);
nand U1901 (N_1901,N_1573,N_1360);
xnor U1902 (N_1902,N_1351,N_1567);
nor U1903 (N_1903,N_1452,N_1439);
nor U1904 (N_1904,N_1232,N_1419);
or U1905 (N_1905,N_1257,N_1266);
or U1906 (N_1906,N_1395,N_1292);
and U1907 (N_1907,N_1584,N_1203);
nor U1908 (N_1908,N_1270,N_1284);
xnor U1909 (N_1909,N_1216,N_1310);
nor U1910 (N_1910,N_1231,N_1294);
xnor U1911 (N_1911,N_1447,N_1329);
nand U1912 (N_1912,N_1312,N_1337);
and U1913 (N_1913,N_1431,N_1509);
and U1914 (N_1914,N_1220,N_1369);
nor U1915 (N_1915,N_1489,N_1491);
or U1916 (N_1916,N_1507,N_1479);
xnor U1917 (N_1917,N_1469,N_1207);
nand U1918 (N_1918,N_1370,N_1525);
and U1919 (N_1919,N_1597,N_1507);
xor U1920 (N_1920,N_1572,N_1384);
nand U1921 (N_1921,N_1422,N_1208);
nor U1922 (N_1922,N_1441,N_1298);
nor U1923 (N_1923,N_1409,N_1245);
nand U1924 (N_1924,N_1424,N_1448);
or U1925 (N_1925,N_1570,N_1542);
nor U1926 (N_1926,N_1236,N_1307);
nor U1927 (N_1927,N_1322,N_1345);
or U1928 (N_1928,N_1335,N_1325);
nand U1929 (N_1929,N_1357,N_1474);
nand U1930 (N_1930,N_1258,N_1481);
and U1931 (N_1931,N_1360,N_1504);
nor U1932 (N_1932,N_1307,N_1300);
nor U1933 (N_1933,N_1375,N_1487);
or U1934 (N_1934,N_1464,N_1341);
nand U1935 (N_1935,N_1303,N_1216);
or U1936 (N_1936,N_1434,N_1400);
xnor U1937 (N_1937,N_1534,N_1468);
and U1938 (N_1938,N_1317,N_1453);
or U1939 (N_1939,N_1358,N_1544);
or U1940 (N_1940,N_1232,N_1244);
nand U1941 (N_1941,N_1287,N_1290);
nor U1942 (N_1942,N_1530,N_1473);
and U1943 (N_1943,N_1578,N_1329);
and U1944 (N_1944,N_1472,N_1509);
or U1945 (N_1945,N_1315,N_1466);
and U1946 (N_1946,N_1334,N_1506);
nand U1947 (N_1947,N_1549,N_1200);
nor U1948 (N_1948,N_1269,N_1379);
nor U1949 (N_1949,N_1496,N_1401);
nor U1950 (N_1950,N_1573,N_1389);
nand U1951 (N_1951,N_1224,N_1241);
or U1952 (N_1952,N_1354,N_1285);
nand U1953 (N_1953,N_1552,N_1516);
xor U1954 (N_1954,N_1408,N_1547);
or U1955 (N_1955,N_1571,N_1451);
or U1956 (N_1956,N_1264,N_1550);
nor U1957 (N_1957,N_1405,N_1455);
nand U1958 (N_1958,N_1523,N_1501);
or U1959 (N_1959,N_1476,N_1512);
and U1960 (N_1960,N_1555,N_1548);
and U1961 (N_1961,N_1202,N_1277);
xor U1962 (N_1962,N_1236,N_1377);
nand U1963 (N_1963,N_1277,N_1405);
xor U1964 (N_1964,N_1587,N_1430);
nand U1965 (N_1965,N_1373,N_1445);
and U1966 (N_1966,N_1590,N_1558);
and U1967 (N_1967,N_1588,N_1432);
nor U1968 (N_1968,N_1472,N_1348);
and U1969 (N_1969,N_1436,N_1367);
and U1970 (N_1970,N_1231,N_1333);
nor U1971 (N_1971,N_1500,N_1230);
nand U1972 (N_1972,N_1419,N_1422);
and U1973 (N_1973,N_1557,N_1490);
nor U1974 (N_1974,N_1279,N_1245);
and U1975 (N_1975,N_1547,N_1302);
and U1976 (N_1976,N_1334,N_1244);
nor U1977 (N_1977,N_1543,N_1482);
nand U1978 (N_1978,N_1304,N_1279);
nor U1979 (N_1979,N_1432,N_1490);
xor U1980 (N_1980,N_1305,N_1395);
and U1981 (N_1981,N_1255,N_1264);
nand U1982 (N_1982,N_1577,N_1372);
nor U1983 (N_1983,N_1211,N_1545);
nor U1984 (N_1984,N_1406,N_1353);
nand U1985 (N_1985,N_1482,N_1428);
or U1986 (N_1986,N_1257,N_1344);
nor U1987 (N_1987,N_1566,N_1323);
and U1988 (N_1988,N_1530,N_1506);
and U1989 (N_1989,N_1292,N_1202);
xnor U1990 (N_1990,N_1304,N_1222);
nor U1991 (N_1991,N_1509,N_1501);
nor U1992 (N_1992,N_1432,N_1429);
nor U1993 (N_1993,N_1588,N_1552);
and U1994 (N_1994,N_1507,N_1217);
nand U1995 (N_1995,N_1543,N_1272);
xor U1996 (N_1996,N_1254,N_1275);
or U1997 (N_1997,N_1243,N_1226);
nand U1998 (N_1998,N_1450,N_1590);
nor U1999 (N_1999,N_1365,N_1537);
and U2000 (N_2000,N_1908,N_1650);
nand U2001 (N_2001,N_1923,N_1994);
xor U2002 (N_2002,N_1892,N_1724);
nand U2003 (N_2003,N_1815,N_1718);
and U2004 (N_2004,N_1922,N_1970);
xnor U2005 (N_2005,N_1877,N_1821);
or U2006 (N_2006,N_1887,N_1961);
nand U2007 (N_2007,N_1969,N_1758);
nor U2008 (N_2008,N_1782,N_1742);
and U2009 (N_2009,N_1940,N_1988);
nor U2010 (N_2010,N_1809,N_1791);
and U2011 (N_2011,N_1703,N_1993);
xor U2012 (N_2012,N_1691,N_1657);
nand U2013 (N_2013,N_1751,N_1654);
or U2014 (N_2014,N_1826,N_1955);
or U2015 (N_2015,N_1768,N_1646);
and U2016 (N_2016,N_1604,N_1671);
xnor U2017 (N_2017,N_1784,N_1824);
and U2018 (N_2018,N_1865,N_1631);
nor U2019 (N_2019,N_1644,N_1800);
and U2020 (N_2020,N_1666,N_1793);
nor U2021 (N_2021,N_1998,N_1948);
nand U2022 (N_2022,N_1947,N_1937);
or U2023 (N_2023,N_1803,N_1856);
nand U2024 (N_2024,N_1950,N_1978);
and U2025 (N_2025,N_1706,N_1665);
nor U2026 (N_2026,N_1959,N_1907);
and U2027 (N_2027,N_1910,N_1629);
nor U2028 (N_2028,N_1769,N_1863);
nand U2029 (N_2029,N_1932,N_1693);
and U2030 (N_2030,N_1726,N_1879);
nand U2031 (N_2031,N_1899,N_1641);
or U2032 (N_2032,N_1684,N_1891);
and U2033 (N_2033,N_1740,N_1913);
or U2034 (N_2034,N_1929,N_1977);
or U2035 (N_2035,N_1674,N_1837);
nor U2036 (N_2036,N_1933,N_1872);
and U2037 (N_2037,N_1976,N_1717);
and U2038 (N_2038,N_1602,N_1788);
and U2039 (N_2039,N_1660,N_1997);
xor U2040 (N_2040,N_1612,N_1886);
and U2041 (N_2041,N_1944,N_1683);
or U2042 (N_2042,N_1920,N_1761);
or U2043 (N_2043,N_1714,N_1668);
nor U2044 (N_2044,N_1888,N_1772);
xor U2045 (N_2045,N_1980,N_1614);
xor U2046 (N_2046,N_1915,N_1607);
or U2047 (N_2047,N_1628,N_1849);
nor U2048 (N_2048,N_1708,N_1797);
and U2049 (N_2049,N_1831,N_1647);
and U2050 (N_2050,N_1799,N_1605);
nor U2051 (N_2051,N_1619,N_1906);
nor U2052 (N_2052,N_1636,N_1852);
xor U2053 (N_2053,N_1720,N_1697);
nand U2054 (N_2054,N_1990,N_1696);
nand U2055 (N_2055,N_1673,N_1971);
xor U2056 (N_2056,N_1652,N_1750);
xor U2057 (N_2057,N_1889,N_1858);
or U2058 (N_2058,N_1973,N_1658);
and U2059 (N_2059,N_1830,N_1667);
xor U2060 (N_2060,N_1918,N_1729);
nand U2061 (N_2061,N_1999,N_1859);
or U2062 (N_2062,N_1618,N_1873);
nand U2063 (N_2063,N_1912,N_1635);
xor U2064 (N_2064,N_1785,N_1651);
nand U2065 (N_2065,N_1956,N_1862);
or U2066 (N_2066,N_1741,N_1765);
nor U2067 (N_2067,N_1927,N_1871);
xor U2068 (N_2068,N_1695,N_1627);
nor U2069 (N_2069,N_1968,N_1883);
nand U2070 (N_2070,N_1848,N_1710);
xnor U2071 (N_2071,N_1952,N_1975);
xor U2072 (N_2072,N_1745,N_1662);
nand U2073 (N_2073,N_1924,N_1818);
and U2074 (N_2074,N_1846,N_1916);
or U2075 (N_2075,N_1960,N_1909);
and U2076 (N_2076,N_1637,N_1656);
and U2077 (N_2077,N_1639,N_1752);
xnor U2078 (N_2078,N_1935,N_1680);
or U2079 (N_2079,N_1953,N_1609);
nand U2080 (N_2080,N_1634,N_1885);
xor U2081 (N_2081,N_1930,N_1640);
or U2082 (N_2082,N_1896,N_1755);
xor U2083 (N_2083,N_1857,N_1806);
or U2084 (N_2084,N_1638,N_1620);
nor U2085 (N_2085,N_1866,N_1672);
nand U2086 (N_2086,N_1825,N_1611);
and U2087 (N_2087,N_1995,N_1814);
or U2088 (N_2088,N_1775,N_1766);
nand U2089 (N_2089,N_1670,N_1794);
or U2090 (N_2090,N_1738,N_1781);
nor U2091 (N_2091,N_1874,N_1748);
xor U2092 (N_2092,N_1867,N_1798);
nand U2093 (N_2093,N_1938,N_1834);
and U2094 (N_2094,N_1942,N_1633);
and U2095 (N_2095,N_1838,N_1880);
or U2096 (N_2096,N_1901,N_1914);
nor U2097 (N_2097,N_1902,N_1664);
or U2098 (N_2098,N_1804,N_1876);
or U2099 (N_2099,N_1931,N_1951);
and U2100 (N_2100,N_1983,N_1965);
nor U2101 (N_2101,N_1987,N_1919);
xor U2102 (N_2102,N_1836,N_1823);
or U2103 (N_2103,N_1796,N_1839);
xor U2104 (N_2104,N_1991,N_1756);
xnor U2105 (N_2105,N_1707,N_1967);
nand U2106 (N_2106,N_1985,N_1686);
xnor U2107 (N_2107,N_1669,N_1810);
xor U2108 (N_2108,N_1763,N_1712);
xnor U2109 (N_2109,N_1648,N_1747);
xnor U2110 (N_2110,N_1685,N_1934);
nand U2111 (N_2111,N_1786,N_1767);
nand U2112 (N_2112,N_1925,N_1676);
nand U2113 (N_2113,N_1954,N_1698);
nor U2114 (N_2114,N_1832,N_1701);
nand U2115 (N_2115,N_1958,N_1939);
and U2116 (N_2116,N_1911,N_1704);
or U2117 (N_2117,N_1816,N_1736);
nor U2118 (N_2118,N_1783,N_1900);
nor U2119 (N_2119,N_1760,N_1805);
and U2120 (N_2120,N_1817,N_1875);
xor U2121 (N_2121,N_1844,N_1904);
nor U2122 (N_2122,N_1600,N_1711);
or U2123 (N_2123,N_1719,N_1715);
nor U2124 (N_2124,N_1770,N_1762);
xor U2125 (N_2125,N_1861,N_1700);
nand U2126 (N_2126,N_1677,N_1655);
xnor U2127 (N_2127,N_1716,N_1776);
or U2128 (N_2128,N_1966,N_1851);
and U2129 (N_2129,N_1835,N_1992);
or U2130 (N_2130,N_1606,N_1820);
and U2131 (N_2131,N_1897,N_1989);
nor U2132 (N_2132,N_1645,N_1709);
or U2133 (N_2133,N_1984,N_1661);
or U2134 (N_2134,N_1903,N_1890);
nand U2135 (N_2135,N_1869,N_1884);
or U2136 (N_2136,N_1898,N_1699);
nor U2137 (N_2137,N_1649,N_1854);
nor U2138 (N_2138,N_1840,N_1790);
nand U2139 (N_2139,N_1653,N_1812);
or U2140 (N_2140,N_1759,N_1739);
nand U2141 (N_2141,N_1822,N_1957);
nor U2142 (N_2142,N_1833,N_1624);
xor U2143 (N_2143,N_1626,N_1829);
nand U2144 (N_2144,N_1981,N_1894);
and U2145 (N_2145,N_1663,N_1705);
and U2146 (N_2146,N_1771,N_1679);
nor U2147 (N_2147,N_1643,N_1725);
nand U2148 (N_2148,N_1690,N_1795);
and U2149 (N_2149,N_1774,N_1789);
xnor U2150 (N_2150,N_1905,N_1949);
nor U2151 (N_2151,N_1630,N_1926);
nand U2152 (N_2152,N_1749,N_1731);
or U2153 (N_2153,N_1728,N_1623);
nand U2154 (N_2154,N_1603,N_1689);
and U2155 (N_2155,N_1855,N_1702);
nor U2156 (N_2156,N_1625,N_1632);
or U2157 (N_2157,N_1675,N_1733);
and U2158 (N_2158,N_1850,N_1737);
or U2159 (N_2159,N_1946,N_1764);
and U2160 (N_2160,N_1746,N_1881);
nor U2161 (N_2161,N_1827,N_1744);
nor U2162 (N_2162,N_1694,N_1882);
nand U2163 (N_2163,N_1681,N_1878);
or U2164 (N_2164,N_1853,N_1687);
nor U2165 (N_2165,N_1610,N_1682);
nor U2166 (N_2166,N_1659,N_1842);
nor U2167 (N_2167,N_1979,N_1678);
and U2168 (N_2168,N_1688,N_1864);
nand U2169 (N_2169,N_1787,N_1895);
and U2170 (N_2170,N_1613,N_1870);
nand U2171 (N_2171,N_1928,N_1847);
or U2172 (N_2172,N_1941,N_1962);
or U2173 (N_2173,N_1811,N_1721);
and U2174 (N_2174,N_1743,N_1779);
and U2175 (N_2175,N_1921,N_1723);
or U2176 (N_2176,N_1843,N_1730);
nor U2177 (N_2177,N_1996,N_1601);
or U2178 (N_2178,N_1828,N_1972);
nor U2179 (N_2179,N_1753,N_1642);
xor U2180 (N_2180,N_1974,N_1792);
nand U2181 (N_2181,N_1964,N_1773);
nand U2182 (N_2182,N_1801,N_1616);
nand U2183 (N_2183,N_1893,N_1917);
nand U2184 (N_2184,N_1986,N_1732);
nand U2185 (N_2185,N_1819,N_1617);
nor U2186 (N_2186,N_1722,N_1735);
nand U2187 (N_2187,N_1802,N_1777);
and U2188 (N_2188,N_1813,N_1780);
or U2189 (N_2189,N_1778,N_1757);
xor U2190 (N_2190,N_1734,N_1868);
nand U2191 (N_2191,N_1807,N_1808);
or U2192 (N_2192,N_1845,N_1622);
and U2193 (N_2193,N_1754,N_1982);
nand U2194 (N_2194,N_1841,N_1860);
xor U2195 (N_2195,N_1727,N_1713);
or U2196 (N_2196,N_1608,N_1945);
nor U2197 (N_2197,N_1936,N_1621);
nand U2198 (N_2198,N_1963,N_1615);
or U2199 (N_2199,N_1692,N_1943);
xnor U2200 (N_2200,N_1642,N_1608);
nand U2201 (N_2201,N_1761,N_1606);
or U2202 (N_2202,N_1632,N_1743);
xor U2203 (N_2203,N_1818,N_1695);
nand U2204 (N_2204,N_1852,N_1912);
nand U2205 (N_2205,N_1924,N_1608);
xor U2206 (N_2206,N_1716,N_1663);
or U2207 (N_2207,N_1733,N_1809);
xnor U2208 (N_2208,N_1650,N_1727);
and U2209 (N_2209,N_1724,N_1986);
nor U2210 (N_2210,N_1947,N_1761);
nand U2211 (N_2211,N_1672,N_1964);
xnor U2212 (N_2212,N_1966,N_1920);
or U2213 (N_2213,N_1634,N_1739);
nand U2214 (N_2214,N_1678,N_1606);
and U2215 (N_2215,N_1745,N_1764);
or U2216 (N_2216,N_1682,N_1605);
or U2217 (N_2217,N_1639,N_1645);
and U2218 (N_2218,N_1709,N_1726);
xor U2219 (N_2219,N_1869,N_1864);
nand U2220 (N_2220,N_1640,N_1629);
xor U2221 (N_2221,N_1726,N_1790);
nor U2222 (N_2222,N_1605,N_1744);
and U2223 (N_2223,N_1956,N_1738);
nor U2224 (N_2224,N_1620,N_1997);
xor U2225 (N_2225,N_1645,N_1882);
or U2226 (N_2226,N_1657,N_1748);
or U2227 (N_2227,N_1799,N_1718);
xnor U2228 (N_2228,N_1944,N_1929);
or U2229 (N_2229,N_1920,N_1646);
nor U2230 (N_2230,N_1645,N_1947);
and U2231 (N_2231,N_1953,N_1924);
or U2232 (N_2232,N_1968,N_1772);
and U2233 (N_2233,N_1891,N_1821);
or U2234 (N_2234,N_1935,N_1803);
nand U2235 (N_2235,N_1716,N_1679);
nand U2236 (N_2236,N_1950,N_1917);
nor U2237 (N_2237,N_1736,N_1937);
nand U2238 (N_2238,N_1630,N_1835);
nand U2239 (N_2239,N_1742,N_1741);
or U2240 (N_2240,N_1635,N_1975);
and U2241 (N_2241,N_1998,N_1681);
or U2242 (N_2242,N_1966,N_1879);
or U2243 (N_2243,N_1602,N_1932);
or U2244 (N_2244,N_1956,N_1960);
xnor U2245 (N_2245,N_1984,N_1641);
and U2246 (N_2246,N_1718,N_1897);
and U2247 (N_2247,N_1670,N_1990);
nor U2248 (N_2248,N_1646,N_1824);
nor U2249 (N_2249,N_1745,N_1655);
nor U2250 (N_2250,N_1672,N_1833);
nor U2251 (N_2251,N_1664,N_1976);
nand U2252 (N_2252,N_1845,N_1631);
or U2253 (N_2253,N_1749,N_1734);
xnor U2254 (N_2254,N_1647,N_1796);
nor U2255 (N_2255,N_1909,N_1756);
nand U2256 (N_2256,N_1684,N_1922);
and U2257 (N_2257,N_1842,N_1674);
or U2258 (N_2258,N_1769,N_1698);
or U2259 (N_2259,N_1792,N_1877);
or U2260 (N_2260,N_1933,N_1713);
nand U2261 (N_2261,N_1822,N_1765);
nor U2262 (N_2262,N_1823,N_1600);
xor U2263 (N_2263,N_1726,N_1985);
or U2264 (N_2264,N_1635,N_1988);
or U2265 (N_2265,N_1828,N_1945);
or U2266 (N_2266,N_1707,N_1684);
and U2267 (N_2267,N_1869,N_1846);
nand U2268 (N_2268,N_1961,N_1699);
or U2269 (N_2269,N_1839,N_1975);
and U2270 (N_2270,N_1880,N_1913);
xnor U2271 (N_2271,N_1937,N_1751);
or U2272 (N_2272,N_1821,N_1758);
nand U2273 (N_2273,N_1620,N_1670);
or U2274 (N_2274,N_1773,N_1833);
xnor U2275 (N_2275,N_1739,N_1669);
nand U2276 (N_2276,N_1891,N_1888);
nand U2277 (N_2277,N_1854,N_1752);
nand U2278 (N_2278,N_1689,N_1679);
xnor U2279 (N_2279,N_1891,N_1885);
or U2280 (N_2280,N_1721,N_1852);
or U2281 (N_2281,N_1997,N_1777);
nor U2282 (N_2282,N_1957,N_1918);
nor U2283 (N_2283,N_1688,N_1790);
xor U2284 (N_2284,N_1634,N_1675);
nand U2285 (N_2285,N_1912,N_1887);
nor U2286 (N_2286,N_1716,N_1738);
or U2287 (N_2287,N_1743,N_1872);
nand U2288 (N_2288,N_1689,N_1919);
nand U2289 (N_2289,N_1783,N_1621);
nand U2290 (N_2290,N_1769,N_1623);
nand U2291 (N_2291,N_1682,N_1831);
or U2292 (N_2292,N_1852,N_1789);
nor U2293 (N_2293,N_1870,N_1673);
or U2294 (N_2294,N_1660,N_1611);
and U2295 (N_2295,N_1823,N_1713);
nor U2296 (N_2296,N_1666,N_1951);
nor U2297 (N_2297,N_1790,N_1686);
nor U2298 (N_2298,N_1662,N_1603);
or U2299 (N_2299,N_1671,N_1632);
and U2300 (N_2300,N_1895,N_1728);
and U2301 (N_2301,N_1805,N_1672);
and U2302 (N_2302,N_1789,N_1848);
xor U2303 (N_2303,N_1775,N_1645);
xor U2304 (N_2304,N_1883,N_1971);
and U2305 (N_2305,N_1694,N_1764);
nand U2306 (N_2306,N_1963,N_1678);
or U2307 (N_2307,N_1840,N_1672);
xor U2308 (N_2308,N_1694,N_1741);
nand U2309 (N_2309,N_1915,N_1688);
nor U2310 (N_2310,N_1969,N_1775);
or U2311 (N_2311,N_1908,N_1990);
and U2312 (N_2312,N_1929,N_1911);
and U2313 (N_2313,N_1645,N_1831);
and U2314 (N_2314,N_1878,N_1613);
xor U2315 (N_2315,N_1780,N_1602);
and U2316 (N_2316,N_1897,N_1769);
and U2317 (N_2317,N_1759,N_1871);
nor U2318 (N_2318,N_1613,N_1833);
nor U2319 (N_2319,N_1965,N_1974);
and U2320 (N_2320,N_1611,N_1759);
xor U2321 (N_2321,N_1820,N_1604);
xor U2322 (N_2322,N_1866,N_1934);
or U2323 (N_2323,N_1905,N_1995);
nand U2324 (N_2324,N_1850,N_1984);
nor U2325 (N_2325,N_1751,N_1744);
nor U2326 (N_2326,N_1992,N_1928);
xnor U2327 (N_2327,N_1976,N_1855);
nor U2328 (N_2328,N_1881,N_1804);
or U2329 (N_2329,N_1691,N_1907);
nor U2330 (N_2330,N_1673,N_1825);
or U2331 (N_2331,N_1704,N_1671);
and U2332 (N_2332,N_1777,N_1978);
and U2333 (N_2333,N_1966,N_1769);
or U2334 (N_2334,N_1923,N_1630);
nand U2335 (N_2335,N_1921,N_1708);
or U2336 (N_2336,N_1909,N_1805);
and U2337 (N_2337,N_1815,N_1950);
or U2338 (N_2338,N_1896,N_1994);
nand U2339 (N_2339,N_1608,N_1903);
nor U2340 (N_2340,N_1939,N_1978);
and U2341 (N_2341,N_1714,N_1813);
and U2342 (N_2342,N_1763,N_1749);
xor U2343 (N_2343,N_1894,N_1672);
or U2344 (N_2344,N_1671,N_1681);
nor U2345 (N_2345,N_1800,N_1871);
xor U2346 (N_2346,N_1766,N_1610);
nand U2347 (N_2347,N_1762,N_1704);
nor U2348 (N_2348,N_1602,N_1962);
and U2349 (N_2349,N_1620,N_1896);
nand U2350 (N_2350,N_1703,N_1730);
nand U2351 (N_2351,N_1862,N_1646);
or U2352 (N_2352,N_1954,N_1616);
and U2353 (N_2353,N_1747,N_1925);
or U2354 (N_2354,N_1795,N_1624);
and U2355 (N_2355,N_1903,N_1869);
and U2356 (N_2356,N_1742,N_1744);
nand U2357 (N_2357,N_1900,N_1838);
or U2358 (N_2358,N_1909,N_1714);
xor U2359 (N_2359,N_1867,N_1718);
and U2360 (N_2360,N_1729,N_1872);
nand U2361 (N_2361,N_1892,N_1646);
xor U2362 (N_2362,N_1853,N_1920);
xor U2363 (N_2363,N_1942,N_1718);
nor U2364 (N_2364,N_1708,N_1986);
xor U2365 (N_2365,N_1798,N_1709);
nand U2366 (N_2366,N_1963,N_1986);
or U2367 (N_2367,N_1835,N_1929);
and U2368 (N_2368,N_1705,N_1700);
or U2369 (N_2369,N_1685,N_1932);
or U2370 (N_2370,N_1910,N_1808);
xnor U2371 (N_2371,N_1650,N_1627);
and U2372 (N_2372,N_1873,N_1901);
nand U2373 (N_2373,N_1888,N_1707);
and U2374 (N_2374,N_1645,N_1779);
and U2375 (N_2375,N_1912,N_1610);
nand U2376 (N_2376,N_1983,N_1629);
nand U2377 (N_2377,N_1830,N_1758);
xnor U2378 (N_2378,N_1945,N_1873);
xnor U2379 (N_2379,N_1728,N_1961);
xor U2380 (N_2380,N_1989,N_1980);
and U2381 (N_2381,N_1975,N_1698);
or U2382 (N_2382,N_1886,N_1993);
nor U2383 (N_2383,N_1709,N_1846);
and U2384 (N_2384,N_1700,N_1701);
nand U2385 (N_2385,N_1962,N_1736);
xor U2386 (N_2386,N_1816,N_1925);
xor U2387 (N_2387,N_1987,N_1989);
nor U2388 (N_2388,N_1952,N_1690);
nand U2389 (N_2389,N_1970,N_1627);
or U2390 (N_2390,N_1627,N_1714);
or U2391 (N_2391,N_1627,N_1721);
or U2392 (N_2392,N_1932,N_1850);
xnor U2393 (N_2393,N_1905,N_1748);
nand U2394 (N_2394,N_1609,N_1704);
nor U2395 (N_2395,N_1986,N_1792);
xnor U2396 (N_2396,N_1933,N_1613);
and U2397 (N_2397,N_1723,N_1717);
nand U2398 (N_2398,N_1619,N_1806);
nor U2399 (N_2399,N_1624,N_1787);
xnor U2400 (N_2400,N_2260,N_2290);
xor U2401 (N_2401,N_2148,N_2326);
nor U2402 (N_2402,N_2024,N_2325);
xor U2403 (N_2403,N_2268,N_2191);
xor U2404 (N_2404,N_2380,N_2309);
nor U2405 (N_2405,N_2033,N_2040);
and U2406 (N_2406,N_2299,N_2264);
xnor U2407 (N_2407,N_2133,N_2188);
or U2408 (N_2408,N_2317,N_2130);
and U2409 (N_2409,N_2289,N_2263);
and U2410 (N_2410,N_2127,N_2386);
or U2411 (N_2411,N_2377,N_2347);
or U2412 (N_2412,N_2054,N_2097);
nand U2413 (N_2413,N_2167,N_2351);
xor U2414 (N_2414,N_2031,N_2261);
or U2415 (N_2415,N_2052,N_2006);
nor U2416 (N_2416,N_2172,N_2275);
nand U2417 (N_2417,N_2335,N_2321);
nor U2418 (N_2418,N_2310,N_2371);
nand U2419 (N_2419,N_2039,N_2147);
nand U2420 (N_2420,N_2233,N_2217);
nand U2421 (N_2421,N_2228,N_2274);
xnor U2422 (N_2422,N_2305,N_2164);
nor U2423 (N_2423,N_2354,N_2041);
and U2424 (N_2424,N_2334,N_2266);
nor U2425 (N_2425,N_2009,N_2062);
and U2426 (N_2426,N_2047,N_2219);
nor U2427 (N_2427,N_2118,N_2091);
nand U2428 (N_2428,N_2243,N_2005);
xnor U2429 (N_2429,N_2012,N_2336);
nand U2430 (N_2430,N_2358,N_2110);
xor U2431 (N_2431,N_2314,N_2270);
and U2432 (N_2432,N_2245,N_2103);
nand U2433 (N_2433,N_2035,N_2315);
nor U2434 (N_2434,N_2066,N_2341);
or U2435 (N_2435,N_2220,N_2144);
and U2436 (N_2436,N_2160,N_2252);
nand U2437 (N_2437,N_2156,N_2124);
nor U2438 (N_2438,N_2286,N_2378);
nor U2439 (N_2439,N_2072,N_2011);
or U2440 (N_2440,N_2185,N_2318);
xnor U2441 (N_2441,N_2203,N_2152);
nor U2442 (N_2442,N_2229,N_2165);
nand U2443 (N_2443,N_2170,N_2368);
nor U2444 (N_2444,N_2319,N_2272);
or U2445 (N_2445,N_2355,N_2149);
and U2446 (N_2446,N_2273,N_2051);
xor U2447 (N_2447,N_2007,N_2365);
xnor U2448 (N_2448,N_2095,N_2308);
nand U2449 (N_2449,N_2253,N_2096);
xnor U2450 (N_2450,N_2232,N_2221);
and U2451 (N_2451,N_2000,N_2019);
nor U2452 (N_2452,N_2028,N_2399);
nand U2453 (N_2453,N_2080,N_2076);
nand U2454 (N_2454,N_2282,N_2171);
and U2455 (N_2455,N_2114,N_2213);
and U2456 (N_2456,N_2364,N_2129);
nand U2457 (N_2457,N_2078,N_2366);
xor U2458 (N_2458,N_2394,N_2269);
or U2459 (N_2459,N_2075,N_2283);
or U2460 (N_2460,N_2117,N_2057);
and U2461 (N_2461,N_2254,N_2257);
or U2462 (N_2462,N_2388,N_2176);
nor U2463 (N_2463,N_2086,N_2045);
or U2464 (N_2464,N_2116,N_2064);
nor U2465 (N_2465,N_2359,N_2175);
xnor U2466 (N_2466,N_2125,N_2048);
nand U2467 (N_2467,N_2251,N_2293);
and U2468 (N_2468,N_2332,N_2145);
nand U2469 (N_2469,N_2242,N_2015);
xnor U2470 (N_2470,N_2003,N_2224);
nand U2471 (N_2471,N_2324,N_2155);
and U2472 (N_2472,N_2139,N_2383);
nand U2473 (N_2473,N_2053,N_2265);
or U2474 (N_2474,N_2025,N_2333);
nor U2475 (N_2475,N_2046,N_2258);
or U2476 (N_2476,N_2250,N_2307);
nand U2477 (N_2477,N_2288,N_2141);
nor U2478 (N_2478,N_2073,N_2234);
or U2479 (N_2479,N_2082,N_2063);
or U2480 (N_2480,N_2302,N_2222);
xnor U2481 (N_2481,N_2236,N_2193);
xnor U2482 (N_2482,N_2043,N_2137);
xor U2483 (N_2483,N_2225,N_2346);
nor U2484 (N_2484,N_2344,N_2140);
and U2485 (N_2485,N_2143,N_2120);
or U2486 (N_2486,N_2036,N_2178);
and U2487 (N_2487,N_2099,N_2104);
xor U2488 (N_2488,N_2074,N_2131);
nand U2489 (N_2489,N_2187,N_2350);
xor U2490 (N_2490,N_2056,N_2259);
xor U2491 (N_2491,N_2026,N_2146);
xor U2492 (N_2492,N_2281,N_2360);
or U2493 (N_2493,N_2018,N_2198);
xor U2494 (N_2494,N_2352,N_2239);
xor U2495 (N_2495,N_2181,N_2055);
xor U2496 (N_2496,N_2134,N_2010);
xor U2497 (N_2497,N_2215,N_2226);
and U2498 (N_2498,N_2372,N_2235);
xnor U2499 (N_2499,N_2398,N_2353);
xnor U2500 (N_2500,N_2022,N_2381);
xor U2501 (N_2501,N_2108,N_2285);
nor U2502 (N_2502,N_2013,N_2295);
nand U2503 (N_2503,N_2238,N_2122);
and U2504 (N_2504,N_2329,N_2162);
and U2505 (N_2505,N_2060,N_2065);
or U2506 (N_2506,N_2348,N_2277);
or U2507 (N_2507,N_2241,N_2397);
nor U2508 (N_2508,N_2304,N_2030);
nor U2509 (N_2509,N_2361,N_2008);
nor U2510 (N_2510,N_2356,N_2159);
or U2511 (N_2511,N_2322,N_2303);
and U2512 (N_2512,N_2231,N_2296);
nor U2513 (N_2513,N_2083,N_2312);
or U2514 (N_2514,N_2115,N_2338);
or U2515 (N_2515,N_2195,N_2100);
xor U2516 (N_2516,N_2330,N_2392);
or U2517 (N_2517,N_2306,N_2343);
or U2518 (N_2518,N_2384,N_2089);
xnor U2519 (N_2519,N_2342,N_2136);
nand U2520 (N_2520,N_2205,N_2262);
and U2521 (N_2521,N_2177,N_2301);
xnor U2522 (N_2522,N_2379,N_2123);
nand U2523 (N_2523,N_2246,N_2363);
or U2524 (N_2524,N_2186,N_2367);
or U2525 (N_2525,N_2339,N_2138);
xor U2526 (N_2526,N_2373,N_2227);
and U2527 (N_2527,N_2151,N_2174);
xor U2528 (N_2528,N_2092,N_2199);
nor U2529 (N_2529,N_2349,N_2284);
or U2530 (N_2530,N_2158,N_2207);
and U2531 (N_2531,N_2393,N_2069);
nor U2532 (N_2532,N_2102,N_2087);
xor U2533 (N_2533,N_2396,N_2044);
nand U2534 (N_2534,N_2316,N_2192);
and U2535 (N_2535,N_2038,N_2276);
nand U2536 (N_2536,N_2369,N_2169);
nand U2537 (N_2537,N_2142,N_2390);
xnor U2538 (N_2538,N_2173,N_2001);
or U2539 (N_2539,N_2020,N_2291);
and U2540 (N_2540,N_2163,N_2294);
nor U2541 (N_2541,N_2328,N_2395);
or U2542 (N_2542,N_2168,N_2027);
or U2543 (N_2543,N_2111,N_2298);
or U2544 (N_2544,N_2204,N_2247);
xnor U2545 (N_2545,N_2340,N_2032);
or U2546 (N_2546,N_2278,N_2081);
nand U2547 (N_2547,N_2128,N_2121);
nor U2548 (N_2548,N_2214,N_2194);
and U2549 (N_2549,N_2202,N_2210);
nor U2550 (N_2550,N_2323,N_2280);
nor U2551 (N_2551,N_2244,N_2300);
nor U2552 (N_2552,N_2077,N_2237);
and U2553 (N_2553,N_2387,N_2119);
or U2554 (N_2554,N_2230,N_2357);
nand U2555 (N_2555,N_2106,N_2098);
xnor U2556 (N_2556,N_2153,N_2068);
nand U2557 (N_2557,N_2211,N_2042);
nor U2558 (N_2558,N_2180,N_2135);
or U2559 (N_2559,N_2201,N_2016);
and U2560 (N_2560,N_2249,N_2161);
and U2561 (N_2561,N_2109,N_2200);
or U2562 (N_2562,N_2154,N_2014);
xor U2563 (N_2563,N_2126,N_2375);
nand U2564 (N_2564,N_2004,N_2132);
or U2565 (N_2565,N_2223,N_2101);
nand U2566 (N_2566,N_2184,N_2088);
or U2567 (N_2567,N_2206,N_2327);
nand U2568 (N_2568,N_2166,N_2034);
or U2569 (N_2569,N_2090,N_2248);
xor U2570 (N_2570,N_2331,N_2362);
nor U2571 (N_2571,N_2391,N_2105);
or U2572 (N_2572,N_2189,N_2113);
or U2573 (N_2573,N_2002,N_2297);
nor U2574 (N_2574,N_2197,N_2029);
and U2575 (N_2575,N_2085,N_2279);
and U2576 (N_2576,N_2093,N_2376);
xor U2577 (N_2577,N_2267,N_2179);
nor U2578 (N_2578,N_2208,N_2079);
xor U2579 (N_2579,N_2382,N_2107);
or U2580 (N_2580,N_2216,N_2374);
and U2581 (N_2581,N_2256,N_2058);
and U2582 (N_2582,N_2017,N_2182);
xnor U2583 (N_2583,N_2313,N_2183);
nor U2584 (N_2584,N_2150,N_2071);
nand U2585 (N_2585,N_2037,N_2112);
and U2586 (N_2586,N_2240,N_2023);
nand U2587 (N_2587,N_2190,N_2070);
or U2588 (N_2588,N_2370,N_2311);
nand U2589 (N_2589,N_2157,N_2345);
xor U2590 (N_2590,N_2271,N_2050);
nor U2591 (N_2591,N_2287,N_2094);
nand U2592 (N_2592,N_2218,N_2212);
nand U2593 (N_2593,N_2337,N_2061);
xnor U2594 (N_2594,N_2084,N_2389);
nor U2595 (N_2595,N_2320,N_2049);
and U2596 (N_2596,N_2021,N_2196);
and U2597 (N_2597,N_2209,N_2385);
nor U2598 (N_2598,N_2067,N_2292);
nor U2599 (N_2599,N_2059,N_2255);
and U2600 (N_2600,N_2269,N_2022);
xnor U2601 (N_2601,N_2365,N_2296);
xor U2602 (N_2602,N_2321,N_2107);
or U2603 (N_2603,N_2223,N_2137);
and U2604 (N_2604,N_2289,N_2361);
and U2605 (N_2605,N_2059,N_2099);
and U2606 (N_2606,N_2093,N_2030);
and U2607 (N_2607,N_2009,N_2199);
or U2608 (N_2608,N_2129,N_2271);
xnor U2609 (N_2609,N_2069,N_2115);
or U2610 (N_2610,N_2190,N_2128);
and U2611 (N_2611,N_2070,N_2292);
xor U2612 (N_2612,N_2308,N_2126);
xor U2613 (N_2613,N_2202,N_2157);
and U2614 (N_2614,N_2319,N_2130);
and U2615 (N_2615,N_2201,N_2248);
nor U2616 (N_2616,N_2076,N_2378);
or U2617 (N_2617,N_2304,N_2116);
nand U2618 (N_2618,N_2190,N_2323);
nor U2619 (N_2619,N_2353,N_2343);
or U2620 (N_2620,N_2181,N_2376);
nor U2621 (N_2621,N_2155,N_2377);
xnor U2622 (N_2622,N_2031,N_2036);
nor U2623 (N_2623,N_2192,N_2107);
nor U2624 (N_2624,N_2144,N_2397);
or U2625 (N_2625,N_2348,N_2312);
and U2626 (N_2626,N_2395,N_2010);
nand U2627 (N_2627,N_2302,N_2255);
nor U2628 (N_2628,N_2217,N_2083);
and U2629 (N_2629,N_2299,N_2214);
and U2630 (N_2630,N_2032,N_2225);
xor U2631 (N_2631,N_2021,N_2017);
xor U2632 (N_2632,N_2127,N_2211);
xnor U2633 (N_2633,N_2185,N_2359);
or U2634 (N_2634,N_2337,N_2204);
xor U2635 (N_2635,N_2365,N_2257);
nand U2636 (N_2636,N_2002,N_2390);
or U2637 (N_2637,N_2108,N_2038);
and U2638 (N_2638,N_2214,N_2287);
and U2639 (N_2639,N_2152,N_2392);
xor U2640 (N_2640,N_2119,N_2320);
xor U2641 (N_2641,N_2006,N_2144);
and U2642 (N_2642,N_2007,N_2215);
nand U2643 (N_2643,N_2342,N_2173);
or U2644 (N_2644,N_2094,N_2306);
nand U2645 (N_2645,N_2282,N_2392);
or U2646 (N_2646,N_2370,N_2378);
or U2647 (N_2647,N_2043,N_2218);
nor U2648 (N_2648,N_2074,N_2174);
xor U2649 (N_2649,N_2392,N_2306);
nand U2650 (N_2650,N_2249,N_2100);
nand U2651 (N_2651,N_2118,N_2277);
or U2652 (N_2652,N_2082,N_2075);
nand U2653 (N_2653,N_2280,N_2143);
nor U2654 (N_2654,N_2280,N_2190);
nand U2655 (N_2655,N_2222,N_2309);
or U2656 (N_2656,N_2070,N_2178);
nand U2657 (N_2657,N_2095,N_2198);
nor U2658 (N_2658,N_2339,N_2040);
or U2659 (N_2659,N_2155,N_2301);
or U2660 (N_2660,N_2390,N_2228);
xnor U2661 (N_2661,N_2136,N_2194);
nand U2662 (N_2662,N_2283,N_2315);
or U2663 (N_2663,N_2027,N_2248);
and U2664 (N_2664,N_2281,N_2017);
xor U2665 (N_2665,N_2363,N_2188);
xor U2666 (N_2666,N_2220,N_2029);
or U2667 (N_2667,N_2182,N_2258);
nand U2668 (N_2668,N_2338,N_2032);
and U2669 (N_2669,N_2037,N_2218);
xor U2670 (N_2670,N_2259,N_2374);
nand U2671 (N_2671,N_2294,N_2149);
nor U2672 (N_2672,N_2035,N_2039);
or U2673 (N_2673,N_2134,N_2394);
nor U2674 (N_2674,N_2307,N_2359);
nand U2675 (N_2675,N_2049,N_2228);
or U2676 (N_2676,N_2115,N_2042);
nand U2677 (N_2677,N_2014,N_2144);
nor U2678 (N_2678,N_2396,N_2042);
nor U2679 (N_2679,N_2248,N_2203);
and U2680 (N_2680,N_2162,N_2123);
nand U2681 (N_2681,N_2053,N_2382);
and U2682 (N_2682,N_2324,N_2218);
and U2683 (N_2683,N_2272,N_2043);
and U2684 (N_2684,N_2277,N_2262);
or U2685 (N_2685,N_2221,N_2047);
xor U2686 (N_2686,N_2374,N_2035);
nor U2687 (N_2687,N_2061,N_2375);
and U2688 (N_2688,N_2063,N_2154);
nor U2689 (N_2689,N_2255,N_2236);
and U2690 (N_2690,N_2274,N_2285);
nand U2691 (N_2691,N_2337,N_2144);
nand U2692 (N_2692,N_2390,N_2185);
or U2693 (N_2693,N_2151,N_2258);
or U2694 (N_2694,N_2276,N_2392);
and U2695 (N_2695,N_2372,N_2123);
nand U2696 (N_2696,N_2141,N_2051);
xnor U2697 (N_2697,N_2240,N_2074);
nor U2698 (N_2698,N_2346,N_2308);
nand U2699 (N_2699,N_2055,N_2317);
nand U2700 (N_2700,N_2068,N_2099);
nand U2701 (N_2701,N_2393,N_2284);
or U2702 (N_2702,N_2228,N_2383);
and U2703 (N_2703,N_2077,N_2145);
nor U2704 (N_2704,N_2231,N_2227);
nor U2705 (N_2705,N_2284,N_2208);
or U2706 (N_2706,N_2280,N_2052);
nand U2707 (N_2707,N_2229,N_2254);
nor U2708 (N_2708,N_2206,N_2398);
and U2709 (N_2709,N_2090,N_2123);
or U2710 (N_2710,N_2229,N_2197);
nor U2711 (N_2711,N_2266,N_2272);
and U2712 (N_2712,N_2127,N_2165);
or U2713 (N_2713,N_2142,N_2048);
or U2714 (N_2714,N_2295,N_2026);
and U2715 (N_2715,N_2146,N_2189);
or U2716 (N_2716,N_2301,N_2241);
xnor U2717 (N_2717,N_2073,N_2282);
or U2718 (N_2718,N_2084,N_2200);
nor U2719 (N_2719,N_2390,N_2241);
xnor U2720 (N_2720,N_2012,N_2342);
nor U2721 (N_2721,N_2024,N_2166);
nand U2722 (N_2722,N_2097,N_2306);
and U2723 (N_2723,N_2216,N_2098);
xnor U2724 (N_2724,N_2390,N_2372);
xor U2725 (N_2725,N_2224,N_2125);
xnor U2726 (N_2726,N_2047,N_2158);
and U2727 (N_2727,N_2256,N_2368);
xor U2728 (N_2728,N_2259,N_2105);
xnor U2729 (N_2729,N_2323,N_2347);
nor U2730 (N_2730,N_2229,N_2048);
or U2731 (N_2731,N_2091,N_2258);
nor U2732 (N_2732,N_2280,N_2028);
nor U2733 (N_2733,N_2241,N_2290);
nor U2734 (N_2734,N_2287,N_2112);
and U2735 (N_2735,N_2317,N_2232);
xor U2736 (N_2736,N_2291,N_2131);
xnor U2737 (N_2737,N_2296,N_2048);
or U2738 (N_2738,N_2096,N_2231);
and U2739 (N_2739,N_2053,N_2259);
xor U2740 (N_2740,N_2157,N_2302);
and U2741 (N_2741,N_2294,N_2212);
xor U2742 (N_2742,N_2213,N_2285);
and U2743 (N_2743,N_2320,N_2193);
nor U2744 (N_2744,N_2201,N_2158);
xnor U2745 (N_2745,N_2174,N_2262);
and U2746 (N_2746,N_2168,N_2196);
or U2747 (N_2747,N_2196,N_2227);
nor U2748 (N_2748,N_2333,N_2198);
nand U2749 (N_2749,N_2235,N_2103);
nand U2750 (N_2750,N_2350,N_2020);
or U2751 (N_2751,N_2192,N_2196);
nand U2752 (N_2752,N_2233,N_2065);
nand U2753 (N_2753,N_2259,N_2395);
nand U2754 (N_2754,N_2332,N_2291);
or U2755 (N_2755,N_2301,N_2278);
and U2756 (N_2756,N_2256,N_2000);
or U2757 (N_2757,N_2241,N_2305);
xor U2758 (N_2758,N_2351,N_2262);
nand U2759 (N_2759,N_2349,N_2081);
or U2760 (N_2760,N_2169,N_2100);
nor U2761 (N_2761,N_2190,N_2024);
xor U2762 (N_2762,N_2003,N_2040);
and U2763 (N_2763,N_2042,N_2071);
and U2764 (N_2764,N_2112,N_2104);
nand U2765 (N_2765,N_2002,N_2374);
or U2766 (N_2766,N_2152,N_2191);
and U2767 (N_2767,N_2101,N_2226);
or U2768 (N_2768,N_2372,N_2180);
nand U2769 (N_2769,N_2081,N_2049);
nand U2770 (N_2770,N_2018,N_2169);
xnor U2771 (N_2771,N_2326,N_2399);
nand U2772 (N_2772,N_2232,N_2173);
xnor U2773 (N_2773,N_2292,N_2060);
xnor U2774 (N_2774,N_2359,N_2067);
nor U2775 (N_2775,N_2120,N_2002);
and U2776 (N_2776,N_2094,N_2270);
or U2777 (N_2777,N_2087,N_2303);
and U2778 (N_2778,N_2378,N_2269);
nand U2779 (N_2779,N_2383,N_2137);
or U2780 (N_2780,N_2190,N_2209);
and U2781 (N_2781,N_2284,N_2241);
xnor U2782 (N_2782,N_2009,N_2314);
nand U2783 (N_2783,N_2095,N_2206);
xor U2784 (N_2784,N_2136,N_2245);
or U2785 (N_2785,N_2130,N_2107);
nand U2786 (N_2786,N_2366,N_2069);
or U2787 (N_2787,N_2384,N_2226);
nand U2788 (N_2788,N_2173,N_2193);
nor U2789 (N_2789,N_2129,N_2226);
xor U2790 (N_2790,N_2228,N_2284);
nor U2791 (N_2791,N_2303,N_2105);
nor U2792 (N_2792,N_2322,N_2024);
nor U2793 (N_2793,N_2323,N_2265);
xnor U2794 (N_2794,N_2341,N_2188);
and U2795 (N_2795,N_2174,N_2276);
xor U2796 (N_2796,N_2237,N_2208);
nand U2797 (N_2797,N_2199,N_2261);
or U2798 (N_2798,N_2377,N_2090);
nand U2799 (N_2799,N_2071,N_2376);
nor U2800 (N_2800,N_2757,N_2700);
nor U2801 (N_2801,N_2785,N_2609);
or U2802 (N_2802,N_2545,N_2527);
or U2803 (N_2803,N_2744,N_2691);
nand U2804 (N_2804,N_2591,N_2606);
nand U2805 (N_2805,N_2650,N_2736);
xnor U2806 (N_2806,N_2665,N_2453);
nand U2807 (N_2807,N_2636,N_2509);
or U2808 (N_2808,N_2641,N_2544);
nand U2809 (N_2809,N_2402,N_2510);
nor U2810 (N_2810,N_2409,N_2783);
or U2811 (N_2811,N_2507,N_2478);
nor U2812 (N_2812,N_2603,N_2717);
nand U2813 (N_2813,N_2612,N_2531);
nor U2814 (N_2814,N_2696,N_2781);
or U2815 (N_2815,N_2726,N_2752);
nor U2816 (N_2816,N_2404,N_2455);
and U2817 (N_2817,N_2487,N_2733);
xor U2818 (N_2818,N_2737,N_2499);
or U2819 (N_2819,N_2642,N_2657);
nand U2820 (N_2820,N_2694,N_2767);
nor U2821 (N_2821,N_2745,N_2461);
and U2822 (N_2822,N_2772,N_2484);
nor U2823 (N_2823,N_2793,N_2723);
or U2824 (N_2824,N_2423,N_2714);
nand U2825 (N_2825,N_2616,N_2607);
or U2826 (N_2826,N_2648,N_2637);
xor U2827 (N_2827,N_2662,N_2787);
or U2828 (N_2828,N_2535,N_2771);
nand U2829 (N_2829,N_2646,N_2673);
xnor U2830 (N_2830,N_2672,N_2569);
xnor U2831 (N_2831,N_2774,N_2652);
nor U2832 (N_2832,N_2795,N_2654);
nand U2833 (N_2833,N_2476,N_2413);
or U2834 (N_2834,N_2460,N_2574);
xnor U2835 (N_2835,N_2469,N_2572);
xor U2836 (N_2836,N_2426,N_2488);
xnor U2837 (N_2837,N_2410,N_2422);
nand U2838 (N_2838,N_2424,N_2494);
nand U2839 (N_2839,N_2605,N_2618);
nand U2840 (N_2840,N_2418,N_2638);
xnor U2841 (N_2841,N_2437,N_2554);
nor U2842 (N_2842,N_2432,N_2506);
and U2843 (N_2843,N_2753,N_2443);
xor U2844 (N_2844,N_2524,N_2634);
nand U2845 (N_2845,N_2441,N_2713);
nand U2846 (N_2846,N_2599,N_2540);
and U2847 (N_2847,N_2762,N_2693);
and U2848 (N_2848,N_2547,N_2649);
xor U2849 (N_2849,N_2595,N_2520);
nor U2850 (N_2850,N_2445,N_2451);
xnor U2851 (N_2851,N_2407,N_2728);
xor U2852 (N_2852,N_2592,N_2589);
xnor U2853 (N_2853,N_2454,N_2565);
nand U2854 (N_2854,N_2770,N_2775);
nor U2855 (N_2855,N_2548,N_2615);
nand U2856 (N_2856,N_2617,N_2695);
nand U2857 (N_2857,N_2663,N_2585);
nor U2858 (N_2858,N_2796,N_2513);
nor U2859 (N_2859,N_2601,N_2579);
xnor U2860 (N_2860,N_2523,N_2439);
xor U2861 (N_2861,N_2556,N_2671);
or U2862 (N_2862,N_2549,N_2707);
nor U2863 (N_2863,N_2756,N_2530);
and U2864 (N_2864,N_2597,N_2558);
nand U2865 (N_2865,N_2715,N_2759);
nor U2866 (N_2866,N_2751,N_2682);
and U2867 (N_2867,N_2765,N_2708);
nor U2868 (N_2868,N_2632,N_2619);
and U2869 (N_2869,N_2496,N_2755);
nand U2870 (N_2870,N_2797,N_2647);
nor U2871 (N_2871,N_2720,N_2406);
nor U2872 (N_2872,N_2446,N_2732);
nor U2873 (N_2873,N_2420,N_2748);
nand U2874 (N_2874,N_2656,N_2552);
or U2875 (N_2875,N_2792,N_2703);
nand U2876 (N_2876,N_2760,N_2676);
nor U2877 (N_2877,N_2639,N_2709);
and U2878 (N_2878,N_2668,N_2697);
and U2879 (N_2879,N_2412,N_2522);
or U2880 (N_2880,N_2500,N_2497);
or U2881 (N_2881,N_2462,N_2746);
xnor U2882 (N_2882,N_2415,N_2456);
nor U2883 (N_2883,N_2575,N_2577);
and U2884 (N_2884,N_2790,N_2479);
or U2885 (N_2885,N_2421,N_2561);
nor U2886 (N_2886,N_2658,N_2722);
nor U2887 (N_2887,N_2623,N_2512);
nor U2888 (N_2888,N_2438,N_2735);
nand U2889 (N_2889,N_2701,N_2777);
nor U2890 (N_2890,N_2434,N_2570);
xor U2891 (N_2891,N_2433,N_2532);
nor U2892 (N_2892,N_2475,N_2564);
nand U2893 (N_2893,N_2780,N_2727);
nor U2894 (N_2894,N_2538,N_2519);
nor U2895 (N_2895,N_2786,N_2403);
and U2896 (N_2896,N_2470,N_2405);
nor U2897 (N_2897,N_2667,N_2675);
nand U2898 (N_2898,N_2425,N_2677);
and U2899 (N_2899,N_2749,N_2583);
nor U2900 (N_2900,N_2710,N_2508);
nor U2901 (N_2901,N_2416,N_2633);
nor U2902 (N_2902,N_2431,N_2679);
or U2903 (N_2903,N_2798,N_2681);
nand U2904 (N_2904,N_2562,N_2624);
xnor U2905 (N_2905,N_2491,N_2536);
nor U2906 (N_2906,N_2498,N_2480);
nand U2907 (N_2907,N_2684,N_2504);
and U2908 (N_2908,N_2690,N_2741);
nor U2909 (N_2909,N_2440,N_2743);
nand U2910 (N_2910,N_2419,N_2576);
xnor U2911 (N_2911,N_2686,N_2529);
nand U2912 (N_2912,N_2429,N_2689);
nor U2913 (N_2913,N_2644,N_2502);
nor U2914 (N_2914,N_2742,N_2468);
or U2915 (N_2915,N_2541,N_2435);
xnor U2916 (N_2916,N_2467,N_2534);
or U2917 (N_2917,N_2430,N_2769);
or U2918 (N_2918,N_2457,N_2761);
or U2919 (N_2919,N_2621,N_2794);
or U2920 (N_2920,N_2763,N_2610);
and U2921 (N_2921,N_2789,N_2537);
nor U2922 (N_2922,N_2640,N_2555);
and U2923 (N_2923,N_2493,N_2628);
nor U2924 (N_2924,N_2501,N_2627);
or U2925 (N_2925,N_2518,N_2517);
nor U2926 (N_2926,N_2593,N_2739);
or U2927 (N_2927,N_2613,N_2731);
xor U2928 (N_2928,N_2670,N_2661);
xor U2929 (N_2929,N_2566,N_2542);
nand U2930 (N_2930,N_2719,N_2669);
nand U2931 (N_2931,N_2614,N_2442);
and U2932 (N_2932,N_2481,N_2448);
xor U2933 (N_2933,N_2573,N_2688);
nor U2934 (N_2934,N_2474,N_2768);
or U2935 (N_2935,N_2465,N_2622);
xor U2936 (N_2936,N_2754,N_2674);
nor U2937 (N_2937,N_2718,N_2666);
or U2938 (N_2938,N_2635,N_2706);
xnor U2939 (N_2939,N_2704,N_2651);
xor U2940 (N_2940,N_2417,N_2664);
and U2941 (N_2941,N_2596,N_2740);
nand U2942 (N_2942,N_2702,N_2764);
nor U2943 (N_2943,N_2631,N_2546);
nor U2944 (N_2944,N_2590,N_2567);
nand U2945 (N_2945,N_2581,N_2678);
nand U2946 (N_2946,N_2643,N_2539);
nand U2947 (N_2947,N_2444,N_2505);
nor U2948 (N_2948,N_2550,N_2463);
or U2949 (N_2949,N_2543,N_2692);
nand U2950 (N_2950,N_2588,N_2799);
xor U2951 (N_2951,N_2471,N_2452);
xor U2952 (N_2952,N_2721,N_2528);
nor U2953 (N_2953,N_2630,N_2482);
and U2954 (N_2954,N_2584,N_2629);
xnor U2955 (N_2955,N_2660,N_2604);
nor U2956 (N_2956,N_2586,N_2791);
and U2957 (N_2957,N_2514,N_2483);
and U2958 (N_2958,N_2408,N_2533);
xor U2959 (N_2959,N_2750,N_2489);
or U2960 (N_2960,N_2427,N_2473);
xor U2961 (N_2961,N_2492,N_2459);
nand U2962 (N_2962,N_2428,N_2788);
or U2963 (N_2963,N_2458,N_2611);
or U2964 (N_2964,N_2776,N_2699);
or U2965 (N_2965,N_2450,N_2626);
nand U2966 (N_2966,N_2725,N_2698);
or U2967 (N_2967,N_2466,N_2683);
and U2968 (N_2968,N_2784,N_2773);
or U2969 (N_2969,N_2414,N_2568);
xnor U2970 (N_2970,N_2521,N_2724);
nor U2971 (N_2971,N_2511,N_2563);
or U2972 (N_2972,N_2447,N_2782);
nor U2973 (N_2973,N_2559,N_2464);
and U2974 (N_2974,N_2716,N_2582);
or U2975 (N_2975,N_2645,N_2600);
and U2976 (N_2976,N_2553,N_2400);
or U2977 (N_2977,N_2490,N_2516);
nand U2978 (N_2978,N_2779,N_2778);
nor U2979 (N_2979,N_2594,N_2578);
nand U2980 (N_2980,N_2449,N_2436);
and U2981 (N_2981,N_2486,N_2598);
nand U2982 (N_2982,N_2477,N_2734);
or U2983 (N_2983,N_2525,N_2602);
nor U2984 (N_2984,N_2625,N_2608);
and U2985 (N_2985,N_2503,N_2655);
or U2986 (N_2986,N_2712,N_2738);
nor U2987 (N_2987,N_2687,N_2747);
or U2988 (N_2988,N_2758,N_2711);
or U2989 (N_2989,N_2659,N_2560);
and U2990 (N_2990,N_2766,N_2401);
or U2991 (N_2991,N_2653,N_2680);
and U2992 (N_2992,N_2485,N_2620);
or U2993 (N_2993,N_2705,N_2580);
xnor U2994 (N_2994,N_2526,N_2557);
nand U2995 (N_2995,N_2730,N_2472);
or U2996 (N_2996,N_2495,N_2551);
or U2997 (N_2997,N_2587,N_2685);
and U2998 (N_2998,N_2515,N_2729);
or U2999 (N_2999,N_2571,N_2411);
and U3000 (N_3000,N_2527,N_2479);
nor U3001 (N_3001,N_2575,N_2616);
nand U3002 (N_3002,N_2787,N_2420);
nor U3003 (N_3003,N_2744,N_2473);
and U3004 (N_3004,N_2716,N_2644);
nand U3005 (N_3005,N_2418,N_2503);
nand U3006 (N_3006,N_2771,N_2498);
or U3007 (N_3007,N_2633,N_2407);
nor U3008 (N_3008,N_2640,N_2546);
and U3009 (N_3009,N_2439,N_2690);
or U3010 (N_3010,N_2434,N_2614);
nor U3011 (N_3011,N_2505,N_2782);
xor U3012 (N_3012,N_2416,N_2598);
nand U3013 (N_3013,N_2599,N_2419);
and U3014 (N_3014,N_2539,N_2680);
xor U3015 (N_3015,N_2798,N_2742);
and U3016 (N_3016,N_2502,N_2774);
nor U3017 (N_3017,N_2658,N_2529);
nand U3018 (N_3018,N_2594,N_2552);
nor U3019 (N_3019,N_2572,N_2492);
xor U3020 (N_3020,N_2464,N_2502);
xnor U3021 (N_3021,N_2585,N_2522);
nor U3022 (N_3022,N_2789,N_2601);
nor U3023 (N_3023,N_2466,N_2611);
nand U3024 (N_3024,N_2793,N_2697);
xnor U3025 (N_3025,N_2632,N_2652);
and U3026 (N_3026,N_2445,N_2465);
or U3027 (N_3027,N_2597,N_2478);
or U3028 (N_3028,N_2508,N_2446);
nand U3029 (N_3029,N_2547,N_2533);
and U3030 (N_3030,N_2597,N_2555);
nor U3031 (N_3031,N_2670,N_2691);
nand U3032 (N_3032,N_2484,N_2795);
nand U3033 (N_3033,N_2696,N_2627);
xnor U3034 (N_3034,N_2708,N_2545);
nand U3035 (N_3035,N_2432,N_2533);
and U3036 (N_3036,N_2430,N_2774);
and U3037 (N_3037,N_2473,N_2785);
or U3038 (N_3038,N_2584,N_2527);
xor U3039 (N_3039,N_2702,N_2537);
nand U3040 (N_3040,N_2509,N_2557);
and U3041 (N_3041,N_2649,N_2530);
and U3042 (N_3042,N_2489,N_2664);
or U3043 (N_3043,N_2419,N_2615);
and U3044 (N_3044,N_2442,N_2511);
and U3045 (N_3045,N_2502,N_2675);
nor U3046 (N_3046,N_2555,N_2425);
nand U3047 (N_3047,N_2532,N_2651);
nor U3048 (N_3048,N_2693,N_2704);
nor U3049 (N_3049,N_2504,N_2716);
or U3050 (N_3050,N_2431,N_2493);
nand U3051 (N_3051,N_2769,N_2713);
nor U3052 (N_3052,N_2785,N_2565);
nand U3053 (N_3053,N_2505,N_2578);
xor U3054 (N_3054,N_2502,N_2522);
xor U3055 (N_3055,N_2710,N_2509);
xor U3056 (N_3056,N_2662,N_2763);
and U3057 (N_3057,N_2682,N_2433);
nor U3058 (N_3058,N_2592,N_2665);
xnor U3059 (N_3059,N_2442,N_2741);
and U3060 (N_3060,N_2724,N_2494);
nand U3061 (N_3061,N_2795,N_2611);
xor U3062 (N_3062,N_2585,N_2691);
and U3063 (N_3063,N_2798,N_2545);
and U3064 (N_3064,N_2433,N_2513);
xor U3065 (N_3065,N_2508,N_2494);
and U3066 (N_3066,N_2750,N_2581);
or U3067 (N_3067,N_2739,N_2531);
nand U3068 (N_3068,N_2632,N_2535);
nor U3069 (N_3069,N_2402,N_2453);
xnor U3070 (N_3070,N_2728,N_2627);
xor U3071 (N_3071,N_2420,N_2513);
or U3072 (N_3072,N_2773,N_2663);
nand U3073 (N_3073,N_2434,N_2727);
nor U3074 (N_3074,N_2498,N_2534);
or U3075 (N_3075,N_2674,N_2481);
nor U3076 (N_3076,N_2775,N_2794);
and U3077 (N_3077,N_2788,N_2725);
and U3078 (N_3078,N_2587,N_2693);
and U3079 (N_3079,N_2577,N_2533);
or U3080 (N_3080,N_2696,N_2788);
and U3081 (N_3081,N_2572,N_2459);
nor U3082 (N_3082,N_2589,N_2778);
nand U3083 (N_3083,N_2648,N_2551);
xnor U3084 (N_3084,N_2772,N_2617);
nand U3085 (N_3085,N_2760,N_2424);
xnor U3086 (N_3086,N_2734,N_2576);
or U3087 (N_3087,N_2659,N_2678);
xnor U3088 (N_3088,N_2564,N_2620);
and U3089 (N_3089,N_2713,N_2538);
or U3090 (N_3090,N_2428,N_2752);
and U3091 (N_3091,N_2519,N_2441);
and U3092 (N_3092,N_2576,N_2501);
xor U3093 (N_3093,N_2645,N_2647);
and U3094 (N_3094,N_2713,N_2744);
nor U3095 (N_3095,N_2505,N_2455);
nand U3096 (N_3096,N_2737,N_2665);
xnor U3097 (N_3097,N_2487,N_2581);
nor U3098 (N_3098,N_2434,N_2553);
or U3099 (N_3099,N_2544,N_2767);
nor U3100 (N_3100,N_2720,N_2757);
xor U3101 (N_3101,N_2484,N_2591);
xnor U3102 (N_3102,N_2591,N_2410);
xnor U3103 (N_3103,N_2744,N_2757);
xor U3104 (N_3104,N_2482,N_2747);
xor U3105 (N_3105,N_2714,N_2420);
and U3106 (N_3106,N_2559,N_2521);
or U3107 (N_3107,N_2710,N_2486);
nor U3108 (N_3108,N_2797,N_2688);
nor U3109 (N_3109,N_2604,N_2401);
nand U3110 (N_3110,N_2572,N_2540);
or U3111 (N_3111,N_2620,N_2407);
nor U3112 (N_3112,N_2650,N_2457);
nor U3113 (N_3113,N_2451,N_2488);
nor U3114 (N_3114,N_2642,N_2507);
nor U3115 (N_3115,N_2558,N_2724);
or U3116 (N_3116,N_2486,N_2498);
and U3117 (N_3117,N_2683,N_2555);
and U3118 (N_3118,N_2762,N_2514);
xnor U3119 (N_3119,N_2684,N_2445);
or U3120 (N_3120,N_2469,N_2520);
xnor U3121 (N_3121,N_2411,N_2738);
xnor U3122 (N_3122,N_2773,N_2465);
nand U3123 (N_3123,N_2674,N_2505);
nand U3124 (N_3124,N_2457,N_2690);
nor U3125 (N_3125,N_2543,N_2542);
and U3126 (N_3126,N_2488,N_2409);
nand U3127 (N_3127,N_2666,N_2590);
nor U3128 (N_3128,N_2764,N_2745);
or U3129 (N_3129,N_2602,N_2642);
nor U3130 (N_3130,N_2518,N_2669);
nand U3131 (N_3131,N_2605,N_2462);
nor U3132 (N_3132,N_2554,N_2771);
xor U3133 (N_3133,N_2409,N_2758);
nor U3134 (N_3134,N_2452,N_2477);
nor U3135 (N_3135,N_2426,N_2677);
or U3136 (N_3136,N_2445,N_2592);
xnor U3137 (N_3137,N_2556,N_2574);
or U3138 (N_3138,N_2712,N_2676);
nand U3139 (N_3139,N_2767,N_2738);
nor U3140 (N_3140,N_2780,N_2496);
and U3141 (N_3141,N_2528,N_2542);
xor U3142 (N_3142,N_2587,N_2522);
nor U3143 (N_3143,N_2555,N_2614);
nand U3144 (N_3144,N_2547,N_2458);
nand U3145 (N_3145,N_2587,N_2411);
or U3146 (N_3146,N_2498,N_2616);
and U3147 (N_3147,N_2430,N_2770);
or U3148 (N_3148,N_2438,N_2451);
nor U3149 (N_3149,N_2418,N_2590);
nor U3150 (N_3150,N_2610,N_2703);
and U3151 (N_3151,N_2497,N_2452);
or U3152 (N_3152,N_2460,N_2599);
and U3153 (N_3153,N_2664,N_2476);
nor U3154 (N_3154,N_2787,N_2687);
nor U3155 (N_3155,N_2457,N_2536);
and U3156 (N_3156,N_2559,N_2788);
or U3157 (N_3157,N_2461,N_2798);
and U3158 (N_3158,N_2541,N_2518);
nand U3159 (N_3159,N_2466,N_2437);
nor U3160 (N_3160,N_2566,N_2649);
or U3161 (N_3161,N_2635,N_2451);
nor U3162 (N_3162,N_2719,N_2695);
or U3163 (N_3163,N_2759,N_2457);
nand U3164 (N_3164,N_2413,N_2710);
or U3165 (N_3165,N_2572,N_2703);
nor U3166 (N_3166,N_2443,N_2580);
nand U3167 (N_3167,N_2668,N_2792);
and U3168 (N_3168,N_2591,N_2453);
or U3169 (N_3169,N_2409,N_2764);
xnor U3170 (N_3170,N_2761,N_2466);
xor U3171 (N_3171,N_2653,N_2478);
xnor U3172 (N_3172,N_2548,N_2464);
or U3173 (N_3173,N_2464,N_2698);
nand U3174 (N_3174,N_2756,N_2402);
nand U3175 (N_3175,N_2652,N_2647);
or U3176 (N_3176,N_2573,N_2402);
or U3177 (N_3177,N_2788,N_2570);
nor U3178 (N_3178,N_2744,N_2614);
or U3179 (N_3179,N_2735,N_2662);
and U3180 (N_3180,N_2561,N_2570);
and U3181 (N_3181,N_2507,N_2623);
nand U3182 (N_3182,N_2603,N_2598);
and U3183 (N_3183,N_2601,N_2722);
and U3184 (N_3184,N_2663,N_2544);
nand U3185 (N_3185,N_2484,N_2642);
xor U3186 (N_3186,N_2692,N_2615);
xnor U3187 (N_3187,N_2468,N_2587);
or U3188 (N_3188,N_2791,N_2579);
xor U3189 (N_3189,N_2797,N_2757);
or U3190 (N_3190,N_2743,N_2477);
nor U3191 (N_3191,N_2768,N_2644);
or U3192 (N_3192,N_2506,N_2773);
nor U3193 (N_3193,N_2728,N_2641);
xnor U3194 (N_3194,N_2592,N_2410);
nor U3195 (N_3195,N_2748,N_2768);
and U3196 (N_3196,N_2771,N_2780);
and U3197 (N_3197,N_2656,N_2795);
xnor U3198 (N_3198,N_2700,N_2734);
nor U3199 (N_3199,N_2664,N_2650);
nand U3200 (N_3200,N_2886,N_2821);
nor U3201 (N_3201,N_2825,N_2954);
nor U3202 (N_3202,N_3110,N_3162);
nor U3203 (N_3203,N_3126,N_2911);
and U3204 (N_3204,N_3112,N_3111);
xnor U3205 (N_3205,N_3180,N_3093);
xnor U3206 (N_3206,N_2939,N_2870);
and U3207 (N_3207,N_3077,N_3047);
nand U3208 (N_3208,N_3082,N_3148);
xnor U3209 (N_3209,N_3069,N_2916);
or U3210 (N_3210,N_3024,N_3163);
xor U3211 (N_3211,N_2882,N_3030);
and U3212 (N_3212,N_3000,N_2927);
or U3213 (N_3213,N_3193,N_3164);
xor U3214 (N_3214,N_2854,N_2915);
xnor U3215 (N_3215,N_2867,N_3139);
and U3216 (N_3216,N_3054,N_2896);
xnor U3217 (N_3217,N_3006,N_2853);
and U3218 (N_3218,N_3130,N_3044);
or U3219 (N_3219,N_3088,N_3142);
xnor U3220 (N_3220,N_3096,N_3166);
or U3221 (N_3221,N_2901,N_3125);
or U3222 (N_3222,N_3115,N_3050);
or U3223 (N_3223,N_3182,N_3133);
xnor U3224 (N_3224,N_2843,N_3091);
and U3225 (N_3225,N_2914,N_3178);
nor U3226 (N_3226,N_2937,N_3056);
nand U3227 (N_3227,N_2877,N_2941);
nor U3228 (N_3228,N_3197,N_3099);
nand U3229 (N_3229,N_3195,N_3022);
xor U3230 (N_3230,N_2864,N_3052);
or U3231 (N_3231,N_2981,N_3114);
or U3232 (N_3232,N_2899,N_3158);
nor U3233 (N_3233,N_2942,N_3068);
nor U3234 (N_3234,N_2921,N_2863);
xnor U3235 (N_3235,N_2988,N_3107);
nand U3236 (N_3236,N_3003,N_2999);
xnor U3237 (N_3237,N_3059,N_3010);
nand U3238 (N_3238,N_3023,N_3161);
or U3239 (N_3239,N_2883,N_3071);
nor U3240 (N_3240,N_2986,N_3150);
nand U3241 (N_3241,N_3080,N_2802);
nor U3242 (N_3242,N_3081,N_3159);
nand U3243 (N_3243,N_3025,N_3045);
nand U3244 (N_3244,N_2991,N_2875);
nor U3245 (N_3245,N_2844,N_2969);
and U3246 (N_3246,N_3097,N_2989);
or U3247 (N_3247,N_2816,N_3145);
and U3248 (N_3248,N_2990,N_2971);
nor U3249 (N_3249,N_2866,N_3013);
and U3250 (N_3250,N_3042,N_2881);
nor U3251 (N_3251,N_3028,N_2823);
nor U3252 (N_3252,N_2849,N_2900);
xnor U3253 (N_3253,N_3043,N_2931);
nor U3254 (N_3254,N_3029,N_3084);
nor U3255 (N_3255,N_3173,N_3175);
xnor U3256 (N_3256,N_2905,N_2839);
xnor U3257 (N_3257,N_2818,N_3035);
or U3258 (N_3258,N_3119,N_2869);
xor U3259 (N_3259,N_2885,N_2830);
and U3260 (N_3260,N_2834,N_3194);
and U3261 (N_3261,N_2878,N_2835);
nand U3262 (N_3262,N_3061,N_3017);
and U3263 (N_3263,N_3118,N_2890);
nor U3264 (N_3264,N_3086,N_2889);
nand U3265 (N_3265,N_3021,N_2928);
or U3266 (N_3266,N_3137,N_3168);
and U3267 (N_3267,N_2959,N_3147);
nor U3268 (N_3268,N_2871,N_3078);
nand U3269 (N_3269,N_3015,N_2933);
and U3270 (N_3270,N_3105,N_2857);
xnor U3271 (N_3271,N_3062,N_2925);
or U3272 (N_3272,N_2862,N_3102);
xnor U3273 (N_3273,N_3160,N_3184);
nor U3274 (N_3274,N_2902,N_3032);
and U3275 (N_3275,N_2836,N_2848);
or U3276 (N_3276,N_3026,N_3014);
nand U3277 (N_3277,N_2811,N_3120);
and U3278 (N_3278,N_3129,N_3034);
or U3279 (N_3279,N_3089,N_2842);
and U3280 (N_3280,N_3183,N_3064);
nand U3281 (N_3281,N_3122,N_2956);
nand U3282 (N_3282,N_2958,N_2934);
nor U3283 (N_3283,N_2963,N_2919);
or U3284 (N_3284,N_3055,N_2822);
and U3285 (N_3285,N_2968,N_2910);
nand U3286 (N_3286,N_3087,N_2838);
nand U3287 (N_3287,N_2984,N_2957);
nand U3288 (N_3288,N_3036,N_3116);
xnor U3289 (N_3289,N_2949,N_2967);
or U3290 (N_3290,N_2922,N_2812);
and U3291 (N_3291,N_3192,N_2966);
xnor U3292 (N_3292,N_3132,N_3004);
xnor U3293 (N_3293,N_3090,N_3037);
or U3294 (N_3294,N_3038,N_2920);
nand U3295 (N_3295,N_3057,N_3020);
xnor U3296 (N_3296,N_2962,N_3108);
and U3297 (N_3297,N_3127,N_3196);
nand U3298 (N_3298,N_2846,N_2831);
and U3299 (N_3299,N_2840,N_2868);
nand U3300 (N_3300,N_2985,N_2918);
or U3301 (N_3301,N_3002,N_3103);
xnor U3302 (N_3302,N_2917,N_2852);
or U3303 (N_3303,N_2826,N_3049);
nor U3304 (N_3304,N_2800,N_3155);
xor U3305 (N_3305,N_3058,N_2924);
xor U3306 (N_3306,N_2809,N_3012);
and U3307 (N_3307,N_2953,N_2837);
and U3308 (N_3308,N_3066,N_3135);
and U3309 (N_3309,N_3011,N_3131);
or U3310 (N_3310,N_2833,N_3151);
nor U3311 (N_3311,N_3016,N_2887);
or U3312 (N_3312,N_2913,N_2879);
xnor U3313 (N_3313,N_2932,N_2992);
or U3314 (N_3314,N_2940,N_2912);
and U3315 (N_3315,N_3157,N_3141);
nor U3316 (N_3316,N_3094,N_2964);
or U3317 (N_3317,N_3001,N_3005);
nor U3318 (N_3318,N_3072,N_2943);
and U3319 (N_3319,N_2814,N_2944);
and U3320 (N_3320,N_3019,N_3191);
nand U3321 (N_3321,N_3143,N_3138);
nor U3322 (N_3322,N_3031,N_2893);
nand U3323 (N_3323,N_3154,N_2998);
nor U3324 (N_3324,N_2960,N_2952);
nor U3325 (N_3325,N_3156,N_2865);
or U3326 (N_3326,N_3189,N_3146);
nor U3327 (N_3327,N_2850,N_2996);
nor U3328 (N_3328,N_3124,N_2815);
nand U3329 (N_3329,N_2858,N_3121);
or U3330 (N_3330,N_3177,N_3092);
nor U3331 (N_3331,N_3046,N_3172);
nand U3332 (N_3332,N_2945,N_3188);
and U3333 (N_3333,N_3152,N_2993);
xnor U3334 (N_3334,N_2923,N_2965);
xnor U3335 (N_3335,N_2892,N_2955);
nand U3336 (N_3336,N_3169,N_2978);
nor U3337 (N_3337,N_2947,N_3104);
nor U3338 (N_3338,N_2860,N_2841);
or U3339 (N_3339,N_2820,N_2894);
nor U3340 (N_3340,N_2813,N_3170);
xor U3341 (N_3341,N_3140,N_2855);
and U3342 (N_3342,N_3100,N_2895);
and U3343 (N_3343,N_2851,N_2926);
xor U3344 (N_3344,N_2977,N_3040);
nand U3345 (N_3345,N_3187,N_3176);
or U3346 (N_3346,N_3174,N_2946);
nor U3347 (N_3347,N_2979,N_2805);
xnor U3348 (N_3348,N_3070,N_2983);
nor U3349 (N_3349,N_3181,N_3167);
nor U3350 (N_3350,N_2801,N_2819);
xnor U3351 (N_3351,N_2859,N_2907);
and U3352 (N_3352,N_3113,N_3185);
and U3353 (N_3353,N_2874,N_3153);
nand U3354 (N_3354,N_2806,N_3079);
or U3355 (N_3355,N_2829,N_3098);
and U3356 (N_3356,N_2982,N_3039);
xor U3357 (N_3357,N_2884,N_3033);
xor U3358 (N_3358,N_2880,N_3123);
xor U3359 (N_3359,N_2891,N_2972);
nand U3360 (N_3360,N_2873,N_3027);
nand U3361 (N_3361,N_2807,N_3149);
or U3362 (N_3362,N_2961,N_3041);
xnor U3363 (N_3363,N_2995,N_2929);
nand U3364 (N_3364,N_2903,N_3179);
xor U3365 (N_3365,N_2994,N_2935);
nor U3366 (N_3366,N_3109,N_2948);
or U3367 (N_3367,N_2804,N_3073);
or U3368 (N_3368,N_3075,N_3009);
nor U3369 (N_3369,N_3165,N_2817);
xor U3370 (N_3370,N_2904,N_2832);
and U3371 (N_3371,N_3065,N_3074);
xnor U3372 (N_3372,N_3083,N_2888);
and U3373 (N_3373,N_3067,N_2906);
or U3374 (N_3374,N_3053,N_2810);
and U3375 (N_3375,N_2973,N_3117);
and U3376 (N_3376,N_2980,N_3101);
or U3377 (N_3377,N_2936,N_3051);
xnor U3378 (N_3378,N_2975,N_2897);
or U3379 (N_3379,N_3095,N_3076);
and U3380 (N_3380,N_2847,N_2970);
and U3381 (N_3381,N_2930,N_3048);
and U3382 (N_3382,N_2803,N_3007);
and U3383 (N_3383,N_3018,N_2987);
and U3384 (N_3384,N_3063,N_2974);
nand U3385 (N_3385,N_3008,N_2824);
xnor U3386 (N_3386,N_2950,N_3144);
nand U3387 (N_3387,N_2872,N_2908);
or U3388 (N_3388,N_2976,N_2845);
nor U3389 (N_3389,N_3136,N_3128);
or U3390 (N_3390,N_3085,N_2808);
nand U3391 (N_3391,N_2827,N_2898);
xnor U3392 (N_3392,N_2951,N_2876);
xnor U3393 (N_3393,N_3186,N_2938);
or U3394 (N_3394,N_2828,N_3171);
xor U3395 (N_3395,N_2856,N_3199);
nor U3396 (N_3396,N_3106,N_3198);
nor U3397 (N_3397,N_3134,N_3190);
and U3398 (N_3398,N_2861,N_3060);
and U3399 (N_3399,N_2909,N_2997);
and U3400 (N_3400,N_2999,N_3079);
or U3401 (N_3401,N_2862,N_3005);
xor U3402 (N_3402,N_3116,N_2830);
nand U3403 (N_3403,N_2990,N_3039);
nor U3404 (N_3404,N_3090,N_3153);
or U3405 (N_3405,N_2901,N_2842);
xor U3406 (N_3406,N_3172,N_2831);
and U3407 (N_3407,N_2960,N_3167);
or U3408 (N_3408,N_3150,N_2828);
nor U3409 (N_3409,N_3175,N_2849);
or U3410 (N_3410,N_2844,N_3166);
xnor U3411 (N_3411,N_3096,N_3095);
and U3412 (N_3412,N_3182,N_3157);
xnor U3413 (N_3413,N_3145,N_3064);
nor U3414 (N_3414,N_3148,N_3004);
nor U3415 (N_3415,N_2924,N_2817);
and U3416 (N_3416,N_2987,N_3054);
nor U3417 (N_3417,N_2943,N_2846);
nand U3418 (N_3418,N_3175,N_3149);
and U3419 (N_3419,N_3074,N_2856);
or U3420 (N_3420,N_2823,N_2812);
and U3421 (N_3421,N_2877,N_3110);
or U3422 (N_3422,N_3051,N_3108);
nor U3423 (N_3423,N_3059,N_3008);
nand U3424 (N_3424,N_3163,N_2971);
nand U3425 (N_3425,N_2933,N_2911);
nand U3426 (N_3426,N_2974,N_3124);
and U3427 (N_3427,N_2817,N_3167);
nor U3428 (N_3428,N_2857,N_2939);
or U3429 (N_3429,N_3159,N_3127);
nor U3430 (N_3430,N_2876,N_3155);
and U3431 (N_3431,N_2857,N_2931);
xnor U3432 (N_3432,N_3098,N_2927);
nor U3433 (N_3433,N_2867,N_3050);
nand U3434 (N_3434,N_2940,N_3108);
xnor U3435 (N_3435,N_3110,N_3181);
nand U3436 (N_3436,N_2913,N_2974);
and U3437 (N_3437,N_2874,N_2872);
and U3438 (N_3438,N_2921,N_3059);
and U3439 (N_3439,N_2984,N_2838);
nand U3440 (N_3440,N_3086,N_3141);
nor U3441 (N_3441,N_2928,N_2920);
nor U3442 (N_3442,N_3002,N_3045);
xor U3443 (N_3443,N_2823,N_2908);
and U3444 (N_3444,N_2879,N_3156);
xor U3445 (N_3445,N_2916,N_2859);
nand U3446 (N_3446,N_3123,N_3093);
or U3447 (N_3447,N_3167,N_3074);
or U3448 (N_3448,N_3145,N_2956);
and U3449 (N_3449,N_3135,N_2924);
xor U3450 (N_3450,N_2903,N_2943);
xor U3451 (N_3451,N_3020,N_3114);
and U3452 (N_3452,N_2859,N_3151);
nand U3453 (N_3453,N_3134,N_2967);
xor U3454 (N_3454,N_3134,N_3125);
and U3455 (N_3455,N_3016,N_2968);
and U3456 (N_3456,N_3046,N_2883);
nor U3457 (N_3457,N_3128,N_2840);
nand U3458 (N_3458,N_3072,N_2815);
nand U3459 (N_3459,N_2954,N_2927);
nor U3460 (N_3460,N_3007,N_2987);
nor U3461 (N_3461,N_2892,N_2824);
nand U3462 (N_3462,N_3187,N_3140);
nor U3463 (N_3463,N_2984,N_2908);
or U3464 (N_3464,N_2944,N_2938);
nor U3465 (N_3465,N_3076,N_2812);
nor U3466 (N_3466,N_2916,N_2971);
and U3467 (N_3467,N_3113,N_2855);
nor U3468 (N_3468,N_3006,N_2968);
or U3469 (N_3469,N_3113,N_2867);
nor U3470 (N_3470,N_2875,N_3171);
and U3471 (N_3471,N_3092,N_3138);
and U3472 (N_3472,N_2818,N_2960);
nor U3473 (N_3473,N_3145,N_2913);
xor U3474 (N_3474,N_2933,N_2900);
nand U3475 (N_3475,N_2832,N_3126);
or U3476 (N_3476,N_2833,N_3013);
xnor U3477 (N_3477,N_2860,N_2856);
and U3478 (N_3478,N_3091,N_2920);
and U3479 (N_3479,N_3079,N_3020);
nand U3480 (N_3480,N_3178,N_2818);
nand U3481 (N_3481,N_3119,N_3025);
nor U3482 (N_3482,N_3004,N_2913);
or U3483 (N_3483,N_2821,N_2977);
and U3484 (N_3484,N_3122,N_3115);
xor U3485 (N_3485,N_2963,N_2923);
or U3486 (N_3486,N_3199,N_3120);
nand U3487 (N_3487,N_3030,N_2881);
xor U3488 (N_3488,N_2814,N_3199);
or U3489 (N_3489,N_2987,N_2898);
nor U3490 (N_3490,N_2982,N_2817);
xnor U3491 (N_3491,N_3019,N_2823);
nor U3492 (N_3492,N_2984,N_3196);
nand U3493 (N_3493,N_3124,N_2912);
xor U3494 (N_3494,N_2947,N_3059);
and U3495 (N_3495,N_3092,N_2894);
and U3496 (N_3496,N_2830,N_2806);
nor U3497 (N_3497,N_3110,N_2966);
or U3498 (N_3498,N_2839,N_3141);
and U3499 (N_3499,N_3135,N_3197);
or U3500 (N_3500,N_2948,N_2807);
xnor U3501 (N_3501,N_3189,N_2971);
or U3502 (N_3502,N_2978,N_3045);
or U3503 (N_3503,N_3108,N_2803);
nor U3504 (N_3504,N_3033,N_2983);
nand U3505 (N_3505,N_2812,N_3153);
nand U3506 (N_3506,N_3101,N_2831);
xor U3507 (N_3507,N_2957,N_2905);
nand U3508 (N_3508,N_2825,N_3149);
xor U3509 (N_3509,N_2868,N_2864);
xnor U3510 (N_3510,N_3159,N_3111);
xor U3511 (N_3511,N_3038,N_3095);
xnor U3512 (N_3512,N_2854,N_2931);
and U3513 (N_3513,N_3032,N_2876);
nand U3514 (N_3514,N_2920,N_3072);
or U3515 (N_3515,N_2800,N_3128);
xnor U3516 (N_3516,N_2822,N_2900);
nand U3517 (N_3517,N_2837,N_3008);
xor U3518 (N_3518,N_3014,N_3078);
nor U3519 (N_3519,N_3181,N_2874);
or U3520 (N_3520,N_2841,N_2984);
nor U3521 (N_3521,N_3098,N_2805);
nand U3522 (N_3522,N_2866,N_3090);
xor U3523 (N_3523,N_2908,N_2892);
nor U3524 (N_3524,N_2927,N_3115);
xnor U3525 (N_3525,N_2816,N_2913);
xor U3526 (N_3526,N_3106,N_3108);
and U3527 (N_3527,N_2984,N_2948);
or U3528 (N_3528,N_3087,N_2819);
nand U3529 (N_3529,N_2879,N_2956);
nand U3530 (N_3530,N_2950,N_3055);
or U3531 (N_3531,N_2909,N_3165);
or U3532 (N_3532,N_2827,N_3111);
nor U3533 (N_3533,N_2897,N_2874);
xor U3534 (N_3534,N_2934,N_3156);
nor U3535 (N_3535,N_3083,N_3159);
xnor U3536 (N_3536,N_2965,N_2831);
nor U3537 (N_3537,N_2994,N_2888);
and U3538 (N_3538,N_2979,N_2987);
nor U3539 (N_3539,N_3017,N_3137);
nor U3540 (N_3540,N_3184,N_2833);
or U3541 (N_3541,N_3118,N_3126);
xor U3542 (N_3542,N_3112,N_3128);
xor U3543 (N_3543,N_2951,N_2954);
and U3544 (N_3544,N_2956,N_2892);
or U3545 (N_3545,N_2802,N_3075);
nand U3546 (N_3546,N_2980,N_2823);
xor U3547 (N_3547,N_3020,N_2885);
and U3548 (N_3548,N_3020,N_2969);
nor U3549 (N_3549,N_2976,N_3089);
nor U3550 (N_3550,N_2889,N_3056);
or U3551 (N_3551,N_3066,N_3147);
nand U3552 (N_3552,N_3106,N_2973);
nor U3553 (N_3553,N_3109,N_2978);
nand U3554 (N_3554,N_2825,N_3186);
nand U3555 (N_3555,N_3114,N_2956);
nor U3556 (N_3556,N_2857,N_3067);
nor U3557 (N_3557,N_2806,N_3184);
or U3558 (N_3558,N_3071,N_2937);
nor U3559 (N_3559,N_3102,N_2941);
nor U3560 (N_3560,N_2861,N_2930);
and U3561 (N_3561,N_3100,N_2874);
xnor U3562 (N_3562,N_3175,N_3065);
and U3563 (N_3563,N_2927,N_2935);
nor U3564 (N_3564,N_3016,N_3184);
nor U3565 (N_3565,N_2939,N_3018);
and U3566 (N_3566,N_3196,N_3071);
or U3567 (N_3567,N_3156,N_3049);
or U3568 (N_3568,N_2904,N_3150);
xor U3569 (N_3569,N_3176,N_2843);
xor U3570 (N_3570,N_2820,N_2922);
and U3571 (N_3571,N_2884,N_3198);
nor U3572 (N_3572,N_3164,N_2843);
and U3573 (N_3573,N_2809,N_3169);
nand U3574 (N_3574,N_2837,N_3187);
and U3575 (N_3575,N_2991,N_2977);
nor U3576 (N_3576,N_3107,N_3095);
nor U3577 (N_3577,N_2856,N_3058);
nor U3578 (N_3578,N_2836,N_2841);
and U3579 (N_3579,N_2969,N_3013);
nand U3580 (N_3580,N_3073,N_3184);
nand U3581 (N_3581,N_2841,N_3124);
nor U3582 (N_3582,N_2968,N_2849);
nand U3583 (N_3583,N_3192,N_3090);
xor U3584 (N_3584,N_3032,N_3177);
nor U3585 (N_3585,N_2983,N_2913);
or U3586 (N_3586,N_2883,N_2967);
nand U3587 (N_3587,N_2858,N_2921);
and U3588 (N_3588,N_3093,N_3055);
xor U3589 (N_3589,N_2981,N_3054);
and U3590 (N_3590,N_3102,N_3007);
xor U3591 (N_3591,N_3146,N_2859);
or U3592 (N_3592,N_3112,N_3049);
xnor U3593 (N_3593,N_2956,N_2927);
nor U3594 (N_3594,N_3147,N_2819);
xnor U3595 (N_3595,N_3041,N_3058);
and U3596 (N_3596,N_3100,N_3065);
nand U3597 (N_3597,N_3068,N_2973);
or U3598 (N_3598,N_2834,N_3083);
and U3599 (N_3599,N_2822,N_2979);
and U3600 (N_3600,N_3309,N_3392);
or U3601 (N_3601,N_3510,N_3304);
xnor U3602 (N_3602,N_3417,N_3519);
nand U3603 (N_3603,N_3327,N_3336);
nor U3604 (N_3604,N_3215,N_3250);
and U3605 (N_3605,N_3216,N_3295);
or U3606 (N_3606,N_3503,N_3213);
nand U3607 (N_3607,N_3361,N_3463);
nand U3608 (N_3608,N_3329,N_3465);
xnor U3609 (N_3609,N_3240,N_3315);
xnor U3610 (N_3610,N_3350,N_3474);
nor U3611 (N_3611,N_3478,N_3439);
and U3612 (N_3612,N_3522,N_3207);
and U3613 (N_3613,N_3449,N_3411);
and U3614 (N_3614,N_3498,N_3460);
xnor U3615 (N_3615,N_3322,N_3370);
or U3616 (N_3616,N_3490,N_3403);
nand U3617 (N_3617,N_3338,N_3367);
or U3618 (N_3618,N_3316,N_3406);
nor U3619 (N_3619,N_3468,N_3530);
and U3620 (N_3620,N_3248,N_3532);
or U3621 (N_3621,N_3223,N_3589);
or U3622 (N_3622,N_3287,N_3337);
and U3623 (N_3623,N_3516,N_3212);
nand U3624 (N_3624,N_3418,N_3475);
xnor U3625 (N_3625,N_3274,N_3257);
or U3626 (N_3626,N_3480,N_3282);
xor U3627 (N_3627,N_3564,N_3552);
nor U3628 (N_3628,N_3229,N_3586);
xor U3629 (N_3629,N_3563,N_3550);
or U3630 (N_3630,N_3587,N_3390);
and U3631 (N_3631,N_3527,N_3515);
and U3632 (N_3632,N_3505,N_3224);
xnor U3633 (N_3633,N_3339,N_3579);
xnor U3634 (N_3634,N_3483,N_3599);
nor U3635 (N_3635,N_3517,N_3397);
nor U3636 (N_3636,N_3299,N_3204);
and U3637 (N_3637,N_3317,N_3412);
and U3638 (N_3638,N_3531,N_3311);
xnor U3639 (N_3639,N_3542,N_3266);
and U3640 (N_3640,N_3259,N_3228);
and U3641 (N_3641,N_3536,N_3497);
nor U3642 (N_3642,N_3584,N_3267);
nand U3643 (N_3643,N_3492,N_3371);
and U3644 (N_3644,N_3328,N_3398);
and U3645 (N_3645,N_3388,N_3422);
and U3646 (N_3646,N_3231,N_3539);
and U3647 (N_3647,N_3400,N_3333);
and U3648 (N_3648,N_3362,N_3500);
xor U3649 (N_3649,N_3445,N_3377);
nor U3650 (N_3650,N_3258,N_3448);
and U3651 (N_3651,N_3383,N_3544);
nand U3652 (N_3652,N_3507,N_3585);
or U3653 (N_3653,N_3344,N_3323);
or U3654 (N_3654,N_3375,N_3293);
and U3655 (N_3655,N_3538,N_3434);
xor U3656 (N_3656,N_3386,N_3302);
nand U3657 (N_3657,N_3238,N_3440);
or U3658 (N_3658,N_3296,N_3473);
xnor U3659 (N_3659,N_3408,N_3308);
and U3660 (N_3660,N_3272,N_3429);
nand U3661 (N_3661,N_3218,N_3312);
nand U3662 (N_3662,N_3413,N_3526);
nand U3663 (N_3663,N_3580,N_3583);
or U3664 (N_3664,N_3470,N_3410);
xor U3665 (N_3665,N_3594,N_3226);
or U3666 (N_3666,N_3358,N_3285);
nor U3667 (N_3667,N_3425,N_3549);
xnor U3668 (N_3668,N_3247,N_3241);
and U3669 (N_3669,N_3235,N_3236);
nand U3670 (N_3670,N_3513,N_3568);
nor U3671 (N_3671,N_3540,N_3442);
nand U3672 (N_3672,N_3225,N_3577);
or U3673 (N_3673,N_3281,N_3276);
and U3674 (N_3674,N_3313,N_3202);
and U3675 (N_3675,N_3331,N_3576);
xor U3676 (N_3676,N_3496,N_3263);
and U3677 (N_3677,N_3464,N_3446);
nor U3678 (N_3678,N_3545,N_3428);
xnor U3679 (N_3679,N_3234,N_3346);
and U3680 (N_3680,N_3501,N_3562);
nand U3681 (N_3681,N_3222,N_3221);
xor U3682 (N_3682,N_3546,N_3591);
nand U3683 (N_3683,N_3488,N_3356);
and U3684 (N_3684,N_3565,N_3363);
nand U3685 (N_3685,N_3399,N_3593);
nand U3686 (N_3686,N_3487,N_3572);
and U3687 (N_3687,N_3255,N_3206);
nand U3688 (N_3688,N_3374,N_3277);
or U3689 (N_3689,N_3220,N_3486);
nand U3690 (N_3690,N_3368,N_3438);
and U3691 (N_3691,N_3479,N_3525);
and U3692 (N_3692,N_3453,N_3376);
nand U3693 (N_3693,N_3462,N_3237);
xor U3694 (N_3694,N_3432,N_3260);
nand U3695 (N_3695,N_3242,N_3269);
and U3696 (N_3696,N_3427,N_3347);
nand U3697 (N_3697,N_3279,N_3431);
or U3698 (N_3698,N_3314,N_3405);
nand U3699 (N_3699,N_3533,N_3203);
xor U3700 (N_3700,N_3265,N_3423);
nand U3701 (N_3701,N_3249,N_3384);
and U3702 (N_3702,N_3205,N_3307);
xnor U3703 (N_3703,N_3320,N_3290);
or U3704 (N_3704,N_3528,N_3401);
and U3705 (N_3705,N_3596,N_3433);
and U3706 (N_3706,N_3289,N_3246);
and U3707 (N_3707,N_3566,N_3381);
or U3708 (N_3708,N_3214,N_3211);
and U3709 (N_3709,N_3209,N_3447);
xor U3710 (N_3710,N_3455,N_3441);
nand U3711 (N_3711,N_3414,N_3430);
nand U3712 (N_3712,N_3556,N_3499);
or U3713 (N_3713,N_3450,N_3387);
and U3714 (N_3714,N_3511,N_3421);
or U3715 (N_3715,N_3286,N_3424);
nand U3716 (N_3716,N_3506,N_3489);
and U3717 (N_3717,N_3553,N_3471);
nor U3718 (N_3718,N_3534,N_3219);
and U3719 (N_3719,N_3523,N_3349);
or U3720 (N_3720,N_3598,N_3554);
xnor U3721 (N_3721,N_3360,N_3491);
or U3722 (N_3722,N_3466,N_3345);
xnor U3723 (N_3723,N_3391,N_3354);
xor U3724 (N_3724,N_3416,N_3404);
or U3725 (N_3725,N_3559,N_3548);
or U3726 (N_3726,N_3458,N_3348);
nor U3727 (N_3727,N_3396,N_3588);
nor U3728 (N_3728,N_3451,N_3210);
and U3729 (N_3729,N_3493,N_3318);
and U3730 (N_3730,N_3292,N_3567);
nand U3731 (N_3731,N_3297,N_3557);
xor U3732 (N_3732,N_3415,N_3504);
or U3733 (N_3733,N_3514,N_3407);
and U3734 (N_3734,N_3341,N_3402);
or U3735 (N_3735,N_3306,N_3590);
nor U3736 (N_3736,N_3570,N_3443);
nor U3737 (N_3737,N_3300,N_3324);
nand U3738 (N_3738,N_3574,N_3420);
and U3739 (N_3739,N_3535,N_3472);
nor U3740 (N_3740,N_3581,N_3230);
or U3741 (N_3741,N_3365,N_3456);
xor U3742 (N_3742,N_3334,N_3294);
xor U3743 (N_3743,N_3518,N_3547);
or U3744 (N_3744,N_3520,N_3254);
or U3745 (N_3745,N_3541,N_3270);
nor U3746 (N_3746,N_3394,N_3325);
or U3747 (N_3747,N_3232,N_3521);
xor U3748 (N_3748,N_3495,N_3342);
and U3749 (N_3749,N_3461,N_3419);
nand U3750 (N_3750,N_3343,N_3571);
nand U3751 (N_3751,N_3459,N_3271);
and U3752 (N_3752,N_3569,N_3597);
xnor U3753 (N_3753,N_3551,N_3382);
xnor U3754 (N_3754,N_3305,N_3366);
and U3755 (N_3755,N_3201,N_3310);
xnor U3756 (N_3756,N_3227,N_3373);
nor U3757 (N_3757,N_3364,N_3273);
xnor U3758 (N_3758,N_3524,N_3200);
and U3759 (N_3759,N_3379,N_3326);
nor U3760 (N_3760,N_3239,N_3351);
and U3761 (N_3761,N_3543,N_3243);
and U3762 (N_3762,N_3359,N_3330);
xnor U3763 (N_3763,N_3537,N_3494);
nor U3764 (N_3764,N_3509,N_3262);
nand U3765 (N_3765,N_3595,N_3357);
or U3766 (N_3766,N_3502,N_3476);
xor U3767 (N_3767,N_3575,N_3508);
nand U3768 (N_3768,N_3284,N_3484);
nand U3769 (N_3769,N_3245,N_3457);
nor U3770 (N_3770,N_3298,N_3409);
or U3771 (N_3771,N_3481,N_3452);
and U3772 (N_3772,N_3444,N_3283);
nand U3773 (N_3773,N_3321,N_3291);
or U3774 (N_3774,N_3301,N_3352);
or U3775 (N_3775,N_3275,N_3512);
nor U3776 (N_3776,N_3426,N_3561);
or U3777 (N_3777,N_3208,N_3319);
xnor U3778 (N_3778,N_3385,N_3454);
xor U3779 (N_3779,N_3485,N_3469);
nand U3780 (N_3780,N_3252,N_3256);
and U3781 (N_3781,N_3482,N_3529);
or U3782 (N_3782,N_3437,N_3592);
and U3783 (N_3783,N_3288,N_3278);
or U3784 (N_3784,N_3393,N_3233);
xnor U3785 (N_3785,N_3251,N_3280);
and U3786 (N_3786,N_3378,N_3335);
xor U3787 (N_3787,N_3369,N_3264);
or U3788 (N_3788,N_3578,N_3573);
or U3789 (N_3789,N_3244,N_3395);
nand U3790 (N_3790,N_3436,N_3332);
xor U3791 (N_3791,N_3355,N_3560);
or U3792 (N_3792,N_3261,N_3467);
or U3793 (N_3793,N_3217,N_3380);
nor U3794 (N_3794,N_3253,N_3372);
nor U3795 (N_3795,N_3555,N_3353);
nor U3796 (N_3796,N_3558,N_3435);
xnor U3797 (N_3797,N_3303,N_3477);
and U3798 (N_3798,N_3582,N_3340);
nand U3799 (N_3799,N_3268,N_3389);
and U3800 (N_3800,N_3217,N_3506);
xnor U3801 (N_3801,N_3447,N_3362);
nand U3802 (N_3802,N_3599,N_3364);
nor U3803 (N_3803,N_3557,N_3580);
or U3804 (N_3804,N_3368,N_3580);
nand U3805 (N_3805,N_3588,N_3444);
nor U3806 (N_3806,N_3347,N_3215);
nor U3807 (N_3807,N_3314,N_3280);
xor U3808 (N_3808,N_3227,N_3393);
nand U3809 (N_3809,N_3516,N_3373);
nor U3810 (N_3810,N_3580,N_3386);
nand U3811 (N_3811,N_3500,N_3491);
nand U3812 (N_3812,N_3452,N_3474);
nand U3813 (N_3813,N_3283,N_3288);
nand U3814 (N_3814,N_3244,N_3299);
nand U3815 (N_3815,N_3517,N_3404);
nand U3816 (N_3816,N_3595,N_3486);
xor U3817 (N_3817,N_3278,N_3205);
and U3818 (N_3818,N_3579,N_3447);
or U3819 (N_3819,N_3509,N_3225);
nor U3820 (N_3820,N_3473,N_3515);
and U3821 (N_3821,N_3572,N_3336);
nand U3822 (N_3822,N_3370,N_3283);
nand U3823 (N_3823,N_3230,N_3338);
nand U3824 (N_3824,N_3596,N_3201);
and U3825 (N_3825,N_3312,N_3511);
or U3826 (N_3826,N_3428,N_3305);
nand U3827 (N_3827,N_3456,N_3206);
or U3828 (N_3828,N_3400,N_3349);
nor U3829 (N_3829,N_3276,N_3581);
and U3830 (N_3830,N_3316,N_3565);
xnor U3831 (N_3831,N_3463,N_3321);
or U3832 (N_3832,N_3348,N_3508);
nor U3833 (N_3833,N_3550,N_3367);
nor U3834 (N_3834,N_3378,N_3372);
nor U3835 (N_3835,N_3568,N_3320);
nor U3836 (N_3836,N_3485,N_3495);
nand U3837 (N_3837,N_3291,N_3560);
xnor U3838 (N_3838,N_3464,N_3254);
or U3839 (N_3839,N_3224,N_3585);
nand U3840 (N_3840,N_3554,N_3227);
nand U3841 (N_3841,N_3533,N_3543);
nand U3842 (N_3842,N_3318,N_3237);
and U3843 (N_3843,N_3581,N_3243);
nor U3844 (N_3844,N_3439,N_3441);
and U3845 (N_3845,N_3363,N_3571);
and U3846 (N_3846,N_3374,N_3398);
nor U3847 (N_3847,N_3252,N_3424);
xor U3848 (N_3848,N_3457,N_3336);
or U3849 (N_3849,N_3336,N_3316);
nand U3850 (N_3850,N_3283,N_3246);
nand U3851 (N_3851,N_3294,N_3272);
nor U3852 (N_3852,N_3454,N_3250);
nor U3853 (N_3853,N_3483,N_3242);
nor U3854 (N_3854,N_3567,N_3230);
and U3855 (N_3855,N_3393,N_3547);
and U3856 (N_3856,N_3441,N_3572);
nand U3857 (N_3857,N_3237,N_3408);
nand U3858 (N_3858,N_3458,N_3582);
nand U3859 (N_3859,N_3546,N_3249);
and U3860 (N_3860,N_3533,N_3252);
or U3861 (N_3861,N_3356,N_3286);
xor U3862 (N_3862,N_3511,N_3591);
and U3863 (N_3863,N_3548,N_3320);
xnor U3864 (N_3864,N_3456,N_3298);
xnor U3865 (N_3865,N_3466,N_3249);
nand U3866 (N_3866,N_3228,N_3598);
nor U3867 (N_3867,N_3590,N_3474);
nor U3868 (N_3868,N_3495,N_3214);
and U3869 (N_3869,N_3284,N_3323);
nor U3870 (N_3870,N_3403,N_3536);
nor U3871 (N_3871,N_3408,N_3258);
and U3872 (N_3872,N_3570,N_3314);
or U3873 (N_3873,N_3229,N_3314);
xor U3874 (N_3874,N_3260,N_3498);
nand U3875 (N_3875,N_3221,N_3220);
and U3876 (N_3876,N_3522,N_3597);
xnor U3877 (N_3877,N_3484,N_3393);
and U3878 (N_3878,N_3336,N_3376);
and U3879 (N_3879,N_3342,N_3316);
and U3880 (N_3880,N_3542,N_3410);
and U3881 (N_3881,N_3274,N_3594);
nand U3882 (N_3882,N_3290,N_3397);
or U3883 (N_3883,N_3552,N_3462);
xnor U3884 (N_3884,N_3575,N_3215);
xnor U3885 (N_3885,N_3290,N_3251);
and U3886 (N_3886,N_3513,N_3417);
or U3887 (N_3887,N_3497,N_3527);
and U3888 (N_3888,N_3499,N_3403);
xor U3889 (N_3889,N_3251,N_3420);
nand U3890 (N_3890,N_3381,N_3400);
xnor U3891 (N_3891,N_3298,N_3414);
xor U3892 (N_3892,N_3564,N_3479);
xor U3893 (N_3893,N_3487,N_3318);
or U3894 (N_3894,N_3238,N_3421);
or U3895 (N_3895,N_3296,N_3435);
or U3896 (N_3896,N_3377,N_3487);
nand U3897 (N_3897,N_3540,N_3364);
nor U3898 (N_3898,N_3304,N_3305);
xor U3899 (N_3899,N_3569,N_3583);
nand U3900 (N_3900,N_3566,N_3398);
or U3901 (N_3901,N_3573,N_3383);
nand U3902 (N_3902,N_3519,N_3551);
xor U3903 (N_3903,N_3350,N_3450);
and U3904 (N_3904,N_3465,N_3504);
and U3905 (N_3905,N_3300,N_3243);
nand U3906 (N_3906,N_3278,N_3214);
or U3907 (N_3907,N_3255,N_3208);
xor U3908 (N_3908,N_3202,N_3535);
nor U3909 (N_3909,N_3430,N_3360);
and U3910 (N_3910,N_3367,N_3427);
or U3911 (N_3911,N_3367,N_3511);
nor U3912 (N_3912,N_3427,N_3213);
and U3913 (N_3913,N_3597,N_3360);
xor U3914 (N_3914,N_3347,N_3404);
xnor U3915 (N_3915,N_3357,N_3252);
or U3916 (N_3916,N_3231,N_3294);
nor U3917 (N_3917,N_3398,N_3570);
nor U3918 (N_3918,N_3467,N_3577);
or U3919 (N_3919,N_3451,N_3458);
xnor U3920 (N_3920,N_3393,N_3474);
and U3921 (N_3921,N_3568,N_3326);
nor U3922 (N_3922,N_3594,N_3393);
or U3923 (N_3923,N_3209,N_3298);
or U3924 (N_3924,N_3350,N_3498);
nand U3925 (N_3925,N_3554,N_3318);
and U3926 (N_3926,N_3303,N_3561);
xor U3927 (N_3927,N_3553,N_3514);
or U3928 (N_3928,N_3475,N_3257);
and U3929 (N_3929,N_3389,N_3513);
nand U3930 (N_3930,N_3407,N_3387);
nor U3931 (N_3931,N_3310,N_3285);
and U3932 (N_3932,N_3217,N_3285);
nand U3933 (N_3933,N_3270,N_3315);
xnor U3934 (N_3934,N_3488,N_3437);
xor U3935 (N_3935,N_3533,N_3318);
xor U3936 (N_3936,N_3300,N_3249);
nor U3937 (N_3937,N_3505,N_3363);
or U3938 (N_3938,N_3425,N_3213);
nor U3939 (N_3939,N_3242,N_3537);
or U3940 (N_3940,N_3318,N_3241);
and U3941 (N_3941,N_3554,N_3205);
nor U3942 (N_3942,N_3521,N_3268);
xor U3943 (N_3943,N_3334,N_3315);
nand U3944 (N_3944,N_3288,N_3355);
or U3945 (N_3945,N_3532,N_3311);
nand U3946 (N_3946,N_3364,N_3244);
or U3947 (N_3947,N_3356,N_3567);
and U3948 (N_3948,N_3213,N_3221);
and U3949 (N_3949,N_3543,N_3425);
nand U3950 (N_3950,N_3504,N_3597);
nor U3951 (N_3951,N_3367,N_3451);
nand U3952 (N_3952,N_3540,N_3535);
nand U3953 (N_3953,N_3562,N_3351);
or U3954 (N_3954,N_3459,N_3441);
nor U3955 (N_3955,N_3543,N_3577);
or U3956 (N_3956,N_3529,N_3461);
xnor U3957 (N_3957,N_3578,N_3385);
and U3958 (N_3958,N_3292,N_3519);
nand U3959 (N_3959,N_3544,N_3489);
xor U3960 (N_3960,N_3212,N_3316);
nand U3961 (N_3961,N_3481,N_3245);
nor U3962 (N_3962,N_3424,N_3418);
and U3963 (N_3963,N_3439,N_3519);
nor U3964 (N_3964,N_3544,N_3297);
and U3965 (N_3965,N_3492,N_3324);
xnor U3966 (N_3966,N_3239,N_3381);
nor U3967 (N_3967,N_3205,N_3436);
xor U3968 (N_3968,N_3567,N_3373);
xnor U3969 (N_3969,N_3238,N_3441);
nor U3970 (N_3970,N_3249,N_3342);
xor U3971 (N_3971,N_3268,N_3292);
nand U3972 (N_3972,N_3433,N_3565);
and U3973 (N_3973,N_3516,N_3387);
nand U3974 (N_3974,N_3308,N_3232);
nor U3975 (N_3975,N_3595,N_3282);
or U3976 (N_3976,N_3310,N_3322);
nor U3977 (N_3977,N_3210,N_3598);
nand U3978 (N_3978,N_3566,N_3241);
and U3979 (N_3979,N_3559,N_3465);
nor U3980 (N_3980,N_3468,N_3347);
or U3981 (N_3981,N_3412,N_3345);
or U3982 (N_3982,N_3452,N_3540);
nand U3983 (N_3983,N_3373,N_3206);
nand U3984 (N_3984,N_3547,N_3272);
or U3985 (N_3985,N_3340,N_3541);
and U3986 (N_3986,N_3316,N_3294);
and U3987 (N_3987,N_3552,N_3478);
nand U3988 (N_3988,N_3461,N_3415);
nand U3989 (N_3989,N_3450,N_3214);
nor U3990 (N_3990,N_3556,N_3276);
xnor U3991 (N_3991,N_3504,N_3526);
nand U3992 (N_3992,N_3381,N_3317);
xnor U3993 (N_3993,N_3210,N_3311);
nand U3994 (N_3994,N_3322,N_3499);
nor U3995 (N_3995,N_3552,N_3481);
and U3996 (N_3996,N_3357,N_3298);
and U3997 (N_3997,N_3475,N_3503);
nor U3998 (N_3998,N_3411,N_3261);
nor U3999 (N_3999,N_3532,N_3546);
or U4000 (N_4000,N_3646,N_3637);
nor U4001 (N_4001,N_3693,N_3781);
xor U4002 (N_4002,N_3645,N_3964);
nor U4003 (N_4003,N_3875,N_3873);
and U4004 (N_4004,N_3634,N_3874);
or U4005 (N_4005,N_3619,N_3881);
and U4006 (N_4006,N_3798,N_3676);
and U4007 (N_4007,N_3754,N_3990);
nand U4008 (N_4008,N_3898,N_3918);
xnor U4009 (N_4009,N_3811,N_3666);
xor U4010 (N_4010,N_3989,N_3616);
xnor U4011 (N_4011,N_3607,N_3952);
nand U4012 (N_4012,N_3924,N_3909);
and U4013 (N_4013,N_3743,N_3677);
xor U4014 (N_4014,N_3672,N_3826);
nand U4015 (N_4015,N_3824,N_3644);
nand U4016 (N_4016,N_3922,N_3911);
nor U4017 (N_4017,N_3617,N_3780);
and U4018 (N_4018,N_3611,N_3707);
xnor U4019 (N_4019,N_3975,N_3769);
and U4020 (N_4020,N_3950,N_3632);
xor U4021 (N_4021,N_3949,N_3795);
nand U4022 (N_4022,N_3937,N_3741);
nor U4023 (N_4023,N_3778,N_3690);
xor U4024 (N_4024,N_3806,N_3804);
nand U4025 (N_4025,N_3731,N_3948);
xnor U4026 (N_4026,N_3863,N_3750);
nand U4027 (N_4027,N_3791,N_3868);
and U4028 (N_4028,N_3794,N_3669);
or U4029 (N_4029,N_3856,N_3932);
xor U4030 (N_4030,N_3788,N_3942);
or U4031 (N_4031,N_3673,N_3879);
or U4032 (N_4032,N_3972,N_3739);
and U4033 (N_4033,N_3810,N_3958);
or U4034 (N_4034,N_3913,N_3774);
xor U4035 (N_4035,N_3653,N_3638);
and U4036 (N_4036,N_3970,N_3947);
and U4037 (N_4037,N_3912,N_3728);
and U4038 (N_4038,N_3887,N_3923);
and U4039 (N_4039,N_3747,N_3738);
nand U4040 (N_4040,N_3792,N_3670);
xnor U4041 (N_4041,N_3822,N_3745);
xnor U4042 (N_4042,N_3787,N_3640);
xor U4043 (N_4043,N_3675,N_3603);
nor U4044 (N_4044,N_3998,N_3997);
nand U4045 (N_4045,N_3901,N_3749);
nor U4046 (N_4046,N_3761,N_3865);
xnor U4047 (N_4047,N_3776,N_3706);
xnor U4048 (N_4048,N_3613,N_3832);
nor U4049 (N_4049,N_3820,N_3725);
nor U4050 (N_4050,N_3680,N_3845);
nor U4051 (N_4051,N_3903,N_3934);
nor U4052 (N_4052,N_3759,N_3860);
nor U4053 (N_4053,N_3762,N_3967);
nor U4054 (N_4054,N_3620,N_3688);
and U4055 (N_4055,N_3930,N_3712);
and U4056 (N_4056,N_3891,N_3622);
and U4057 (N_4057,N_3662,N_3809);
or U4058 (N_4058,N_3940,N_3831);
nand U4059 (N_4059,N_3612,N_3757);
and U4060 (N_4060,N_3877,N_3803);
nor U4061 (N_4061,N_3604,N_3816);
nand U4062 (N_4062,N_3805,N_3802);
or U4063 (N_4063,N_3984,N_3827);
nand U4064 (N_4064,N_3661,N_3818);
or U4065 (N_4065,N_3734,N_3713);
nand U4066 (N_4066,N_3627,N_3751);
xnor U4067 (N_4067,N_3800,N_3855);
nor U4068 (N_4068,N_3629,N_3657);
xor U4069 (N_4069,N_3876,N_3847);
nor U4070 (N_4070,N_3885,N_3609);
xor U4071 (N_4071,N_3777,N_3862);
and U4072 (N_4072,N_3872,N_3718);
and U4073 (N_4073,N_3702,N_3758);
xor U4074 (N_4074,N_3878,N_3850);
nand U4075 (N_4075,N_3753,N_3605);
nand U4076 (N_4076,N_3819,N_3689);
nand U4077 (N_4077,N_3674,N_3900);
nand U4078 (N_4078,N_3601,N_3602);
or U4079 (N_4079,N_3721,N_3740);
or U4080 (N_4080,N_3985,N_3695);
nor U4081 (N_4081,N_3766,N_3708);
and U4082 (N_4082,N_3719,N_3987);
xnor U4083 (N_4083,N_3659,N_3821);
and U4084 (N_4084,N_3710,N_3973);
nand U4085 (N_4085,N_3732,N_3767);
and U4086 (N_4086,N_3969,N_3957);
and U4087 (N_4087,N_3979,N_3935);
xnor U4088 (N_4088,N_3928,N_3641);
nor U4089 (N_4089,N_3834,N_3894);
nor U4090 (N_4090,N_3848,N_3853);
nor U4091 (N_4091,N_3889,N_3796);
and U4092 (N_4092,N_3882,N_3807);
xnor U4093 (N_4093,N_3859,N_3699);
or U4094 (N_4094,N_3737,N_3765);
nand U4095 (N_4095,N_3888,N_3663);
or U4096 (N_4096,N_3671,N_3647);
xor U4097 (N_4097,N_3905,N_3775);
nor U4098 (N_4098,N_3956,N_3823);
nor U4099 (N_4099,N_3830,N_3698);
xnor U4100 (N_4100,N_3615,N_3733);
nor U4101 (N_4101,N_3782,N_3624);
nand U4102 (N_4102,N_3681,N_3991);
nor U4103 (N_4103,N_3814,N_3929);
xnor U4104 (N_4104,N_3880,N_3829);
xnor U4105 (N_4105,N_3944,N_3655);
and U4106 (N_4106,N_3927,N_3630);
nor U4107 (N_4107,N_3864,N_3633);
xor U4108 (N_4108,N_3919,N_3703);
or U4109 (N_4109,N_3883,N_3960);
xor U4110 (N_4110,N_3770,N_3892);
nand U4111 (N_4111,N_3628,N_3784);
xor U4112 (N_4112,N_3692,N_3642);
nor U4113 (N_4113,N_3705,N_3908);
nor U4114 (N_4114,N_3665,N_3768);
nor U4115 (N_4115,N_3682,N_3906);
nor U4116 (N_4116,N_3925,N_3623);
xnor U4117 (N_4117,N_3606,N_3939);
nor U4118 (N_4118,N_3686,N_3697);
or U4119 (N_4119,N_3684,N_3799);
nand U4120 (N_4120,N_3600,N_3717);
or U4121 (N_4121,N_3843,N_3771);
nor U4122 (N_4122,N_3841,N_3895);
xnor U4123 (N_4123,N_3654,N_3650);
nand U4124 (N_4124,N_3610,N_3978);
nand U4125 (N_4125,N_3700,N_3683);
and U4126 (N_4126,N_3730,N_3993);
nand U4127 (N_4127,N_3755,N_3696);
nand U4128 (N_4128,N_3965,N_3994);
xor U4129 (N_4129,N_3926,N_3722);
nand U4130 (N_4130,N_3854,N_3812);
nor U4131 (N_4131,N_3773,N_3867);
and U4132 (N_4132,N_3621,N_3961);
or U4133 (N_4133,N_3779,N_3667);
nor U4134 (N_4134,N_3954,N_3763);
or U4135 (N_4135,N_3715,N_3825);
nor U4136 (N_4136,N_3760,N_3846);
and U4137 (N_4137,N_3968,N_3723);
and U4138 (N_4138,N_3917,N_3836);
nand U4139 (N_4139,N_3742,N_3735);
nand U4140 (N_4140,N_3996,N_3959);
nand U4141 (N_4141,N_3983,N_3789);
or U4142 (N_4142,N_3720,N_3813);
and U4143 (N_4143,N_3636,N_3678);
nand U4144 (N_4144,N_3711,N_3986);
nor U4145 (N_4145,N_3904,N_3946);
and U4146 (N_4146,N_3910,N_3727);
nand U4147 (N_4147,N_3963,N_3691);
or U4148 (N_4148,N_3694,N_3614);
or U4149 (N_4149,N_3988,N_3902);
or U4150 (N_4150,N_3649,N_3943);
or U4151 (N_4151,N_3833,N_3941);
xnor U4152 (N_4152,N_3744,N_3842);
nand U4153 (N_4153,N_3626,N_3999);
xnor U4154 (N_4154,N_3899,N_3815);
xor U4155 (N_4155,N_3953,N_3938);
and U4156 (N_4156,N_3992,N_3658);
or U4157 (N_4157,N_3648,N_3748);
and U4158 (N_4158,N_3772,N_3783);
or U4159 (N_4159,N_3790,N_3982);
xnor U4160 (N_4160,N_3752,N_3651);
nand U4161 (N_4161,N_3668,N_3664);
nand U4162 (N_4162,N_3916,N_3709);
nor U4163 (N_4163,N_3980,N_3870);
or U4164 (N_4164,N_3652,N_3660);
xnor U4165 (N_4165,N_3951,N_3838);
nand U4166 (N_4166,N_3945,N_3851);
nand U4167 (N_4167,N_3840,N_3716);
nor U4168 (N_4168,N_3726,N_3955);
and U4169 (N_4169,N_3801,N_3890);
and U4170 (N_4170,N_3871,N_3835);
or U4171 (N_4171,N_3746,N_3995);
and U4172 (N_4172,N_3736,N_3962);
xor U4173 (N_4173,N_3921,N_3685);
or U4174 (N_4174,N_3724,N_3679);
and U4175 (N_4175,N_3974,N_3635);
xnor U4176 (N_4176,N_3785,N_3618);
nand U4177 (N_4177,N_3896,N_3861);
nor U4178 (N_4178,N_3849,N_3808);
nand U4179 (N_4179,N_3893,N_3852);
or U4180 (N_4180,N_3839,N_3966);
nand U4181 (N_4181,N_3976,N_3933);
nor U4182 (N_4182,N_3797,N_3857);
xor U4183 (N_4183,N_3687,N_3858);
nand U4184 (N_4184,N_3817,N_3793);
or U4185 (N_4185,N_3936,N_3625);
and U4186 (N_4186,N_3866,N_3608);
nor U4187 (N_4187,N_3756,N_3704);
or U4188 (N_4188,N_3786,N_3897);
or U4189 (N_4189,N_3631,N_3656);
nand U4190 (N_4190,N_3837,N_3714);
or U4191 (N_4191,N_3931,N_3884);
or U4192 (N_4192,N_3914,N_3764);
or U4193 (N_4193,N_3977,N_3844);
xor U4194 (N_4194,N_3828,N_3729);
nand U4195 (N_4195,N_3981,N_3907);
nor U4196 (N_4196,N_3643,N_3920);
or U4197 (N_4197,N_3869,N_3886);
xnor U4198 (N_4198,N_3639,N_3915);
xnor U4199 (N_4199,N_3701,N_3971);
xor U4200 (N_4200,N_3918,N_3672);
xnor U4201 (N_4201,N_3844,N_3707);
nor U4202 (N_4202,N_3713,N_3950);
nand U4203 (N_4203,N_3641,N_3924);
and U4204 (N_4204,N_3888,N_3814);
nand U4205 (N_4205,N_3890,N_3614);
nand U4206 (N_4206,N_3616,N_3961);
nor U4207 (N_4207,N_3977,N_3885);
nand U4208 (N_4208,N_3915,N_3662);
or U4209 (N_4209,N_3983,N_3630);
xor U4210 (N_4210,N_3891,N_3691);
nor U4211 (N_4211,N_3613,N_3699);
xor U4212 (N_4212,N_3606,N_3724);
and U4213 (N_4213,N_3851,N_3975);
nand U4214 (N_4214,N_3922,N_3883);
xor U4215 (N_4215,N_3776,N_3819);
xor U4216 (N_4216,N_3668,N_3843);
nor U4217 (N_4217,N_3956,N_3675);
and U4218 (N_4218,N_3794,N_3820);
nor U4219 (N_4219,N_3979,N_3700);
nand U4220 (N_4220,N_3908,N_3646);
nor U4221 (N_4221,N_3844,N_3831);
nand U4222 (N_4222,N_3767,N_3682);
and U4223 (N_4223,N_3702,N_3756);
xnor U4224 (N_4224,N_3823,N_3804);
and U4225 (N_4225,N_3727,N_3641);
nand U4226 (N_4226,N_3907,N_3650);
xnor U4227 (N_4227,N_3852,N_3844);
nand U4228 (N_4228,N_3614,N_3858);
nand U4229 (N_4229,N_3760,N_3894);
nand U4230 (N_4230,N_3807,N_3697);
nand U4231 (N_4231,N_3773,N_3690);
or U4232 (N_4232,N_3638,N_3770);
or U4233 (N_4233,N_3767,N_3891);
nand U4234 (N_4234,N_3836,N_3950);
xor U4235 (N_4235,N_3676,N_3880);
xnor U4236 (N_4236,N_3642,N_3687);
xor U4237 (N_4237,N_3919,N_3866);
nor U4238 (N_4238,N_3764,N_3803);
or U4239 (N_4239,N_3928,N_3741);
or U4240 (N_4240,N_3735,N_3931);
or U4241 (N_4241,N_3689,N_3745);
xnor U4242 (N_4242,N_3727,N_3681);
nand U4243 (N_4243,N_3965,N_3800);
nor U4244 (N_4244,N_3613,N_3964);
or U4245 (N_4245,N_3863,N_3622);
or U4246 (N_4246,N_3870,N_3795);
nor U4247 (N_4247,N_3995,N_3738);
nor U4248 (N_4248,N_3914,N_3744);
and U4249 (N_4249,N_3997,N_3729);
xor U4250 (N_4250,N_3663,N_3954);
and U4251 (N_4251,N_3681,N_3777);
nor U4252 (N_4252,N_3852,N_3756);
xor U4253 (N_4253,N_3914,N_3711);
nor U4254 (N_4254,N_3692,N_3992);
or U4255 (N_4255,N_3904,N_3871);
nor U4256 (N_4256,N_3845,N_3957);
nand U4257 (N_4257,N_3895,N_3941);
or U4258 (N_4258,N_3926,N_3810);
nor U4259 (N_4259,N_3714,N_3754);
or U4260 (N_4260,N_3626,N_3705);
and U4261 (N_4261,N_3687,N_3635);
or U4262 (N_4262,N_3655,N_3857);
nand U4263 (N_4263,N_3736,N_3906);
and U4264 (N_4264,N_3957,N_3733);
or U4265 (N_4265,N_3924,N_3801);
nor U4266 (N_4266,N_3814,N_3625);
or U4267 (N_4267,N_3847,N_3623);
nand U4268 (N_4268,N_3738,N_3678);
xor U4269 (N_4269,N_3816,N_3880);
nor U4270 (N_4270,N_3719,N_3936);
nand U4271 (N_4271,N_3681,N_3840);
and U4272 (N_4272,N_3874,N_3883);
nand U4273 (N_4273,N_3939,N_3851);
xnor U4274 (N_4274,N_3940,N_3612);
nand U4275 (N_4275,N_3997,N_3935);
nor U4276 (N_4276,N_3717,N_3928);
nor U4277 (N_4277,N_3920,N_3980);
and U4278 (N_4278,N_3924,N_3769);
xor U4279 (N_4279,N_3952,N_3646);
or U4280 (N_4280,N_3803,N_3824);
and U4281 (N_4281,N_3938,N_3929);
or U4282 (N_4282,N_3723,N_3733);
nand U4283 (N_4283,N_3879,N_3947);
xnor U4284 (N_4284,N_3709,N_3614);
xnor U4285 (N_4285,N_3678,N_3856);
nor U4286 (N_4286,N_3708,N_3919);
xor U4287 (N_4287,N_3878,N_3615);
nor U4288 (N_4288,N_3875,N_3928);
or U4289 (N_4289,N_3864,N_3714);
xor U4290 (N_4290,N_3741,N_3705);
or U4291 (N_4291,N_3698,N_3603);
nor U4292 (N_4292,N_3867,N_3634);
and U4293 (N_4293,N_3823,N_3833);
nand U4294 (N_4294,N_3721,N_3724);
and U4295 (N_4295,N_3618,N_3666);
and U4296 (N_4296,N_3977,N_3949);
or U4297 (N_4297,N_3605,N_3680);
or U4298 (N_4298,N_3994,N_3770);
nor U4299 (N_4299,N_3672,N_3971);
or U4300 (N_4300,N_3750,N_3872);
xnor U4301 (N_4301,N_3847,N_3783);
or U4302 (N_4302,N_3933,N_3928);
or U4303 (N_4303,N_3983,N_3857);
nand U4304 (N_4304,N_3686,N_3986);
nor U4305 (N_4305,N_3746,N_3993);
xnor U4306 (N_4306,N_3970,N_3705);
and U4307 (N_4307,N_3888,N_3612);
or U4308 (N_4308,N_3796,N_3644);
nand U4309 (N_4309,N_3645,N_3991);
nand U4310 (N_4310,N_3686,N_3749);
nand U4311 (N_4311,N_3896,N_3805);
nor U4312 (N_4312,N_3684,N_3806);
nand U4313 (N_4313,N_3768,N_3800);
or U4314 (N_4314,N_3612,N_3639);
xnor U4315 (N_4315,N_3876,N_3850);
nor U4316 (N_4316,N_3765,N_3773);
xor U4317 (N_4317,N_3878,N_3920);
xor U4318 (N_4318,N_3708,N_3993);
and U4319 (N_4319,N_3952,N_3631);
xor U4320 (N_4320,N_3946,N_3764);
and U4321 (N_4321,N_3858,N_3647);
nor U4322 (N_4322,N_3854,N_3888);
and U4323 (N_4323,N_3732,N_3844);
or U4324 (N_4324,N_3844,N_3690);
and U4325 (N_4325,N_3703,N_3972);
xor U4326 (N_4326,N_3928,N_3756);
nor U4327 (N_4327,N_3913,N_3936);
or U4328 (N_4328,N_3920,N_3669);
and U4329 (N_4329,N_3827,N_3657);
nand U4330 (N_4330,N_3709,N_3681);
or U4331 (N_4331,N_3812,N_3984);
xnor U4332 (N_4332,N_3694,N_3902);
and U4333 (N_4333,N_3717,N_3666);
and U4334 (N_4334,N_3977,N_3648);
xnor U4335 (N_4335,N_3864,N_3926);
or U4336 (N_4336,N_3635,N_3913);
xor U4337 (N_4337,N_3648,N_3763);
nor U4338 (N_4338,N_3910,N_3931);
xnor U4339 (N_4339,N_3894,N_3824);
nand U4340 (N_4340,N_3911,N_3956);
and U4341 (N_4341,N_3683,N_3618);
nand U4342 (N_4342,N_3729,N_3985);
or U4343 (N_4343,N_3822,N_3851);
and U4344 (N_4344,N_3853,N_3929);
and U4345 (N_4345,N_3815,N_3797);
and U4346 (N_4346,N_3887,N_3893);
xnor U4347 (N_4347,N_3923,N_3874);
xnor U4348 (N_4348,N_3831,N_3783);
nand U4349 (N_4349,N_3995,N_3980);
xor U4350 (N_4350,N_3863,N_3716);
and U4351 (N_4351,N_3914,N_3877);
nor U4352 (N_4352,N_3894,N_3613);
nor U4353 (N_4353,N_3814,N_3755);
nand U4354 (N_4354,N_3760,N_3863);
nand U4355 (N_4355,N_3737,N_3917);
nor U4356 (N_4356,N_3689,N_3601);
nor U4357 (N_4357,N_3851,N_3900);
or U4358 (N_4358,N_3669,N_3741);
nor U4359 (N_4359,N_3608,N_3800);
nand U4360 (N_4360,N_3858,N_3857);
nand U4361 (N_4361,N_3699,N_3606);
xor U4362 (N_4362,N_3659,N_3691);
and U4363 (N_4363,N_3936,N_3604);
or U4364 (N_4364,N_3854,N_3677);
nor U4365 (N_4365,N_3671,N_3879);
and U4366 (N_4366,N_3938,N_3650);
and U4367 (N_4367,N_3643,N_3839);
and U4368 (N_4368,N_3740,N_3613);
xnor U4369 (N_4369,N_3651,N_3833);
nand U4370 (N_4370,N_3659,N_3843);
nor U4371 (N_4371,N_3700,N_3609);
nor U4372 (N_4372,N_3837,N_3911);
nor U4373 (N_4373,N_3904,N_3680);
and U4374 (N_4374,N_3858,N_3887);
xor U4375 (N_4375,N_3853,N_3927);
and U4376 (N_4376,N_3632,N_3910);
or U4377 (N_4377,N_3698,N_3976);
nor U4378 (N_4378,N_3862,N_3802);
nand U4379 (N_4379,N_3948,N_3699);
or U4380 (N_4380,N_3845,N_3828);
or U4381 (N_4381,N_3872,N_3998);
and U4382 (N_4382,N_3887,N_3826);
or U4383 (N_4383,N_3844,N_3655);
or U4384 (N_4384,N_3835,N_3806);
nand U4385 (N_4385,N_3624,N_3757);
or U4386 (N_4386,N_3600,N_3946);
xnor U4387 (N_4387,N_3961,N_3639);
nand U4388 (N_4388,N_3839,N_3763);
nand U4389 (N_4389,N_3827,N_3688);
or U4390 (N_4390,N_3960,N_3813);
and U4391 (N_4391,N_3707,N_3678);
nand U4392 (N_4392,N_3780,N_3984);
xnor U4393 (N_4393,N_3732,N_3613);
xnor U4394 (N_4394,N_3783,N_3603);
and U4395 (N_4395,N_3908,N_3970);
or U4396 (N_4396,N_3699,N_3716);
nor U4397 (N_4397,N_3622,N_3844);
or U4398 (N_4398,N_3827,N_3766);
nor U4399 (N_4399,N_3633,N_3616);
nand U4400 (N_4400,N_4208,N_4192);
or U4401 (N_4401,N_4075,N_4132);
or U4402 (N_4402,N_4303,N_4153);
nand U4403 (N_4403,N_4367,N_4291);
xnor U4404 (N_4404,N_4321,N_4210);
xnor U4405 (N_4405,N_4378,N_4341);
or U4406 (N_4406,N_4113,N_4056);
or U4407 (N_4407,N_4123,N_4306);
nor U4408 (N_4408,N_4252,N_4081);
nand U4409 (N_4409,N_4028,N_4147);
or U4410 (N_4410,N_4246,N_4371);
nand U4411 (N_4411,N_4307,N_4216);
nand U4412 (N_4412,N_4296,N_4279);
xnor U4413 (N_4413,N_4396,N_4323);
nand U4414 (N_4414,N_4036,N_4095);
xor U4415 (N_4415,N_4100,N_4399);
nand U4416 (N_4416,N_4394,N_4373);
nand U4417 (N_4417,N_4333,N_4227);
nand U4418 (N_4418,N_4012,N_4005);
or U4419 (N_4419,N_4156,N_4034);
nand U4420 (N_4420,N_4224,N_4327);
nor U4421 (N_4421,N_4070,N_4173);
nor U4422 (N_4422,N_4236,N_4003);
xnor U4423 (N_4423,N_4043,N_4335);
nor U4424 (N_4424,N_4151,N_4134);
and U4425 (N_4425,N_4127,N_4266);
xnor U4426 (N_4426,N_4154,N_4260);
nand U4427 (N_4427,N_4242,N_4239);
nand U4428 (N_4428,N_4118,N_4128);
and U4429 (N_4429,N_4293,N_4365);
or U4430 (N_4430,N_4097,N_4200);
nand U4431 (N_4431,N_4361,N_4244);
nor U4432 (N_4432,N_4344,N_4355);
or U4433 (N_4433,N_4018,N_4363);
nor U4434 (N_4434,N_4025,N_4146);
and U4435 (N_4435,N_4276,N_4179);
or U4436 (N_4436,N_4073,N_4368);
nand U4437 (N_4437,N_4275,N_4250);
nor U4438 (N_4438,N_4254,N_4330);
and U4439 (N_4439,N_4105,N_4141);
or U4440 (N_4440,N_4129,N_4230);
or U4441 (N_4441,N_4271,N_4196);
xor U4442 (N_4442,N_4114,N_4088);
nor U4443 (N_4443,N_4176,N_4274);
and U4444 (N_4444,N_4352,N_4382);
nand U4445 (N_4445,N_4066,N_4152);
nor U4446 (N_4446,N_4009,N_4305);
xnor U4447 (N_4447,N_4150,N_4169);
nand U4448 (N_4448,N_4071,N_4063);
xor U4449 (N_4449,N_4002,N_4024);
or U4450 (N_4450,N_4353,N_4023);
or U4451 (N_4451,N_4051,N_4162);
or U4452 (N_4452,N_4389,N_4313);
or U4453 (N_4453,N_4297,N_4261);
nand U4454 (N_4454,N_4186,N_4046);
nand U4455 (N_4455,N_4057,N_4386);
or U4456 (N_4456,N_4052,N_4331);
nor U4457 (N_4457,N_4388,N_4161);
nand U4458 (N_4458,N_4251,N_4093);
nor U4459 (N_4459,N_4229,N_4283);
nor U4460 (N_4460,N_4272,N_4112);
or U4461 (N_4461,N_4326,N_4245);
or U4462 (N_4462,N_4180,N_4017);
nand U4463 (N_4463,N_4101,N_4202);
nor U4464 (N_4464,N_4064,N_4302);
or U4465 (N_4465,N_4068,N_4050);
or U4466 (N_4466,N_4354,N_4234);
nor U4467 (N_4467,N_4304,N_4339);
nor U4468 (N_4468,N_4285,N_4155);
or U4469 (N_4469,N_4164,N_4182);
nand U4470 (N_4470,N_4092,N_4022);
and U4471 (N_4471,N_4026,N_4011);
or U4472 (N_4472,N_4243,N_4209);
or U4473 (N_4473,N_4054,N_4312);
nor U4474 (N_4474,N_4139,N_4178);
nand U4475 (N_4475,N_4048,N_4165);
xor U4476 (N_4476,N_4122,N_4084);
or U4477 (N_4477,N_4265,N_4356);
and U4478 (N_4478,N_4079,N_4387);
and U4479 (N_4479,N_4248,N_4171);
or U4480 (N_4480,N_4351,N_4278);
or U4481 (N_4481,N_4294,N_4223);
xor U4482 (N_4482,N_4309,N_4348);
nand U4483 (N_4483,N_4350,N_4393);
and U4484 (N_4484,N_4383,N_4201);
xor U4485 (N_4485,N_4019,N_4374);
xor U4486 (N_4486,N_4035,N_4332);
or U4487 (N_4487,N_4214,N_4218);
and U4488 (N_4488,N_4044,N_4148);
and U4489 (N_4489,N_4379,N_4119);
or U4490 (N_4490,N_4108,N_4299);
nand U4491 (N_4491,N_4189,N_4238);
xnor U4492 (N_4492,N_4130,N_4167);
xnor U4493 (N_4493,N_4170,N_4172);
nand U4494 (N_4494,N_4256,N_4083);
xnor U4495 (N_4495,N_4324,N_4264);
xnor U4496 (N_4496,N_4049,N_4174);
xor U4497 (N_4497,N_4273,N_4194);
and U4498 (N_4498,N_4398,N_4337);
nor U4499 (N_4499,N_4377,N_4041);
xor U4500 (N_4500,N_4329,N_4006);
xnor U4501 (N_4501,N_4369,N_4376);
and U4502 (N_4502,N_4007,N_4366);
nor U4503 (N_4503,N_4221,N_4163);
xor U4504 (N_4504,N_4397,N_4072);
xor U4505 (N_4505,N_4298,N_4077);
nor U4506 (N_4506,N_4149,N_4027);
nor U4507 (N_4507,N_4222,N_4203);
nand U4508 (N_4508,N_4207,N_4029);
nor U4509 (N_4509,N_4267,N_4395);
or U4510 (N_4510,N_4342,N_4287);
or U4511 (N_4511,N_4020,N_4080);
xnor U4512 (N_4512,N_4257,N_4136);
nor U4513 (N_4513,N_4206,N_4219);
or U4514 (N_4514,N_4037,N_4262);
or U4515 (N_4515,N_4258,N_4142);
and U4516 (N_4516,N_4385,N_4059);
or U4517 (N_4517,N_4199,N_4381);
xor U4518 (N_4518,N_4177,N_4082);
nor U4519 (N_4519,N_4021,N_4269);
nand U4520 (N_4520,N_4340,N_4008);
nand U4521 (N_4521,N_4213,N_4345);
xor U4522 (N_4522,N_4187,N_4282);
and U4523 (N_4523,N_4181,N_4107);
xnor U4524 (N_4524,N_4133,N_4362);
xnor U4525 (N_4525,N_4175,N_4033);
nand U4526 (N_4526,N_4109,N_4315);
nor U4527 (N_4527,N_4228,N_4085);
nor U4528 (N_4528,N_4065,N_4268);
and U4529 (N_4529,N_4058,N_4288);
and U4530 (N_4530,N_4010,N_4115);
and U4531 (N_4531,N_4074,N_4205);
or U4532 (N_4532,N_4126,N_4241);
nand U4533 (N_4533,N_4193,N_4295);
or U4534 (N_4534,N_4102,N_4322);
nand U4535 (N_4535,N_4137,N_4391);
and U4536 (N_4536,N_4184,N_4053);
xnor U4537 (N_4537,N_4259,N_4096);
nand U4538 (N_4538,N_4121,N_4131);
or U4539 (N_4539,N_4346,N_4380);
xnor U4540 (N_4540,N_4042,N_4031);
or U4541 (N_4541,N_4292,N_4090);
or U4542 (N_4542,N_4231,N_4078);
nand U4543 (N_4543,N_4325,N_4370);
xor U4544 (N_4544,N_4240,N_4125);
and U4545 (N_4545,N_4349,N_4390);
nor U4546 (N_4546,N_4098,N_4392);
and U4547 (N_4547,N_4328,N_4076);
nand U4548 (N_4548,N_4284,N_4289);
xnor U4549 (N_4549,N_4040,N_4117);
and U4550 (N_4550,N_4166,N_4168);
and U4551 (N_4551,N_4357,N_4045);
nor U4552 (N_4552,N_4138,N_4384);
nor U4553 (N_4553,N_4318,N_4300);
nor U4554 (N_4554,N_4232,N_4310);
or U4555 (N_4555,N_4198,N_4067);
xor U4556 (N_4556,N_4111,N_4220);
nor U4557 (N_4557,N_4217,N_4336);
or U4558 (N_4558,N_4016,N_4091);
xor U4559 (N_4559,N_4104,N_4110);
nor U4560 (N_4560,N_4343,N_4060);
and U4561 (N_4561,N_4185,N_4347);
xnor U4562 (N_4562,N_4233,N_4263);
xnor U4563 (N_4563,N_4281,N_4145);
nor U4564 (N_4564,N_4247,N_4124);
nand U4565 (N_4565,N_4094,N_4055);
xnor U4566 (N_4566,N_4069,N_4249);
and U4567 (N_4567,N_4160,N_4375);
and U4568 (N_4568,N_4372,N_4211);
nand U4569 (N_4569,N_4195,N_4225);
or U4570 (N_4570,N_4099,N_4191);
nor U4571 (N_4571,N_4237,N_4158);
nand U4572 (N_4572,N_4197,N_4030);
nor U4573 (N_4573,N_4212,N_4159);
nand U4574 (N_4574,N_4140,N_4280);
or U4575 (N_4575,N_4061,N_4047);
xnor U4576 (N_4576,N_4062,N_4314);
xor U4577 (N_4577,N_4286,N_4014);
or U4578 (N_4578,N_4204,N_4039);
or U4579 (N_4579,N_4270,N_4135);
nand U4580 (N_4580,N_4255,N_4215);
xnor U4581 (N_4581,N_4277,N_4317);
nor U4582 (N_4582,N_4290,N_4226);
nand U4583 (N_4583,N_4120,N_4143);
xor U4584 (N_4584,N_4360,N_4364);
or U4585 (N_4585,N_4338,N_4103);
and U4586 (N_4586,N_4183,N_4308);
and U4587 (N_4587,N_4157,N_4320);
or U4588 (N_4588,N_4188,N_4316);
or U4589 (N_4589,N_4089,N_4087);
nor U4590 (N_4590,N_4106,N_4015);
nor U4591 (N_4591,N_4358,N_4190);
nor U4592 (N_4592,N_4000,N_4038);
or U4593 (N_4593,N_4004,N_4001);
or U4594 (N_4594,N_4311,N_4013);
nor U4595 (N_4595,N_4086,N_4032);
and U4596 (N_4596,N_4235,N_4359);
nor U4597 (N_4597,N_4334,N_4319);
or U4598 (N_4598,N_4116,N_4253);
xor U4599 (N_4599,N_4301,N_4144);
or U4600 (N_4600,N_4353,N_4379);
xor U4601 (N_4601,N_4174,N_4165);
nand U4602 (N_4602,N_4088,N_4308);
nor U4603 (N_4603,N_4011,N_4141);
nor U4604 (N_4604,N_4069,N_4173);
nand U4605 (N_4605,N_4142,N_4178);
and U4606 (N_4606,N_4087,N_4159);
nand U4607 (N_4607,N_4015,N_4112);
nand U4608 (N_4608,N_4240,N_4150);
xnor U4609 (N_4609,N_4016,N_4064);
nand U4610 (N_4610,N_4011,N_4342);
xor U4611 (N_4611,N_4284,N_4278);
or U4612 (N_4612,N_4157,N_4082);
nand U4613 (N_4613,N_4080,N_4179);
nor U4614 (N_4614,N_4322,N_4356);
and U4615 (N_4615,N_4127,N_4384);
xnor U4616 (N_4616,N_4012,N_4094);
nand U4617 (N_4617,N_4386,N_4255);
and U4618 (N_4618,N_4073,N_4319);
xnor U4619 (N_4619,N_4036,N_4164);
nor U4620 (N_4620,N_4005,N_4032);
xor U4621 (N_4621,N_4298,N_4378);
xor U4622 (N_4622,N_4192,N_4246);
or U4623 (N_4623,N_4037,N_4148);
nand U4624 (N_4624,N_4334,N_4367);
and U4625 (N_4625,N_4054,N_4332);
or U4626 (N_4626,N_4079,N_4075);
and U4627 (N_4627,N_4086,N_4275);
nor U4628 (N_4628,N_4179,N_4140);
nor U4629 (N_4629,N_4124,N_4258);
or U4630 (N_4630,N_4004,N_4281);
or U4631 (N_4631,N_4116,N_4159);
and U4632 (N_4632,N_4392,N_4356);
or U4633 (N_4633,N_4034,N_4330);
xor U4634 (N_4634,N_4034,N_4235);
nor U4635 (N_4635,N_4216,N_4372);
nand U4636 (N_4636,N_4011,N_4198);
nor U4637 (N_4637,N_4124,N_4251);
nand U4638 (N_4638,N_4232,N_4392);
or U4639 (N_4639,N_4010,N_4390);
nand U4640 (N_4640,N_4297,N_4262);
xor U4641 (N_4641,N_4373,N_4062);
and U4642 (N_4642,N_4149,N_4329);
xnor U4643 (N_4643,N_4224,N_4185);
nor U4644 (N_4644,N_4171,N_4223);
xor U4645 (N_4645,N_4284,N_4169);
nand U4646 (N_4646,N_4365,N_4061);
xnor U4647 (N_4647,N_4038,N_4173);
or U4648 (N_4648,N_4250,N_4170);
nor U4649 (N_4649,N_4089,N_4034);
nand U4650 (N_4650,N_4317,N_4081);
nor U4651 (N_4651,N_4336,N_4282);
xnor U4652 (N_4652,N_4227,N_4117);
nor U4653 (N_4653,N_4250,N_4355);
and U4654 (N_4654,N_4323,N_4232);
and U4655 (N_4655,N_4255,N_4077);
nand U4656 (N_4656,N_4051,N_4155);
nor U4657 (N_4657,N_4087,N_4138);
xnor U4658 (N_4658,N_4060,N_4199);
xor U4659 (N_4659,N_4347,N_4079);
and U4660 (N_4660,N_4397,N_4196);
or U4661 (N_4661,N_4258,N_4350);
nor U4662 (N_4662,N_4135,N_4046);
xnor U4663 (N_4663,N_4064,N_4009);
xor U4664 (N_4664,N_4123,N_4003);
nand U4665 (N_4665,N_4011,N_4335);
nand U4666 (N_4666,N_4110,N_4009);
nand U4667 (N_4667,N_4174,N_4145);
xnor U4668 (N_4668,N_4347,N_4311);
nor U4669 (N_4669,N_4299,N_4310);
or U4670 (N_4670,N_4346,N_4190);
nand U4671 (N_4671,N_4089,N_4020);
and U4672 (N_4672,N_4220,N_4387);
or U4673 (N_4673,N_4044,N_4110);
xor U4674 (N_4674,N_4264,N_4086);
nor U4675 (N_4675,N_4398,N_4340);
or U4676 (N_4676,N_4181,N_4021);
xnor U4677 (N_4677,N_4337,N_4154);
or U4678 (N_4678,N_4071,N_4179);
or U4679 (N_4679,N_4391,N_4132);
nand U4680 (N_4680,N_4104,N_4076);
xor U4681 (N_4681,N_4248,N_4276);
nand U4682 (N_4682,N_4174,N_4327);
or U4683 (N_4683,N_4193,N_4014);
or U4684 (N_4684,N_4067,N_4118);
nor U4685 (N_4685,N_4250,N_4351);
nor U4686 (N_4686,N_4182,N_4015);
and U4687 (N_4687,N_4152,N_4226);
and U4688 (N_4688,N_4295,N_4119);
or U4689 (N_4689,N_4259,N_4172);
nor U4690 (N_4690,N_4112,N_4254);
and U4691 (N_4691,N_4314,N_4261);
nand U4692 (N_4692,N_4253,N_4161);
nand U4693 (N_4693,N_4061,N_4298);
or U4694 (N_4694,N_4128,N_4094);
nand U4695 (N_4695,N_4178,N_4392);
or U4696 (N_4696,N_4257,N_4154);
or U4697 (N_4697,N_4150,N_4039);
and U4698 (N_4698,N_4347,N_4030);
nor U4699 (N_4699,N_4357,N_4291);
nor U4700 (N_4700,N_4168,N_4254);
and U4701 (N_4701,N_4151,N_4248);
nor U4702 (N_4702,N_4261,N_4137);
or U4703 (N_4703,N_4195,N_4028);
xnor U4704 (N_4704,N_4130,N_4088);
nand U4705 (N_4705,N_4321,N_4265);
xnor U4706 (N_4706,N_4365,N_4298);
or U4707 (N_4707,N_4335,N_4137);
and U4708 (N_4708,N_4028,N_4319);
and U4709 (N_4709,N_4162,N_4085);
nor U4710 (N_4710,N_4313,N_4304);
or U4711 (N_4711,N_4191,N_4087);
nand U4712 (N_4712,N_4194,N_4087);
xor U4713 (N_4713,N_4109,N_4191);
and U4714 (N_4714,N_4293,N_4393);
nor U4715 (N_4715,N_4002,N_4277);
nand U4716 (N_4716,N_4280,N_4301);
nand U4717 (N_4717,N_4125,N_4157);
xnor U4718 (N_4718,N_4155,N_4238);
xor U4719 (N_4719,N_4131,N_4263);
nor U4720 (N_4720,N_4368,N_4060);
and U4721 (N_4721,N_4070,N_4184);
and U4722 (N_4722,N_4280,N_4094);
or U4723 (N_4723,N_4052,N_4232);
nand U4724 (N_4724,N_4243,N_4248);
xnor U4725 (N_4725,N_4176,N_4261);
or U4726 (N_4726,N_4218,N_4391);
and U4727 (N_4727,N_4383,N_4117);
nor U4728 (N_4728,N_4372,N_4046);
and U4729 (N_4729,N_4098,N_4048);
or U4730 (N_4730,N_4309,N_4289);
nor U4731 (N_4731,N_4074,N_4375);
or U4732 (N_4732,N_4220,N_4138);
or U4733 (N_4733,N_4022,N_4352);
xnor U4734 (N_4734,N_4243,N_4336);
xor U4735 (N_4735,N_4266,N_4324);
nor U4736 (N_4736,N_4131,N_4074);
nor U4737 (N_4737,N_4364,N_4215);
or U4738 (N_4738,N_4073,N_4235);
xor U4739 (N_4739,N_4067,N_4216);
or U4740 (N_4740,N_4296,N_4205);
and U4741 (N_4741,N_4376,N_4005);
nand U4742 (N_4742,N_4086,N_4076);
or U4743 (N_4743,N_4280,N_4285);
or U4744 (N_4744,N_4037,N_4368);
xnor U4745 (N_4745,N_4360,N_4376);
or U4746 (N_4746,N_4052,N_4136);
and U4747 (N_4747,N_4005,N_4331);
xor U4748 (N_4748,N_4260,N_4100);
xnor U4749 (N_4749,N_4326,N_4031);
xnor U4750 (N_4750,N_4036,N_4067);
xor U4751 (N_4751,N_4208,N_4274);
and U4752 (N_4752,N_4068,N_4186);
or U4753 (N_4753,N_4195,N_4387);
nor U4754 (N_4754,N_4271,N_4249);
xnor U4755 (N_4755,N_4390,N_4301);
nor U4756 (N_4756,N_4236,N_4398);
nor U4757 (N_4757,N_4201,N_4310);
nor U4758 (N_4758,N_4108,N_4188);
nand U4759 (N_4759,N_4121,N_4059);
nand U4760 (N_4760,N_4198,N_4350);
or U4761 (N_4761,N_4028,N_4269);
and U4762 (N_4762,N_4298,N_4271);
nand U4763 (N_4763,N_4187,N_4006);
xnor U4764 (N_4764,N_4359,N_4273);
nor U4765 (N_4765,N_4124,N_4005);
or U4766 (N_4766,N_4221,N_4344);
and U4767 (N_4767,N_4198,N_4259);
and U4768 (N_4768,N_4214,N_4008);
and U4769 (N_4769,N_4052,N_4389);
or U4770 (N_4770,N_4144,N_4320);
nand U4771 (N_4771,N_4266,N_4164);
nand U4772 (N_4772,N_4216,N_4338);
and U4773 (N_4773,N_4380,N_4229);
xor U4774 (N_4774,N_4182,N_4230);
and U4775 (N_4775,N_4027,N_4068);
and U4776 (N_4776,N_4276,N_4022);
xor U4777 (N_4777,N_4386,N_4139);
or U4778 (N_4778,N_4107,N_4206);
xor U4779 (N_4779,N_4176,N_4109);
xor U4780 (N_4780,N_4192,N_4074);
and U4781 (N_4781,N_4027,N_4342);
or U4782 (N_4782,N_4185,N_4020);
nand U4783 (N_4783,N_4336,N_4032);
nand U4784 (N_4784,N_4139,N_4217);
or U4785 (N_4785,N_4190,N_4394);
or U4786 (N_4786,N_4093,N_4201);
xnor U4787 (N_4787,N_4316,N_4337);
nand U4788 (N_4788,N_4377,N_4025);
nand U4789 (N_4789,N_4037,N_4063);
xnor U4790 (N_4790,N_4218,N_4217);
and U4791 (N_4791,N_4373,N_4007);
and U4792 (N_4792,N_4179,N_4043);
or U4793 (N_4793,N_4337,N_4168);
and U4794 (N_4794,N_4135,N_4254);
xor U4795 (N_4795,N_4262,N_4059);
nor U4796 (N_4796,N_4298,N_4257);
nor U4797 (N_4797,N_4308,N_4336);
nor U4798 (N_4798,N_4125,N_4319);
xnor U4799 (N_4799,N_4200,N_4125);
xnor U4800 (N_4800,N_4661,N_4400);
nor U4801 (N_4801,N_4535,N_4500);
or U4802 (N_4802,N_4692,N_4673);
nand U4803 (N_4803,N_4480,N_4577);
xor U4804 (N_4804,N_4620,N_4617);
nand U4805 (N_4805,N_4537,N_4656);
nor U4806 (N_4806,N_4791,N_4531);
or U4807 (N_4807,N_4686,N_4787);
and U4808 (N_4808,N_4514,N_4748);
nor U4809 (N_4809,N_4666,N_4770);
nand U4810 (N_4810,N_4676,N_4754);
xor U4811 (N_4811,N_4483,N_4688);
xnor U4812 (N_4812,N_4516,N_4684);
and U4813 (N_4813,N_4559,N_4543);
or U4814 (N_4814,N_4469,N_4546);
xor U4815 (N_4815,N_4716,N_4722);
and U4816 (N_4816,N_4486,N_4455);
and U4817 (N_4817,N_4721,N_4547);
and U4818 (N_4818,N_4578,N_4653);
or U4819 (N_4819,N_4654,N_4513);
and U4820 (N_4820,N_4752,N_4565);
nor U4821 (N_4821,N_4541,N_4408);
and U4822 (N_4822,N_4439,N_4471);
xor U4823 (N_4823,N_4574,N_4583);
nor U4824 (N_4824,N_4570,N_4689);
xnor U4825 (N_4825,N_4773,N_4639);
xor U4826 (N_4826,N_4587,N_4490);
nand U4827 (N_4827,N_4644,N_4498);
nor U4828 (N_4828,N_4586,N_4781);
nand U4829 (N_4829,N_4517,N_4563);
or U4830 (N_4830,N_4777,N_4709);
xnor U4831 (N_4831,N_4691,N_4718);
or U4832 (N_4832,N_4618,N_4645);
nand U4833 (N_4833,N_4599,N_4790);
nand U4834 (N_4834,N_4562,N_4590);
and U4835 (N_4835,N_4479,N_4706);
or U4836 (N_4836,N_4637,N_4534);
xor U4837 (N_4837,N_4602,N_4726);
and U4838 (N_4838,N_4506,N_4521);
nand U4839 (N_4839,N_4774,N_4433);
and U4840 (N_4840,N_4452,N_4663);
or U4841 (N_4841,N_4621,N_4643);
nor U4842 (N_4842,N_4404,N_4446);
nor U4843 (N_4843,N_4738,N_4609);
nor U4844 (N_4844,N_4613,N_4734);
nand U4845 (N_4845,N_4536,N_4557);
nand U4846 (N_4846,N_4789,N_4667);
nor U4847 (N_4847,N_4509,N_4550);
or U4848 (N_4848,N_4607,N_4788);
nor U4849 (N_4849,N_4711,N_4473);
xnor U4850 (N_4850,N_4730,N_4679);
nand U4851 (N_4851,N_4647,N_4792);
or U4852 (N_4852,N_4527,N_4674);
xor U4853 (N_4853,N_4407,N_4410);
or U4854 (N_4854,N_4717,N_4725);
nor U4855 (N_4855,N_4459,N_4572);
nor U4856 (N_4856,N_4603,N_4489);
nand U4857 (N_4857,N_4705,N_4488);
and U4858 (N_4858,N_4524,N_4727);
nor U4859 (N_4859,N_4427,N_4735);
or U4860 (N_4860,N_4780,N_4438);
and U4861 (N_4861,N_4454,N_4403);
and U4862 (N_4862,N_4551,N_4478);
xor U4863 (N_4863,N_4652,N_4693);
or U4864 (N_4864,N_4704,N_4405);
and U4865 (N_4865,N_4712,N_4542);
and U4866 (N_4866,N_4458,N_4464);
xor U4867 (N_4867,N_4423,N_4659);
or U4868 (N_4868,N_4751,N_4503);
nor U4869 (N_4869,N_4682,N_4675);
nor U4870 (N_4870,N_4462,N_4664);
xor U4871 (N_4871,N_4418,N_4756);
nor U4872 (N_4872,N_4625,N_4669);
and U4873 (N_4873,N_4648,N_4495);
nand U4874 (N_4874,N_4622,N_4635);
nand U4875 (N_4875,N_4651,N_4745);
xnor U4876 (N_4876,N_4591,N_4461);
nand U4877 (N_4877,N_4604,N_4515);
nand U4878 (N_4878,N_4581,N_4614);
xor U4879 (N_4879,N_4786,N_4589);
xnor U4880 (N_4880,N_4782,N_4573);
or U4881 (N_4881,N_4434,N_4494);
nor U4882 (N_4882,N_4470,N_4508);
or U4883 (N_4883,N_4576,N_4561);
nor U4884 (N_4884,N_4525,N_4594);
nand U4885 (N_4885,N_4548,N_4641);
xnor U4886 (N_4886,N_4595,N_4799);
nand U4887 (N_4887,N_4448,N_4475);
and U4888 (N_4888,N_4698,N_4678);
or U4889 (N_4889,N_4593,N_4680);
xor U4890 (N_4890,N_4632,N_4526);
nand U4891 (N_4891,N_4624,N_4768);
xor U4892 (N_4892,N_4504,N_4747);
or U4893 (N_4893,N_4700,N_4539);
or U4894 (N_4894,N_4755,N_4511);
xor U4895 (N_4895,N_4775,N_4665);
nor U4896 (N_4896,N_4568,N_4660);
or U4897 (N_4897,N_4638,N_4450);
nand U4898 (N_4898,N_4797,N_4715);
nand U4899 (N_4899,N_4484,N_4736);
and U4900 (N_4900,N_4796,N_4558);
nand U4901 (N_4901,N_4762,N_4611);
and U4902 (N_4902,N_4491,N_4630);
nand U4903 (N_4903,N_4646,N_4487);
and U4904 (N_4904,N_4420,N_4720);
or U4905 (N_4905,N_4507,N_4662);
xor U4906 (N_4906,N_4642,N_4552);
and U4907 (N_4907,N_4695,N_4671);
and U4908 (N_4908,N_4690,N_4428);
or U4909 (N_4909,N_4406,N_4477);
and U4910 (N_4910,N_4465,N_4556);
xor U4911 (N_4911,N_4426,N_4633);
nor U4912 (N_4912,N_4655,N_4566);
nand U4913 (N_4913,N_4744,N_4723);
and U4914 (N_4914,N_4401,N_4794);
nand U4915 (N_4915,N_4584,N_4657);
or U4916 (N_4916,N_4615,N_4746);
nand U4917 (N_4917,N_4766,N_4442);
nor U4918 (N_4918,N_4415,N_4417);
and U4919 (N_4919,N_4592,N_4757);
or U4920 (N_4920,N_4710,N_4650);
xnor U4921 (N_4921,N_4636,N_4419);
nor U4922 (N_4922,N_4598,N_4416);
or U4923 (N_4923,N_4554,N_4668);
and U4924 (N_4924,N_4749,N_4610);
nor U4925 (N_4925,N_4596,N_4430);
nand U4926 (N_4926,N_4619,N_4560);
nor U4927 (N_4927,N_4532,N_4545);
nor U4928 (N_4928,N_4697,N_4585);
nand U4929 (N_4929,N_4658,N_4764);
and U4930 (N_4930,N_4449,N_4582);
or U4931 (N_4931,N_4694,N_4441);
and U4932 (N_4932,N_4743,N_4606);
nand U4933 (N_4933,N_4413,N_4776);
xnor U4934 (N_4934,N_4579,N_4758);
and U4935 (N_4935,N_4771,N_4778);
or U4936 (N_4936,N_4785,N_4729);
and U4937 (N_4937,N_4699,N_4608);
nor U4938 (N_4938,N_4409,N_4519);
and U4939 (N_4939,N_4798,N_4402);
or U4940 (N_4940,N_4476,N_4685);
or U4941 (N_4941,N_4580,N_4493);
and U4942 (N_4942,N_4518,N_4451);
nand U4943 (N_4943,N_4424,N_4701);
or U4944 (N_4944,N_4444,N_4763);
nor U4945 (N_4945,N_4767,N_4411);
xor U4946 (N_4946,N_4421,N_4540);
or U4947 (N_4947,N_4623,N_4567);
xnor U4948 (N_4948,N_4772,N_4728);
nand U4949 (N_4949,N_4670,N_4779);
or U4950 (N_4950,N_4457,N_4485);
or U4951 (N_4951,N_4629,N_4522);
or U4952 (N_4952,N_4425,N_4520);
xor U4953 (N_4953,N_4683,N_4528);
and U4954 (N_4954,N_4708,N_4492);
nand U4955 (N_4955,N_4553,N_4482);
xnor U4956 (N_4956,N_4443,N_4497);
nor U4957 (N_4957,N_4714,N_4703);
xnor U4958 (N_4958,N_4634,N_4436);
xor U4959 (N_4959,N_4737,N_4742);
and U4960 (N_4960,N_4719,N_4765);
xor U4961 (N_4961,N_4505,N_4523);
and U4962 (N_4962,N_4753,N_4440);
nor U4963 (N_4963,N_4741,N_4456);
and U4964 (N_4964,N_4733,N_4453);
nor U4965 (N_4965,N_4713,N_4571);
xnor U4966 (N_4966,N_4575,N_4628);
nor U4967 (N_4967,N_4696,N_4588);
nor U4968 (N_4968,N_4422,N_4463);
or U4969 (N_4969,N_4672,N_4414);
xor U4970 (N_4970,N_4468,N_4732);
and U4971 (N_4971,N_4501,N_4445);
nor U4972 (N_4972,N_4499,N_4512);
nand U4973 (N_4973,N_4481,N_4597);
or U4974 (N_4974,N_4460,N_4739);
xnor U4975 (N_4975,N_4472,N_4564);
or U4976 (N_4976,N_4412,N_4533);
or U4977 (N_4977,N_4496,N_4544);
nand U4978 (N_4978,N_4759,N_4760);
nor U4979 (N_4979,N_4761,N_4784);
nand U4980 (N_4980,N_4769,N_4681);
nand U4981 (N_4981,N_4601,N_4626);
and U4982 (N_4982,N_4447,N_4467);
or U4983 (N_4983,N_4549,N_4750);
or U4984 (N_4984,N_4783,N_4432);
nand U4985 (N_4985,N_4795,N_4502);
xor U4986 (N_4986,N_4435,N_4793);
xnor U4987 (N_4987,N_4731,N_4740);
nor U4988 (N_4988,N_4724,N_4431);
and U4989 (N_4989,N_4510,N_4640);
or U4990 (N_4990,N_4429,N_4612);
and U4991 (N_4991,N_4605,N_4600);
xnor U4992 (N_4992,N_4529,N_4530);
xor U4993 (N_4993,N_4677,N_4649);
and U4994 (N_4994,N_4627,N_4707);
nor U4995 (N_4995,N_4569,N_4555);
xor U4996 (N_4996,N_4687,N_4474);
or U4997 (N_4997,N_4702,N_4437);
and U4998 (N_4998,N_4538,N_4466);
nand U4999 (N_4999,N_4631,N_4616);
xor U5000 (N_5000,N_4661,N_4468);
or U5001 (N_5001,N_4585,N_4465);
nand U5002 (N_5002,N_4584,N_4416);
or U5003 (N_5003,N_4404,N_4778);
and U5004 (N_5004,N_4724,N_4641);
and U5005 (N_5005,N_4571,N_4724);
nor U5006 (N_5006,N_4718,N_4537);
or U5007 (N_5007,N_4586,N_4708);
xnor U5008 (N_5008,N_4498,N_4621);
xnor U5009 (N_5009,N_4762,N_4480);
xor U5010 (N_5010,N_4567,N_4494);
xor U5011 (N_5011,N_4446,N_4458);
nor U5012 (N_5012,N_4553,N_4461);
or U5013 (N_5013,N_4668,N_4420);
nand U5014 (N_5014,N_4462,N_4706);
xor U5015 (N_5015,N_4508,N_4612);
or U5016 (N_5016,N_4486,N_4570);
or U5017 (N_5017,N_4545,N_4723);
or U5018 (N_5018,N_4584,N_4410);
and U5019 (N_5019,N_4794,N_4569);
and U5020 (N_5020,N_4416,N_4406);
and U5021 (N_5021,N_4741,N_4521);
nand U5022 (N_5022,N_4441,N_4781);
or U5023 (N_5023,N_4514,N_4589);
and U5024 (N_5024,N_4406,N_4660);
xor U5025 (N_5025,N_4698,N_4567);
or U5026 (N_5026,N_4491,N_4647);
xor U5027 (N_5027,N_4637,N_4612);
or U5028 (N_5028,N_4433,N_4645);
and U5029 (N_5029,N_4786,N_4764);
xnor U5030 (N_5030,N_4689,N_4762);
or U5031 (N_5031,N_4558,N_4414);
nor U5032 (N_5032,N_4780,N_4762);
nor U5033 (N_5033,N_4559,N_4490);
and U5034 (N_5034,N_4427,N_4716);
nand U5035 (N_5035,N_4482,N_4738);
xnor U5036 (N_5036,N_4656,N_4464);
or U5037 (N_5037,N_4545,N_4743);
or U5038 (N_5038,N_4581,N_4554);
xnor U5039 (N_5039,N_4432,N_4505);
or U5040 (N_5040,N_4770,N_4537);
nor U5041 (N_5041,N_4547,N_4433);
or U5042 (N_5042,N_4652,N_4644);
or U5043 (N_5043,N_4762,N_4520);
and U5044 (N_5044,N_4616,N_4508);
nand U5045 (N_5045,N_4576,N_4616);
nand U5046 (N_5046,N_4427,N_4585);
nor U5047 (N_5047,N_4766,N_4492);
or U5048 (N_5048,N_4585,N_4495);
xor U5049 (N_5049,N_4462,N_4602);
nor U5050 (N_5050,N_4696,N_4673);
nor U5051 (N_5051,N_4780,N_4590);
or U5052 (N_5052,N_4410,N_4590);
nor U5053 (N_5053,N_4506,N_4551);
nor U5054 (N_5054,N_4497,N_4732);
nor U5055 (N_5055,N_4645,N_4590);
and U5056 (N_5056,N_4716,N_4551);
and U5057 (N_5057,N_4490,N_4600);
nor U5058 (N_5058,N_4668,N_4721);
and U5059 (N_5059,N_4566,N_4755);
xor U5060 (N_5060,N_4797,N_4595);
xnor U5061 (N_5061,N_4508,N_4623);
nor U5062 (N_5062,N_4772,N_4400);
nor U5063 (N_5063,N_4751,N_4685);
and U5064 (N_5064,N_4651,N_4557);
or U5065 (N_5065,N_4598,N_4655);
and U5066 (N_5066,N_4555,N_4614);
or U5067 (N_5067,N_4546,N_4607);
nand U5068 (N_5068,N_4525,N_4429);
xnor U5069 (N_5069,N_4659,N_4517);
or U5070 (N_5070,N_4776,N_4667);
nor U5071 (N_5071,N_4437,N_4430);
nand U5072 (N_5072,N_4443,N_4561);
and U5073 (N_5073,N_4720,N_4482);
and U5074 (N_5074,N_4517,N_4730);
nor U5075 (N_5075,N_4672,N_4513);
and U5076 (N_5076,N_4567,N_4535);
nand U5077 (N_5077,N_4535,N_4498);
xor U5078 (N_5078,N_4750,N_4738);
and U5079 (N_5079,N_4778,N_4529);
nor U5080 (N_5080,N_4672,N_4784);
or U5081 (N_5081,N_4558,N_4574);
or U5082 (N_5082,N_4688,N_4647);
and U5083 (N_5083,N_4497,N_4558);
xor U5084 (N_5084,N_4438,N_4474);
nor U5085 (N_5085,N_4545,N_4680);
and U5086 (N_5086,N_4799,N_4797);
nand U5087 (N_5087,N_4744,N_4682);
and U5088 (N_5088,N_4551,N_4793);
and U5089 (N_5089,N_4413,N_4708);
xnor U5090 (N_5090,N_4735,N_4785);
xnor U5091 (N_5091,N_4411,N_4725);
nand U5092 (N_5092,N_4710,N_4757);
nand U5093 (N_5093,N_4449,N_4785);
or U5094 (N_5094,N_4731,N_4637);
or U5095 (N_5095,N_4685,N_4740);
and U5096 (N_5096,N_4668,N_4534);
or U5097 (N_5097,N_4467,N_4566);
and U5098 (N_5098,N_4544,N_4611);
nor U5099 (N_5099,N_4525,N_4418);
nand U5100 (N_5100,N_4759,N_4705);
and U5101 (N_5101,N_4729,N_4697);
and U5102 (N_5102,N_4667,N_4609);
and U5103 (N_5103,N_4411,N_4670);
or U5104 (N_5104,N_4704,N_4606);
and U5105 (N_5105,N_4479,N_4471);
and U5106 (N_5106,N_4789,N_4499);
or U5107 (N_5107,N_4433,N_4527);
nor U5108 (N_5108,N_4549,N_4475);
xor U5109 (N_5109,N_4660,N_4586);
nor U5110 (N_5110,N_4700,N_4552);
xnor U5111 (N_5111,N_4774,N_4435);
nand U5112 (N_5112,N_4756,N_4451);
nand U5113 (N_5113,N_4642,N_4431);
and U5114 (N_5114,N_4402,N_4648);
nor U5115 (N_5115,N_4647,N_4789);
and U5116 (N_5116,N_4582,N_4543);
nor U5117 (N_5117,N_4755,N_4580);
and U5118 (N_5118,N_4526,N_4687);
and U5119 (N_5119,N_4499,N_4430);
nor U5120 (N_5120,N_4628,N_4509);
and U5121 (N_5121,N_4455,N_4439);
nand U5122 (N_5122,N_4452,N_4425);
and U5123 (N_5123,N_4474,N_4655);
or U5124 (N_5124,N_4589,N_4542);
nand U5125 (N_5125,N_4735,N_4606);
nor U5126 (N_5126,N_4630,N_4721);
nor U5127 (N_5127,N_4409,N_4556);
nor U5128 (N_5128,N_4577,N_4600);
nor U5129 (N_5129,N_4648,N_4567);
or U5130 (N_5130,N_4684,N_4415);
and U5131 (N_5131,N_4568,N_4424);
xnor U5132 (N_5132,N_4734,N_4729);
nand U5133 (N_5133,N_4713,N_4530);
or U5134 (N_5134,N_4558,N_4509);
or U5135 (N_5135,N_4789,N_4606);
nand U5136 (N_5136,N_4678,N_4761);
xnor U5137 (N_5137,N_4798,N_4562);
and U5138 (N_5138,N_4586,N_4644);
xor U5139 (N_5139,N_4579,N_4780);
and U5140 (N_5140,N_4651,N_4714);
xor U5141 (N_5141,N_4563,N_4499);
or U5142 (N_5142,N_4456,N_4433);
nand U5143 (N_5143,N_4719,N_4588);
or U5144 (N_5144,N_4658,N_4449);
and U5145 (N_5145,N_4545,N_4584);
xor U5146 (N_5146,N_4527,N_4675);
xnor U5147 (N_5147,N_4591,N_4471);
and U5148 (N_5148,N_4662,N_4677);
and U5149 (N_5149,N_4749,N_4418);
xnor U5150 (N_5150,N_4640,N_4427);
nand U5151 (N_5151,N_4755,N_4564);
nor U5152 (N_5152,N_4651,N_4782);
and U5153 (N_5153,N_4731,N_4649);
and U5154 (N_5154,N_4757,N_4443);
or U5155 (N_5155,N_4482,N_4717);
or U5156 (N_5156,N_4695,N_4546);
xnor U5157 (N_5157,N_4665,N_4529);
and U5158 (N_5158,N_4659,N_4696);
xnor U5159 (N_5159,N_4607,N_4682);
xnor U5160 (N_5160,N_4742,N_4720);
and U5161 (N_5161,N_4611,N_4753);
nand U5162 (N_5162,N_4657,N_4452);
xnor U5163 (N_5163,N_4415,N_4554);
nor U5164 (N_5164,N_4416,N_4508);
nand U5165 (N_5165,N_4538,N_4463);
and U5166 (N_5166,N_4656,N_4610);
nor U5167 (N_5167,N_4407,N_4772);
and U5168 (N_5168,N_4732,N_4428);
xnor U5169 (N_5169,N_4708,N_4719);
or U5170 (N_5170,N_4718,N_4769);
or U5171 (N_5171,N_4511,N_4498);
nor U5172 (N_5172,N_4779,N_4753);
or U5173 (N_5173,N_4769,N_4784);
nor U5174 (N_5174,N_4781,N_4515);
and U5175 (N_5175,N_4613,N_4578);
or U5176 (N_5176,N_4419,N_4544);
nor U5177 (N_5177,N_4553,N_4563);
and U5178 (N_5178,N_4711,N_4507);
nand U5179 (N_5179,N_4600,N_4437);
and U5180 (N_5180,N_4580,N_4645);
xnor U5181 (N_5181,N_4491,N_4553);
nand U5182 (N_5182,N_4465,N_4408);
nor U5183 (N_5183,N_4605,N_4615);
and U5184 (N_5184,N_4645,N_4620);
and U5185 (N_5185,N_4782,N_4619);
xnor U5186 (N_5186,N_4554,N_4708);
nand U5187 (N_5187,N_4445,N_4719);
xnor U5188 (N_5188,N_4669,N_4520);
nor U5189 (N_5189,N_4403,N_4446);
or U5190 (N_5190,N_4452,N_4640);
xor U5191 (N_5191,N_4619,N_4786);
nor U5192 (N_5192,N_4639,N_4721);
and U5193 (N_5193,N_4685,N_4688);
or U5194 (N_5194,N_4440,N_4607);
xnor U5195 (N_5195,N_4403,N_4630);
nand U5196 (N_5196,N_4561,N_4559);
xnor U5197 (N_5197,N_4722,N_4622);
nor U5198 (N_5198,N_4411,N_4553);
and U5199 (N_5199,N_4644,N_4545);
nor U5200 (N_5200,N_5064,N_5159);
nor U5201 (N_5201,N_4863,N_5176);
xor U5202 (N_5202,N_4965,N_4937);
nand U5203 (N_5203,N_4885,N_4829);
xnor U5204 (N_5204,N_4903,N_4913);
nand U5205 (N_5205,N_4822,N_4897);
or U5206 (N_5206,N_5073,N_5184);
or U5207 (N_5207,N_5095,N_5045);
nand U5208 (N_5208,N_4874,N_4813);
xnor U5209 (N_5209,N_5134,N_5167);
nor U5210 (N_5210,N_5088,N_5149);
or U5211 (N_5211,N_4986,N_5032);
xor U5212 (N_5212,N_4925,N_5086);
xor U5213 (N_5213,N_5166,N_5078);
xor U5214 (N_5214,N_4981,N_4988);
or U5215 (N_5215,N_5070,N_4892);
and U5216 (N_5216,N_4815,N_5007);
nor U5217 (N_5217,N_5173,N_4875);
xnor U5218 (N_5218,N_5116,N_4802);
xnor U5219 (N_5219,N_4873,N_5139);
nor U5220 (N_5220,N_4915,N_5191);
nor U5221 (N_5221,N_5113,N_5006);
nor U5222 (N_5222,N_5172,N_4804);
or U5223 (N_5223,N_5024,N_4984);
xnor U5224 (N_5224,N_5158,N_4806);
nand U5225 (N_5225,N_4890,N_4834);
nand U5226 (N_5226,N_5089,N_5133);
nand U5227 (N_5227,N_4974,N_5187);
or U5228 (N_5228,N_5147,N_5143);
and U5229 (N_5229,N_5084,N_4831);
xnor U5230 (N_5230,N_4976,N_5196);
xor U5231 (N_5231,N_4816,N_5194);
or U5232 (N_5232,N_4911,N_4868);
nor U5233 (N_5233,N_5115,N_5002);
nor U5234 (N_5234,N_5192,N_5059);
nor U5235 (N_5235,N_4920,N_4879);
nor U5236 (N_5236,N_4844,N_5021);
nand U5237 (N_5237,N_4803,N_4832);
nor U5238 (N_5238,N_5195,N_5055);
and U5239 (N_5239,N_4809,N_4852);
and U5240 (N_5240,N_4961,N_5018);
xor U5241 (N_5241,N_4871,N_5010);
nand U5242 (N_5242,N_5051,N_4870);
or U5243 (N_5243,N_5156,N_4837);
or U5244 (N_5244,N_5044,N_4891);
nor U5245 (N_5245,N_4881,N_5092);
and U5246 (N_5246,N_4973,N_4898);
xnor U5247 (N_5247,N_4939,N_4833);
or U5248 (N_5248,N_4956,N_5154);
xnor U5249 (N_5249,N_5065,N_4884);
xor U5250 (N_5250,N_5123,N_4841);
and U5251 (N_5251,N_5058,N_5129);
nand U5252 (N_5252,N_4880,N_5015);
or U5253 (N_5253,N_5011,N_4906);
nor U5254 (N_5254,N_4995,N_5128);
and U5255 (N_5255,N_4845,N_5074);
and U5256 (N_5256,N_5008,N_5110);
nand U5257 (N_5257,N_5186,N_4894);
or U5258 (N_5258,N_5132,N_4846);
or U5259 (N_5259,N_4872,N_4889);
nand U5260 (N_5260,N_5124,N_4955);
xor U5261 (N_5261,N_5103,N_5035);
nand U5262 (N_5262,N_4825,N_4991);
xnor U5263 (N_5263,N_5081,N_5020);
nor U5264 (N_5264,N_5041,N_5104);
or U5265 (N_5265,N_4824,N_5190);
nor U5266 (N_5266,N_4912,N_5109);
or U5267 (N_5267,N_4975,N_5130);
and U5268 (N_5268,N_5049,N_5171);
nand U5269 (N_5269,N_5122,N_4848);
nor U5270 (N_5270,N_4967,N_4946);
nor U5271 (N_5271,N_4923,N_4908);
and U5272 (N_5272,N_4882,N_5183);
nor U5273 (N_5273,N_4859,N_4836);
or U5274 (N_5274,N_5025,N_4944);
nand U5275 (N_5275,N_4926,N_5004);
nand U5276 (N_5276,N_4977,N_4985);
xnor U5277 (N_5277,N_4817,N_4993);
or U5278 (N_5278,N_4971,N_4917);
or U5279 (N_5279,N_5189,N_5105);
xnor U5280 (N_5280,N_4933,N_4962);
or U5281 (N_5281,N_4867,N_4919);
nor U5282 (N_5282,N_5131,N_5097);
nand U5283 (N_5283,N_4930,N_4830);
xor U5284 (N_5284,N_5151,N_5188);
or U5285 (N_5285,N_5162,N_4843);
or U5286 (N_5286,N_4948,N_5034);
or U5287 (N_5287,N_4929,N_4945);
or U5288 (N_5288,N_5180,N_4969);
xor U5289 (N_5289,N_4978,N_4847);
nor U5290 (N_5290,N_5111,N_4954);
nor U5291 (N_5291,N_4861,N_5168);
xnor U5292 (N_5292,N_5150,N_4805);
nand U5293 (N_5293,N_5135,N_4998);
nand U5294 (N_5294,N_4900,N_4916);
or U5295 (N_5295,N_4992,N_5155);
xor U5296 (N_5296,N_5146,N_5069);
xnor U5297 (N_5297,N_4850,N_5157);
xor U5298 (N_5298,N_5031,N_4950);
nand U5299 (N_5299,N_4990,N_4869);
nand U5300 (N_5300,N_4996,N_5145);
nand U5301 (N_5301,N_4957,N_4932);
or U5302 (N_5302,N_4970,N_4949);
or U5303 (N_5303,N_5026,N_5057);
and U5304 (N_5304,N_4936,N_5164);
nand U5305 (N_5305,N_5077,N_5013);
or U5306 (N_5306,N_4994,N_5096);
or U5307 (N_5307,N_4959,N_4800);
and U5308 (N_5308,N_5062,N_4819);
or U5309 (N_5309,N_4856,N_4952);
or U5310 (N_5310,N_5193,N_4812);
nand U5311 (N_5311,N_4828,N_5056);
or U5312 (N_5312,N_4857,N_4983);
or U5313 (N_5313,N_5170,N_4835);
xnor U5314 (N_5314,N_5136,N_5100);
xnor U5315 (N_5315,N_4943,N_4940);
and U5316 (N_5316,N_5120,N_5048);
or U5317 (N_5317,N_5152,N_4877);
or U5318 (N_5318,N_4826,N_4855);
nand U5319 (N_5319,N_4941,N_4927);
xnor U5320 (N_5320,N_4960,N_4909);
nor U5321 (N_5321,N_5112,N_5165);
nand U5322 (N_5322,N_5185,N_5108);
nand U5323 (N_5323,N_5079,N_5153);
and U5324 (N_5324,N_5005,N_5001);
nor U5325 (N_5325,N_4921,N_5102);
nand U5326 (N_5326,N_5117,N_5175);
or U5327 (N_5327,N_4910,N_4887);
and U5328 (N_5328,N_5101,N_5029);
and U5329 (N_5329,N_5037,N_5106);
nor U5330 (N_5330,N_5082,N_4934);
nand U5331 (N_5331,N_4808,N_5038);
and U5332 (N_5332,N_4997,N_5163);
nand U5333 (N_5333,N_5148,N_5090);
nor U5334 (N_5334,N_4807,N_5125);
xnor U5335 (N_5335,N_5043,N_4935);
and U5336 (N_5336,N_5030,N_5174);
nor U5337 (N_5337,N_4901,N_4858);
nand U5338 (N_5338,N_5071,N_5076);
nor U5339 (N_5339,N_4951,N_5138);
and U5340 (N_5340,N_4902,N_5072);
nor U5341 (N_5341,N_4982,N_4914);
or U5342 (N_5342,N_4905,N_5039);
nand U5343 (N_5343,N_4989,N_5068);
or U5344 (N_5344,N_5000,N_4922);
nand U5345 (N_5345,N_4842,N_5107);
nor U5346 (N_5346,N_4814,N_5182);
nand U5347 (N_5347,N_4853,N_5142);
nor U5348 (N_5348,N_5141,N_5053);
nor U5349 (N_5349,N_5161,N_5023);
or U5350 (N_5350,N_5197,N_4883);
and U5351 (N_5351,N_5098,N_4864);
or U5352 (N_5352,N_5014,N_4980);
and U5353 (N_5353,N_5169,N_4999);
nand U5354 (N_5354,N_4823,N_5119);
xor U5355 (N_5355,N_5060,N_5027);
and U5356 (N_5356,N_4953,N_4876);
nor U5357 (N_5357,N_4979,N_5199);
xnor U5358 (N_5358,N_4818,N_4849);
nand U5359 (N_5359,N_5160,N_5003);
and U5360 (N_5360,N_4928,N_5040);
nor U5361 (N_5361,N_5046,N_4963);
nor U5362 (N_5362,N_5093,N_5019);
or U5363 (N_5363,N_5198,N_5091);
xnor U5364 (N_5364,N_4968,N_4931);
or U5365 (N_5365,N_5137,N_4851);
nor U5366 (N_5366,N_4972,N_5181);
xor U5367 (N_5367,N_4860,N_4821);
and U5368 (N_5368,N_5118,N_5179);
xnor U5369 (N_5369,N_5061,N_5126);
or U5370 (N_5370,N_5022,N_5085);
and U5371 (N_5371,N_5052,N_5094);
and U5372 (N_5372,N_4888,N_4896);
nor U5373 (N_5373,N_5099,N_4862);
and U5374 (N_5374,N_4942,N_4907);
nor U5375 (N_5375,N_5012,N_5036);
and U5376 (N_5376,N_4895,N_4801);
xor U5377 (N_5377,N_4839,N_5066);
nor U5378 (N_5378,N_4964,N_4827);
nor U5379 (N_5379,N_4966,N_4810);
and U5380 (N_5380,N_4854,N_5083);
nand U5381 (N_5381,N_5177,N_5067);
and U5382 (N_5382,N_5114,N_5033);
nand U5383 (N_5383,N_5050,N_4811);
or U5384 (N_5384,N_5063,N_4865);
xor U5385 (N_5385,N_4878,N_5009);
or U5386 (N_5386,N_5047,N_4904);
and U5387 (N_5387,N_5042,N_5017);
nor U5388 (N_5388,N_5080,N_4958);
or U5389 (N_5389,N_4918,N_4886);
and U5390 (N_5390,N_5087,N_4838);
xor U5391 (N_5391,N_4820,N_5144);
or U5392 (N_5392,N_5140,N_5127);
nand U5393 (N_5393,N_4987,N_5121);
nand U5394 (N_5394,N_4947,N_4866);
and U5395 (N_5395,N_5016,N_5178);
nand U5396 (N_5396,N_4893,N_4938);
nor U5397 (N_5397,N_4840,N_5075);
nor U5398 (N_5398,N_5028,N_4924);
and U5399 (N_5399,N_5054,N_4899);
nor U5400 (N_5400,N_5004,N_4949);
nor U5401 (N_5401,N_4805,N_5122);
or U5402 (N_5402,N_4966,N_4878);
and U5403 (N_5403,N_4958,N_5151);
nand U5404 (N_5404,N_4918,N_5167);
and U5405 (N_5405,N_5060,N_5070);
xor U5406 (N_5406,N_5105,N_4906);
nor U5407 (N_5407,N_5019,N_5046);
nor U5408 (N_5408,N_4859,N_5182);
nand U5409 (N_5409,N_5133,N_5076);
or U5410 (N_5410,N_4986,N_5116);
nor U5411 (N_5411,N_4823,N_5028);
xor U5412 (N_5412,N_4964,N_4801);
nor U5413 (N_5413,N_4966,N_5017);
nor U5414 (N_5414,N_5147,N_4860);
nor U5415 (N_5415,N_4880,N_5189);
nor U5416 (N_5416,N_4855,N_4829);
and U5417 (N_5417,N_5156,N_5027);
nor U5418 (N_5418,N_4992,N_5021);
nand U5419 (N_5419,N_4948,N_4879);
nor U5420 (N_5420,N_5074,N_4917);
or U5421 (N_5421,N_4853,N_4927);
nor U5422 (N_5422,N_5165,N_4974);
nor U5423 (N_5423,N_5103,N_4923);
nand U5424 (N_5424,N_5051,N_5118);
and U5425 (N_5425,N_5084,N_5151);
xnor U5426 (N_5426,N_5035,N_4894);
and U5427 (N_5427,N_5166,N_5098);
or U5428 (N_5428,N_5024,N_4914);
or U5429 (N_5429,N_4942,N_5042);
nor U5430 (N_5430,N_5046,N_4934);
and U5431 (N_5431,N_4932,N_5034);
nor U5432 (N_5432,N_5117,N_5001);
or U5433 (N_5433,N_4891,N_5074);
nor U5434 (N_5434,N_5151,N_5144);
xnor U5435 (N_5435,N_5157,N_5171);
and U5436 (N_5436,N_5074,N_4910);
nor U5437 (N_5437,N_4907,N_5107);
nor U5438 (N_5438,N_4912,N_5110);
and U5439 (N_5439,N_4915,N_5067);
and U5440 (N_5440,N_5182,N_5030);
xnor U5441 (N_5441,N_5142,N_4894);
xnor U5442 (N_5442,N_4987,N_5128);
xnor U5443 (N_5443,N_5061,N_4985);
or U5444 (N_5444,N_4821,N_4829);
and U5445 (N_5445,N_5199,N_4879);
nor U5446 (N_5446,N_5112,N_5182);
nand U5447 (N_5447,N_5128,N_4828);
nand U5448 (N_5448,N_4947,N_5169);
nor U5449 (N_5449,N_4804,N_5090);
nor U5450 (N_5450,N_4896,N_4886);
and U5451 (N_5451,N_5024,N_5001);
nand U5452 (N_5452,N_5184,N_5150);
nor U5453 (N_5453,N_5104,N_5063);
and U5454 (N_5454,N_4963,N_5143);
xnor U5455 (N_5455,N_5016,N_5185);
and U5456 (N_5456,N_4800,N_5039);
nand U5457 (N_5457,N_4923,N_5028);
nand U5458 (N_5458,N_4844,N_4881);
and U5459 (N_5459,N_4906,N_4905);
nor U5460 (N_5460,N_4800,N_4862);
and U5461 (N_5461,N_5169,N_4910);
and U5462 (N_5462,N_4833,N_5007);
or U5463 (N_5463,N_4854,N_5008);
nand U5464 (N_5464,N_4944,N_5153);
or U5465 (N_5465,N_5048,N_4942);
and U5466 (N_5466,N_5075,N_4849);
xnor U5467 (N_5467,N_5147,N_5011);
xnor U5468 (N_5468,N_4898,N_4963);
nand U5469 (N_5469,N_5115,N_5051);
and U5470 (N_5470,N_4941,N_5185);
nand U5471 (N_5471,N_4959,N_5111);
and U5472 (N_5472,N_5006,N_4986);
xor U5473 (N_5473,N_4858,N_4808);
nor U5474 (N_5474,N_5140,N_5039);
nand U5475 (N_5475,N_4939,N_5072);
and U5476 (N_5476,N_4818,N_4816);
xnor U5477 (N_5477,N_5001,N_4960);
nor U5478 (N_5478,N_5186,N_4945);
nor U5479 (N_5479,N_4825,N_4952);
nand U5480 (N_5480,N_5060,N_5128);
and U5481 (N_5481,N_4806,N_5019);
nand U5482 (N_5482,N_4919,N_4986);
nor U5483 (N_5483,N_5134,N_4806);
or U5484 (N_5484,N_4867,N_5004);
xor U5485 (N_5485,N_4892,N_5107);
or U5486 (N_5486,N_4802,N_5022);
and U5487 (N_5487,N_5070,N_5170);
or U5488 (N_5488,N_5045,N_5190);
nand U5489 (N_5489,N_5095,N_4956);
and U5490 (N_5490,N_4917,N_5156);
nor U5491 (N_5491,N_4831,N_4940);
or U5492 (N_5492,N_4955,N_5119);
nor U5493 (N_5493,N_5182,N_5009);
nand U5494 (N_5494,N_4824,N_5145);
nor U5495 (N_5495,N_4883,N_5108);
nor U5496 (N_5496,N_4941,N_4969);
nand U5497 (N_5497,N_5066,N_5028);
and U5498 (N_5498,N_5188,N_5042);
nand U5499 (N_5499,N_4867,N_4856);
xor U5500 (N_5500,N_5020,N_4949);
nor U5501 (N_5501,N_5016,N_4954);
xor U5502 (N_5502,N_5047,N_4846);
xor U5503 (N_5503,N_4855,N_4945);
nor U5504 (N_5504,N_4808,N_4992);
nor U5505 (N_5505,N_4955,N_4951);
nor U5506 (N_5506,N_4941,N_4973);
nor U5507 (N_5507,N_4865,N_4880);
nor U5508 (N_5508,N_4885,N_5142);
and U5509 (N_5509,N_5049,N_5063);
and U5510 (N_5510,N_5016,N_4918);
nor U5511 (N_5511,N_4840,N_5124);
or U5512 (N_5512,N_4951,N_5140);
and U5513 (N_5513,N_5026,N_5102);
nand U5514 (N_5514,N_5085,N_5079);
xor U5515 (N_5515,N_4965,N_4988);
nand U5516 (N_5516,N_4998,N_5122);
nor U5517 (N_5517,N_4961,N_5046);
or U5518 (N_5518,N_5110,N_4872);
xor U5519 (N_5519,N_4898,N_5019);
nor U5520 (N_5520,N_4914,N_4945);
nor U5521 (N_5521,N_5077,N_5005);
or U5522 (N_5522,N_5145,N_4817);
or U5523 (N_5523,N_5106,N_5132);
nor U5524 (N_5524,N_4961,N_4826);
nand U5525 (N_5525,N_4924,N_5007);
nand U5526 (N_5526,N_4949,N_5014);
and U5527 (N_5527,N_5152,N_4929);
and U5528 (N_5528,N_4914,N_4980);
nand U5529 (N_5529,N_4863,N_4862);
or U5530 (N_5530,N_4962,N_5037);
and U5531 (N_5531,N_5186,N_5161);
xnor U5532 (N_5532,N_5085,N_4937);
and U5533 (N_5533,N_4872,N_5195);
and U5534 (N_5534,N_5188,N_5085);
or U5535 (N_5535,N_4852,N_5163);
or U5536 (N_5536,N_5049,N_4891);
or U5537 (N_5537,N_4975,N_5139);
xor U5538 (N_5538,N_4904,N_5173);
nor U5539 (N_5539,N_4984,N_4994);
xor U5540 (N_5540,N_5180,N_4945);
nor U5541 (N_5541,N_5131,N_4942);
xor U5542 (N_5542,N_4918,N_4900);
and U5543 (N_5543,N_4819,N_4859);
nor U5544 (N_5544,N_4994,N_4871);
nor U5545 (N_5545,N_5091,N_4987);
nor U5546 (N_5546,N_5064,N_4804);
and U5547 (N_5547,N_5173,N_4922);
nand U5548 (N_5548,N_5178,N_4840);
and U5549 (N_5549,N_4839,N_5172);
nand U5550 (N_5550,N_5149,N_5137);
nor U5551 (N_5551,N_5023,N_5154);
nand U5552 (N_5552,N_4989,N_4920);
nor U5553 (N_5553,N_4951,N_5028);
nor U5554 (N_5554,N_4925,N_4814);
or U5555 (N_5555,N_4974,N_4955);
and U5556 (N_5556,N_4968,N_5047);
nor U5557 (N_5557,N_5199,N_4947);
xor U5558 (N_5558,N_4922,N_4961);
nand U5559 (N_5559,N_4834,N_5008);
or U5560 (N_5560,N_5110,N_4926);
or U5561 (N_5561,N_4976,N_4965);
nand U5562 (N_5562,N_4913,N_4935);
xnor U5563 (N_5563,N_5023,N_4979);
xnor U5564 (N_5564,N_4899,N_4952);
nand U5565 (N_5565,N_4907,N_4971);
xnor U5566 (N_5566,N_4976,N_5080);
or U5567 (N_5567,N_5175,N_5104);
and U5568 (N_5568,N_5084,N_4980);
nand U5569 (N_5569,N_4831,N_4880);
xor U5570 (N_5570,N_5195,N_4972);
nand U5571 (N_5571,N_4862,N_5173);
or U5572 (N_5572,N_5024,N_5112);
nand U5573 (N_5573,N_5169,N_5067);
and U5574 (N_5574,N_5038,N_5164);
or U5575 (N_5575,N_4899,N_4826);
nand U5576 (N_5576,N_4965,N_4888);
xor U5577 (N_5577,N_5136,N_4889);
nor U5578 (N_5578,N_5011,N_5194);
nor U5579 (N_5579,N_4987,N_5081);
or U5580 (N_5580,N_5041,N_4951);
xor U5581 (N_5581,N_4865,N_4995);
nor U5582 (N_5582,N_4857,N_4888);
nor U5583 (N_5583,N_4812,N_4899);
nor U5584 (N_5584,N_4987,N_5114);
nor U5585 (N_5585,N_5141,N_5098);
and U5586 (N_5586,N_5129,N_5041);
and U5587 (N_5587,N_4986,N_5129);
or U5588 (N_5588,N_5131,N_5070);
nand U5589 (N_5589,N_4971,N_4912);
xnor U5590 (N_5590,N_5086,N_5122);
and U5591 (N_5591,N_5083,N_4944);
and U5592 (N_5592,N_4820,N_4921);
xor U5593 (N_5593,N_5092,N_5029);
or U5594 (N_5594,N_5185,N_4929);
xor U5595 (N_5595,N_5190,N_4949);
or U5596 (N_5596,N_5046,N_4900);
or U5597 (N_5597,N_4904,N_4968);
and U5598 (N_5598,N_4993,N_5172);
nand U5599 (N_5599,N_5037,N_4938);
or U5600 (N_5600,N_5388,N_5421);
and U5601 (N_5601,N_5531,N_5265);
nand U5602 (N_5602,N_5343,N_5237);
xor U5603 (N_5603,N_5319,N_5363);
or U5604 (N_5604,N_5377,N_5520);
nand U5605 (N_5605,N_5386,N_5438);
nor U5606 (N_5606,N_5532,N_5518);
and U5607 (N_5607,N_5381,N_5496);
nand U5608 (N_5608,N_5544,N_5457);
and U5609 (N_5609,N_5311,N_5346);
nor U5610 (N_5610,N_5399,N_5272);
xor U5611 (N_5611,N_5347,N_5546);
nand U5612 (N_5612,N_5474,N_5368);
and U5613 (N_5613,N_5390,N_5461);
xor U5614 (N_5614,N_5226,N_5414);
and U5615 (N_5615,N_5261,N_5203);
xor U5616 (N_5616,N_5396,N_5374);
nor U5617 (N_5617,N_5331,N_5511);
xnor U5618 (N_5618,N_5538,N_5507);
or U5619 (N_5619,N_5528,N_5455);
and U5620 (N_5620,N_5301,N_5249);
nor U5621 (N_5621,N_5254,N_5587);
xnor U5622 (N_5622,N_5584,N_5269);
nor U5623 (N_5623,N_5371,N_5534);
nand U5624 (N_5624,N_5586,N_5597);
nor U5625 (N_5625,N_5250,N_5333);
and U5626 (N_5626,N_5354,N_5380);
xnor U5627 (N_5627,N_5452,N_5306);
and U5628 (N_5628,N_5418,N_5530);
nor U5629 (N_5629,N_5458,N_5335);
xnor U5630 (N_5630,N_5425,N_5562);
and U5631 (N_5631,N_5238,N_5566);
nand U5632 (N_5632,N_5324,N_5208);
nand U5633 (N_5633,N_5495,N_5524);
nor U5634 (N_5634,N_5204,N_5393);
xnor U5635 (N_5635,N_5304,N_5353);
nor U5636 (N_5636,N_5283,N_5310);
nor U5637 (N_5637,N_5594,N_5257);
nor U5638 (N_5638,N_5296,N_5579);
or U5639 (N_5639,N_5561,N_5305);
nor U5640 (N_5640,N_5357,N_5423);
nor U5641 (N_5641,N_5350,N_5475);
nor U5642 (N_5642,N_5378,N_5401);
and U5643 (N_5643,N_5448,N_5300);
xnor U5644 (N_5644,N_5504,N_5573);
nor U5645 (N_5645,N_5485,N_5361);
nor U5646 (N_5646,N_5293,N_5429);
xor U5647 (N_5647,N_5451,N_5280);
nor U5648 (N_5648,N_5494,N_5271);
xnor U5649 (N_5649,N_5539,N_5221);
or U5650 (N_5650,N_5405,N_5466);
nand U5651 (N_5651,N_5411,N_5270);
and U5652 (N_5652,N_5246,N_5591);
nor U5653 (N_5653,N_5403,N_5336);
nor U5654 (N_5654,N_5235,N_5574);
nand U5655 (N_5655,N_5444,N_5486);
nor U5656 (N_5656,N_5576,N_5211);
and U5657 (N_5657,N_5223,N_5456);
nor U5658 (N_5658,N_5541,N_5442);
nand U5659 (N_5659,N_5510,N_5351);
xnor U5660 (N_5660,N_5503,N_5500);
xor U5661 (N_5661,N_5537,N_5542);
or U5662 (N_5662,N_5206,N_5345);
xor U5663 (N_5663,N_5329,N_5536);
or U5664 (N_5664,N_5218,N_5327);
nor U5665 (N_5665,N_5598,N_5552);
nor U5666 (N_5666,N_5326,N_5366);
or U5667 (N_5667,N_5593,N_5572);
or U5668 (N_5668,N_5207,N_5568);
and U5669 (N_5669,N_5328,N_5286);
nand U5670 (N_5670,N_5325,N_5323);
or U5671 (N_5671,N_5290,N_5316);
xor U5672 (N_5672,N_5342,N_5404);
xnor U5673 (N_5673,N_5549,N_5557);
nand U5674 (N_5674,N_5349,N_5428);
or U5675 (N_5675,N_5493,N_5372);
nand U5676 (N_5676,N_5288,N_5449);
or U5677 (N_5677,N_5525,N_5558);
nor U5678 (N_5678,N_5416,N_5577);
nand U5679 (N_5679,N_5420,N_5565);
nor U5680 (N_5680,N_5513,N_5295);
nor U5681 (N_5681,N_5468,N_5232);
nor U5682 (N_5682,N_5266,N_5433);
nor U5683 (N_5683,N_5464,N_5337);
nor U5684 (N_5684,N_5364,N_5419);
nand U5685 (N_5685,N_5545,N_5341);
xor U5686 (N_5686,N_5356,N_5596);
and U5687 (N_5687,N_5445,N_5330);
or U5688 (N_5688,N_5589,N_5370);
nand U5689 (N_5689,N_5297,N_5225);
xnor U5690 (N_5690,N_5437,N_5523);
or U5691 (N_5691,N_5369,N_5375);
xnor U5692 (N_5692,N_5450,N_5473);
nor U5693 (N_5693,N_5563,N_5412);
nand U5694 (N_5694,N_5580,N_5459);
nand U5695 (N_5695,N_5321,N_5533);
nand U5696 (N_5696,N_5282,N_5248);
nor U5697 (N_5697,N_5583,N_5240);
xor U5698 (N_5698,N_5505,N_5340);
nor U5699 (N_5699,N_5294,N_5287);
or U5700 (N_5700,N_5317,N_5564);
or U5701 (N_5701,N_5529,N_5307);
or U5702 (N_5702,N_5467,N_5259);
xnor U5703 (N_5703,N_5521,N_5434);
nor U5704 (N_5704,N_5268,N_5365);
xnor U5705 (N_5705,N_5360,N_5263);
and U5706 (N_5706,N_5209,N_5488);
nand U5707 (N_5707,N_5314,N_5383);
nand U5708 (N_5708,N_5410,N_5278);
or U5709 (N_5709,N_5522,N_5230);
nor U5710 (N_5710,N_5277,N_5526);
xnor U5711 (N_5711,N_5470,N_5479);
nand U5712 (N_5712,N_5490,N_5476);
nand U5713 (N_5713,N_5447,N_5373);
or U5714 (N_5714,N_5519,N_5540);
or U5715 (N_5715,N_5400,N_5391);
and U5716 (N_5716,N_5582,N_5251);
or U5717 (N_5717,N_5216,N_5567);
xor U5718 (N_5718,N_5469,N_5492);
nor U5719 (N_5719,N_5432,N_5236);
nand U5720 (N_5720,N_5430,N_5367);
nor U5721 (N_5721,N_5478,N_5590);
and U5722 (N_5722,N_5506,N_5312);
or U5723 (N_5723,N_5385,N_5313);
and U5724 (N_5724,N_5426,N_5202);
xor U5725 (N_5725,N_5348,N_5392);
nor U5726 (N_5726,N_5309,N_5227);
or U5727 (N_5727,N_5344,N_5484);
or U5728 (N_5728,N_5220,N_5440);
nor U5729 (N_5729,N_5446,N_5424);
and U5730 (N_5730,N_5571,N_5441);
or U5731 (N_5731,N_5548,N_5355);
xor U5732 (N_5732,N_5535,N_5436);
nand U5733 (N_5733,N_5508,N_5217);
nand U5734 (N_5734,N_5352,N_5570);
xor U5735 (N_5735,N_5481,N_5554);
or U5736 (N_5736,N_5384,N_5402);
xor U5737 (N_5737,N_5415,N_5581);
nand U5738 (N_5738,N_5210,N_5233);
and U5739 (N_5739,N_5243,N_5362);
xor U5740 (N_5740,N_5422,N_5483);
xnor U5741 (N_5741,N_5359,N_5480);
nand U5742 (N_5742,N_5595,N_5334);
xor U5743 (N_5743,N_5273,N_5245);
and U5744 (N_5744,N_5560,N_5315);
nor U5745 (N_5745,N_5219,N_5276);
and U5746 (N_5746,N_5454,N_5213);
or U5747 (N_5747,N_5244,N_5289);
nand U5748 (N_5748,N_5298,N_5253);
or U5749 (N_5749,N_5275,N_5200);
or U5750 (N_5750,N_5379,N_5252);
xnor U5751 (N_5751,N_5382,N_5499);
nand U5752 (N_5752,N_5527,N_5201);
or U5753 (N_5753,N_5453,N_5575);
xor U5754 (N_5754,N_5222,N_5395);
or U5755 (N_5755,N_5256,N_5241);
and U5756 (N_5756,N_5292,N_5376);
nand U5757 (N_5757,N_5299,N_5515);
xor U5758 (N_5758,N_5212,N_5555);
nor U5759 (N_5759,N_5264,N_5578);
or U5760 (N_5760,N_5215,N_5409);
xnor U5761 (N_5761,N_5543,N_5407);
or U5762 (N_5762,N_5398,N_5205);
nor U5763 (N_5763,N_5258,N_5431);
xor U5764 (N_5764,N_5556,N_5599);
nor U5765 (N_5765,N_5477,N_5260);
nor U5766 (N_5766,N_5284,N_5231);
nor U5767 (N_5767,N_5338,N_5285);
nor U5768 (N_5768,N_5585,N_5413);
and U5769 (N_5769,N_5491,N_5439);
or U5770 (N_5770,N_5592,N_5322);
or U5771 (N_5771,N_5242,N_5427);
xor U5772 (N_5772,N_5267,N_5463);
or U5773 (N_5773,N_5239,N_5318);
nand U5774 (N_5774,N_5358,N_5406);
and U5775 (N_5775,N_5417,N_5435);
xnor U5776 (N_5776,N_5588,N_5394);
xnor U5777 (N_5777,N_5247,N_5443);
nor U5778 (N_5778,N_5547,N_5501);
or U5779 (N_5779,N_5229,N_5502);
nor U5780 (N_5780,N_5234,N_5489);
or U5781 (N_5781,N_5559,N_5339);
nand U5782 (N_5782,N_5262,N_5465);
nor U5783 (N_5783,N_5472,N_5214);
nand U5784 (N_5784,N_5387,N_5553);
and U5785 (N_5785,N_5497,N_5462);
nand U5786 (N_5786,N_5487,N_5569);
nand U5787 (N_5787,N_5255,N_5397);
xor U5788 (N_5788,N_5303,N_5460);
nand U5789 (N_5789,N_5308,N_5550);
and U5790 (N_5790,N_5498,N_5281);
and U5791 (N_5791,N_5320,N_5389);
nor U5792 (N_5792,N_5509,N_5279);
or U5793 (N_5793,N_5291,N_5302);
nand U5794 (N_5794,N_5482,N_5517);
and U5795 (N_5795,N_5551,N_5512);
nor U5796 (N_5796,N_5274,N_5332);
nor U5797 (N_5797,N_5408,N_5471);
and U5798 (N_5798,N_5228,N_5516);
xnor U5799 (N_5799,N_5224,N_5514);
nor U5800 (N_5800,N_5587,N_5279);
nor U5801 (N_5801,N_5385,N_5375);
xor U5802 (N_5802,N_5544,N_5568);
and U5803 (N_5803,N_5387,N_5599);
or U5804 (N_5804,N_5324,N_5335);
nand U5805 (N_5805,N_5543,N_5344);
nor U5806 (N_5806,N_5242,N_5527);
xnor U5807 (N_5807,N_5347,N_5313);
xor U5808 (N_5808,N_5207,N_5284);
nor U5809 (N_5809,N_5238,N_5483);
nor U5810 (N_5810,N_5377,N_5495);
and U5811 (N_5811,N_5379,N_5293);
and U5812 (N_5812,N_5320,N_5583);
nor U5813 (N_5813,N_5464,N_5392);
and U5814 (N_5814,N_5207,N_5259);
or U5815 (N_5815,N_5403,N_5392);
nor U5816 (N_5816,N_5244,N_5433);
and U5817 (N_5817,N_5227,N_5204);
and U5818 (N_5818,N_5313,N_5375);
and U5819 (N_5819,N_5455,N_5286);
and U5820 (N_5820,N_5247,N_5523);
xor U5821 (N_5821,N_5438,N_5504);
xor U5822 (N_5822,N_5251,N_5563);
or U5823 (N_5823,N_5247,N_5517);
nand U5824 (N_5824,N_5354,N_5319);
xor U5825 (N_5825,N_5490,N_5353);
and U5826 (N_5826,N_5342,N_5272);
or U5827 (N_5827,N_5403,N_5247);
nand U5828 (N_5828,N_5535,N_5362);
nor U5829 (N_5829,N_5317,N_5436);
xor U5830 (N_5830,N_5582,N_5272);
and U5831 (N_5831,N_5583,N_5478);
nor U5832 (N_5832,N_5501,N_5237);
nor U5833 (N_5833,N_5443,N_5363);
or U5834 (N_5834,N_5243,N_5549);
nand U5835 (N_5835,N_5562,N_5522);
and U5836 (N_5836,N_5285,N_5586);
xnor U5837 (N_5837,N_5430,N_5404);
nor U5838 (N_5838,N_5341,N_5500);
xnor U5839 (N_5839,N_5369,N_5218);
xnor U5840 (N_5840,N_5261,N_5546);
and U5841 (N_5841,N_5571,N_5370);
nand U5842 (N_5842,N_5409,N_5591);
nand U5843 (N_5843,N_5576,N_5453);
nand U5844 (N_5844,N_5332,N_5343);
xnor U5845 (N_5845,N_5466,N_5301);
or U5846 (N_5846,N_5519,N_5571);
and U5847 (N_5847,N_5526,N_5350);
xnor U5848 (N_5848,N_5379,N_5349);
and U5849 (N_5849,N_5514,N_5367);
nand U5850 (N_5850,N_5467,N_5554);
xnor U5851 (N_5851,N_5492,N_5233);
or U5852 (N_5852,N_5484,N_5515);
nand U5853 (N_5853,N_5296,N_5499);
or U5854 (N_5854,N_5291,N_5203);
nor U5855 (N_5855,N_5550,N_5442);
xnor U5856 (N_5856,N_5479,N_5202);
nand U5857 (N_5857,N_5358,N_5306);
nand U5858 (N_5858,N_5487,N_5208);
or U5859 (N_5859,N_5532,N_5268);
and U5860 (N_5860,N_5409,N_5460);
nand U5861 (N_5861,N_5346,N_5253);
or U5862 (N_5862,N_5244,N_5205);
and U5863 (N_5863,N_5238,N_5365);
or U5864 (N_5864,N_5484,N_5457);
or U5865 (N_5865,N_5579,N_5527);
xor U5866 (N_5866,N_5300,N_5595);
nor U5867 (N_5867,N_5363,N_5579);
or U5868 (N_5868,N_5366,N_5413);
nand U5869 (N_5869,N_5376,N_5431);
and U5870 (N_5870,N_5242,N_5223);
nor U5871 (N_5871,N_5474,N_5248);
xor U5872 (N_5872,N_5518,N_5432);
nand U5873 (N_5873,N_5221,N_5446);
xnor U5874 (N_5874,N_5433,N_5457);
or U5875 (N_5875,N_5363,N_5520);
xnor U5876 (N_5876,N_5304,N_5398);
xnor U5877 (N_5877,N_5381,N_5475);
or U5878 (N_5878,N_5396,N_5475);
xnor U5879 (N_5879,N_5396,N_5299);
and U5880 (N_5880,N_5544,N_5440);
or U5881 (N_5881,N_5598,N_5329);
nor U5882 (N_5882,N_5203,N_5574);
xor U5883 (N_5883,N_5249,N_5265);
nand U5884 (N_5884,N_5239,N_5463);
nor U5885 (N_5885,N_5582,N_5403);
nor U5886 (N_5886,N_5384,N_5448);
xor U5887 (N_5887,N_5558,N_5336);
and U5888 (N_5888,N_5558,N_5449);
and U5889 (N_5889,N_5252,N_5212);
nand U5890 (N_5890,N_5548,N_5553);
and U5891 (N_5891,N_5235,N_5252);
nor U5892 (N_5892,N_5428,N_5570);
nand U5893 (N_5893,N_5553,N_5399);
and U5894 (N_5894,N_5419,N_5457);
nand U5895 (N_5895,N_5308,N_5259);
nand U5896 (N_5896,N_5204,N_5249);
nor U5897 (N_5897,N_5217,N_5415);
nor U5898 (N_5898,N_5549,N_5224);
and U5899 (N_5899,N_5339,N_5491);
or U5900 (N_5900,N_5273,N_5433);
or U5901 (N_5901,N_5291,N_5208);
nand U5902 (N_5902,N_5442,N_5361);
and U5903 (N_5903,N_5233,N_5592);
nand U5904 (N_5904,N_5374,N_5438);
nand U5905 (N_5905,N_5447,N_5570);
xor U5906 (N_5906,N_5307,N_5558);
or U5907 (N_5907,N_5221,N_5323);
nor U5908 (N_5908,N_5583,N_5422);
nand U5909 (N_5909,N_5412,N_5481);
xor U5910 (N_5910,N_5241,N_5200);
nor U5911 (N_5911,N_5386,N_5207);
or U5912 (N_5912,N_5350,N_5456);
and U5913 (N_5913,N_5552,N_5555);
nand U5914 (N_5914,N_5548,N_5306);
or U5915 (N_5915,N_5540,N_5336);
nor U5916 (N_5916,N_5258,N_5328);
nand U5917 (N_5917,N_5349,N_5212);
nor U5918 (N_5918,N_5494,N_5374);
nand U5919 (N_5919,N_5414,N_5560);
xnor U5920 (N_5920,N_5288,N_5415);
nor U5921 (N_5921,N_5535,N_5361);
nor U5922 (N_5922,N_5294,N_5312);
xor U5923 (N_5923,N_5528,N_5467);
nand U5924 (N_5924,N_5261,N_5298);
nand U5925 (N_5925,N_5244,N_5542);
nor U5926 (N_5926,N_5464,N_5470);
xor U5927 (N_5927,N_5331,N_5409);
or U5928 (N_5928,N_5592,N_5553);
xnor U5929 (N_5929,N_5414,N_5594);
xnor U5930 (N_5930,N_5205,N_5296);
or U5931 (N_5931,N_5534,N_5470);
and U5932 (N_5932,N_5298,N_5394);
or U5933 (N_5933,N_5491,N_5247);
nor U5934 (N_5934,N_5576,N_5273);
or U5935 (N_5935,N_5449,N_5515);
nor U5936 (N_5936,N_5222,N_5590);
or U5937 (N_5937,N_5428,N_5333);
or U5938 (N_5938,N_5273,N_5222);
xnor U5939 (N_5939,N_5502,N_5409);
nand U5940 (N_5940,N_5458,N_5447);
nand U5941 (N_5941,N_5256,N_5245);
xor U5942 (N_5942,N_5260,N_5230);
nor U5943 (N_5943,N_5303,N_5317);
nand U5944 (N_5944,N_5211,N_5382);
or U5945 (N_5945,N_5445,N_5511);
and U5946 (N_5946,N_5540,N_5573);
xnor U5947 (N_5947,N_5552,N_5255);
nand U5948 (N_5948,N_5463,N_5298);
and U5949 (N_5949,N_5593,N_5278);
nor U5950 (N_5950,N_5421,N_5351);
xnor U5951 (N_5951,N_5411,N_5405);
or U5952 (N_5952,N_5398,N_5492);
nor U5953 (N_5953,N_5470,N_5305);
xor U5954 (N_5954,N_5437,N_5326);
and U5955 (N_5955,N_5511,N_5491);
nand U5956 (N_5956,N_5328,N_5311);
and U5957 (N_5957,N_5247,N_5281);
or U5958 (N_5958,N_5351,N_5516);
nor U5959 (N_5959,N_5394,N_5375);
xnor U5960 (N_5960,N_5399,N_5318);
nor U5961 (N_5961,N_5406,N_5473);
nor U5962 (N_5962,N_5414,N_5203);
and U5963 (N_5963,N_5510,N_5545);
nor U5964 (N_5964,N_5502,N_5473);
nand U5965 (N_5965,N_5444,N_5252);
xnor U5966 (N_5966,N_5383,N_5549);
nor U5967 (N_5967,N_5544,N_5204);
nand U5968 (N_5968,N_5383,N_5385);
or U5969 (N_5969,N_5359,N_5571);
nor U5970 (N_5970,N_5389,N_5576);
xor U5971 (N_5971,N_5595,N_5264);
and U5972 (N_5972,N_5278,N_5351);
or U5973 (N_5973,N_5426,N_5402);
or U5974 (N_5974,N_5401,N_5431);
or U5975 (N_5975,N_5209,N_5548);
or U5976 (N_5976,N_5522,N_5435);
xor U5977 (N_5977,N_5511,N_5412);
xnor U5978 (N_5978,N_5542,N_5444);
nor U5979 (N_5979,N_5367,N_5489);
or U5980 (N_5980,N_5433,N_5437);
nor U5981 (N_5981,N_5337,N_5212);
xnor U5982 (N_5982,N_5312,N_5409);
nor U5983 (N_5983,N_5232,N_5231);
and U5984 (N_5984,N_5300,N_5263);
and U5985 (N_5985,N_5290,N_5238);
or U5986 (N_5986,N_5508,N_5323);
or U5987 (N_5987,N_5308,N_5219);
or U5988 (N_5988,N_5258,N_5220);
xor U5989 (N_5989,N_5422,N_5527);
or U5990 (N_5990,N_5466,N_5546);
xnor U5991 (N_5991,N_5203,N_5283);
nand U5992 (N_5992,N_5250,N_5462);
or U5993 (N_5993,N_5281,N_5368);
nor U5994 (N_5994,N_5301,N_5294);
xor U5995 (N_5995,N_5292,N_5328);
and U5996 (N_5996,N_5204,N_5223);
nand U5997 (N_5997,N_5455,N_5376);
nor U5998 (N_5998,N_5331,N_5351);
and U5999 (N_5999,N_5334,N_5438);
or U6000 (N_6000,N_5985,N_5767);
and U6001 (N_6001,N_5826,N_5788);
xor U6002 (N_6002,N_5827,N_5951);
nor U6003 (N_6003,N_5706,N_5792);
nor U6004 (N_6004,N_5714,N_5682);
nand U6005 (N_6005,N_5881,N_5806);
nand U6006 (N_6006,N_5915,N_5815);
or U6007 (N_6007,N_5898,N_5833);
xor U6008 (N_6008,N_5908,N_5777);
nand U6009 (N_6009,N_5784,N_5984);
and U6010 (N_6010,N_5997,N_5846);
nor U6011 (N_6011,N_5701,N_5916);
xor U6012 (N_6012,N_5606,N_5691);
nand U6013 (N_6013,N_5905,N_5889);
nand U6014 (N_6014,N_5938,N_5628);
or U6015 (N_6015,N_5869,N_5974);
nand U6016 (N_6016,N_5931,N_5883);
nand U6017 (N_6017,N_5808,N_5862);
xor U6018 (N_6018,N_5977,N_5865);
and U6019 (N_6019,N_5635,N_5939);
nor U6020 (N_6020,N_5677,N_5825);
or U6021 (N_6021,N_5947,N_5769);
xor U6022 (N_6022,N_5885,N_5958);
and U6023 (N_6023,N_5992,N_5854);
or U6024 (N_6024,N_5617,N_5936);
or U6025 (N_6025,N_5659,N_5751);
nand U6026 (N_6026,N_5824,N_5671);
nand U6027 (N_6027,N_5819,N_5723);
xor U6028 (N_6028,N_5796,N_5741);
and U6029 (N_6029,N_5674,N_5952);
xor U6030 (N_6030,N_5948,N_5725);
xor U6031 (N_6031,N_5790,N_5717);
xor U6032 (N_6032,N_5721,N_5665);
nand U6033 (N_6033,N_5868,N_5861);
xnor U6034 (N_6034,N_5837,N_5849);
or U6035 (N_6035,N_5660,N_5716);
and U6036 (N_6036,N_5633,N_5732);
xnor U6037 (N_6037,N_5904,N_5967);
nor U6038 (N_6038,N_5686,N_5656);
and U6039 (N_6039,N_5911,N_5787);
nand U6040 (N_6040,N_5776,N_5630);
and U6041 (N_6041,N_5745,N_5711);
xnor U6042 (N_6042,N_5965,N_5636);
nand U6043 (N_6043,N_5813,N_5744);
nand U6044 (N_6044,N_5839,N_5774);
xnor U6045 (N_6045,N_5964,N_5834);
or U6046 (N_6046,N_5900,N_5983);
or U6047 (N_6047,N_5734,N_5971);
or U6048 (N_6048,N_5622,N_5782);
or U6049 (N_6049,N_5903,N_5728);
and U6050 (N_6050,N_5654,N_5828);
or U6051 (N_6051,N_5852,N_5795);
or U6052 (N_6052,N_5949,N_5912);
xor U6053 (N_6053,N_5888,N_5611);
nand U6054 (N_6054,N_5731,N_5803);
nor U6055 (N_6055,N_5830,N_5943);
nor U6056 (N_6056,N_5764,N_5978);
nor U6057 (N_6057,N_5661,N_5797);
or U6058 (N_6058,N_5755,N_5627);
xor U6059 (N_6059,N_5609,N_5866);
nor U6060 (N_6060,N_5876,N_5894);
or U6061 (N_6061,N_5968,N_5634);
nor U6062 (N_6062,N_5873,N_5812);
xor U6063 (N_6063,N_5793,N_5919);
nand U6064 (N_6064,N_5874,N_5648);
nand U6065 (N_6065,N_5637,N_5644);
or U6066 (N_6066,N_5791,N_5831);
nor U6067 (N_6067,N_5647,N_5690);
nand U6068 (N_6068,N_5749,N_5698);
xnor U6069 (N_6069,N_5932,N_5937);
nand U6070 (N_6070,N_5884,N_5618);
xor U6071 (N_6071,N_5859,N_5925);
or U6072 (N_6072,N_5941,N_5853);
xor U6073 (N_6073,N_5961,N_5867);
or U6074 (N_6074,N_5973,N_5653);
or U6075 (N_6075,N_5991,N_5928);
xor U6076 (N_6076,N_5929,N_5705);
nor U6077 (N_6077,N_5707,N_5680);
nor U6078 (N_6078,N_5718,N_5761);
and U6079 (N_6079,N_5724,N_5935);
nor U6080 (N_6080,N_5993,N_5641);
or U6081 (N_6081,N_5989,N_5838);
nand U6082 (N_6082,N_5766,N_5614);
and U6083 (N_6083,N_5802,N_5959);
nand U6084 (N_6084,N_5902,N_5730);
nand U6085 (N_6085,N_5799,N_5986);
and U6086 (N_6086,N_5963,N_5639);
xnor U6087 (N_6087,N_5969,N_5804);
and U6088 (N_6088,N_5768,N_5794);
or U6089 (N_6089,N_5844,N_5673);
nand U6090 (N_6090,N_5652,N_5856);
nand U6091 (N_6091,N_5818,N_5783);
and U6092 (N_6092,N_5860,N_5956);
nor U6093 (N_6093,N_5798,N_5603);
xnor U6094 (N_6094,N_5891,N_5920);
nand U6095 (N_6095,N_5650,N_5922);
nor U6096 (N_6096,N_5886,N_5763);
and U6097 (N_6097,N_5944,N_5981);
xor U6098 (N_6098,N_5709,N_5923);
nand U6099 (N_6099,N_5785,N_5924);
and U6100 (N_6100,N_5610,N_5693);
or U6101 (N_6101,N_5942,N_5684);
or U6102 (N_6102,N_5613,N_5700);
or U6103 (N_6103,N_5835,N_5770);
nand U6104 (N_6104,N_5821,N_5695);
nand U6105 (N_6105,N_5845,N_5623);
or U6106 (N_6106,N_5664,N_5934);
nor U6107 (N_6107,N_5737,N_5913);
and U6108 (N_6108,N_5829,N_5990);
nand U6109 (N_6109,N_5864,N_5762);
or U6110 (N_6110,N_5672,N_5820);
nor U6111 (N_6111,N_5739,N_5616);
and U6112 (N_6112,N_5870,N_5918);
nor U6113 (N_6113,N_5608,N_5748);
and U6114 (N_6114,N_5712,N_5950);
xnor U6115 (N_6115,N_5926,N_5980);
xor U6116 (N_6116,N_5987,N_5675);
and U6117 (N_6117,N_5962,N_5863);
nand U6118 (N_6118,N_5921,N_5676);
or U6119 (N_6119,N_5933,N_5740);
or U6120 (N_6120,N_5893,N_5946);
nor U6121 (N_6121,N_5708,N_5955);
or U6122 (N_6122,N_5880,N_5996);
xnor U6123 (N_6123,N_5729,N_5697);
and U6124 (N_6124,N_5800,N_5779);
and U6125 (N_6125,N_5607,N_5927);
or U6126 (N_6126,N_5687,N_5836);
xor U6127 (N_6127,N_5759,N_5688);
nand U6128 (N_6128,N_5786,N_5643);
and U6129 (N_6129,N_5663,N_5662);
nand U6130 (N_6130,N_5752,N_5601);
nor U6131 (N_6131,N_5851,N_5757);
xor U6132 (N_6132,N_5638,N_5624);
nor U6133 (N_6133,N_5976,N_5954);
xor U6134 (N_6134,N_5668,N_5625);
xor U6135 (N_6135,N_5892,N_5602);
xor U6136 (N_6136,N_5979,N_5720);
nand U6137 (N_6137,N_5970,N_5896);
xor U6138 (N_6138,N_5906,N_5754);
or U6139 (N_6139,N_5899,N_5667);
nand U6140 (N_6140,N_5909,N_5907);
xor U6141 (N_6141,N_5817,N_5940);
and U6142 (N_6142,N_5738,N_5649);
and U6143 (N_6143,N_5887,N_5679);
xnor U6144 (N_6144,N_5736,N_5771);
xnor U6145 (N_6145,N_5890,N_5789);
or U6146 (N_6146,N_5850,N_5685);
nor U6147 (N_6147,N_5760,N_5620);
xor U6148 (N_6148,N_5841,N_5972);
xnor U6149 (N_6149,N_5692,N_5914);
xnor U6150 (N_6150,N_5742,N_5683);
or U6151 (N_6151,N_5678,N_5681);
nand U6152 (N_6152,N_5722,N_5758);
xor U6153 (N_6153,N_5703,N_5966);
nand U6154 (N_6154,N_5823,N_5957);
and U6155 (N_6155,N_5995,N_5848);
nor U6156 (N_6156,N_5619,N_5726);
nand U6157 (N_6157,N_5651,N_5612);
nand U6158 (N_6158,N_5811,N_5832);
nand U6159 (N_6159,N_5882,N_5646);
nor U6160 (N_6160,N_5810,N_5901);
xor U6161 (N_6161,N_5805,N_5999);
nor U6162 (N_6162,N_5666,N_5855);
xor U6163 (N_6163,N_5746,N_5753);
nor U6164 (N_6164,N_5975,N_5632);
and U6165 (N_6165,N_5843,N_5840);
xnor U6166 (N_6166,N_5878,N_5604);
nand U6167 (N_6167,N_5822,N_5998);
nor U6168 (N_6168,N_5772,N_5858);
and U6169 (N_6169,N_5696,N_5719);
nor U6170 (N_6170,N_5775,N_5655);
nand U6171 (N_6171,N_5756,N_5715);
xnor U6172 (N_6172,N_5988,N_5930);
and U6173 (N_6173,N_5626,N_5877);
and U6174 (N_6174,N_5642,N_5733);
or U6175 (N_6175,N_5750,N_5872);
or U6176 (N_6176,N_5699,N_5743);
and U6177 (N_6177,N_5658,N_5640);
nor U6178 (N_6178,N_5945,N_5765);
nor U6179 (N_6179,N_5727,N_5689);
xor U6180 (N_6180,N_5694,N_5857);
and U6181 (N_6181,N_5600,N_5910);
and U6182 (N_6182,N_5702,N_5895);
or U6183 (N_6183,N_5747,N_5875);
and U6184 (N_6184,N_5629,N_5960);
nor U6185 (N_6185,N_5816,N_5780);
and U6186 (N_6186,N_5842,N_5704);
and U6187 (N_6187,N_5615,N_5631);
or U6188 (N_6188,N_5982,N_5781);
nor U6189 (N_6189,N_5645,N_5713);
nand U6190 (N_6190,N_5710,N_5871);
nand U6191 (N_6191,N_5994,N_5917);
nand U6192 (N_6192,N_5605,N_5621);
nor U6193 (N_6193,N_5809,N_5847);
nand U6194 (N_6194,N_5657,N_5670);
and U6195 (N_6195,N_5801,N_5953);
nand U6196 (N_6196,N_5814,N_5669);
or U6197 (N_6197,N_5879,N_5778);
nand U6198 (N_6198,N_5735,N_5773);
nor U6199 (N_6199,N_5897,N_5807);
or U6200 (N_6200,N_5974,N_5719);
nor U6201 (N_6201,N_5898,N_5952);
or U6202 (N_6202,N_5797,N_5863);
xnor U6203 (N_6203,N_5937,N_5638);
nand U6204 (N_6204,N_5645,N_5917);
or U6205 (N_6205,N_5815,N_5718);
nand U6206 (N_6206,N_5970,N_5669);
xor U6207 (N_6207,N_5624,N_5718);
xnor U6208 (N_6208,N_5983,N_5661);
or U6209 (N_6209,N_5985,N_5911);
and U6210 (N_6210,N_5667,N_5959);
nand U6211 (N_6211,N_5980,N_5692);
nand U6212 (N_6212,N_5606,N_5926);
or U6213 (N_6213,N_5602,N_5709);
nand U6214 (N_6214,N_5764,N_5964);
nand U6215 (N_6215,N_5658,N_5971);
or U6216 (N_6216,N_5810,N_5768);
or U6217 (N_6217,N_5627,N_5811);
nor U6218 (N_6218,N_5674,N_5775);
and U6219 (N_6219,N_5750,N_5797);
or U6220 (N_6220,N_5653,N_5824);
xnor U6221 (N_6221,N_5638,N_5666);
nor U6222 (N_6222,N_5890,N_5956);
and U6223 (N_6223,N_5715,N_5691);
nand U6224 (N_6224,N_5891,N_5675);
or U6225 (N_6225,N_5908,N_5647);
nand U6226 (N_6226,N_5871,N_5657);
or U6227 (N_6227,N_5785,N_5635);
and U6228 (N_6228,N_5801,N_5778);
nand U6229 (N_6229,N_5830,N_5985);
or U6230 (N_6230,N_5745,N_5830);
nand U6231 (N_6231,N_5853,N_5646);
or U6232 (N_6232,N_5776,N_5794);
nor U6233 (N_6233,N_5857,N_5948);
xor U6234 (N_6234,N_5832,N_5776);
nand U6235 (N_6235,N_5822,N_5914);
nor U6236 (N_6236,N_5800,N_5766);
xnor U6237 (N_6237,N_5894,N_5753);
nor U6238 (N_6238,N_5863,N_5770);
nor U6239 (N_6239,N_5851,N_5940);
or U6240 (N_6240,N_5853,N_5720);
or U6241 (N_6241,N_5922,N_5624);
nor U6242 (N_6242,N_5643,N_5860);
nand U6243 (N_6243,N_5604,N_5781);
or U6244 (N_6244,N_5681,N_5626);
nand U6245 (N_6245,N_5637,N_5792);
and U6246 (N_6246,N_5924,N_5774);
and U6247 (N_6247,N_5848,N_5704);
xnor U6248 (N_6248,N_5928,N_5652);
nand U6249 (N_6249,N_5753,N_5827);
and U6250 (N_6250,N_5834,N_5890);
nor U6251 (N_6251,N_5727,N_5975);
nand U6252 (N_6252,N_5926,N_5899);
and U6253 (N_6253,N_5713,N_5773);
and U6254 (N_6254,N_5820,N_5960);
and U6255 (N_6255,N_5937,N_5731);
or U6256 (N_6256,N_5840,N_5689);
nor U6257 (N_6257,N_5687,N_5633);
or U6258 (N_6258,N_5654,N_5883);
nor U6259 (N_6259,N_5940,N_5761);
xor U6260 (N_6260,N_5941,N_5862);
and U6261 (N_6261,N_5669,N_5694);
and U6262 (N_6262,N_5607,N_5769);
nor U6263 (N_6263,N_5932,N_5680);
or U6264 (N_6264,N_5705,N_5779);
nor U6265 (N_6265,N_5719,N_5936);
or U6266 (N_6266,N_5609,N_5995);
xnor U6267 (N_6267,N_5938,N_5646);
xnor U6268 (N_6268,N_5760,N_5976);
and U6269 (N_6269,N_5946,N_5825);
or U6270 (N_6270,N_5620,N_5730);
xor U6271 (N_6271,N_5981,N_5707);
xnor U6272 (N_6272,N_5649,N_5750);
xor U6273 (N_6273,N_5872,N_5685);
and U6274 (N_6274,N_5665,N_5650);
nand U6275 (N_6275,N_5600,N_5606);
nor U6276 (N_6276,N_5961,N_5770);
and U6277 (N_6277,N_5791,N_5653);
or U6278 (N_6278,N_5911,N_5758);
and U6279 (N_6279,N_5920,N_5738);
xor U6280 (N_6280,N_5843,N_5889);
nor U6281 (N_6281,N_5955,N_5933);
and U6282 (N_6282,N_5953,N_5885);
xor U6283 (N_6283,N_5988,N_5644);
and U6284 (N_6284,N_5763,N_5836);
and U6285 (N_6285,N_5808,N_5687);
and U6286 (N_6286,N_5692,N_5722);
nor U6287 (N_6287,N_5777,N_5713);
nor U6288 (N_6288,N_5767,N_5733);
xnor U6289 (N_6289,N_5974,N_5981);
nand U6290 (N_6290,N_5746,N_5987);
nand U6291 (N_6291,N_5733,N_5654);
or U6292 (N_6292,N_5792,N_5997);
or U6293 (N_6293,N_5745,N_5884);
nand U6294 (N_6294,N_5888,N_5760);
and U6295 (N_6295,N_5660,N_5817);
nand U6296 (N_6296,N_5857,N_5674);
or U6297 (N_6297,N_5867,N_5697);
nor U6298 (N_6298,N_5755,N_5882);
and U6299 (N_6299,N_5918,N_5928);
and U6300 (N_6300,N_5885,N_5949);
xnor U6301 (N_6301,N_5835,N_5796);
or U6302 (N_6302,N_5648,N_5687);
and U6303 (N_6303,N_5805,N_5681);
and U6304 (N_6304,N_5612,N_5891);
nand U6305 (N_6305,N_5832,N_5756);
xnor U6306 (N_6306,N_5625,N_5916);
nand U6307 (N_6307,N_5602,N_5898);
nand U6308 (N_6308,N_5714,N_5825);
and U6309 (N_6309,N_5662,N_5623);
and U6310 (N_6310,N_5855,N_5637);
nor U6311 (N_6311,N_5747,N_5759);
nor U6312 (N_6312,N_5652,N_5745);
nand U6313 (N_6313,N_5884,N_5856);
nand U6314 (N_6314,N_5626,N_5796);
xor U6315 (N_6315,N_5812,N_5841);
or U6316 (N_6316,N_5962,N_5654);
and U6317 (N_6317,N_5682,N_5903);
xor U6318 (N_6318,N_5642,N_5980);
xor U6319 (N_6319,N_5627,N_5723);
nand U6320 (N_6320,N_5630,N_5759);
nor U6321 (N_6321,N_5956,N_5871);
xnor U6322 (N_6322,N_5901,N_5900);
nand U6323 (N_6323,N_5982,N_5749);
nand U6324 (N_6324,N_5620,N_5767);
and U6325 (N_6325,N_5616,N_5679);
nand U6326 (N_6326,N_5669,N_5982);
or U6327 (N_6327,N_5888,N_5913);
and U6328 (N_6328,N_5936,N_5833);
and U6329 (N_6329,N_5680,N_5976);
nor U6330 (N_6330,N_5810,N_5722);
or U6331 (N_6331,N_5912,N_5725);
nand U6332 (N_6332,N_5705,N_5772);
or U6333 (N_6333,N_5858,N_5953);
nand U6334 (N_6334,N_5760,N_5761);
nor U6335 (N_6335,N_5811,N_5769);
or U6336 (N_6336,N_5923,N_5831);
nor U6337 (N_6337,N_5666,N_5635);
nor U6338 (N_6338,N_5673,N_5996);
or U6339 (N_6339,N_5917,N_5996);
and U6340 (N_6340,N_5880,N_5957);
nand U6341 (N_6341,N_5738,N_5626);
xor U6342 (N_6342,N_5601,N_5970);
and U6343 (N_6343,N_5737,N_5748);
xor U6344 (N_6344,N_5718,N_5613);
nand U6345 (N_6345,N_5993,N_5740);
and U6346 (N_6346,N_5964,N_5922);
xnor U6347 (N_6347,N_5855,N_5840);
nor U6348 (N_6348,N_5934,N_5639);
and U6349 (N_6349,N_5639,N_5891);
and U6350 (N_6350,N_5884,N_5712);
or U6351 (N_6351,N_5720,N_5611);
and U6352 (N_6352,N_5999,N_5786);
nor U6353 (N_6353,N_5916,N_5620);
nor U6354 (N_6354,N_5783,N_5732);
and U6355 (N_6355,N_5934,N_5699);
or U6356 (N_6356,N_5793,N_5716);
xnor U6357 (N_6357,N_5874,N_5756);
and U6358 (N_6358,N_5976,N_5675);
xnor U6359 (N_6359,N_5928,N_5832);
xor U6360 (N_6360,N_5876,N_5972);
nand U6361 (N_6361,N_5919,N_5886);
nand U6362 (N_6362,N_5685,N_5855);
or U6363 (N_6363,N_5993,N_5868);
xor U6364 (N_6364,N_5942,N_5743);
xor U6365 (N_6365,N_5651,N_5898);
nor U6366 (N_6366,N_5730,N_5839);
and U6367 (N_6367,N_5758,N_5749);
nand U6368 (N_6368,N_5679,N_5961);
nand U6369 (N_6369,N_5801,N_5623);
xor U6370 (N_6370,N_5711,N_5847);
and U6371 (N_6371,N_5809,N_5902);
nand U6372 (N_6372,N_5753,N_5701);
and U6373 (N_6373,N_5989,N_5968);
or U6374 (N_6374,N_5638,N_5703);
and U6375 (N_6375,N_5917,N_5833);
or U6376 (N_6376,N_5639,N_5878);
nor U6377 (N_6377,N_5775,N_5838);
xnor U6378 (N_6378,N_5727,N_5712);
nand U6379 (N_6379,N_5881,N_5836);
or U6380 (N_6380,N_5846,N_5660);
nor U6381 (N_6381,N_5602,N_5699);
and U6382 (N_6382,N_5885,N_5733);
nand U6383 (N_6383,N_5712,N_5889);
and U6384 (N_6384,N_5898,N_5646);
and U6385 (N_6385,N_5749,N_5754);
nand U6386 (N_6386,N_5863,N_5761);
nand U6387 (N_6387,N_5633,N_5765);
and U6388 (N_6388,N_5825,N_5978);
xor U6389 (N_6389,N_5892,N_5693);
and U6390 (N_6390,N_5851,N_5859);
xor U6391 (N_6391,N_5993,N_5746);
nor U6392 (N_6392,N_5604,N_5629);
nor U6393 (N_6393,N_5630,N_5956);
or U6394 (N_6394,N_5964,N_5657);
nor U6395 (N_6395,N_5726,N_5673);
xor U6396 (N_6396,N_5679,N_5983);
xor U6397 (N_6397,N_5872,N_5726);
nand U6398 (N_6398,N_5604,N_5609);
and U6399 (N_6399,N_5930,N_5802);
nand U6400 (N_6400,N_6194,N_6002);
and U6401 (N_6401,N_6377,N_6089);
or U6402 (N_6402,N_6282,N_6143);
xor U6403 (N_6403,N_6385,N_6199);
or U6404 (N_6404,N_6230,N_6388);
xor U6405 (N_6405,N_6149,N_6390);
nand U6406 (N_6406,N_6139,N_6387);
and U6407 (N_6407,N_6093,N_6075);
nor U6408 (N_6408,N_6115,N_6320);
xor U6409 (N_6409,N_6142,N_6195);
nor U6410 (N_6410,N_6361,N_6373);
nand U6411 (N_6411,N_6008,N_6267);
xor U6412 (N_6412,N_6040,N_6256);
nand U6413 (N_6413,N_6109,N_6290);
xnor U6414 (N_6414,N_6277,N_6317);
nand U6415 (N_6415,N_6127,N_6119);
nand U6416 (N_6416,N_6296,N_6244);
or U6417 (N_6417,N_6322,N_6196);
or U6418 (N_6418,N_6270,N_6327);
nand U6419 (N_6419,N_6017,N_6177);
and U6420 (N_6420,N_6105,N_6031);
nand U6421 (N_6421,N_6355,N_6088);
nand U6422 (N_6422,N_6281,N_6333);
xor U6423 (N_6423,N_6259,N_6136);
or U6424 (N_6424,N_6133,N_6353);
xor U6425 (N_6425,N_6231,N_6280);
or U6426 (N_6426,N_6248,N_6135);
nor U6427 (N_6427,N_6058,N_6092);
or U6428 (N_6428,N_6329,N_6313);
nor U6429 (N_6429,N_6396,N_6225);
nand U6430 (N_6430,N_6399,N_6162);
or U6431 (N_6431,N_6336,N_6069);
and U6432 (N_6432,N_6125,N_6309);
and U6433 (N_6433,N_6180,N_6352);
nand U6434 (N_6434,N_6154,N_6386);
xnor U6435 (N_6435,N_6001,N_6156);
or U6436 (N_6436,N_6351,N_6184);
or U6437 (N_6437,N_6182,N_6150);
nor U6438 (N_6438,N_6090,N_6397);
nand U6439 (N_6439,N_6024,N_6272);
nand U6440 (N_6440,N_6011,N_6203);
and U6441 (N_6441,N_6219,N_6208);
or U6442 (N_6442,N_6275,N_6384);
and U6443 (N_6443,N_6285,N_6269);
nor U6444 (N_6444,N_6077,N_6114);
or U6445 (N_6445,N_6273,N_6026);
nand U6446 (N_6446,N_6021,N_6066);
nor U6447 (N_6447,N_6006,N_6094);
nand U6448 (N_6448,N_6237,N_6205);
or U6449 (N_6449,N_6372,N_6364);
nand U6450 (N_6450,N_6249,N_6144);
and U6451 (N_6451,N_6048,N_6350);
or U6452 (N_6452,N_6212,N_6246);
nor U6453 (N_6453,N_6147,N_6032);
nor U6454 (N_6454,N_6044,N_6170);
and U6455 (N_6455,N_6095,N_6016);
nor U6456 (N_6456,N_6153,N_6383);
nor U6457 (N_6457,N_6247,N_6347);
nor U6458 (N_6458,N_6028,N_6227);
nand U6459 (N_6459,N_6302,N_6071);
xnor U6460 (N_6460,N_6356,N_6067);
nand U6461 (N_6461,N_6348,N_6254);
xnor U6462 (N_6462,N_6366,N_6202);
and U6463 (N_6463,N_6264,N_6191);
nand U6464 (N_6464,N_6365,N_6051);
or U6465 (N_6465,N_6297,N_6304);
or U6466 (N_6466,N_6039,N_6164);
nor U6467 (N_6467,N_6286,N_6243);
or U6468 (N_6468,N_6229,N_6197);
nor U6469 (N_6469,N_6129,N_6371);
and U6470 (N_6470,N_6014,N_6060);
or U6471 (N_6471,N_6370,N_6165);
nand U6472 (N_6472,N_6343,N_6107);
nor U6473 (N_6473,N_6151,N_6326);
and U6474 (N_6474,N_6027,N_6068);
nor U6475 (N_6475,N_6260,N_6284);
nand U6476 (N_6476,N_6301,N_6158);
nor U6477 (N_6477,N_6221,N_6188);
or U6478 (N_6478,N_6220,N_6111);
nor U6479 (N_6479,N_6303,N_6190);
or U6480 (N_6480,N_6233,N_6339);
or U6481 (N_6481,N_6344,N_6314);
nand U6482 (N_6482,N_6321,N_6086);
nand U6483 (N_6483,N_6148,N_6187);
or U6484 (N_6484,N_6210,N_6169);
and U6485 (N_6485,N_6342,N_6228);
or U6486 (N_6486,N_6161,N_6185);
nor U6487 (N_6487,N_6157,N_6192);
and U6488 (N_6488,N_6059,N_6193);
xnor U6489 (N_6489,N_6263,N_6116);
or U6490 (N_6490,N_6003,N_6382);
xor U6491 (N_6491,N_6084,N_6065);
nor U6492 (N_6492,N_6106,N_6393);
nand U6493 (N_6493,N_6056,N_6181);
and U6494 (N_6494,N_6380,N_6070);
or U6495 (N_6495,N_6152,N_6074);
xnor U6496 (N_6496,N_6018,N_6323);
or U6497 (N_6497,N_6292,N_6015);
nor U6498 (N_6498,N_6389,N_6020);
nor U6499 (N_6499,N_6045,N_6214);
xor U6500 (N_6500,N_6341,N_6005);
nand U6501 (N_6501,N_6076,N_6101);
nand U6502 (N_6502,N_6236,N_6010);
nor U6503 (N_6503,N_6340,N_6080);
nand U6504 (N_6504,N_6337,N_6168);
xor U6505 (N_6505,N_6310,N_6346);
nor U6506 (N_6506,N_6207,N_6271);
nand U6507 (N_6507,N_6175,N_6038);
xor U6508 (N_6508,N_6091,N_6118);
nor U6509 (N_6509,N_6315,N_6345);
and U6510 (N_6510,N_6369,N_6265);
xnor U6511 (N_6511,N_6025,N_6007);
and U6512 (N_6512,N_6166,N_6122);
nand U6513 (N_6513,N_6183,N_6335);
nand U6514 (N_6514,N_6253,N_6287);
and U6515 (N_6515,N_6251,N_6103);
nor U6516 (N_6516,N_6201,N_6121);
nor U6517 (N_6517,N_6167,N_6100);
and U6518 (N_6518,N_6087,N_6223);
or U6519 (N_6519,N_6252,N_6022);
nor U6520 (N_6520,N_6288,N_6216);
or U6521 (N_6521,N_6206,N_6030);
nor U6522 (N_6522,N_6000,N_6368);
nand U6523 (N_6523,N_6173,N_6276);
nand U6524 (N_6524,N_6359,N_6261);
nand U6525 (N_6525,N_6037,N_6174);
or U6526 (N_6526,N_6360,N_6262);
nor U6527 (N_6527,N_6033,N_6374);
xor U6528 (N_6528,N_6307,N_6198);
and U6529 (N_6529,N_6041,N_6300);
or U6530 (N_6530,N_6160,N_6395);
nor U6531 (N_6531,N_6137,N_6306);
nor U6532 (N_6532,N_6305,N_6062);
xor U6533 (N_6533,N_6034,N_6312);
nand U6534 (N_6534,N_6283,N_6132);
and U6535 (N_6535,N_6117,N_6126);
nand U6536 (N_6536,N_6381,N_6078);
nor U6537 (N_6537,N_6330,N_6113);
nand U6538 (N_6538,N_6036,N_6053);
xnor U6539 (N_6539,N_6325,N_6104);
nand U6540 (N_6540,N_6042,N_6072);
nor U6541 (N_6541,N_6004,N_6391);
xnor U6542 (N_6542,N_6145,N_6061);
nand U6543 (N_6543,N_6081,N_6082);
nand U6544 (N_6544,N_6064,N_6289);
nand U6545 (N_6545,N_6134,N_6367);
and U6546 (N_6546,N_6099,N_6049);
and U6547 (N_6547,N_6200,N_6311);
xnor U6548 (N_6548,N_6146,N_6124);
nand U6549 (N_6549,N_6217,N_6238);
nor U6550 (N_6550,N_6332,N_6226);
or U6551 (N_6551,N_6354,N_6108);
and U6552 (N_6552,N_6130,N_6338);
or U6553 (N_6553,N_6023,N_6172);
and U6554 (N_6554,N_6138,N_6159);
nand U6555 (N_6555,N_6394,N_6375);
and U6556 (N_6556,N_6308,N_6178);
and U6557 (N_6557,N_6291,N_6097);
nand U6558 (N_6558,N_6363,N_6234);
nand U6559 (N_6559,N_6224,N_6057);
nor U6560 (N_6560,N_6029,N_6128);
and U6561 (N_6561,N_6055,N_6241);
xnor U6562 (N_6562,N_6073,N_6123);
xnor U6563 (N_6563,N_6046,N_6163);
and U6564 (N_6564,N_6398,N_6102);
nor U6565 (N_6565,N_6293,N_6098);
nor U6566 (N_6566,N_6050,N_6019);
and U6567 (N_6567,N_6112,N_6141);
nand U6568 (N_6568,N_6186,N_6096);
nor U6569 (N_6569,N_6179,N_6328);
nor U6570 (N_6570,N_6392,N_6250);
nor U6571 (N_6571,N_6035,N_6268);
nor U6572 (N_6572,N_6318,N_6215);
and U6573 (N_6573,N_6295,N_6211);
nor U6574 (N_6574,N_6245,N_6140);
or U6575 (N_6575,N_6043,N_6209);
or U6576 (N_6576,N_6120,N_6012);
nor U6577 (N_6577,N_6299,N_6298);
nor U6578 (N_6578,N_6047,N_6278);
or U6579 (N_6579,N_6255,N_6063);
xor U6580 (N_6580,N_6331,N_6213);
xor U6581 (N_6581,N_6218,N_6085);
nand U6582 (N_6582,N_6274,N_6232);
or U6583 (N_6583,N_6009,N_6358);
nor U6584 (N_6584,N_6235,N_6362);
nand U6585 (N_6585,N_6240,N_6013);
nand U6586 (N_6586,N_6083,N_6171);
xnor U6587 (N_6587,N_6316,N_6294);
or U6588 (N_6588,N_6349,N_6279);
nand U6589 (N_6589,N_6189,N_6324);
xnor U6590 (N_6590,N_6054,N_6376);
nor U6591 (N_6591,N_6176,N_6242);
nand U6592 (N_6592,N_6131,N_6222);
or U6593 (N_6593,N_6378,N_6379);
xor U6594 (N_6594,N_6319,N_6204);
nand U6595 (N_6595,N_6239,N_6155);
xnor U6596 (N_6596,N_6110,N_6052);
nor U6597 (N_6597,N_6257,N_6079);
and U6598 (N_6598,N_6357,N_6266);
nor U6599 (N_6599,N_6258,N_6334);
nor U6600 (N_6600,N_6052,N_6036);
nand U6601 (N_6601,N_6149,N_6146);
and U6602 (N_6602,N_6157,N_6036);
xor U6603 (N_6603,N_6046,N_6086);
or U6604 (N_6604,N_6108,N_6140);
nand U6605 (N_6605,N_6196,N_6107);
nor U6606 (N_6606,N_6383,N_6347);
or U6607 (N_6607,N_6100,N_6177);
or U6608 (N_6608,N_6099,N_6223);
xor U6609 (N_6609,N_6325,N_6176);
and U6610 (N_6610,N_6328,N_6383);
xnor U6611 (N_6611,N_6038,N_6170);
nor U6612 (N_6612,N_6080,N_6181);
xnor U6613 (N_6613,N_6326,N_6171);
nand U6614 (N_6614,N_6307,N_6352);
and U6615 (N_6615,N_6379,N_6036);
or U6616 (N_6616,N_6259,N_6168);
or U6617 (N_6617,N_6351,N_6186);
nor U6618 (N_6618,N_6375,N_6332);
nor U6619 (N_6619,N_6290,N_6012);
nand U6620 (N_6620,N_6008,N_6158);
nand U6621 (N_6621,N_6156,N_6049);
xor U6622 (N_6622,N_6307,N_6134);
or U6623 (N_6623,N_6363,N_6359);
nand U6624 (N_6624,N_6223,N_6185);
and U6625 (N_6625,N_6378,N_6166);
xnor U6626 (N_6626,N_6162,N_6202);
and U6627 (N_6627,N_6003,N_6036);
xnor U6628 (N_6628,N_6300,N_6180);
nor U6629 (N_6629,N_6380,N_6105);
xor U6630 (N_6630,N_6308,N_6009);
xor U6631 (N_6631,N_6157,N_6073);
and U6632 (N_6632,N_6148,N_6059);
nand U6633 (N_6633,N_6092,N_6330);
nor U6634 (N_6634,N_6204,N_6099);
xor U6635 (N_6635,N_6107,N_6090);
and U6636 (N_6636,N_6094,N_6372);
xor U6637 (N_6637,N_6055,N_6311);
nand U6638 (N_6638,N_6061,N_6359);
nand U6639 (N_6639,N_6334,N_6385);
nand U6640 (N_6640,N_6090,N_6094);
and U6641 (N_6641,N_6190,N_6291);
nor U6642 (N_6642,N_6152,N_6261);
nor U6643 (N_6643,N_6330,N_6109);
nand U6644 (N_6644,N_6201,N_6324);
nor U6645 (N_6645,N_6087,N_6017);
xor U6646 (N_6646,N_6343,N_6235);
nand U6647 (N_6647,N_6275,N_6199);
xor U6648 (N_6648,N_6294,N_6214);
or U6649 (N_6649,N_6356,N_6197);
or U6650 (N_6650,N_6086,N_6113);
and U6651 (N_6651,N_6265,N_6039);
nand U6652 (N_6652,N_6395,N_6352);
nor U6653 (N_6653,N_6248,N_6359);
nand U6654 (N_6654,N_6006,N_6141);
xor U6655 (N_6655,N_6397,N_6343);
or U6656 (N_6656,N_6124,N_6046);
nand U6657 (N_6657,N_6285,N_6329);
and U6658 (N_6658,N_6199,N_6146);
nor U6659 (N_6659,N_6324,N_6264);
nand U6660 (N_6660,N_6141,N_6194);
nor U6661 (N_6661,N_6308,N_6204);
nor U6662 (N_6662,N_6028,N_6201);
nor U6663 (N_6663,N_6368,N_6151);
nand U6664 (N_6664,N_6274,N_6006);
and U6665 (N_6665,N_6258,N_6314);
nand U6666 (N_6666,N_6159,N_6188);
nand U6667 (N_6667,N_6228,N_6295);
and U6668 (N_6668,N_6354,N_6134);
nand U6669 (N_6669,N_6373,N_6010);
xnor U6670 (N_6670,N_6232,N_6373);
xnor U6671 (N_6671,N_6242,N_6185);
or U6672 (N_6672,N_6349,N_6196);
and U6673 (N_6673,N_6069,N_6061);
xnor U6674 (N_6674,N_6201,N_6251);
xor U6675 (N_6675,N_6357,N_6210);
and U6676 (N_6676,N_6362,N_6087);
and U6677 (N_6677,N_6381,N_6399);
or U6678 (N_6678,N_6383,N_6229);
or U6679 (N_6679,N_6278,N_6204);
or U6680 (N_6680,N_6382,N_6236);
or U6681 (N_6681,N_6338,N_6298);
xor U6682 (N_6682,N_6135,N_6098);
nand U6683 (N_6683,N_6288,N_6213);
and U6684 (N_6684,N_6001,N_6164);
or U6685 (N_6685,N_6178,N_6391);
or U6686 (N_6686,N_6339,N_6078);
nor U6687 (N_6687,N_6141,N_6245);
and U6688 (N_6688,N_6045,N_6289);
nand U6689 (N_6689,N_6193,N_6279);
nand U6690 (N_6690,N_6369,N_6261);
nor U6691 (N_6691,N_6337,N_6141);
and U6692 (N_6692,N_6001,N_6324);
nand U6693 (N_6693,N_6205,N_6216);
xor U6694 (N_6694,N_6196,N_6381);
nand U6695 (N_6695,N_6282,N_6215);
nand U6696 (N_6696,N_6343,N_6060);
nor U6697 (N_6697,N_6032,N_6072);
or U6698 (N_6698,N_6383,N_6218);
nand U6699 (N_6699,N_6262,N_6315);
xnor U6700 (N_6700,N_6096,N_6040);
or U6701 (N_6701,N_6345,N_6172);
nor U6702 (N_6702,N_6129,N_6287);
nand U6703 (N_6703,N_6304,N_6033);
xor U6704 (N_6704,N_6031,N_6318);
nor U6705 (N_6705,N_6112,N_6232);
xor U6706 (N_6706,N_6218,N_6138);
or U6707 (N_6707,N_6241,N_6343);
and U6708 (N_6708,N_6233,N_6168);
xor U6709 (N_6709,N_6300,N_6326);
and U6710 (N_6710,N_6039,N_6276);
or U6711 (N_6711,N_6182,N_6356);
nand U6712 (N_6712,N_6273,N_6251);
nor U6713 (N_6713,N_6071,N_6326);
xor U6714 (N_6714,N_6222,N_6012);
and U6715 (N_6715,N_6351,N_6249);
xnor U6716 (N_6716,N_6084,N_6232);
and U6717 (N_6717,N_6112,N_6279);
nor U6718 (N_6718,N_6242,N_6033);
and U6719 (N_6719,N_6170,N_6199);
and U6720 (N_6720,N_6080,N_6141);
or U6721 (N_6721,N_6035,N_6229);
xor U6722 (N_6722,N_6184,N_6113);
and U6723 (N_6723,N_6255,N_6136);
xor U6724 (N_6724,N_6130,N_6364);
xor U6725 (N_6725,N_6352,N_6164);
nand U6726 (N_6726,N_6246,N_6351);
or U6727 (N_6727,N_6117,N_6334);
xor U6728 (N_6728,N_6376,N_6399);
and U6729 (N_6729,N_6252,N_6200);
nand U6730 (N_6730,N_6255,N_6289);
or U6731 (N_6731,N_6350,N_6369);
xor U6732 (N_6732,N_6111,N_6121);
xnor U6733 (N_6733,N_6256,N_6308);
nor U6734 (N_6734,N_6357,N_6293);
and U6735 (N_6735,N_6233,N_6113);
nor U6736 (N_6736,N_6075,N_6067);
nor U6737 (N_6737,N_6091,N_6082);
and U6738 (N_6738,N_6247,N_6221);
nor U6739 (N_6739,N_6368,N_6332);
or U6740 (N_6740,N_6056,N_6154);
xor U6741 (N_6741,N_6284,N_6184);
nor U6742 (N_6742,N_6358,N_6128);
nor U6743 (N_6743,N_6333,N_6043);
or U6744 (N_6744,N_6091,N_6023);
xnor U6745 (N_6745,N_6222,N_6233);
xor U6746 (N_6746,N_6229,N_6233);
nor U6747 (N_6747,N_6390,N_6264);
xnor U6748 (N_6748,N_6347,N_6023);
nor U6749 (N_6749,N_6024,N_6321);
and U6750 (N_6750,N_6099,N_6040);
or U6751 (N_6751,N_6110,N_6107);
nor U6752 (N_6752,N_6236,N_6198);
nand U6753 (N_6753,N_6070,N_6287);
or U6754 (N_6754,N_6035,N_6037);
nor U6755 (N_6755,N_6094,N_6386);
xnor U6756 (N_6756,N_6191,N_6165);
nor U6757 (N_6757,N_6318,N_6084);
nand U6758 (N_6758,N_6022,N_6113);
nand U6759 (N_6759,N_6178,N_6145);
or U6760 (N_6760,N_6252,N_6230);
or U6761 (N_6761,N_6056,N_6130);
xor U6762 (N_6762,N_6319,N_6294);
and U6763 (N_6763,N_6243,N_6190);
xor U6764 (N_6764,N_6048,N_6052);
and U6765 (N_6765,N_6192,N_6324);
xor U6766 (N_6766,N_6070,N_6166);
nor U6767 (N_6767,N_6337,N_6328);
and U6768 (N_6768,N_6089,N_6381);
and U6769 (N_6769,N_6188,N_6279);
nand U6770 (N_6770,N_6083,N_6346);
and U6771 (N_6771,N_6333,N_6233);
nor U6772 (N_6772,N_6372,N_6061);
and U6773 (N_6773,N_6366,N_6255);
and U6774 (N_6774,N_6276,N_6284);
xnor U6775 (N_6775,N_6102,N_6152);
nand U6776 (N_6776,N_6330,N_6300);
nand U6777 (N_6777,N_6061,N_6346);
nor U6778 (N_6778,N_6293,N_6208);
xnor U6779 (N_6779,N_6324,N_6195);
nor U6780 (N_6780,N_6385,N_6179);
nand U6781 (N_6781,N_6095,N_6212);
xnor U6782 (N_6782,N_6112,N_6201);
xnor U6783 (N_6783,N_6054,N_6107);
and U6784 (N_6784,N_6094,N_6258);
or U6785 (N_6785,N_6131,N_6340);
and U6786 (N_6786,N_6096,N_6116);
nor U6787 (N_6787,N_6096,N_6335);
and U6788 (N_6788,N_6372,N_6388);
xor U6789 (N_6789,N_6390,N_6059);
xnor U6790 (N_6790,N_6295,N_6129);
nand U6791 (N_6791,N_6069,N_6259);
xor U6792 (N_6792,N_6057,N_6144);
nor U6793 (N_6793,N_6208,N_6136);
and U6794 (N_6794,N_6090,N_6258);
nor U6795 (N_6795,N_6271,N_6326);
xor U6796 (N_6796,N_6216,N_6141);
or U6797 (N_6797,N_6025,N_6362);
or U6798 (N_6798,N_6222,N_6261);
or U6799 (N_6799,N_6393,N_6221);
or U6800 (N_6800,N_6498,N_6525);
nor U6801 (N_6801,N_6503,N_6576);
nand U6802 (N_6802,N_6603,N_6476);
xor U6803 (N_6803,N_6638,N_6514);
or U6804 (N_6804,N_6686,N_6552);
or U6805 (N_6805,N_6414,N_6444);
xor U6806 (N_6806,N_6559,N_6736);
nor U6807 (N_6807,N_6690,N_6483);
xnor U6808 (N_6808,N_6474,N_6642);
or U6809 (N_6809,N_6423,N_6458);
nand U6810 (N_6810,N_6779,N_6705);
and U6811 (N_6811,N_6477,N_6534);
nor U6812 (N_6812,N_6785,N_6738);
xor U6813 (N_6813,N_6568,N_6680);
nor U6814 (N_6814,N_6772,N_6502);
nand U6815 (N_6815,N_6693,N_6600);
xnor U6816 (N_6816,N_6595,N_6405);
xor U6817 (N_6817,N_6701,N_6530);
nor U6818 (N_6818,N_6579,N_6465);
or U6819 (N_6819,N_6520,N_6415);
xnor U6820 (N_6820,N_6636,N_6781);
or U6821 (N_6821,N_6623,N_6577);
and U6822 (N_6822,N_6681,N_6728);
or U6823 (N_6823,N_6448,N_6446);
or U6824 (N_6824,N_6644,N_6777);
nor U6825 (N_6825,N_6723,N_6548);
nor U6826 (N_6826,N_6511,N_6765);
or U6827 (N_6827,N_6541,N_6729);
xnor U6828 (N_6828,N_6584,N_6747);
nor U6829 (N_6829,N_6773,N_6687);
nor U6830 (N_6830,N_6794,N_6641);
xor U6831 (N_6831,N_6594,N_6732);
nand U6832 (N_6832,N_6752,N_6433);
nor U6833 (N_6833,N_6704,N_6570);
and U6834 (N_6834,N_6425,N_6484);
xor U6835 (N_6835,N_6434,N_6572);
nor U6836 (N_6836,N_6697,N_6605);
and U6837 (N_6837,N_6791,N_6413);
xor U6838 (N_6838,N_6418,N_6515);
or U6839 (N_6839,N_6657,N_6717);
and U6840 (N_6840,N_6479,N_6497);
or U6841 (N_6841,N_6507,N_6582);
and U6842 (N_6842,N_6678,N_6599);
or U6843 (N_6843,N_6506,N_6424);
nand U6844 (N_6844,N_6420,N_6560);
or U6845 (N_6845,N_6755,N_6626);
nor U6846 (N_6846,N_6661,N_6406);
and U6847 (N_6847,N_6537,N_6770);
or U6848 (N_6848,N_6422,N_6783);
and U6849 (N_6849,N_6533,N_6691);
or U6850 (N_6850,N_6574,N_6618);
nor U6851 (N_6851,N_6632,N_6432);
or U6852 (N_6852,N_6653,N_6412);
xnor U6853 (N_6853,N_6768,N_6470);
nand U6854 (N_6854,N_6667,N_6712);
or U6855 (N_6855,N_6524,N_6714);
and U6856 (N_6856,N_6788,N_6656);
xnor U6857 (N_6857,N_6786,N_6513);
nor U6858 (N_6858,N_6663,N_6567);
and U6859 (N_6859,N_6716,N_6437);
and U6860 (N_6860,N_6543,N_6436);
nand U6861 (N_6861,N_6496,N_6692);
nor U6862 (N_6862,N_6608,N_6666);
nand U6863 (N_6863,N_6401,N_6580);
nand U6864 (N_6864,N_6550,N_6419);
and U6865 (N_6865,N_6538,N_6442);
and U6866 (N_6866,N_6759,N_6737);
xor U6867 (N_6867,N_6555,N_6672);
and U6868 (N_6868,N_6761,N_6659);
xor U6869 (N_6869,N_6633,N_6628);
nor U6870 (N_6870,N_6535,N_6492);
xor U6871 (N_6871,N_6546,N_6440);
nor U6872 (N_6872,N_6671,N_6494);
nor U6873 (N_6873,N_6542,N_6665);
or U6874 (N_6874,N_6583,N_6725);
and U6875 (N_6875,N_6733,N_6435);
nor U6876 (N_6876,N_6766,N_6517);
nor U6877 (N_6877,N_6493,N_6673);
nand U6878 (N_6878,N_6464,N_6519);
and U6879 (N_6879,N_6554,N_6764);
nor U6880 (N_6880,N_6463,N_6426);
xor U6881 (N_6881,N_6718,N_6689);
nor U6882 (N_6882,N_6763,N_6526);
or U6883 (N_6883,N_6708,N_6707);
and U6884 (N_6884,N_6604,N_6468);
nand U6885 (N_6885,N_6473,N_6649);
xnor U6886 (N_6886,N_6449,N_6557);
and U6887 (N_6887,N_6450,N_6640);
nor U6888 (N_6888,N_6715,N_6696);
xor U6889 (N_6889,N_6551,N_6549);
and U6890 (N_6890,N_6482,N_6427);
nor U6891 (N_6891,N_6586,N_6590);
and U6892 (N_6892,N_6527,N_6719);
xor U6893 (N_6893,N_6521,N_6578);
or U6894 (N_6894,N_6466,N_6409);
and U6895 (N_6895,N_6411,N_6711);
and U6896 (N_6896,N_6553,N_6784);
xnor U6897 (N_6897,N_6529,N_6795);
or U6898 (N_6898,N_6683,N_6792);
or U6899 (N_6899,N_6778,N_6487);
xnor U6900 (N_6900,N_6634,N_6430);
or U6901 (N_6901,N_6581,N_6695);
nand U6902 (N_6902,N_6756,N_6481);
and U6903 (N_6903,N_6743,N_6652);
xor U6904 (N_6904,N_6757,N_6735);
or U6905 (N_6905,N_6726,N_6565);
nand U6906 (N_6906,N_6739,N_6621);
nand U6907 (N_6907,N_6601,N_6655);
nand U6908 (N_6908,N_6528,N_6563);
and U6909 (N_6909,N_6585,N_6475);
and U6910 (N_6910,N_6721,N_6611);
and U6911 (N_6911,N_6460,N_6616);
and U6912 (N_6912,N_6539,N_6703);
nand U6913 (N_6913,N_6713,N_6421);
and U6914 (N_6914,N_6631,N_6547);
and U6915 (N_6915,N_6485,N_6780);
xor U6916 (N_6916,N_6403,N_6588);
or U6917 (N_6917,N_6540,N_6688);
xor U6918 (N_6918,N_6602,N_6499);
nand U6919 (N_6919,N_6402,N_6461);
or U6920 (N_6920,N_6610,N_6682);
and U6921 (N_6921,N_6478,N_6455);
or U6922 (N_6922,N_6587,N_6769);
nor U6923 (N_6923,N_6408,N_6662);
nor U6924 (N_6924,N_6544,N_6650);
xor U6925 (N_6925,N_6495,N_6531);
nand U6926 (N_6926,N_6516,N_6518);
or U6927 (N_6927,N_6647,N_6431);
or U6928 (N_6928,N_6658,N_6564);
nor U6929 (N_6929,N_6676,N_6654);
and U6930 (N_6930,N_6619,N_6648);
xnor U6931 (N_6931,N_6573,N_6651);
xnor U6932 (N_6932,N_6700,N_6612);
or U6933 (N_6933,N_6740,N_6500);
or U6934 (N_6934,N_6536,N_6722);
nor U6935 (N_6935,N_6710,N_6558);
or U6936 (N_6936,N_6720,N_6767);
or U6937 (N_6937,N_6698,N_6760);
nand U6938 (N_6938,N_6637,N_6614);
and U6939 (N_6939,N_6668,N_6504);
nor U6940 (N_6940,N_6630,N_6694);
and U6941 (N_6941,N_6699,N_6509);
and U6942 (N_6942,N_6569,N_6751);
xnor U6943 (N_6943,N_6742,N_6727);
or U6944 (N_6944,N_6627,N_6645);
nor U6945 (N_6945,N_6472,N_6545);
xnor U6946 (N_6946,N_6488,N_6561);
nand U6947 (N_6947,N_6798,N_6439);
nor U6948 (N_6948,N_6615,N_6684);
nor U6949 (N_6949,N_6454,N_6776);
xnor U6950 (N_6950,N_6591,N_6489);
nor U6951 (N_6951,N_6775,N_6452);
nor U6952 (N_6952,N_6598,N_6746);
or U6953 (N_6953,N_6669,N_6467);
or U6954 (N_6954,N_6753,N_6407);
and U6955 (N_6955,N_6622,N_6575);
or U6956 (N_6956,N_6429,N_6505);
nor U6957 (N_6957,N_6624,N_6709);
or U6958 (N_6958,N_6787,N_6660);
and U6959 (N_6959,N_6731,N_6749);
nor U6960 (N_6960,N_6782,N_6491);
xnor U6961 (N_6961,N_6670,N_6702);
xnor U6962 (N_6962,N_6643,N_6674);
nand U6963 (N_6963,N_6522,N_6750);
xnor U6964 (N_6964,N_6556,N_6571);
xor U6965 (N_6965,N_6469,N_6457);
and U6966 (N_6966,N_6706,N_6593);
nor U6967 (N_6967,N_6617,N_6428);
or U6968 (N_6968,N_6486,N_6607);
and U6969 (N_6969,N_6456,N_6748);
and U6970 (N_6970,N_6620,N_6451);
and U6971 (N_6971,N_6625,N_6741);
nor U6972 (N_6972,N_6532,N_6685);
or U6973 (N_6973,N_6480,N_6459);
nand U6974 (N_6974,N_6445,N_6566);
xor U6975 (N_6975,N_6471,N_6789);
xor U6976 (N_6976,N_6609,N_6562);
nand U6977 (N_6977,N_6416,N_6730);
and U6978 (N_6978,N_6400,N_6596);
xor U6979 (N_6979,N_6597,N_6677);
xnor U6980 (N_6980,N_6510,N_6501);
or U6981 (N_6981,N_6734,N_6724);
xor U6982 (N_6982,N_6675,N_6758);
or U6983 (N_6983,N_6404,N_6438);
nor U6984 (N_6984,N_6797,N_6744);
nor U6985 (N_6985,N_6417,N_6679);
nand U6986 (N_6986,N_6606,N_6441);
xor U6987 (N_6987,N_6646,N_6664);
and U6988 (N_6988,N_6745,N_6774);
nor U6989 (N_6989,N_6613,N_6790);
and U6990 (N_6990,N_6447,N_6754);
xnor U6991 (N_6991,N_6799,N_6490);
and U6992 (N_6992,N_6635,N_6796);
nand U6993 (N_6993,N_6629,N_6592);
nand U6994 (N_6994,N_6512,N_6462);
and U6995 (N_6995,N_6793,N_6508);
nor U6996 (N_6996,N_6639,N_6410);
or U6997 (N_6997,N_6771,N_6589);
nand U6998 (N_6998,N_6453,N_6443);
and U6999 (N_6999,N_6523,N_6762);
nand U7000 (N_7000,N_6789,N_6765);
and U7001 (N_7001,N_6651,N_6654);
nor U7002 (N_7002,N_6595,N_6717);
xor U7003 (N_7003,N_6572,N_6611);
nand U7004 (N_7004,N_6583,N_6655);
nor U7005 (N_7005,N_6743,N_6785);
nor U7006 (N_7006,N_6406,N_6666);
nand U7007 (N_7007,N_6619,N_6471);
nor U7008 (N_7008,N_6460,N_6475);
or U7009 (N_7009,N_6796,N_6716);
or U7010 (N_7010,N_6753,N_6770);
or U7011 (N_7011,N_6659,N_6678);
nand U7012 (N_7012,N_6557,N_6556);
nor U7013 (N_7013,N_6604,N_6608);
nand U7014 (N_7014,N_6699,N_6578);
and U7015 (N_7015,N_6718,N_6694);
xnor U7016 (N_7016,N_6627,N_6780);
or U7017 (N_7017,N_6579,N_6701);
or U7018 (N_7018,N_6410,N_6513);
and U7019 (N_7019,N_6419,N_6490);
nand U7020 (N_7020,N_6773,N_6676);
or U7021 (N_7021,N_6421,N_6753);
and U7022 (N_7022,N_6706,N_6798);
and U7023 (N_7023,N_6684,N_6521);
nand U7024 (N_7024,N_6790,N_6432);
and U7025 (N_7025,N_6415,N_6557);
nor U7026 (N_7026,N_6614,N_6499);
nand U7027 (N_7027,N_6570,N_6525);
or U7028 (N_7028,N_6604,N_6662);
or U7029 (N_7029,N_6609,N_6579);
nor U7030 (N_7030,N_6575,N_6512);
xor U7031 (N_7031,N_6563,N_6668);
nor U7032 (N_7032,N_6640,N_6647);
or U7033 (N_7033,N_6660,N_6466);
and U7034 (N_7034,N_6622,N_6685);
and U7035 (N_7035,N_6680,N_6793);
or U7036 (N_7036,N_6408,N_6570);
nor U7037 (N_7037,N_6718,N_6725);
nand U7038 (N_7038,N_6555,N_6726);
nor U7039 (N_7039,N_6661,N_6667);
or U7040 (N_7040,N_6417,N_6701);
or U7041 (N_7041,N_6627,N_6617);
xnor U7042 (N_7042,N_6520,N_6694);
nand U7043 (N_7043,N_6633,N_6539);
and U7044 (N_7044,N_6741,N_6713);
nand U7045 (N_7045,N_6595,N_6688);
nand U7046 (N_7046,N_6484,N_6691);
nand U7047 (N_7047,N_6455,N_6608);
nor U7048 (N_7048,N_6785,N_6580);
and U7049 (N_7049,N_6464,N_6454);
and U7050 (N_7050,N_6435,N_6713);
nand U7051 (N_7051,N_6688,N_6505);
xor U7052 (N_7052,N_6527,N_6556);
or U7053 (N_7053,N_6525,N_6666);
nor U7054 (N_7054,N_6605,N_6495);
nand U7055 (N_7055,N_6444,N_6630);
or U7056 (N_7056,N_6533,N_6545);
or U7057 (N_7057,N_6752,N_6582);
or U7058 (N_7058,N_6598,N_6769);
nor U7059 (N_7059,N_6441,N_6591);
nor U7060 (N_7060,N_6453,N_6568);
nand U7061 (N_7061,N_6746,N_6626);
and U7062 (N_7062,N_6570,N_6465);
nor U7063 (N_7063,N_6653,N_6455);
xnor U7064 (N_7064,N_6653,N_6663);
nand U7065 (N_7065,N_6713,N_6778);
and U7066 (N_7066,N_6474,N_6490);
nor U7067 (N_7067,N_6695,N_6611);
and U7068 (N_7068,N_6459,N_6493);
nor U7069 (N_7069,N_6714,N_6505);
nand U7070 (N_7070,N_6771,N_6483);
and U7071 (N_7071,N_6704,N_6629);
xnor U7072 (N_7072,N_6773,N_6445);
and U7073 (N_7073,N_6453,N_6629);
or U7074 (N_7074,N_6412,N_6749);
xor U7075 (N_7075,N_6519,N_6521);
xor U7076 (N_7076,N_6768,N_6535);
and U7077 (N_7077,N_6497,N_6491);
nand U7078 (N_7078,N_6634,N_6566);
and U7079 (N_7079,N_6669,N_6786);
nor U7080 (N_7080,N_6643,N_6484);
xor U7081 (N_7081,N_6670,N_6654);
or U7082 (N_7082,N_6606,N_6785);
xor U7083 (N_7083,N_6645,N_6459);
nand U7084 (N_7084,N_6499,N_6506);
or U7085 (N_7085,N_6504,N_6746);
nor U7086 (N_7086,N_6683,N_6426);
nand U7087 (N_7087,N_6648,N_6465);
or U7088 (N_7088,N_6757,N_6510);
nand U7089 (N_7089,N_6787,N_6731);
nor U7090 (N_7090,N_6542,N_6509);
or U7091 (N_7091,N_6729,N_6517);
nor U7092 (N_7092,N_6485,N_6553);
xnor U7093 (N_7093,N_6400,N_6771);
nand U7094 (N_7094,N_6654,N_6644);
nor U7095 (N_7095,N_6599,N_6625);
nor U7096 (N_7096,N_6448,N_6580);
and U7097 (N_7097,N_6709,N_6496);
or U7098 (N_7098,N_6456,N_6729);
xnor U7099 (N_7099,N_6704,N_6681);
and U7100 (N_7100,N_6735,N_6718);
or U7101 (N_7101,N_6702,N_6430);
or U7102 (N_7102,N_6513,N_6750);
nor U7103 (N_7103,N_6573,N_6687);
or U7104 (N_7104,N_6444,N_6652);
and U7105 (N_7105,N_6699,N_6681);
nor U7106 (N_7106,N_6698,N_6706);
nand U7107 (N_7107,N_6634,N_6474);
xnor U7108 (N_7108,N_6700,N_6707);
and U7109 (N_7109,N_6678,N_6469);
xor U7110 (N_7110,N_6457,N_6775);
or U7111 (N_7111,N_6518,N_6689);
xnor U7112 (N_7112,N_6526,N_6747);
or U7113 (N_7113,N_6542,N_6408);
xor U7114 (N_7114,N_6466,N_6491);
nor U7115 (N_7115,N_6646,N_6783);
xor U7116 (N_7116,N_6534,N_6771);
and U7117 (N_7117,N_6571,N_6400);
nand U7118 (N_7118,N_6595,N_6494);
xnor U7119 (N_7119,N_6467,N_6782);
xor U7120 (N_7120,N_6468,N_6493);
or U7121 (N_7121,N_6775,N_6436);
nand U7122 (N_7122,N_6503,N_6773);
or U7123 (N_7123,N_6798,N_6742);
and U7124 (N_7124,N_6596,N_6587);
nor U7125 (N_7125,N_6499,N_6799);
or U7126 (N_7126,N_6668,N_6673);
or U7127 (N_7127,N_6564,N_6543);
or U7128 (N_7128,N_6538,N_6532);
xor U7129 (N_7129,N_6504,N_6530);
nor U7130 (N_7130,N_6461,N_6611);
and U7131 (N_7131,N_6610,N_6650);
nor U7132 (N_7132,N_6658,N_6770);
nand U7133 (N_7133,N_6494,N_6629);
nand U7134 (N_7134,N_6764,N_6502);
or U7135 (N_7135,N_6642,N_6610);
nor U7136 (N_7136,N_6722,N_6681);
nor U7137 (N_7137,N_6401,N_6706);
and U7138 (N_7138,N_6764,N_6624);
xor U7139 (N_7139,N_6714,N_6632);
nor U7140 (N_7140,N_6793,N_6499);
and U7141 (N_7141,N_6678,N_6764);
or U7142 (N_7142,N_6430,N_6669);
xnor U7143 (N_7143,N_6530,N_6471);
xnor U7144 (N_7144,N_6657,N_6532);
and U7145 (N_7145,N_6472,N_6491);
or U7146 (N_7146,N_6527,N_6771);
and U7147 (N_7147,N_6537,N_6442);
xnor U7148 (N_7148,N_6515,N_6679);
xor U7149 (N_7149,N_6736,N_6510);
nand U7150 (N_7150,N_6484,N_6435);
nor U7151 (N_7151,N_6567,N_6619);
nor U7152 (N_7152,N_6511,N_6736);
xor U7153 (N_7153,N_6701,N_6422);
nand U7154 (N_7154,N_6623,N_6637);
nand U7155 (N_7155,N_6627,N_6497);
nor U7156 (N_7156,N_6688,N_6753);
xor U7157 (N_7157,N_6433,N_6703);
nand U7158 (N_7158,N_6462,N_6788);
nor U7159 (N_7159,N_6547,N_6448);
nor U7160 (N_7160,N_6448,N_6404);
xor U7161 (N_7161,N_6573,N_6743);
and U7162 (N_7162,N_6433,N_6693);
xor U7163 (N_7163,N_6619,N_6479);
and U7164 (N_7164,N_6521,N_6568);
nor U7165 (N_7165,N_6410,N_6566);
xor U7166 (N_7166,N_6504,N_6732);
xnor U7167 (N_7167,N_6736,N_6560);
or U7168 (N_7168,N_6635,N_6719);
nor U7169 (N_7169,N_6490,N_6592);
or U7170 (N_7170,N_6777,N_6622);
xnor U7171 (N_7171,N_6452,N_6720);
and U7172 (N_7172,N_6622,N_6551);
and U7173 (N_7173,N_6453,N_6465);
or U7174 (N_7174,N_6595,N_6751);
and U7175 (N_7175,N_6660,N_6544);
xnor U7176 (N_7176,N_6716,N_6525);
nor U7177 (N_7177,N_6637,N_6691);
nor U7178 (N_7178,N_6515,N_6408);
nand U7179 (N_7179,N_6702,N_6766);
or U7180 (N_7180,N_6608,N_6737);
nor U7181 (N_7181,N_6431,N_6776);
xnor U7182 (N_7182,N_6665,N_6797);
nand U7183 (N_7183,N_6666,N_6643);
or U7184 (N_7184,N_6436,N_6526);
nor U7185 (N_7185,N_6607,N_6521);
nand U7186 (N_7186,N_6573,N_6414);
and U7187 (N_7187,N_6603,N_6447);
and U7188 (N_7188,N_6434,N_6588);
nand U7189 (N_7189,N_6513,N_6639);
xnor U7190 (N_7190,N_6488,N_6645);
nor U7191 (N_7191,N_6611,N_6421);
or U7192 (N_7192,N_6413,N_6585);
nor U7193 (N_7193,N_6523,N_6437);
nor U7194 (N_7194,N_6590,N_6663);
or U7195 (N_7195,N_6496,N_6539);
nand U7196 (N_7196,N_6501,N_6482);
nor U7197 (N_7197,N_6435,N_6575);
xor U7198 (N_7198,N_6741,N_6673);
nand U7199 (N_7199,N_6551,N_6649);
xor U7200 (N_7200,N_7166,N_7136);
and U7201 (N_7201,N_7110,N_6885);
nand U7202 (N_7202,N_7133,N_6858);
or U7203 (N_7203,N_7080,N_7098);
nand U7204 (N_7204,N_7118,N_7053);
nor U7205 (N_7205,N_7026,N_7087);
nand U7206 (N_7206,N_6897,N_6844);
and U7207 (N_7207,N_6963,N_7031);
or U7208 (N_7208,N_6909,N_7059);
nand U7209 (N_7209,N_7153,N_6908);
xnor U7210 (N_7210,N_7109,N_7086);
xor U7211 (N_7211,N_6834,N_7128);
or U7212 (N_7212,N_7065,N_6875);
and U7213 (N_7213,N_7008,N_7150);
nand U7214 (N_7214,N_7124,N_7077);
or U7215 (N_7215,N_6949,N_6914);
and U7216 (N_7216,N_7130,N_6887);
nor U7217 (N_7217,N_7148,N_6876);
xnor U7218 (N_7218,N_6978,N_7137);
nor U7219 (N_7219,N_6999,N_7082);
or U7220 (N_7220,N_7127,N_6955);
nand U7221 (N_7221,N_7058,N_6935);
or U7222 (N_7222,N_6830,N_6966);
nand U7223 (N_7223,N_6950,N_6918);
nor U7224 (N_7224,N_6925,N_6855);
and U7225 (N_7225,N_6873,N_6919);
nand U7226 (N_7226,N_6939,N_7171);
and U7227 (N_7227,N_6981,N_6936);
nand U7228 (N_7228,N_7009,N_7186);
nand U7229 (N_7229,N_7091,N_6943);
xor U7230 (N_7230,N_6930,N_7067);
and U7231 (N_7231,N_6849,N_7168);
xnor U7232 (N_7232,N_6945,N_7084);
or U7233 (N_7233,N_7001,N_6920);
xor U7234 (N_7234,N_7043,N_6888);
xor U7235 (N_7235,N_7023,N_7006);
or U7236 (N_7236,N_7047,N_7060);
nand U7237 (N_7237,N_6942,N_7174);
and U7238 (N_7238,N_7126,N_6992);
nor U7239 (N_7239,N_7192,N_7050);
or U7240 (N_7240,N_7167,N_6972);
xnor U7241 (N_7241,N_6804,N_6941);
nand U7242 (N_7242,N_7040,N_6946);
and U7243 (N_7243,N_7030,N_7129);
xor U7244 (N_7244,N_7041,N_6890);
xnor U7245 (N_7245,N_6901,N_6997);
or U7246 (N_7246,N_7072,N_6838);
nand U7247 (N_7247,N_6837,N_7123);
and U7248 (N_7248,N_6889,N_7063);
and U7249 (N_7249,N_6868,N_7048);
or U7250 (N_7250,N_7143,N_6974);
xnor U7251 (N_7251,N_7119,N_7177);
and U7252 (N_7252,N_6952,N_6884);
nand U7253 (N_7253,N_7070,N_6987);
nor U7254 (N_7254,N_6977,N_7011);
xnor U7255 (N_7255,N_7120,N_7134);
nand U7256 (N_7256,N_7022,N_7079);
xor U7257 (N_7257,N_7151,N_7176);
nor U7258 (N_7258,N_6816,N_6864);
and U7259 (N_7259,N_6944,N_6959);
or U7260 (N_7260,N_7092,N_6903);
and U7261 (N_7261,N_6917,N_6988);
and U7262 (N_7262,N_6927,N_6851);
xor U7263 (N_7263,N_7131,N_7090);
xor U7264 (N_7264,N_6926,N_7025);
nor U7265 (N_7265,N_7034,N_7158);
or U7266 (N_7266,N_7096,N_6979);
and U7267 (N_7267,N_6869,N_6835);
nand U7268 (N_7268,N_6986,N_6900);
and U7269 (N_7269,N_7056,N_6863);
xnor U7270 (N_7270,N_6895,N_7154);
xnor U7271 (N_7271,N_6825,N_7042);
and U7272 (N_7272,N_7159,N_7198);
nor U7273 (N_7273,N_7139,N_6847);
nor U7274 (N_7274,N_7036,N_7113);
or U7275 (N_7275,N_6983,N_6993);
and U7276 (N_7276,N_6877,N_6915);
nand U7277 (N_7277,N_6861,N_7175);
nor U7278 (N_7278,N_6848,N_6802);
or U7279 (N_7279,N_7140,N_7102);
or U7280 (N_7280,N_7162,N_7196);
and U7281 (N_7281,N_7097,N_6817);
nand U7282 (N_7282,N_7108,N_6843);
xor U7283 (N_7283,N_6800,N_6934);
and U7284 (N_7284,N_6990,N_7014);
xnor U7285 (N_7285,N_6985,N_6867);
nand U7286 (N_7286,N_7054,N_6836);
xor U7287 (N_7287,N_7019,N_7135);
or U7288 (N_7288,N_7061,N_6961);
xnor U7289 (N_7289,N_6829,N_7142);
nor U7290 (N_7290,N_6809,N_7003);
nor U7291 (N_7291,N_7149,N_6902);
xor U7292 (N_7292,N_7156,N_7094);
or U7293 (N_7293,N_7170,N_6832);
nor U7294 (N_7294,N_7172,N_6883);
xnor U7295 (N_7295,N_6956,N_6938);
and U7296 (N_7296,N_7007,N_7112);
or U7297 (N_7297,N_6906,N_7066);
nor U7298 (N_7298,N_7029,N_6905);
and U7299 (N_7299,N_6904,N_7164);
nor U7300 (N_7300,N_7002,N_6991);
or U7301 (N_7301,N_7138,N_6911);
and U7302 (N_7302,N_6931,N_6968);
nor U7303 (N_7303,N_7116,N_7191);
xor U7304 (N_7304,N_7046,N_6996);
and U7305 (N_7305,N_6912,N_6929);
nand U7306 (N_7306,N_6824,N_7173);
xnor U7307 (N_7307,N_7188,N_7163);
xor U7308 (N_7308,N_6973,N_6880);
or U7309 (N_7309,N_7179,N_7028);
nor U7310 (N_7310,N_6921,N_7106);
and U7311 (N_7311,N_7017,N_6916);
nor U7312 (N_7312,N_6886,N_7044);
xnor U7313 (N_7313,N_7157,N_7181);
nand U7314 (N_7314,N_7012,N_7194);
xnor U7315 (N_7315,N_6962,N_7189);
xnor U7316 (N_7316,N_7104,N_6923);
or U7317 (N_7317,N_7193,N_6805);
nand U7318 (N_7318,N_6913,N_6937);
nor U7319 (N_7319,N_7075,N_7004);
nand U7320 (N_7320,N_6841,N_7085);
or U7321 (N_7321,N_7105,N_7052);
xnor U7322 (N_7322,N_6907,N_7078);
or U7323 (N_7323,N_6980,N_6957);
nand U7324 (N_7324,N_7197,N_7146);
and U7325 (N_7325,N_7184,N_6899);
nand U7326 (N_7326,N_7013,N_6964);
and U7327 (N_7327,N_6967,N_6823);
and U7328 (N_7328,N_6954,N_7101);
nor U7329 (N_7329,N_7027,N_6994);
or U7330 (N_7330,N_6826,N_7111);
xor U7331 (N_7331,N_6860,N_6982);
or U7332 (N_7332,N_7089,N_6828);
or U7333 (N_7333,N_7161,N_7195);
xor U7334 (N_7334,N_6808,N_6958);
nand U7335 (N_7335,N_7064,N_6818);
or U7336 (N_7336,N_6846,N_6928);
and U7337 (N_7337,N_7035,N_7160);
nand U7338 (N_7338,N_7010,N_6839);
xnor U7339 (N_7339,N_7005,N_6821);
nor U7340 (N_7340,N_6891,N_6801);
or U7341 (N_7341,N_7199,N_6813);
nor U7342 (N_7342,N_6810,N_7185);
or U7343 (N_7343,N_6998,N_6984);
xor U7344 (N_7344,N_7055,N_6833);
nor U7345 (N_7345,N_6893,N_6910);
and U7346 (N_7346,N_7093,N_6976);
or U7347 (N_7347,N_7107,N_7016);
nor U7348 (N_7348,N_6862,N_7068);
xnor U7349 (N_7349,N_7057,N_6866);
nand U7350 (N_7350,N_6953,N_6857);
nor U7351 (N_7351,N_7178,N_7121);
or U7352 (N_7352,N_7020,N_6853);
or U7353 (N_7353,N_6940,N_6859);
or U7354 (N_7354,N_6819,N_7018);
nor U7355 (N_7355,N_6881,N_6814);
nor U7356 (N_7356,N_6995,N_6827);
and U7357 (N_7357,N_6822,N_6882);
nor U7358 (N_7358,N_7122,N_6850);
xor U7359 (N_7359,N_7076,N_7147);
xnor U7360 (N_7360,N_6879,N_7152);
nand U7361 (N_7361,N_6871,N_7169);
nand U7362 (N_7362,N_6806,N_6845);
nor U7363 (N_7363,N_6856,N_7038);
and U7364 (N_7364,N_7190,N_6870);
nor U7365 (N_7365,N_7039,N_7095);
and U7366 (N_7366,N_7037,N_6807);
or U7367 (N_7367,N_7081,N_6922);
or U7368 (N_7368,N_6989,N_7132);
xnor U7369 (N_7369,N_7144,N_6803);
nand U7370 (N_7370,N_6820,N_6947);
nand U7371 (N_7371,N_7099,N_7115);
nor U7372 (N_7372,N_6896,N_7141);
or U7373 (N_7373,N_6894,N_6812);
xnor U7374 (N_7374,N_7083,N_6960);
nand U7375 (N_7375,N_6840,N_6951);
or U7376 (N_7376,N_7074,N_7145);
and U7377 (N_7377,N_7187,N_6852);
and U7378 (N_7378,N_7103,N_6811);
nand U7379 (N_7379,N_6965,N_7049);
nand U7380 (N_7380,N_6898,N_7021);
or U7381 (N_7381,N_6975,N_6969);
and U7382 (N_7382,N_7114,N_7183);
and U7383 (N_7383,N_6878,N_7033);
nor U7384 (N_7384,N_6872,N_6932);
xnor U7385 (N_7385,N_7062,N_6933);
or U7386 (N_7386,N_7015,N_6970);
or U7387 (N_7387,N_6971,N_7100);
nor U7388 (N_7388,N_6892,N_7155);
xnor U7389 (N_7389,N_7071,N_6842);
nor U7390 (N_7390,N_7069,N_6948);
xor U7391 (N_7391,N_7117,N_7165);
xnor U7392 (N_7392,N_7088,N_6865);
nand U7393 (N_7393,N_6854,N_7051);
or U7394 (N_7394,N_7000,N_6815);
nor U7395 (N_7395,N_6874,N_7024);
nand U7396 (N_7396,N_6924,N_7032);
xor U7397 (N_7397,N_7125,N_6831);
or U7398 (N_7398,N_7073,N_7180);
xor U7399 (N_7399,N_7182,N_7045);
nor U7400 (N_7400,N_7171,N_6912);
and U7401 (N_7401,N_6849,N_6982);
xor U7402 (N_7402,N_7095,N_7156);
nor U7403 (N_7403,N_7102,N_7101);
nor U7404 (N_7404,N_7194,N_6954);
nor U7405 (N_7405,N_7149,N_6891);
and U7406 (N_7406,N_6853,N_7156);
xnor U7407 (N_7407,N_7054,N_6893);
or U7408 (N_7408,N_7137,N_6911);
xor U7409 (N_7409,N_7146,N_7193);
and U7410 (N_7410,N_6826,N_6971);
or U7411 (N_7411,N_6883,N_6863);
xnor U7412 (N_7412,N_7008,N_7028);
or U7413 (N_7413,N_7057,N_7012);
nor U7414 (N_7414,N_7126,N_7156);
nand U7415 (N_7415,N_7099,N_6836);
and U7416 (N_7416,N_6921,N_7143);
nor U7417 (N_7417,N_6867,N_7176);
xor U7418 (N_7418,N_7072,N_6874);
nor U7419 (N_7419,N_7016,N_7141);
and U7420 (N_7420,N_6900,N_7138);
or U7421 (N_7421,N_6936,N_6925);
nand U7422 (N_7422,N_6918,N_6969);
or U7423 (N_7423,N_7091,N_6956);
and U7424 (N_7424,N_6944,N_7124);
and U7425 (N_7425,N_7019,N_7156);
nand U7426 (N_7426,N_6851,N_6921);
or U7427 (N_7427,N_6852,N_7137);
nor U7428 (N_7428,N_6909,N_7115);
nor U7429 (N_7429,N_6897,N_7000);
nand U7430 (N_7430,N_7029,N_7193);
nand U7431 (N_7431,N_6977,N_6976);
nand U7432 (N_7432,N_7007,N_7170);
nor U7433 (N_7433,N_6832,N_7115);
and U7434 (N_7434,N_7147,N_7009);
or U7435 (N_7435,N_6986,N_7151);
xor U7436 (N_7436,N_6998,N_6876);
nand U7437 (N_7437,N_7136,N_6884);
and U7438 (N_7438,N_6856,N_7063);
or U7439 (N_7439,N_7199,N_6954);
or U7440 (N_7440,N_6817,N_6851);
nand U7441 (N_7441,N_6959,N_7183);
xor U7442 (N_7442,N_6904,N_6868);
or U7443 (N_7443,N_7130,N_7098);
nand U7444 (N_7444,N_6965,N_6816);
xor U7445 (N_7445,N_7120,N_7140);
and U7446 (N_7446,N_6981,N_6865);
or U7447 (N_7447,N_7172,N_7197);
xnor U7448 (N_7448,N_7001,N_6901);
nor U7449 (N_7449,N_6949,N_6992);
or U7450 (N_7450,N_6927,N_7195);
and U7451 (N_7451,N_6937,N_7002);
or U7452 (N_7452,N_6861,N_6959);
and U7453 (N_7453,N_7016,N_6955);
nor U7454 (N_7454,N_7186,N_7135);
nand U7455 (N_7455,N_6964,N_6991);
and U7456 (N_7456,N_7057,N_6954);
or U7457 (N_7457,N_7031,N_7159);
and U7458 (N_7458,N_7084,N_6911);
and U7459 (N_7459,N_6955,N_7177);
or U7460 (N_7460,N_7022,N_7151);
xnor U7461 (N_7461,N_6828,N_7067);
and U7462 (N_7462,N_6800,N_7188);
nand U7463 (N_7463,N_7189,N_7023);
nor U7464 (N_7464,N_6833,N_6929);
and U7465 (N_7465,N_7073,N_6936);
nand U7466 (N_7466,N_6973,N_7018);
nor U7467 (N_7467,N_7030,N_7193);
nor U7468 (N_7468,N_7108,N_6978);
nand U7469 (N_7469,N_6952,N_7051);
nand U7470 (N_7470,N_6875,N_6819);
or U7471 (N_7471,N_7026,N_7013);
xnor U7472 (N_7472,N_7173,N_7012);
xor U7473 (N_7473,N_6844,N_7142);
xnor U7474 (N_7474,N_6863,N_7097);
nor U7475 (N_7475,N_6898,N_7042);
or U7476 (N_7476,N_6809,N_6808);
or U7477 (N_7477,N_6905,N_6930);
and U7478 (N_7478,N_7042,N_7029);
nor U7479 (N_7479,N_6983,N_7068);
or U7480 (N_7480,N_7136,N_7062);
nor U7481 (N_7481,N_6953,N_7024);
nand U7482 (N_7482,N_7080,N_6916);
xnor U7483 (N_7483,N_7073,N_7000);
nor U7484 (N_7484,N_6880,N_6848);
xnor U7485 (N_7485,N_6909,N_7175);
nand U7486 (N_7486,N_7012,N_6883);
or U7487 (N_7487,N_7016,N_6971);
and U7488 (N_7488,N_7070,N_6912);
nor U7489 (N_7489,N_7139,N_7179);
or U7490 (N_7490,N_7170,N_6843);
nor U7491 (N_7491,N_7110,N_6900);
and U7492 (N_7492,N_6890,N_7054);
xnor U7493 (N_7493,N_6905,N_6980);
xnor U7494 (N_7494,N_6805,N_6860);
nand U7495 (N_7495,N_6945,N_7103);
or U7496 (N_7496,N_6897,N_6809);
and U7497 (N_7497,N_6922,N_7054);
and U7498 (N_7498,N_6932,N_7150);
xor U7499 (N_7499,N_6857,N_7003);
nor U7500 (N_7500,N_7118,N_7005);
nand U7501 (N_7501,N_6828,N_7127);
nor U7502 (N_7502,N_6947,N_6955);
nor U7503 (N_7503,N_6955,N_7010);
and U7504 (N_7504,N_7176,N_7199);
and U7505 (N_7505,N_6934,N_7019);
xnor U7506 (N_7506,N_7002,N_7198);
and U7507 (N_7507,N_6806,N_6890);
and U7508 (N_7508,N_7124,N_7123);
nor U7509 (N_7509,N_6816,N_7073);
nor U7510 (N_7510,N_7066,N_7027);
xor U7511 (N_7511,N_7061,N_7104);
nand U7512 (N_7512,N_7064,N_7022);
nor U7513 (N_7513,N_7055,N_7115);
nor U7514 (N_7514,N_6953,N_6811);
or U7515 (N_7515,N_7031,N_7044);
nor U7516 (N_7516,N_6834,N_6925);
xor U7517 (N_7517,N_6809,N_7094);
nand U7518 (N_7518,N_6829,N_7092);
xnor U7519 (N_7519,N_6829,N_7007);
nand U7520 (N_7520,N_7124,N_6976);
or U7521 (N_7521,N_6902,N_7198);
nor U7522 (N_7522,N_6903,N_6998);
or U7523 (N_7523,N_7120,N_6833);
nand U7524 (N_7524,N_6996,N_6857);
nor U7525 (N_7525,N_7149,N_6984);
nand U7526 (N_7526,N_7044,N_6931);
xnor U7527 (N_7527,N_7085,N_7055);
or U7528 (N_7528,N_7197,N_6826);
and U7529 (N_7529,N_6863,N_6845);
or U7530 (N_7530,N_6860,N_6960);
xor U7531 (N_7531,N_6969,N_7032);
or U7532 (N_7532,N_7021,N_7111);
and U7533 (N_7533,N_6827,N_7159);
and U7534 (N_7534,N_7172,N_7103);
xor U7535 (N_7535,N_7153,N_6854);
or U7536 (N_7536,N_7174,N_7156);
or U7537 (N_7537,N_7110,N_6952);
and U7538 (N_7538,N_6919,N_7190);
or U7539 (N_7539,N_6831,N_6839);
and U7540 (N_7540,N_6860,N_6884);
or U7541 (N_7541,N_6873,N_6888);
or U7542 (N_7542,N_7072,N_6815);
or U7543 (N_7543,N_7007,N_7197);
and U7544 (N_7544,N_6993,N_6937);
nor U7545 (N_7545,N_7120,N_7090);
nor U7546 (N_7546,N_7191,N_7172);
nor U7547 (N_7547,N_6958,N_7083);
and U7548 (N_7548,N_6873,N_7016);
or U7549 (N_7549,N_6824,N_6889);
nand U7550 (N_7550,N_7053,N_7189);
xnor U7551 (N_7551,N_7140,N_6893);
nor U7552 (N_7552,N_6847,N_7181);
or U7553 (N_7553,N_6987,N_7017);
and U7554 (N_7554,N_7123,N_7026);
nand U7555 (N_7555,N_7108,N_6970);
xnor U7556 (N_7556,N_6902,N_6846);
xor U7557 (N_7557,N_6883,N_7001);
and U7558 (N_7558,N_6945,N_7198);
nand U7559 (N_7559,N_6811,N_6980);
xor U7560 (N_7560,N_7192,N_7079);
or U7561 (N_7561,N_7166,N_6971);
or U7562 (N_7562,N_7011,N_7064);
nor U7563 (N_7563,N_7089,N_7127);
nand U7564 (N_7564,N_6821,N_7176);
nor U7565 (N_7565,N_7112,N_7012);
nor U7566 (N_7566,N_7082,N_6823);
and U7567 (N_7567,N_7008,N_7016);
or U7568 (N_7568,N_7000,N_7123);
and U7569 (N_7569,N_7032,N_7156);
and U7570 (N_7570,N_7036,N_6835);
or U7571 (N_7571,N_6847,N_6916);
and U7572 (N_7572,N_6806,N_7108);
xor U7573 (N_7573,N_7021,N_6850);
nand U7574 (N_7574,N_7079,N_6935);
nor U7575 (N_7575,N_6822,N_6808);
and U7576 (N_7576,N_6909,N_6938);
xor U7577 (N_7577,N_7157,N_6930);
or U7578 (N_7578,N_7186,N_6836);
xor U7579 (N_7579,N_6820,N_6929);
or U7580 (N_7580,N_6802,N_7173);
nand U7581 (N_7581,N_7161,N_6853);
nand U7582 (N_7582,N_7136,N_7038);
xor U7583 (N_7583,N_6866,N_7030);
and U7584 (N_7584,N_7044,N_7003);
nand U7585 (N_7585,N_6902,N_6913);
or U7586 (N_7586,N_7066,N_7050);
xnor U7587 (N_7587,N_7127,N_6819);
nor U7588 (N_7588,N_6994,N_6827);
nand U7589 (N_7589,N_6935,N_7080);
xor U7590 (N_7590,N_7066,N_6805);
xnor U7591 (N_7591,N_6924,N_7184);
nor U7592 (N_7592,N_6955,N_7017);
and U7593 (N_7593,N_6854,N_7182);
xnor U7594 (N_7594,N_7146,N_7144);
and U7595 (N_7595,N_6899,N_6910);
xnor U7596 (N_7596,N_7135,N_7198);
xnor U7597 (N_7597,N_7134,N_6822);
nor U7598 (N_7598,N_7053,N_6810);
and U7599 (N_7599,N_6867,N_7011);
xnor U7600 (N_7600,N_7275,N_7413);
and U7601 (N_7601,N_7415,N_7438);
nor U7602 (N_7602,N_7260,N_7297);
xor U7603 (N_7603,N_7398,N_7435);
or U7604 (N_7604,N_7540,N_7311);
nand U7605 (N_7605,N_7556,N_7344);
or U7606 (N_7606,N_7478,N_7386);
and U7607 (N_7607,N_7256,N_7347);
nand U7608 (N_7608,N_7566,N_7425);
and U7609 (N_7609,N_7531,N_7414);
nand U7610 (N_7610,N_7244,N_7302);
and U7611 (N_7611,N_7561,N_7591);
nand U7612 (N_7612,N_7376,N_7358);
xor U7613 (N_7613,N_7221,N_7384);
nand U7614 (N_7614,N_7286,N_7322);
nand U7615 (N_7615,N_7563,N_7545);
or U7616 (N_7616,N_7580,N_7465);
nand U7617 (N_7617,N_7573,N_7250);
nand U7618 (N_7618,N_7208,N_7459);
xor U7619 (N_7619,N_7220,N_7292);
xor U7620 (N_7620,N_7535,N_7536);
nand U7621 (N_7621,N_7254,N_7530);
and U7622 (N_7622,N_7417,N_7326);
and U7623 (N_7623,N_7330,N_7232);
and U7624 (N_7624,N_7258,N_7323);
nand U7625 (N_7625,N_7419,N_7240);
xnor U7626 (N_7626,N_7389,N_7225);
and U7627 (N_7627,N_7441,N_7482);
and U7628 (N_7628,N_7215,N_7248);
and U7629 (N_7629,N_7271,N_7495);
nand U7630 (N_7630,N_7255,N_7328);
xnor U7631 (N_7631,N_7372,N_7367);
nor U7632 (N_7632,N_7557,N_7310);
and U7633 (N_7633,N_7370,N_7381);
xnor U7634 (N_7634,N_7309,N_7498);
or U7635 (N_7635,N_7444,N_7526);
xor U7636 (N_7636,N_7568,N_7351);
nand U7637 (N_7637,N_7385,N_7296);
nand U7638 (N_7638,N_7513,N_7587);
or U7639 (N_7639,N_7393,N_7507);
nand U7640 (N_7640,N_7265,N_7246);
and U7641 (N_7641,N_7518,N_7219);
nor U7642 (N_7642,N_7598,N_7327);
nand U7643 (N_7643,N_7445,N_7333);
xor U7644 (N_7644,N_7509,N_7424);
or U7645 (N_7645,N_7457,N_7592);
or U7646 (N_7646,N_7234,N_7289);
and U7647 (N_7647,N_7453,N_7353);
xor U7648 (N_7648,N_7581,N_7588);
nand U7649 (N_7649,N_7325,N_7269);
nand U7650 (N_7650,N_7470,N_7456);
xnor U7651 (N_7651,N_7510,N_7348);
nand U7652 (N_7652,N_7550,N_7437);
xnor U7653 (N_7653,N_7501,N_7368);
xor U7654 (N_7654,N_7516,N_7281);
xor U7655 (N_7655,N_7253,N_7524);
nor U7656 (N_7656,N_7489,N_7318);
nor U7657 (N_7657,N_7541,N_7506);
nor U7658 (N_7658,N_7469,N_7231);
nor U7659 (N_7659,N_7484,N_7412);
nor U7660 (N_7660,N_7223,N_7446);
xnor U7661 (N_7661,N_7512,N_7373);
or U7662 (N_7662,N_7502,N_7527);
or U7663 (N_7663,N_7483,N_7547);
xor U7664 (N_7664,N_7418,N_7555);
nor U7665 (N_7665,N_7490,N_7500);
nand U7666 (N_7666,N_7316,N_7324);
and U7667 (N_7667,N_7434,N_7369);
nor U7668 (N_7668,N_7451,N_7543);
nor U7669 (N_7669,N_7315,N_7411);
xor U7670 (N_7670,N_7525,N_7241);
xor U7671 (N_7671,N_7596,N_7280);
or U7672 (N_7672,N_7522,N_7511);
nand U7673 (N_7673,N_7577,N_7239);
xor U7674 (N_7674,N_7338,N_7494);
nor U7675 (N_7675,N_7242,N_7421);
nor U7676 (N_7676,N_7211,N_7546);
and U7677 (N_7677,N_7339,N_7493);
and U7678 (N_7678,N_7397,N_7375);
nand U7679 (N_7679,N_7554,N_7464);
or U7680 (N_7680,N_7475,N_7204);
nand U7681 (N_7681,N_7343,N_7477);
xor U7682 (N_7682,N_7593,N_7450);
nand U7683 (N_7683,N_7471,N_7481);
xor U7684 (N_7684,N_7340,N_7583);
and U7685 (N_7685,N_7491,N_7431);
or U7686 (N_7686,N_7449,N_7523);
xnor U7687 (N_7687,N_7294,N_7274);
or U7688 (N_7688,N_7429,N_7301);
nor U7689 (N_7689,N_7436,N_7420);
xnor U7690 (N_7690,N_7261,N_7224);
and U7691 (N_7691,N_7454,N_7564);
nor U7692 (N_7692,N_7277,N_7486);
and U7693 (N_7693,N_7589,N_7216);
xor U7694 (N_7694,N_7466,N_7217);
and U7695 (N_7695,N_7538,N_7395);
xnor U7696 (N_7696,N_7503,N_7366);
nor U7697 (N_7697,N_7440,N_7514);
nand U7698 (N_7698,N_7562,N_7226);
xor U7699 (N_7699,N_7342,N_7262);
xor U7700 (N_7700,N_7350,N_7205);
or U7701 (N_7701,N_7227,N_7291);
nor U7702 (N_7702,N_7505,N_7213);
and U7703 (N_7703,N_7359,N_7508);
and U7704 (N_7704,N_7365,N_7249);
nand U7705 (N_7705,N_7480,N_7448);
nor U7706 (N_7706,N_7492,N_7442);
and U7707 (N_7707,N_7408,N_7474);
and U7708 (N_7708,N_7599,N_7243);
nand U7709 (N_7709,N_7569,N_7409);
xor U7710 (N_7710,N_7559,N_7595);
nor U7711 (N_7711,N_7264,N_7357);
or U7712 (N_7712,N_7214,N_7218);
or U7713 (N_7713,N_7272,N_7594);
xor U7714 (N_7714,N_7346,N_7496);
or U7715 (N_7715,N_7430,N_7364);
nand U7716 (N_7716,N_7273,N_7532);
nand U7717 (N_7717,N_7497,N_7251);
or U7718 (N_7718,N_7206,N_7553);
nor U7719 (N_7719,N_7304,N_7293);
xnor U7720 (N_7720,N_7319,N_7299);
or U7721 (N_7721,N_7487,N_7352);
and U7722 (N_7722,N_7401,N_7383);
xor U7723 (N_7723,N_7229,N_7537);
and U7724 (N_7724,N_7329,N_7499);
nor U7725 (N_7725,N_7578,N_7377);
xnor U7726 (N_7726,N_7282,N_7228);
and U7727 (N_7727,N_7472,N_7290);
and U7728 (N_7728,N_7402,N_7378);
nand U7729 (N_7729,N_7267,N_7485);
nand U7730 (N_7730,N_7300,N_7572);
xor U7731 (N_7731,N_7355,N_7519);
nand U7732 (N_7732,N_7288,N_7374);
xnor U7733 (N_7733,N_7207,N_7461);
nand U7734 (N_7734,N_7576,N_7257);
nand U7735 (N_7735,N_7210,N_7529);
nor U7736 (N_7736,N_7548,N_7400);
and U7737 (N_7737,N_7458,N_7387);
and U7738 (N_7738,N_7380,N_7321);
xnor U7739 (N_7739,N_7452,N_7287);
or U7740 (N_7740,N_7590,N_7479);
nand U7741 (N_7741,N_7520,N_7295);
xor U7742 (N_7742,N_7201,N_7468);
or U7743 (N_7743,N_7432,N_7423);
nand U7744 (N_7744,N_7396,N_7579);
nor U7745 (N_7745,N_7200,N_7575);
xnor U7746 (N_7746,N_7504,N_7570);
xnor U7747 (N_7747,N_7305,N_7433);
and U7748 (N_7748,N_7574,N_7331);
and U7749 (N_7749,N_7391,N_7533);
or U7750 (N_7750,N_7382,N_7460);
xnor U7751 (N_7751,N_7335,N_7360);
nor U7752 (N_7752,N_7404,N_7422);
and U7753 (N_7753,N_7266,N_7317);
or U7754 (N_7754,N_7259,N_7416);
nor U7755 (N_7755,N_7515,N_7551);
or U7756 (N_7756,N_7586,N_7285);
or U7757 (N_7757,N_7361,N_7270);
or U7758 (N_7758,N_7447,N_7332);
nor U7759 (N_7759,N_7263,N_7279);
and U7760 (N_7760,N_7276,N_7582);
and U7761 (N_7761,N_7426,N_7284);
nor U7762 (N_7762,N_7356,N_7209);
or U7763 (N_7763,N_7394,N_7565);
and U7764 (N_7764,N_7307,N_7406);
and U7765 (N_7765,N_7467,N_7403);
and U7766 (N_7766,N_7283,N_7390);
and U7767 (N_7767,N_7410,N_7462);
xnor U7768 (N_7768,N_7363,N_7362);
or U7769 (N_7769,N_7314,N_7354);
nor U7770 (N_7770,N_7236,N_7476);
nor U7771 (N_7771,N_7528,N_7407);
nor U7772 (N_7772,N_7312,N_7571);
and U7773 (N_7773,N_7298,N_7203);
nor U7774 (N_7774,N_7278,N_7245);
xor U7775 (N_7775,N_7560,N_7534);
or U7776 (N_7776,N_7371,N_7345);
xnor U7777 (N_7777,N_7388,N_7230);
or U7778 (N_7778,N_7336,N_7584);
or U7779 (N_7779,N_7399,N_7549);
and U7780 (N_7780,N_7268,N_7567);
or U7781 (N_7781,N_7334,N_7558);
xnor U7782 (N_7782,N_7379,N_7544);
xor U7783 (N_7783,N_7222,N_7542);
nor U7784 (N_7784,N_7585,N_7443);
nor U7785 (N_7785,N_7463,N_7439);
and U7786 (N_7786,N_7337,N_7247);
and U7787 (N_7787,N_7517,N_7552);
nor U7788 (N_7788,N_7473,N_7212);
or U7789 (N_7789,N_7303,N_7235);
or U7790 (N_7790,N_7488,N_7320);
and U7791 (N_7791,N_7237,N_7308);
and U7792 (N_7792,N_7597,N_7539);
and U7793 (N_7793,N_7428,N_7427);
or U7794 (N_7794,N_7392,N_7349);
nor U7795 (N_7795,N_7455,N_7405);
nor U7796 (N_7796,N_7521,N_7341);
nand U7797 (N_7797,N_7202,N_7233);
nand U7798 (N_7798,N_7306,N_7238);
or U7799 (N_7799,N_7313,N_7252);
xor U7800 (N_7800,N_7232,N_7372);
nand U7801 (N_7801,N_7514,N_7422);
nand U7802 (N_7802,N_7469,N_7447);
xor U7803 (N_7803,N_7314,N_7279);
xnor U7804 (N_7804,N_7314,N_7455);
nor U7805 (N_7805,N_7519,N_7526);
xor U7806 (N_7806,N_7412,N_7303);
nand U7807 (N_7807,N_7392,N_7227);
and U7808 (N_7808,N_7367,N_7566);
nor U7809 (N_7809,N_7344,N_7358);
xnor U7810 (N_7810,N_7364,N_7524);
nor U7811 (N_7811,N_7317,N_7254);
or U7812 (N_7812,N_7548,N_7498);
nor U7813 (N_7813,N_7366,N_7484);
xnor U7814 (N_7814,N_7519,N_7201);
nand U7815 (N_7815,N_7470,N_7366);
and U7816 (N_7816,N_7299,N_7434);
or U7817 (N_7817,N_7246,N_7596);
or U7818 (N_7818,N_7403,N_7517);
nor U7819 (N_7819,N_7444,N_7454);
nand U7820 (N_7820,N_7222,N_7583);
nand U7821 (N_7821,N_7424,N_7477);
nor U7822 (N_7822,N_7321,N_7489);
xnor U7823 (N_7823,N_7423,N_7404);
and U7824 (N_7824,N_7358,N_7521);
and U7825 (N_7825,N_7406,N_7440);
xnor U7826 (N_7826,N_7535,N_7581);
or U7827 (N_7827,N_7479,N_7276);
xnor U7828 (N_7828,N_7312,N_7215);
and U7829 (N_7829,N_7247,N_7410);
nor U7830 (N_7830,N_7535,N_7334);
nand U7831 (N_7831,N_7279,N_7216);
and U7832 (N_7832,N_7206,N_7366);
nor U7833 (N_7833,N_7311,N_7442);
or U7834 (N_7834,N_7209,N_7316);
nor U7835 (N_7835,N_7286,N_7366);
xor U7836 (N_7836,N_7398,N_7552);
nand U7837 (N_7837,N_7444,N_7285);
nor U7838 (N_7838,N_7354,N_7523);
or U7839 (N_7839,N_7442,N_7374);
nor U7840 (N_7840,N_7410,N_7221);
xnor U7841 (N_7841,N_7472,N_7309);
or U7842 (N_7842,N_7317,N_7544);
nand U7843 (N_7843,N_7375,N_7441);
nor U7844 (N_7844,N_7324,N_7467);
and U7845 (N_7845,N_7342,N_7261);
nor U7846 (N_7846,N_7568,N_7488);
nor U7847 (N_7847,N_7541,N_7210);
and U7848 (N_7848,N_7287,N_7464);
and U7849 (N_7849,N_7508,N_7376);
and U7850 (N_7850,N_7380,N_7356);
nor U7851 (N_7851,N_7202,N_7278);
nor U7852 (N_7852,N_7310,N_7416);
nand U7853 (N_7853,N_7479,N_7580);
xnor U7854 (N_7854,N_7384,N_7406);
nor U7855 (N_7855,N_7278,N_7350);
nor U7856 (N_7856,N_7353,N_7228);
nand U7857 (N_7857,N_7418,N_7500);
or U7858 (N_7858,N_7269,N_7555);
nand U7859 (N_7859,N_7508,N_7588);
xnor U7860 (N_7860,N_7248,N_7276);
nand U7861 (N_7861,N_7404,N_7582);
or U7862 (N_7862,N_7316,N_7491);
nand U7863 (N_7863,N_7550,N_7312);
and U7864 (N_7864,N_7284,N_7353);
xnor U7865 (N_7865,N_7565,N_7287);
nand U7866 (N_7866,N_7531,N_7570);
and U7867 (N_7867,N_7585,N_7209);
xor U7868 (N_7868,N_7572,N_7514);
xnor U7869 (N_7869,N_7294,N_7450);
and U7870 (N_7870,N_7575,N_7492);
nand U7871 (N_7871,N_7330,N_7514);
or U7872 (N_7872,N_7264,N_7439);
xor U7873 (N_7873,N_7430,N_7394);
xor U7874 (N_7874,N_7365,N_7414);
xor U7875 (N_7875,N_7556,N_7310);
nor U7876 (N_7876,N_7225,N_7449);
nor U7877 (N_7877,N_7249,N_7302);
xnor U7878 (N_7878,N_7495,N_7242);
or U7879 (N_7879,N_7244,N_7355);
and U7880 (N_7880,N_7570,N_7518);
and U7881 (N_7881,N_7241,N_7461);
xor U7882 (N_7882,N_7239,N_7291);
nor U7883 (N_7883,N_7247,N_7294);
xnor U7884 (N_7884,N_7254,N_7393);
and U7885 (N_7885,N_7263,N_7492);
nor U7886 (N_7886,N_7420,N_7504);
nor U7887 (N_7887,N_7207,N_7405);
xnor U7888 (N_7888,N_7382,N_7395);
and U7889 (N_7889,N_7549,N_7447);
nor U7890 (N_7890,N_7402,N_7502);
xnor U7891 (N_7891,N_7470,N_7494);
and U7892 (N_7892,N_7478,N_7512);
or U7893 (N_7893,N_7407,N_7380);
xor U7894 (N_7894,N_7229,N_7571);
nand U7895 (N_7895,N_7335,N_7292);
or U7896 (N_7896,N_7204,N_7353);
nand U7897 (N_7897,N_7218,N_7342);
xor U7898 (N_7898,N_7586,N_7569);
and U7899 (N_7899,N_7477,N_7599);
or U7900 (N_7900,N_7308,N_7344);
nor U7901 (N_7901,N_7553,N_7494);
nor U7902 (N_7902,N_7201,N_7246);
nand U7903 (N_7903,N_7206,N_7497);
nand U7904 (N_7904,N_7263,N_7252);
xor U7905 (N_7905,N_7356,N_7491);
nor U7906 (N_7906,N_7365,N_7517);
or U7907 (N_7907,N_7284,N_7263);
or U7908 (N_7908,N_7421,N_7314);
nand U7909 (N_7909,N_7206,N_7260);
or U7910 (N_7910,N_7283,N_7296);
nand U7911 (N_7911,N_7403,N_7339);
and U7912 (N_7912,N_7483,N_7300);
and U7913 (N_7913,N_7410,N_7238);
or U7914 (N_7914,N_7512,N_7405);
nor U7915 (N_7915,N_7358,N_7292);
nand U7916 (N_7916,N_7420,N_7448);
and U7917 (N_7917,N_7385,N_7325);
xor U7918 (N_7918,N_7203,N_7347);
xnor U7919 (N_7919,N_7556,N_7228);
or U7920 (N_7920,N_7288,N_7471);
xor U7921 (N_7921,N_7230,N_7460);
nor U7922 (N_7922,N_7527,N_7238);
nor U7923 (N_7923,N_7296,N_7343);
xor U7924 (N_7924,N_7475,N_7566);
nor U7925 (N_7925,N_7318,N_7471);
xor U7926 (N_7926,N_7468,N_7205);
nor U7927 (N_7927,N_7339,N_7473);
nand U7928 (N_7928,N_7452,N_7461);
nand U7929 (N_7929,N_7372,N_7373);
nor U7930 (N_7930,N_7548,N_7237);
and U7931 (N_7931,N_7578,N_7328);
xor U7932 (N_7932,N_7392,N_7515);
or U7933 (N_7933,N_7444,N_7321);
nand U7934 (N_7934,N_7275,N_7420);
nor U7935 (N_7935,N_7395,N_7497);
or U7936 (N_7936,N_7375,N_7369);
nand U7937 (N_7937,N_7205,N_7483);
xor U7938 (N_7938,N_7207,N_7282);
or U7939 (N_7939,N_7381,N_7341);
nand U7940 (N_7940,N_7275,N_7255);
nor U7941 (N_7941,N_7426,N_7385);
nor U7942 (N_7942,N_7255,N_7341);
or U7943 (N_7943,N_7462,N_7598);
and U7944 (N_7944,N_7454,N_7403);
or U7945 (N_7945,N_7440,N_7436);
nor U7946 (N_7946,N_7552,N_7313);
and U7947 (N_7947,N_7289,N_7319);
nor U7948 (N_7948,N_7366,N_7526);
nor U7949 (N_7949,N_7523,N_7349);
or U7950 (N_7950,N_7205,N_7509);
nor U7951 (N_7951,N_7279,N_7360);
or U7952 (N_7952,N_7533,N_7420);
nand U7953 (N_7953,N_7548,N_7230);
and U7954 (N_7954,N_7282,N_7592);
nand U7955 (N_7955,N_7314,N_7374);
xor U7956 (N_7956,N_7597,N_7391);
and U7957 (N_7957,N_7494,N_7211);
and U7958 (N_7958,N_7242,N_7314);
xnor U7959 (N_7959,N_7481,N_7380);
and U7960 (N_7960,N_7461,N_7380);
xnor U7961 (N_7961,N_7480,N_7201);
and U7962 (N_7962,N_7204,N_7208);
nand U7963 (N_7963,N_7560,N_7380);
nand U7964 (N_7964,N_7374,N_7557);
and U7965 (N_7965,N_7222,N_7379);
nand U7966 (N_7966,N_7305,N_7579);
nand U7967 (N_7967,N_7568,N_7200);
nor U7968 (N_7968,N_7388,N_7368);
or U7969 (N_7969,N_7413,N_7231);
xor U7970 (N_7970,N_7291,N_7580);
nor U7971 (N_7971,N_7532,N_7449);
and U7972 (N_7972,N_7424,N_7580);
and U7973 (N_7973,N_7423,N_7338);
xor U7974 (N_7974,N_7518,N_7315);
xor U7975 (N_7975,N_7369,N_7249);
and U7976 (N_7976,N_7596,N_7275);
xor U7977 (N_7977,N_7278,N_7257);
xnor U7978 (N_7978,N_7497,N_7526);
xnor U7979 (N_7979,N_7577,N_7590);
and U7980 (N_7980,N_7544,N_7497);
nor U7981 (N_7981,N_7212,N_7452);
xor U7982 (N_7982,N_7472,N_7278);
xnor U7983 (N_7983,N_7331,N_7467);
and U7984 (N_7984,N_7447,N_7342);
nand U7985 (N_7985,N_7373,N_7308);
nor U7986 (N_7986,N_7255,N_7310);
nand U7987 (N_7987,N_7261,N_7266);
and U7988 (N_7988,N_7251,N_7213);
xor U7989 (N_7989,N_7558,N_7595);
and U7990 (N_7990,N_7473,N_7262);
or U7991 (N_7991,N_7209,N_7468);
and U7992 (N_7992,N_7484,N_7534);
nor U7993 (N_7993,N_7364,N_7408);
nor U7994 (N_7994,N_7255,N_7366);
or U7995 (N_7995,N_7218,N_7225);
or U7996 (N_7996,N_7227,N_7257);
nand U7997 (N_7997,N_7375,N_7464);
nor U7998 (N_7998,N_7335,N_7287);
xor U7999 (N_7999,N_7302,N_7465);
nor U8000 (N_8000,N_7997,N_7689);
nand U8001 (N_8001,N_7921,N_7703);
nor U8002 (N_8002,N_7826,N_7701);
and U8003 (N_8003,N_7851,N_7927);
xor U8004 (N_8004,N_7632,N_7678);
xor U8005 (N_8005,N_7892,N_7923);
or U8006 (N_8006,N_7849,N_7875);
nor U8007 (N_8007,N_7957,N_7772);
nor U8008 (N_8008,N_7977,N_7971);
nand U8009 (N_8009,N_7958,N_7746);
and U8010 (N_8010,N_7634,N_7866);
xor U8011 (N_8011,N_7685,N_7613);
and U8012 (N_8012,N_7918,N_7872);
or U8013 (N_8013,N_7982,N_7965);
nand U8014 (N_8014,N_7687,N_7868);
nor U8015 (N_8015,N_7920,N_7908);
and U8016 (N_8016,N_7814,N_7843);
nand U8017 (N_8017,N_7691,N_7718);
nor U8018 (N_8018,N_7641,N_7804);
nand U8019 (N_8019,N_7650,N_7943);
xnor U8020 (N_8020,N_7963,N_7615);
nand U8021 (N_8021,N_7754,N_7862);
and U8022 (N_8022,N_7706,N_7616);
xor U8023 (N_8023,N_7792,N_7626);
xnor U8024 (N_8024,N_7759,N_7993);
and U8025 (N_8025,N_7838,N_7713);
and U8026 (N_8026,N_7812,N_7708);
xnor U8027 (N_8027,N_7952,N_7854);
xor U8028 (N_8028,N_7954,N_7635);
or U8029 (N_8029,N_7960,N_7933);
nor U8030 (N_8030,N_7979,N_7704);
or U8031 (N_8031,N_7797,N_7999);
nand U8032 (N_8032,N_7828,N_7765);
nand U8033 (N_8033,N_7643,N_7646);
and U8034 (N_8034,N_7939,N_7707);
xnor U8035 (N_8035,N_7837,N_7739);
xor U8036 (N_8036,N_7865,N_7863);
xnor U8037 (N_8037,N_7767,N_7919);
nand U8038 (N_8038,N_7833,N_7916);
nor U8039 (N_8039,N_7947,N_7897);
xnor U8040 (N_8040,N_7606,N_7747);
nor U8041 (N_8041,N_7751,N_7905);
xnor U8042 (N_8042,N_7624,N_7877);
xor U8043 (N_8043,N_7727,N_7755);
nand U8044 (N_8044,N_7961,N_7645);
nand U8045 (N_8045,N_7675,N_7612);
and U8046 (N_8046,N_7839,N_7667);
nand U8047 (N_8047,N_7787,N_7909);
and U8048 (N_8048,N_7693,N_7700);
nor U8049 (N_8049,N_7903,N_7842);
nor U8050 (N_8050,N_7625,N_7978);
and U8051 (N_8051,N_7815,N_7976);
xor U8052 (N_8052,N_7912,N_7980);
nand U8053 (N_8053,N_7734,N_7663);
xor U8054 (N_8054,N_7941,N_7763);
nand U8055 (N_8055,N_7768,N_7834);
nand U8056 (N_8056,N_7848,N_7855);
xnor U8057 (N_8057,N_7924,N_7955);
xnor U8058 (N_8058,N_7741,N_7984);
nand U8059 (N_8059,N_7789,N_7884);
and U8060 (N_8060,N_7620,N_7853);
nor U8061 (N_8061,N_7657,N_7989);
or U8062 (N_8062,N_7761,N_7896);
nor U8063 (N_8063,N_7609,N_7680);
nor U8064 (N_8064,N_7686,N_7944);
and U8065 (N_8065,N_7934,N_7795);
and U8066 (N_8066,N_7864,N_7770);
xnor U8067 (N_8067,N_7659,N_7887);
xnor U8068 (N_8068,N_7990,N_7845);
nor U8069 (N_8069,N_7720,N_7983);
and U8070 (N_8070,N_7758,N_7820);
or U8071 (N_8071,N_7723,N_7810);
xnor U8072 (N_8072,N_7835,N_7968);
xnor U8073 (N_8073,N_7827,N_7604);
nand U8074 (N_8074,N_7935,N_7931);
nor U8075 (N_8075,N_7651,N_7817);
nor U8076 (N_8076,N_7679,N_7942);
nand U8077 (N_8077,N_7779,N_7750);
xnor U8078 (N_8078,N_7981,N_7946);
or U8079 (N_8079,N_7695,N_7959);
or U8080 (N_8080,N_7873,N_7859);
xnor U8081 (N_8081,N_7882,N_7682);
nand U8082 (N_8082,N_7860,N_7986);
nor U8083 (N_8083,N_7743,N_7647);
nor U8084 (N_8084,N_7953,N_7972);
xnor U8085 (N_8085,N_7825,N_7846);
or U8086 (N_8086,N_7658,N_7627);
or U8087 (N_8087,N_7736,N_7614);
and U8088 (N_8088,N_7794,N_7926);
nand U8089 (N_8089,N_7760,N_7890);
or U8090 (N_8090,N_7867,N_7660);
nand U8091 (N_8091,N_7692,N_7777);
nor U8092 (N_8092,N_7824,N_7781);
and U8093 (N_8093,N_7840,N_7748);
nor U8094 (N_8094,N_7726,N_7662);
xor U8095 (N_8095,N_7816,N_7813);
nand U8096 (N_8096,N_7893,N_7936);
nand U8097 (N_8097,N_7642,N_7948);
xor U8098 (N_8098,N_7889,N_7841);
nor U8099 (N_8099,N_7764,N_7638);
nand U8100 (N_8100,N_7898,N_7880);
or U8101 (N_8101,N_7610,N_7929);
or U8102 (N_8102,N_7785,N_7805);
xor U8103 (N_8103,N_7987,N_7652);
nor U8104 (N_8104,N_7661,N_7871);
xnor U8105 (N_8105,N_7605,N_7907);
nor U8106 (N_8106,N_7698,N_7911);
and U8107 (N_8107,N_7684,N_7883);
and U8108 (N_8108,N_7823,N_7966);
nand U8109 (N_8109,N_7636,N_7631);
and U8110 (N_8110,N_7670,N_7829);
and U8111 (N_8111,N_7910,N_7822);
nand U8112 (N_8112,N_7915,N_7717);
nor U8113 (N_8113,N_7722,N_7697);
or U8114 (N_8114,N_7611,N_7702);
and U8115 (N_8115,N_7836,N_7696);
or U8116 (N_8116,N_7728,N_7742);
xor U8117 (N_8117,N_7786,N_7694);
and U8118 (N_8118,N_7886,N_7962);
nor U8119 (N_8119,N_7811,N_7874);
and U8120 (N_8120,N_7895,N_7628);
xor U8121 (N_8121,N_7821,N_7830);
and U8122 (N_8122,N_7637,N_7803);
xnor U8123 (N_8123,N_7753,N_7802);
nand U8124 (N_8124,N_7745,N_7623);
xor U8125 (N_8125,N_7608,N_7749);
nand U8126 (N_8126,N_7809,N_7964);
or U8127 (N_8127,N_7683,N_7668);
nand U8128 (N_8128,N_7975,N_7858);
nor U8129 (N_8129,N_7856,N_7644);
xor U8130 (N_8130,N_7629,N_7656);
or U8131 (N_8131,N_7688,N_7998);
nor U8132 (N_8132,N_7806,N_7681);
nand U8133 (N_8133,N_7714,N_7653);
nand U8134 (N_8134,N_7699,N_7819);
xnor U8135 (N_8135,N_7956,N_7666);
and U8136 (N_8136,N_7901,N_7807);
nand U8137 (N_8137,N_7640,N_7974);
nand U8138 (N_8138,N_7818,N_7994);
nor U8139 (N_8139,N_7729,N_7672);
and U8140 (N_8140,N_7607,N_7917);
xnor U8141 (N_8141,N_7783,N_7664);
and U8142 (N_8142,N_7951,N_7676);
nand U8143 (N_8143,N_7602,N_7735);
nor U8144 (N_8144,N_7861,N_7832);
nor U8145 (N_8145,N_7850,N_7949);
or U8146 (N_8146,N_7793,N_7796);
or U8147 (N_8147,N_7940,N_7885);
and U8148 (N_8148,N_7857,N_7879);
or U8149 (N_8149,N_7674,N_7639);
nor U8150 (N_8150,N_7721,N_7782);
nor U8151 (N_8151,N_7967,N_7771);
and U8152 (N_8152,N_7788,N_7891);
and U8153 (N_8153,N_7970,N_7669);
or U8154 (N_8154,N_7938,N_7709);
xnor U8155 (N_8155,N_7799,N_7894);
nand U8156 (N_8156,N_7791,N_7902);
nor U8157 (N_8157,N_7844,N_7775);
xnor U8158 (N_8158,N_7800,N_7690);
nand U8159 (N_8159,N_7730,N_7878);
or U8160 (N_8160,N_7622,N_7869);
nand U8161 (N_8161,N_7731,N_7985);
nor U8162 (N_8162,N_7600,N_7945);
nand U8163 (N_8163,N_7665,N_7724);
or U8164 (N_8164,N_7773,N_7888);
or U8165 (N_8165,N_7633,N_7712);
xnor U8166 (N_8166,N_7715,N_7619);
xnor U8167 (N_8167,N_7995,N_7769);
xor U8168 (N_8168,N_7601,N_7950);
or U8169 (N_8169,N_7617,N_7870);
and U8170 (N_8170,N_7603,N_7928);
and U8171 (N_8171,N_7649,N_7992);
and U8172 (N_8172,N_7737,N_7937);
and U8173 (N_8173,N_7798,N_7801);
nor U8174 (N_8174,N_7876,N_7881);
nor U8175 (N_8175,N_7932,N_7710);
or U8176 (N_8176,N_7744,N_7756);
nand U8177 (N_8177,N_7719,N_7725);
nor U8178 (N_8178,N_7677,N_7988);
nand U8179 (N_8179,N_7925,N_7790);
nor U8180 (N_8180,N_7732,N_7904);
or U8181 (N_8181,N_7648,N_7762);
and U8182 (N_8182,N_7996,N_7654);
and U8183 (N_8183,N_7705,N_7831);
nand U8184 (N_8184,N_7673,N_7973);
xor U8185 (N_8185,N_7906,N_7808);
and U8186 (N_8186,N_7766,N_7774);
and U8187 (N_8187,N_7716,N_7969);
xnor U8188 (N_8188,N_7733,N_7655);
or U8189 (N_8189,N_7991,N_7757);
and U8190 (N_8190,N_7922,N_7630);
xor U8191 (N_8191,N_7913,N_7778);
xor U8192 (N_8192,N_7899,N_7621);
and U8193 (N_8193,N_7852,N_7847);
nor U8194 (N_8194,N_7671,N_7618);
and U8195 (N_8195,N_7784,N_7740);
or U8196 (N_8196,N_7914,N_7780);
or U8197 (N_8197,N_7776,N_7752);
nor U8198 (N_8198,N_7738,N_7711);
xor U8199 (N_8199,N_7900,N_7930);
nand U8200 (N_8200,N_7896,N_7950);
nor U8201 (N_8201,N_7629,N_7832);
xor U8202 (N_8202,N_7806,N_7643);
and U8203 (N_8203,N_7952,N_7758);
nor U8204 (N_8204,N_7658,N_7984);
or U8205 (N_8205,N_7670,N_7774);
or U8206 (N_8206,N_7998,N_7801);
xor U8207 (N_8207,N_7857,N_7764);
xor U8208 (N_8208,N_7938,N_7903);
nor U8209 (N_8209,N_7747,N_7800);
or U8210 (N_8210,N_7623,N_7812);
nor U8211 (N_8211,N_7870,N_7601);
nor U8212 (N_8212,N_7672,N_7983);
xnor U8213 (N_8213,N_7683,N_7785);
and U8214 (N_8214,N_7853,N_7837);
and U8215 (N_8215,N_7741,N_7730);
xor U8216 (N_8216,N_7907,N_7633);
and U8217 (N_8217,N_7990,N_7804);
nor U8218 (N_8218,N_7691,N_7704);
xnor U8219 (N_8219,N_7609,N_7779);
and U8220 (N_8220,N_7908,N_7864);
or U8221 (N_8221,N_7942,N_7805);
xor U8222 (N_8222,N_7730,N_7757);
nand U8223 (N_8223,N_7644,N_7832);
nand U8224 (N_8224,N_7748,N_7958);
and U8225 (N_8225,N_7816,N_7620);
nor U8226 (N_8226,N_7743,N_7872);
or U8227 (N_8227,N_7969,N_7748);
and U8228 (N_8228,N_7822,N_7991);
nand U8229 (N_8229,N_7885,N_7636);
nand U8230 (N_8230,N_7756,N_7669);
or U8231 (N_8231,N_7656,N_7735);
or U8232 (N_8232,N_7610,N_7949);
or U8233 (N_8233,N_7648,N_7637);
or U8234 (N_8234,N_7606,N_7786);
or U8235 (N_8235,N_7831,N_7914);
and U8236 (N_8236,N_7752,N_7801);
or U8237 (N_8237,N_7811,N_7729);
and U8238 (N_8238,N_7934,N_7781);
nor U8239 (N_8239,N_7656,N_7831);
and U8240 (N_8240,N_7848,N_7940);
nor U8241 (N_8241,N_7844,N_7601);
and U8242 (N_8242,N_7814,N_7922);
and U8243 (N_8243,N_7905,N_7973);
xor U8244 (N_8244,N_7766,N_7677);
or U8245 (N_8245,N_7923,N_7791);
and U8246 (N_8246,N_7708,N_7619);
nor U8247 (N_8247,N_7954,N_7784);
nand U8248 (N_8248,N_7864,N_7603);
xor U8249 (N_8249,N_7876,N_7784);
nor U8250 (N_8250,N_7897,N_7918);
or U8251 (N_8251,N_7958,N_7858);
or U8252 (N_8252,N_7688,N_7702);
nor U8253 (N_8253,N_7887,N_7639);
or U8254 (N_8254,N_7612,N_7665);
and U8255 (N_8255,N_7849,N_7800);
nor U8256 (N_8256,N_7861,N_7820);
xor U8257 (N_8257,N_7830,N_7925);
nor U8258 (N_8258,N_7658,N_7871);
nand U8259 (N_8259,N_7866,N_7757);
and U8260 (N_8260,N_7635,N_7810);
nand U8261 (N_8261,N_7638,N_7707);
xor U8262 (N_8262,N_7758,N_7768);
xor U8263 (N_8263,N_7918,N_7601);
nor U8264 (N_8264,N_7633,N_7652);
or U8265 (N_8265,N_7816,N_7774);
xor U8266 (N_8266,N_7933,N_7829);
nor U8267 (N_8267,N_7718,N_7706);
or U8268 (N_8268,N_7648,N_7764);
nand U8269 (N_8269,N_7989,N_7890);
nand U8270 (N_8270,N_7995,N_7966);
and U8271 (N_8271,N_7931,N_7853);
nor U8272 (N_8272,N_7819,N_7931);
xnor U8273 (N_8273,N_7748,N_7672);
or U8274 (N_8274,N_7837,N_7975);
nand U8275 (N_8275,N_7909,N_7927);
xnor U8276 (N_8276,N_7953,N_7796);
xor U8277 (N_8277,N_7888,N_7685);
or U8278 (N_8278,N_7761,N_7934);
nand U8279 (N_8279,N_7698,N_7631);
and U8280 (N_8280,N_7693,N_7607);
and U8281 (N_8281,N_7704,N_7797);
xor U8282 (N_8282,N_7874,N_7747);
nand U8283 (N_8283,N_7845,N_7742);
nand U8284 (N_8284,N_7607,N_7679);
and U8285 (N_8285,N_7654,N_7676);
nand U8286 (N_8286,N_7651,N_7675);
nand U8287 (N_8287,N_7928,N_7978);
nor U8288 (N_8288,N_7766,N_7711);
or U8289 (N_8289,N_7973,N_7684);
and U8290 (N_8290,N_7856,N_7624);
nand U8291 (N_8291,N_7818,N_7697);
nand U8292 (N_8292,N_7744,N_7712);
or U8293 (N_8293,N_7693,N_7751);
xor U8294 (N_8294,N_7674,N_7625);
or U8295 (N_8295,N_7750,N_7637);
nor U8296 (N_8296,N_7628,N_7655);
nand U8297 (N_8297,N_7901,N_7836);
nor U8298 (N_8298,N_7688,N_7726);
nor U8299 (N_8299,N_7918,N_7678);
nand U8300 (N_8300,N_7813,N_7767);
nor U8301 (N_8301,N_7614,N_7639);
nor U8302 (N_8302,N_7886,N_7884);
or U8303 (N_8303,N_7648,N_7630);
or U8304 (N_8304,N_7743,N_7988);
nand U8305 (N_8305,N_7629,N_7833);
nor U8306 (N_8306,N_7600,N_7988);
nor U8307 (N_8307,N_7737,N_7770);
xor U8308 (N_8308,N_7846,N_7871);
nand U8309 (N_8309,N_7762,N_7894);
and U8310 (N_8310,N_7832,N_7691);
xnor U8311 (N_8311,N_7820,N_7608);
and U8312 (N_8312,N_7747,N_7812);
xnor U8313 (N_8313,N_7776,N_7701);
xnor U8314 (N_8314,N_7855,N_7777);
or U8315 (N_8315,N_7818,N_7742);
nand U8316 (N_8316,N_7725,N_7941);
nand U8317 (N_8317,N_7824,N_7640);
nor U8318 (N_8318,N_7861,N_7731);
and U8319 (N_8319,N_7676,N_7631);
nand U8320 (N_8320,N_7943,N_7805);
nand U8321 (N_8321,N_7761,N_7889);
nor U8322 (N_8322,N_7965,N_7883);
nor U8323 (N_8323,N_7958,N_7948);
nand U8324 (N_8324,N_7709,N_7810);
xor U8325 (N_8325,N_7643,N_7941);
xor U8326 (N_8326,N_7717,N_7773);
and U8327 (N_8327,N_7833,N_7861);
nor U8328 (N_8328,N_7810,N_7777);
or U8329 (N_8329,N_7854,N_7865);
nor U8330 (N_8330,N_7915,N_7839);
xor U8331 (N_8331,N_7973,N_7649);
nand U8332 (N_8332,N_7838,N_7625);
nor U8333 (N_8333,N_7881,N_7966);
and U8334 (N_8334,N_7632,N_7614);
nor U8335 (N_8335,N_7655,N_7747);
xor U8336 (N_8336,N_7991,N_7890);
nand U8337 (N_8337,N_7684,N_7611);
xor U8338 (N_8338,N_7810,N_7758);
or U8339 (N_8339,N_7857,N_7646);
nor U8340 (N_8340,N_7627,N_7693);
nand U8341 (N_8341,N_7638,N_7865);
or U8342 (N_8342,N_7848,N_7904);
nor U8343 (N_8343,N_7932,N_7951);
or U8344 (N_8344,N_7707,N_7924);
and U8345 (N_8345,N_7780,N_7672);
xor U8346 (N_8346,N_7781,N_7639);
nand U8347 (N_8347,N_7899,N_7632);
or U8348 (N_8348,N_7992,N_7932);
nand U8349 (N_8349,N_7708,N_7662);
and U8350 (N_8350,N_7614,N_7666);
xnor U8351 (N_8351,N_7733,N_7777);
or U8352 (N_8352,N_7971,N_7746);
nand U8353 (N_8353,N_7817,N_7778);
and U8354 (N_8354,N_7789,N_7680);
nand U8355 (N_8355,N_7617,N_7914);
and U8356 (N_8356,N_7615,N_7761);
nor U8357 (N_8357,N_7705,N_7975);
and U8358 (N_8358,N_7805,N_7715);
nor U8359 (N_8359,N_7982,N_7665);
xnor U8360 (N_8360,N_7925,N_7980);
or U8361 (N_8361,N_7939,N_7634);
xnor U8362 (N_8362,N_7811,N_7910);
nor U8363 (N_8363,N_7672,N_7791);
nor U8364 (N_8364,N_7835,N_7850);
or U8365 (N_8365,N_7920,N_7965);
nor U8366 (N_8366,N_7883,N_7602);
or U8367 (N_8367,N_7782,N_7985);
or U8368 (N_8368,N_7814,N_7657);
nand U8369 (N_8369,N_7761,N_7620);
nand U8370 (N_8370,N_7641,N_7837);
nor U8371 (N_8371,N_7636,N_7845);
nand U8372 (N_8372,N_7717,N_7835);
or U8373 (N_8373,N_7851,N_7871);
nand U8374 (N_8374,N_7877,N_7772);
nor U8375 (N_8375,N_7798,N_7885);
nand U8376 (N_8376,N_7737,N_7700);
nand U8377 (N_8377,N_7865,N_7952);
nor U8378 (N_8378,N_7828,N_7863);
nor U8379 (N_8379,N_7817,N_7723);
nand U8380 (N_8380,N_7669,N_7931);
or U8381 (N_8381,N_7774,N_7906);
or U8382 (N_8382,N_7690,N_7783);
nand U8383 (N_8383,N_7622,N_7768);
nor U8384 (N_8384,N_7758,N_7784);
nor U8385 (N_8385,N_7794,N_7731);
and U8386 (N_8386,N_7874,N_7829);
or U8387 (N_8387,N_7777,N_7785);
nand U8388 (N_8388,N_7997,N_7910);
and U8389 (N_8389,N_7609,N_7917);
or U8390 (N_8390,N_7870,N_7904);
nand U8391 (N_8391,N_7609,N_7700);
xnor U8392 (N_8392,N_7753,N_7781);
and U8393 (N_8393,N_7720,N_7996);
nor U8394 (N_8394,N_7666,N_7632);
nand U8395 (N_8395,N_7730,N_7798);
nor U8396 (N_8396,N_7702,N_7750);
and U8397 (N_8397,N_7724,N_7645);
or U8398 (N_8398,N_7802,N_7797);
nor U8399 (N_8399,N_7879,N_7672);
or U8400 (N_8400,N_8181,N_8201);
and U8401 (N_8401,N_8095,N_8256);
and U8402 (N_8402,N_8145,N_8363);
nand U8403 (N_8403,N_8069,N_8073);
nand U8404 (N_8404,N_8184,N_8066);
nand U8405 (N_8405,N_8165,N_8376);
and U8406 (N_8406,N_8253,N_8299);
or U8407 (N_8407,N_8268,N_8242);
and U8408 (N_8408,N_8250,N_8124);
xnor U8409 (N_8409,N_8150,N_8000);
and U8410 (N_8410,N_8009,N_8125);
nor U8411 (N_8411,N_8086,N_8016);
and U8412 (N_8412,N_8334,N_8198);
or U8413 (N_8413,N_8378,N_8007);
nor U8414 (N_8414,N_8075,N_8336);
xor U8415 (N_8415,N_8266,N_8079);
xor U8416 (N_8416,N_8282,N_8032);
and U8417 (N_8417,N_8313,N_8135);
or U8418 (N_8418,N_8239,N_8084);
nand U8419 (N_8419,N_8333,N_8331);
or U8420 (N_8420,N_8352,N_8301);
or U8421 (N_8421,N_8104,N_8248);
and U8422 (N_8422,N_8312,N_8288);
nor U8423 (N_8423,N_8296,N_8329);
nand U8424 (N_8424,N_8044,N_8056);
nand U8425 (N_8425,N_8099,N_8219);
or U8426 (N_8426,N_8136,N_8121);
xnor U8427 (N_8427,N_8081,N_8223);
xnor U8428 (N_8428,N_8259,N_8311);
nand U8429 (N_8429,N_8089,N_8055);
nor U8430 (N_8430,N_8207,N_8300);
or U8431 (N_8431,N_8083,N_8255);
nor U8432 (N_8432,N_8241,N_8019);
nand U8433 (N_8433,N_8152,N_8391);
xor U8434 (N_8434,N_8225,N_8074);
or U8435 (N_8435,N_8130,N_8309);
xnor U8436 (N_8436,N_8271,N_8214);
nor U8437 (N_8437,N_8036,N_8330);
or U8438 (N_8438,N_8180,N_8353);
xnor U8439 (N_8439,N_8062,N_8210);
or U8440 (N_8440,N_8090,N_8398);
and U8441 (N_8441,N_8321,N_8211);
or U8442 (N_8442,N_8120,N_8097);
and U8443 (N_8443,N_8339,N_8295);
nand U8444 (N_8444,N_8341,N_8366);
nor U8445 (N_8445,N_8149,N_8316);
or U8446 (N_8446,N_8098,N_8160);
xor U8447 (N_8447,N_8108,N_8008);
xnor U8448 (N_8448,N_8292,N_8272);
nor U8449 (N_8449,N_8174,N_8025);
or U8450 (N_8450,N_8251,N_8085);
xnor U8451 (N_8451,N_8020,N_8034);
nor U8452 (N_8452,N_8050,N_8328);
xor U8453 (N_8453,N_8018,N_8208);
xnor U8454 (N_8454,N_8162,N_8118);
nor U8455 (N_8455,N_8023,N_8171);
xor U8456 (N_8456,N_8355,N_8358);
nand U8457 (N_8457,N_8059,N_8123);
and U8458 (N_8458,N_8220,N_8063);
xor U8459 (N_8459,N_8322,N_8384);
or U8460 (N_8460,N_8240,N_8371);
xnor U8461 (N_8461,N_8040,N_8033);
nor U8462 (N_8462,N_8116,N_8192);
and U8463 (N_8463,N_8230,N_8191);
and U8464 (N_8464,N_8027,N_8183);
xnor U8465 (N_8465,N_8289,N_8068);
nor U8466 (N_8466,N_8260,N_8164);
and U8467 (N_8467,N_8045,N_8013);
nor U8468 (N_8468,N_8237,N_8350);
and U8469 (N_8469,N_8148,N_8014);
nand U8470 (N_8470,N_8325,N_8115);
and U8471 (N_8471,N_8235,N_8394);
nor U8472 (N_8472,N_8269,N_8395);
nand U8473 (N_8473,N_8129,N_8206);
and U8474 (N_8474,N_8113,N_8274);
and U8475 (N_8475,N_8356,N_8385);
nand U8476 (N_8476,N_8182,N_8303);
and U8477 (N_8477,N_8302,N_8314);
and U8478 (N_8478,N_8047,N_8332);
or U8479 (N_8479,N_8367,N_8179);
nand U8480 (N_8480,N_8388,N_8270);
nand U8481 (N_8481,N_8111,N_8243);
nor U8482 (N_8482,N_8380,N_8067);
or U8483 (N_8483,N_8375,N_8317);
or U8484 (N_8484,N_8012,N_8138);
or U8485 (N_8485,N_8131,N_8058);
xnor U8486 (N_8486,N_8053,N_8003);
and U8487 (N_8487,N_8344,N_8258);
nand U8488 (N_8488,N_8185,N_8277);
nor U8489 (N_8489,N_8107,N_8163);
and U8490 (N_8490,N_8305,N_8140);
xnor U8491 (N_8491,N_8194,N_8080);
nor U8492 (N_8492,N_8369,N_8114);
or U8493 (N_8493,N_8028,N_8263);
or U8494 (N_8494,N_8372,N_8335);
nor U8495 (N_8495,N_8294,N_8026);
nand U8496 (N_8496,N_8228,N_8222);
nand U8497 (N_8497,N_8134,N_8373);
and U8498 (N_8498,N_8196,N_8381);
or U8499 (N_8499,N_8158,N_8061);
or U8500 (N_8500,N_8199,N_8257);
nand U8501 (N_8501,N_8147,N_8117);
xor U8502 (N_8502,N_8168,N_8049);
and U8503 (N_8503,N_8057,N_8362);
and U8504 (N_8504,N_8320,N_8261);
nor U8505 (N_8505,N_8155,N_8357);
nand U8506 (N_8506,N_8342,N_8024);
nor U8507 (N_8507,N_8188,N_8153);
or U8508 (N_8508,N_8232,N_8318);
nand U8509 (N_8509,N_8374,N_8015);
xnor U8510 (N_8510,N_8054,N_8340);
and U8511 (N_8511,N_8159,N_8209);
or U8512 (N_8512,N_8349,N_8389);
nand U8513 (N_8513,N_8151,N_8200);
or U8514 (N_8514,N_8324,N_8285);
nand U8515 (N_8515,N_8254,N_8143);
and U8516 (N_8516,N_8154,N_8133);
nor U8517 (N_8517,N_8010,N_8071);
or U8518 (N_8518,N_8106,N_8144);
nor U8519 (N_8519,N_8139,N_8137);
or U8520 (N_8520,N_8382,N_8283);
or U8521 (N_8521,N_8119,N_8190);
or U8522 (N_8522,N_8397,N_8100);
nand U8523 (N_8523,N_8052,N_8203);
xor U8524 (N_8524,N_8177,N_8002);
nand U8525 (N_8525,N_8166,N_8364);
or U8526 (N_8526,N_8310,N_8102);
nor U8527 (N_8527,N_8379,N_8234);
xnor U8528 (N_8528,N_8038,N_8078);
nand U8529 (N_8529,N_8005,N_8286);
and U8530 (N_8530,N_8216,N_8246);
xor U8531 (N_8531,N_8326,N_8264);
nand U8532 (N_8532,N_8105,N_8226);
nor U8533 (N_8533,N_8193,N_8224);
or U8534 (N_8534,N_8244,N_8146);
or U8535 (N_8535,N_8279,N_8187);
nand U8536 (N_8536,N_8094,N_8161);
nor U8537 (N_8537,N_8278,N_8315);
nand U8538 (N_8538,N_8267,N_8360);
or U8539 (N_8539,N_8287,N_8291);
xnor U8540 (N_8540,N_8354,N_8029);
xor U8541 (N_8541,N_8204,N_8060);
and U8542 (N_8542,N_8186,N_8396);
xor U8543 (N_8543,N_8039,N_8276);
nor U8544 (N_8544,N_8077,N_8281);
nand U8545 (N_8545,N_8127,N_8215);
nor U8546 (N_8546,N_8370,N_8070);
xnor U8547 (N_8547,N_8172,N_8399);
nor U8548 (N_8548,N_8368,N_8280);
nor U8549 (N_8549,N_8393,N_8087);
and U8550 (N_8550,N_8293,N_8017);
or U8551 (N_8551,N_8043,N_8297);
or U8552 (N_8552,N_8212,N_8175);
or U8553 (N_8553,N_8323,N_8343);
and U8554 (N_8554,N_8103,N_8217);
and U8555 (N_8555,N_8122,N_8327);
and U8556 (N_8556,N_8319,N_8189);
nor U8557 (N_8557,N_8390,N_8233);
nand U8558 (N_8558,N_8169,N_8361);
or U8559 (N_8559,N_8262,N_8245);
nand U8560 (N_8560,N_8064,N_8132);
xnor U8561 (N_8561,N_8048,N_8167);
nor U8562 (N_8562,N_8392,N_8157);
nand U8563 (N_8563,N_8006,N_8001);
xor U8564 (N_8564,N_8377,N_8273);
xor U8565 (N_8565,N_8101,N_8156);
nor U8566 (N_8566,N_8141,N_8093);
or U8567 (N_8567,N_8021,N_8359);
nand U8568 (N_8568,N_8227,N_8337);
and U8569 (N_8569,N_8076,N_8035);
nand U8570 (N_8570,N_8197,N_8298);
nand U8571 (N_8571,N_8128,N_8037);
nor U8572 (N_8572,N_8022,N_8091);
and U8573 (N_8573,N_8365,N_8275);
or U8574 (N_8574,N_8348,N_8092);
or U8575 (N_8575,N_8347,N_8307);
and U8576 (N_8576,N_8249,N_8351);
or U8577 (N_8577,N_8088,N_8247);
nor U8578 (N_8578,N_8051,N_8221);
nand U8579 (N_8579,N_8112,N_8072);
or U8580 (N_8580,N_8173,N_8041);
xor U8581 (N_8581,N_8030,N_8011);
nand U8582 (N_8582,N_8290,N_8031);
nand U8583 (N_8583,N_8231,N_8042);
and U8584 (N_8584,N_8065,N_8345);
nand U8585 (N_8585,N_8306,N_8238);
or U8586 (N_8586,N_8284,N_8205);
and U8587 (N_8587,N_8176,N_8110);
nor U8588 (N_8588,N_8386,N_8304);
and U8589 (N_8589,N_8170,N_8387);
and U8590 (N_8590,N_8229,N_8202);
or U8591 (N_8591,N_8346,N_8109);
xnor U8592 (N_8592,N_8383,N_8142);
and U8593 (N_8593,N_8082,N_8252);
or U8594 (N_8594,N_8046,N_8004);
xor U8595 (N_8595,N_8126,N_8265);
and U8596 (N_8596,N_8178,N_8338);
nor U8597 (N_8597,N_8213,N_8308);
xnor U8598 (N_8598,N_8218,N_8096);
or U8599 (N_8599,N_8195,N_8236);
nand U8600 (N_8600,N_8356,N_8138);
nor U8601 (N_8601,N_8359,N_8302);
nor U8602 (N_8602,N_8098,N_8230);
or U8603 (N_8603,N_8330,N_8002);
nor U8604 (N_8604,N_8291,N_8255);
xor U8605 (N_8605,N_8078,N_8246);
nor U8606 (N_8606,N_8124,N_8190);
xnor U8607 (N_8607,N_8212,N_8348);
and U8608 (N_8608,N_8357,N_8158);
nor U8609 (N_8609,N_8026,N_8292);
and U8610 (N_8610,N_8232,N_8072);
nand U8611 (N_8611,N_8258,N_8024);
nor U8612 (N_8612,N_8287,N_8386);
nor U8613 (N_8613,N_8371,N_8049);
and U8614 (N_8614,N_8052,N_8164);
nor U8615 (N_8615,N_8191,N_8258);
nor U8616 (N_8616,N_8063,N_8050);
or U8617 (N_8617,N_8063,N_8075);
xnor U8618 (N_8618,N_8066,N_8260);
and U8619 (N_8619,N_8219,N_8086);
nor U8620 (N_8620,N_8324,N_8024);
xnor U8621 (N_8621,N_8021,N_8200);
or U8622 (N_8622,N_8025,N_8294);
nand U8623 (N_8623,N_8263,N_8319);
nand U8624 (N_8624,N_8031,N_8171);
and U8625 (N_8625,N_8096,N_8243);
nand U8626 (N_8626,N_8294,N_8219);
xnor U8627 (N_8627,N_8290,N_8191);
nand U8628 (N_8628,N_8335,N_8143);
nor U8629 (N_8629,N_8189,N_8226);
and U8630 (N_8630,N_8024,N_8065);
nor U8631 (N_8631,N_8069,N_8232);
nor U8632 (N_8632,N_8384,N_8124);
and U8633 (N_8633,N_8202,N_8104);
nand U8634 (N_8634,N_8036,N_8049);
and U8635 (N_8635,N_8021,N_8157);
nor U8636 (N_8636,N_8302,N_8224);
or U8637 (N_8637,N_8000,N_8163);
or U8638 (N_8638,N_8393,N_8001);
or U8639 (N_8639,N_8358,N_8129);
and U8640 (N_8640,N_8184,N_8182);
nand U8641 (N_8641,N_8194,N_8017);
xor U8642 (N_8642,N_8200,N_8139);
and U8643 (N_8643,N_8291,N_8182);
nand U8644 (N_8644,N_8218,N_8314);
nor U8645 (N_8645,N_8191,N_8235);
xor U8646 (N_8646,N_8170,N_8159);
xnor U8647 (N_8647,N_8002,N_8057);
nor U8648 (N_8648,N_8048,N_8128);
or U8649 (N_8649,N_8396,N_8398);
xor U8650 (N_8650,N_8171,N_8380);
nand U8651 (N_8651,N_8033,N_8183);
or U8652 (N_8652,N_8144,N_8009);
nand U8653 (N_8653,N_8193,N_8038);
nor U8654 (N_8654,N_8126,N_8178);
and U8655 (N_8655,N_8203,N_8299);
and U8656 (N_8656,N_8020,N_8044);
nand U8657 (N_8657,N_8205,N_8076);
and U8658 (N_8658,N_8119,N_8378);
nor U8659 (N_8659,N_8102,N_8263);
and U8660 (N_8660,N_8172,N_8112);
nand U8661 (N_8661,N_8270,N_8244);
nand U8662 (N_8662,N_8145,N_8062);
and U8663 (N_8663,N_8338,N_8352);
and U8664 (N_8664,N_8182,N_8144);
or U8665 (N_8665,N_8093,N_8163);
xnor U8666 (N_8666,N_8035,N_8384);
or U8667 (N_8667,N_8253,N_8313);
or U8668 (N_8668,N_8092,N_8160);
or U8669 (N_8669,N_8236,N_8298);
nand U8670 (N_8670,N_8336,N_8212);
and U8671 (N_8671,N_8347,N_8109);
nand U8672 (N_8672,N_8292,N_8094);
nor U8673 (N_8673,N_8339,N_8394);
nor U8674 (N_8674,N_8133,N_8030);
nor U8675 (N_8675,N_8352,N_8047);
nand U8676 (N_8676,N_8313,N_8136);
and U8677 (N_8677,N_8131,N_8052);
or U8678 (N_8678,N_8042,N_8391);
nor U8679 (N_8679,N_8152,N_8031);
and U8680 (N_8680,N_8082,N_8010);
and U8681 (N_8681,N_8392,N_8323);
nor U8682 (N_8682,N_8258,N_8348);
xor U8683 (N_8683,N_8238,N_8216);
and U8684 (N_8684,N_8221,N_8200);
or U8685 (N_8685,N_8248,N_8314);
or U8686 (N_8686,N_8398,N_8128);
xor U8687 (N_8687,N_8318,N_8183);
nand U8688 (N_8688,N_8387,N_8389);
nor U8689 (N_8689,N_8214,N_8286);
or U8690 (N_8690,N_8043,N_8095);
nand U8691 (N_8691,N_8059,N_8014);
xnor U8692 (N_8692,N_8172,N_8029);
xor U8693 (N_8693,N_8294,N_8159);
xnor U8694 (N_8694,N_8121,N_8000);
or U8695 (N_8695,N_8261,N_8331);
nor U8696 (N_8696,N_8000,N_8012);
or U8697 (N_8697,N_8112,N_8274);
xnor U8698 (N_8698,N_8102,N_8179);
nor U8699 (N_8699,N_8336,N_8169);
or U8700 (N_8700,N_8214,N_8081);
xor U8701 (N_8701,N_8079,N_8294);
and U8702 (N_8702,N_8284,N_8292);
nand U8703 (N_8703,N_8274,N_8322);
and U8704 (N_8704,N_8369,N_8097);
xnor U8705 (N_8705,N_8216,N_8067);
xnor U8706 (N_8706,N_8110,N_8358);
nand U8707 (N_8707,N_8061,N_8396);
nand U8708 (N_8708,N_8133,N_8285);
and U8709 (N_8709,N_8223,N_8327);
or U8710 (N_8710,N_8365,N_8351);
nand U8711 (N_8711,N_8102,N_8071);
nor U8712 (N_8712,N_8219,N_8088);
nand U8713 (N_8713,N_8053,N_8234);
nand U8714 (N_8714,N_8037,N_8153);
and U8715 (N_8715,N_8029,N_8165);
nand U8716 (N_8716,N_8249,N_8122);
nand U8717 (N_8717,N_8304,N_8135);
and U8718 (N_8718,N_8156,N_8380);
and U8719 (N_8719,N_8189,N_8337);
and U8720 (N_8720,N_8156,N_8035);
and U8721 (N_8721,N_8152,N_8159);
nor U8722 (N_8722,N_8069,N_8291);
nand U8723 (N_8723,N_8058,N_8079);
and U8724 (N_8724,N_8344,N_8342);
or U8725 (N_8725,N_8032,N_8335);
and U8726 (N_8726,N_8342,N_8244);
nand U8727 (N_8727,N_8019,N_8126);
or U8728 (N_8728,N_8077,N_8160);
and U8729 (N_8729,N_8135,N_8239);
and U8730 (N_8730,N_8134,N_8033);
nand U8731 (N_8731,N_8124,N_8014);
or U8732 (N_8732,N_8152,N_8259);
and U8733 (N_8733,N_8070,N_8208);
nor U8734 (N_8734,N_8370,N_8032);
and U8735 (N_8735,N_8317,N_8383);
xnor U8736 (N_8736,N_8206,N_8173);
and U8737 (N_8737,N_8129,N_8029);
or U8738 (N_8738,N_8105,N_8205);
nor U8739 (N_8739,N_8049,N_8313);
or U8740 (N_8740,N_8151,N_8240);
nor U8741 (N_8741,N_8372,N_8262);
or U8742 (N_8742,N_8023,N_8283);
or U8743 (N_8743,N_8067,N_8037);
nand U8744 (N_8744,N_8396,N_8279);
or U8745 (N_8745,N_8329,N_8299);
nor U8746 (N_8746,N_8282,N_8065);
nor U8747 (N_8747,N_8301,N_8097);
xnor U8748 (N_8748,N_8194,N_8156);
or U8749 (N_8749,N_8374,N_8346);
or U8750 (N_8750,N_8349,N_8330);
or U8751 (N_8751,N_8250,N_8004);
or U8752 (N_8752,N_8094,N_8174);
or U8753 (N_8753,N_8236,N_8331);
nor U8754 (N_8754,N_8286,N_8148);
nor U8755 (N_8755,N_8366,N_8347);
xnor U8756 (N_8756,N_8162,N_8246);
and U8757 (N_8757,N_8130,N_8002);
nor U8758 (N_8758,N_8146,N_8174);
or U8759 (N_8759,N_8179,N_8096);
nand U8760 (N_8760,N_8045,N_8393);
nand U8761 (N_8761,N_8218,N_8123);
nand U8762 (N_8762,N_8021,N_8100);
nor U8763 (N_8763,N_8330,N_8039);
and U8764 (N_8764,N_8197,N_8318);
or U8765 (N_8765,N_8308,N_8131);
nor U8766 (N_8766,N_8187,N_8392);
nor U8767 (N_8767,N_8038,N_8183);
nand U8768 (N_8768,N_8351,N_8301);
nand U8769 (N_8769,N_8310,N_8203);
nor U8770 (N_8770,N_8292,N_8075);
or U8771 (N_8771,N_8326,N_8185);
nand U8772 (N_8772,N_8394,N_8325);
or U8773 (N_8773,N_8267,N_8395);
nand U8774 (N_8774,N_8043,N_8224);
nand U8775 (N_8775,N_8360,N_8197);
xnor U8776 (N_8776,N_8192,N_8126);
or U8777 (N_8777,N_8098,N_8185);
nand U8778 (N_8778,N_8006,N_8204);
or U8779 (N_8779,N_8110,N_8352);
xnor U8780 (N_8780,N_8252,N_8195);
or U8781 (N_8781,N_8240,N_8083);
xnor U8782 (N_8782,N_8218,N_8339);
nor U8783 (N_8783,N_8099,N_8000);
nand U8784 (N_8784,N_8247,N_8254);
or U8785 (N_8785,N_8149,N_8370);
or U8786 (N_8786,N_8335,N_8288);
nor U8787 (N_8787,N_8192,N_8148);
xor U8788 (N_8788,N_8045,N_8367);
nand U8789 (N_8789,N_8260,N_8101);
nand U8790 (N_8790,N_8087,N_8121);
nand U8791 (N_8791,N_8364,N_8365);
and U8792 (N_8792,N_8050,N_8258);
nand U8793 (N_8793,N_8065,N_8347);
and U8794 (N_8794,N_8201,N_8066);
nand U8795 (N_8795,N_8365,N_8139);
nor U8796 (N_8796,N_8236,N_8304);
nor U8797 (N_8797,N_8059,N_8339);
xor U8798 (N_8798,N_8311,N_8339);
and U8799 (N_8799,N_8175,N_8046);
or U8800 (N_8800,N_8709,N_8421);
nand U8801 (N_8801,N_8573,N_8589);
or U8802 (N_8802,N_8682,N_8492);
or U8803 (N_8803,N_8595,N_8488);
nand U8804 (N_8804,N_8522,N_8455);
or U8805 (N_8805,N_8648,N_8440);
nand U8806 (N_8806,N_8763,N_8732);
and U8807 (N_8807,N_8627,N_8783);
nand U8808 (N_8808,N_8694,N_8592);
and U8809 (N_8809,N_8442,N_8727);
and U8810 (N_8810,N_8553,N_8643);
xnor U8811 (N_8811,N_8497,N_8425);
and U8812 (N_8812,N_8608,N_8700);
xor U8813 (N_8813,N_8435,N_8605);
nand U8814 (N_8814,N_8529,N_8565);
nor U8815 (N_8815,N_8438,N_8656);
or U8816 (N_8816,N_8427,N_8730);
xnor U8817 (N_8817,N_8658,N_8657);
or U8818 (N_8818,N_8786,N_8638);
nor U8819 (N_8819,N_8487,N_8717);
xnor U8820 (N_8820,N_8702,N_8422);
nand U8821 (N_8821,N_8517,N_8486);
and U8822 (N_8822,N_8527,N_8654);
nand U8823 (N_8823,N_8568,N_8646);
and U8824 (N_8824,N_8647,N_8613);
nor U8825 (N_8825,N_8535,N_8621);
and U8826 (N_8826,N_8401,N_8687);
and U8827 (N_8827,N_8408,N_8799);
and U8828 (N_8828,N_8505,N_8411);
nor U8829 (N_8829,N_8521,N_8728);
nand U8830 (N_8830,N_8641,N_8457);
nand U8831 (N_8831,N_8432,N_8630);
or U8832 (N_8832,N_8499,N_8580);
or U8833 (N_8833,N_8752,N_8761);
and U8834 (N_8834,N_8746,N_8731);
or U8835 (N_8835,N_8566,N_8669);
xor U8836 (N_8836,N_8779,N_8410);
xnor U8837 (N_8837,N_8426,N_8644);
and U8838 (N_8838,N_8631,N_8675);
or U8839 (N_8839,N_8639,N_8788);
xnor U8840 (N_8840,N_8551,N_8526);
xor U8841 (N_8841,N_8473,N_8636);
nor U8842 (N_8842,N_8528,N_8572);
nor U8843 (N_8843,N_8453,N_8742);
nor U8844 (N_8844,N_8692,N_8478);
xor U8845 (N_8845,N_8449,N_8718);
nand U8846 (N_8846,N_8691,N_8650);
nand U8847 (N_8847,N_8753,N_8738);
xor U8848 (N_8848,N_8481,N_8543);
xnor U8849 (N_8849,N_8663,N_8744);
xor U8850 (N_8850,N_8604,N_8445);
nor U8851 (N_8851,N_8689,N_8634);
or U8852 (N_8852,N_8587,N_8405);
and U8853 (N_8853,N_8552,N_8433);
xnor U8854 (N_8854,N_8520,N_8768);
nand U8855 (N_8855,N_8640,N_8791);
and U8856 (N_8856,N_8655,N_8705);
or U8857 (N_8857,N_8671,N_8429);
nor U8858 (N_8858,N_8450,N_8562);
nand U8859 (N_8859,N_8780,N_8794);
nand U8860 (N_8860,N_8414,N_8620);
or U8861 (N_8861,N_8710,N_8515);
or U8862 (N_8862,N_8494,N_8476);
nor U8863 (N_8863,N_8574,N_8769);
or U8864 (N_8864,N_8696,N_8525);
xnor U8865 (N_8865,N_8510,N_8558);
and U8866 (N_8866,N_8404,N_8496);
and U8867 (N_8867,N_8623,N_8512);
nand U8868 (N_8868,N_8632,N_8725);
or U8869 (N_8869,N_8561,N_8706);
and U8870 (N_8870,N_8452,N_8614);
and U8871 (N_8871,N_8578,N_8424);
nand U8872 (N_8872,N_8686,N_8491);
and U8873 (N_8873,N_8795,N_8609);
or U8874 (N_8874,N_8617,N_8736);
nand U8875 (N_8875,N_8420,N_8530);
nand U8876 (N_8876,N_8628,N_8431);
and U8877 (N_8877,N_8653,N_8774);
and U8878 (N_8878,N_8518,N_8667);
or U8879 (N_8879,N_8743,N_8511);
or U8880 (N_8880,N_8550,N_8524);
nor U8881 (N_8881,N_8469,N_8498);
and U8882 (N_8882,N_8541,N_8575);
or U8883 (N_8883,N_8747,N_8724);
and U8884 (N_8884,N_8439,N_8461);
nand U8885 (N_8885,N_8721,N_8502);
or U8886 (N_8886,N_8619,N_8597);
or U8887 (N_8887,N_8489,N_8599);
nor U8888 (N_8888,N_8423,N_8602);
nand U8889 (N_8889,N_8600,N_8436);
or U8890 (N_8890,N_8661,N_8665);
xnor U8891 (N_8891,N_8538,N_8585);
xnor U8892 (N_8892,N_8466,N_8635);
or U8893 (N_8893,N_8737,N_8506);
and U8894 (N_8894,N_8775,N_8699);
xnor U8895 (N_8895,N_8790,N_8548);
and U8896 (N_8896,N_8662,N_8701);
and U8897 (N_8897,N_8674,N_8723);
nand U8898 (N_8898,N_8468,N_8485);
nand U8899 (N_8899,N_8570,N_8523);
nand U8900 (N_8900,N_8680,N_8633);
or U8901 (N_8901,N_8428,N_8733);
xnor U8902 (N_8902,N_8532,N_8475);
and U8903 (N_8903,N_8579,N_8772);
nand U8904 (N_8904,N_8569,N_8765);
nor U8905 (N_8905,N_8516,N_8584);
and U8906 (N_8906,N_8708,N_8479);
or U8907 (N_8907,N_8666,N_8484);
nand U8908 (N_8908,N_8659,N_8500);
nand U8909 (N_8909,N_8531,N_8714);
xnor U8910 (N_8910,N_8402,N_8451);
or U8911 (N_8911,N_8734,N_8465);
or U8912 (N_8912,N_8622,N_8651);
xnor U8913 (N_8913,N_8434,N_8764);
nor U8914 (N_8914,N_8509,N_8537);
nor U8915 (N_8915,N_8698,N_8462);
and U8916 (N_8916,N_8787,N_8582);
xnor U8917 (N_8917,N_8754,N_8618);
or U8918 (N_8918,N_8418,N_8467);
and U8919 (N_8919,N_8480,N_8777);
xnor U8920 (N_8920,N_8493,N_8782);
nand U8921 (N_8921,N_8715,N_8773);
xor U8922 (N_8922,N_8611,N_8626);
nor U8923 (N_8923,N_8472,N_8759);
nor U8924 (N_8924,N_8533,N_8456);
and U8925 (N_8925,N_8606,N_8771);
xor U8926 (N_8926,N_8668,N_8751);
xnor U8927 (N_8927,N_8474,N_8583);
nor U8928 (N_8928,N_8697,N_8564);
and U8929 (N_8929,N_8546,N_8762);
or U8930 (N_8930,N_8798,N_8625);
xor U8931 (N_8931,N_8704,N_8495);
and U8932 (N_8932,N_8792,N_8660);
and U8933 (N_8933,N_8471,N_8672);
xor U8934 (N_8934,N_8598,N_8610);
xor U8935 (N_8935,N_8707,N_8403);
xor U8936 (N_8936,N_8588,N_8560);
xor U8937 (N_8937,N_8416,N_8735);
nand U8938 (N_8938,N_8557,N_8693);
nor U8939 (N_8939,N_8603,N_8419);
xnor U8940 (N_8940,N_8415,N_8748);
nand U8941 (N_8941,N_8470,N_8785);
nand U8942 (N_8942,N_8591,N_8417);
xor U8943 (N_8943,N_8757,N_8464);
nor U8944 (N_8944,N_8454,N_8594);
nor U8945 (N_8945,N_8616,N_8784);
xor U8946 (N_8946,N_8443,N_8673);
nor U8947 (N_8947,N_8571,N_8463);
or U8948 (N_8948,N_8750,N_8596);
and U8949 (N_8949,N_8519,N_8712);
or U8950 (N_8950,N_8615,N_8501);
or U8951 (N_8951,N_8676,N_8679);
nand U8952 (N_8952,N_8760,N_8504);
and U8953 (N_8953,N_8776,N_8683);
nor U8954 (N_8954,N_8444,N_8503);
and U8955 (N_8955,N_8581,N_8545);
xor U8956 (N_8956,N_8720,N_8690);
nand U8957 (N_8957,N_8678,N_8547);
nand U8958 (N_8958,N_8601,N_8586);
xnor U8959 (N_8959,N_8756,N_8745);
or U8960 (N_8960,N_8577,N_8593);
nor U8961 (N_8961,N_8446,N_8448);
xnor U8962 (N_8962,N_8607,N_8508);
or U8963 (N_8963,N_8685,N_8441);
xor U8964 (N_8964,N_8749,N_8739);
or U8965 (N_8965,N_8797,N_8576);
and U8966 (N_8966,N_8536,N_8719);
xor U8967 (N_8967,N_8629,N_8540);
xor U8968 (N_8968,N_8766,N_8758);
xor U8969 (N_8969,N_8555,N_8729);
or U8970 (N_8970,N_8649,N_8437);
xnor U8971 (N_8971,N_8755,N_8483);
xor U8972 (N_8972,N_8534,N_8612);
or U8973 (N_8973,N_8460,N_8514);
xnor U8974 (N_8974,N_8695,N_8624);
and U8975 (N_8975,N_8507,N_8430);
xor U8976 (N_8976,N_8740,N_8590);
or U8977 (N_8977,N_8664,N_8767);
and U8978 (N_8978,N_8645,N_8781);
xnor U8979 (N_8979,N_8793,N_8482);
nor U8980 (N_8980,N_8703,N_8458);
xnor U8981 (N_8981,N_8770,N_8567);
nor U8982 (N_8982,N_8741,N_8711);
and U8983 (N_8983,N_8559,N_8652);
nand U8984 (N_8984,N_8513,N_8677);
or U8985 (N_8985,N_8722,N_8539);
or U8986 (N_8986,N_8400,N_8477);
and U8987 (N_8987,N_8789,N_8542);
and U8988 (N_8988,N_8447,N_8554);
nand U8989 (N_8989,N_8796,N_8406);
and U8990 (N_8990,N_8556,N_8713);
nand U8991 (N_8991,N_8716,N_8642);
and U8992 (N_8992,N_8490,N_8407);
nand U8993 (N_8993,N_8670,N_8688);
and U8994 (N_8994,N_8778,N_8637);
nand U8995 (N_8995,N_8684,N_8459);
or U8996 (N_8996,N_8413,N_8409);
xor U8997 (N_8997,N_8412,N_8549);
nor U8998 (N_8998,N_8544,N_8681);
or U8999 (N_8999,N_8726,N_8563);
xor U9000 (N_9000,N_8507,N_8547);
nor U9001 (N_9001,N_8582,N_8621);
xor U9002 (N_9002,N_8511,N_8643);
or U9003 (N_9003,N_8561,N_8440);
or U9004 (N_9004,N_8748,N_8518);
nor U9005 (N_9005,N_8523,N_8455);
or U9006 (N_9006,N_8665,N_8790);
xor U9007 (N_9007,N_8512,N_8555);
nand U9008 (N_9008,N_8624,N_8731);
and U9009 (N_9009,N_8660,N_8615);
nand U9010 (N_9010,N_8446,N_8631);
xor U9011 (N_9011,N_8584,N_8427);
xnor U9012 (N_9012,N_8661,N_8571);
nand U9013 (N_9013,N_8570,N_8711);
or U9014 (N_9014,N_8691,N_8615);
or U9015 (N_9015,N_8749,N_8459);
or U9016 (N_9016,N_8432,N_8733);
xor U9017 (N_9017,N_8789,N_8796);
xor U9018 (N_9018,N_8502,N_8707);
nand U9019 (N_9019,N_8540,N_8544);
or U9020 (N_9020,N_8473,N_8647);
or U9021 (N_9021,N_8536,N_8433);
or U9022 (N_9022,N_8651,N_8702);
or U9023 (N_9023,N_8539,N_8532);
or U9024 (N_9024,N_8759,N_8487);
nand U9025 (N_9025,N_8773,N_8630);
or U9026 (N_9026,N_8421,N_8768);
xnor U9027 (N_9027,N_8492,N_8416);
or U9028 (N_9028,N_8775,N_8646);
or U9029 (N_9029,N_8404,N_8599);
nor U9030 (N_9030,N_8408,N_8459);
xnor U9031 (N_9031,N_8746,N_8516);
xor U9032 (N_9032,N_8484,N_8727);
nand U9033 (N_9033,N_8658,N_8520);
xor U9034 (N_9034,N_8452,N_8573);
xnor U9035 (N_9035,N_8615,N_8552);
and U9036 (N_9036,N_8661,N_8401);
xnor U9037 (N_9037,N_8409,N_8608);
or U9038 (N_9038,N_8703,N_8552);
or U9039 (N_9039,N_8688,N_8501);
or U9040 (N_9040,N_8418,N_8443);
and U9041 (N_9041,N_8627,N_8433);
or U9042 (N_9042,N_8619,N_8564);
or U9043 (N_9043,N_8424,N_8701);
xnor U9044 (N_9044,N_8728,N_8425);
xor U9045 (N_9045,N_8657,N_8529);
and U9046 (N_9046,N_8767,N_8558);
and U9047 (N_9047,N_8636,N_8630);
or U9048 (N_9048,N_8474,N_8492);
nand U9049 (N_9049,N_8502,N_8407);
and U9050 (N_9050,N_8415,N_8703);
and U9051 (N_9051,N_8561,N_8549);
or U9052 (N_9052,N_8453,N_8669);
xor U9053 (N_9053,N_8472,N_8753);
xor U9054 (N_9054,N_8459,N_8528);
and U9055 (N_9055,N_8607,N_8789);
nand U9056 (N_9056,N_8474,N_8452);
or U9057 (N_9057,N_8520,N_8798);
or U9058 (N_9058,N_8488,N_8493);
and U9059 (N_9059,N_8709,N_8693);
nor U9060 (N_9060,N_8470,N_8460);
or U9061 (N_9061,N_8790,N_8624);
and U9062 (N_9062,N_8520,N_8611);
xnor U9063 (N_9063,N_8684,N_8786);
nand U9064 (N_9064,N_8596,N_8513);
xor U9065 (N_9065,N_8627,N_8647);
xnor U9066 (N_9066,N_8524,N_8655);
or U9067 (N_9067,N_8462,N_8426);
nor U9068 (N_9068,N_8761,N_8732);
or U9069 (N_9069,N_8607,N_8458);
nor U9070 (N_9070,N_8546,N_8424);
xor U9071 (N_9071,N_8713,N_8580);
or U9072 (N_9072,N_8574,N_8787);
nand U9073 (N_9073,N_8665,N_8436);
nor U9074 (N_9074,N_8545,N_8593);
and U9075 (N_9075,N_8720,N_8739);
xnor U9076 (N_9076,N_8622,N_8613);
xor U9077 (N_9077,N_8406,N_8427);
or U9078 (N_9078,N_8647,N_8617);
and U9079 (N_9079,N_8706,N_8743);
nand U9080 (N_9080,N_8720,N_8608);
nand U9081 (N_9081,N_8558,N_8692);
and U9082 (N_9082,N_8585,N_8441);
or U9083 (N_9083,N_8785,N_8701);
xor U9084 (N_9084,N_8455,N_8741);
xnor U9085 (N_9085,N_8595,N_8481);
and U9086 (N_9086,N_8753,N_8797);
and U9087 (N_9087,N_8643,N_8733);
nand U9088 (N_9088,N_8777,N_8674);
nor U9089 (N_9089,N_8619,N_8423);
or U9090 (N_9090,N_8667,N_8541);
and U9091 (N_9091,N_8410,N_8686);
xnor U9092 (N_9092,N_8480,N_8672);
xnor U9093 (N_9093,N_8526,N_8453);
or U9094 (N_9094,N_8515,N_8745);
or U9095 (N_9095,N_8778,N_8699);
and U9096 (N_9096,N_8787,N_8509);
nand U9097 (N_9097,N_8660,N_8661);
or U9098 (N_9098,N_8723,N_8489);
nor U9099 (N_9099,N_8418,N_8608);
nor U9100 (N_9100,N_8701,N_8570);
xnor U9101 (N_9101,N_8693,N_8691);
xor U9102 (N_9102,N_8706,N_8587);
or U9103 (N_9103,N_8562,N_8771);
nor U9104 (N_9104,N_8775,N_8616);
and U9105 (N_9105,N_8741,N_8740);
or U9106 (N_9106,N_8770,N_8455);
nand U9107 (N_9107,N_8734,N_8613);
xnor U9108 (N_9108,N_8440,N_8419);
xor U9109 (N_9109,N_8769,N_8633);
nor U9110 (N_9110,N_8530,N_8725);
nor U9111 (N_9111,N_8523,N_8498);
and U9112 (N_9112,N_8607,N_8643);
xnor U9113 (N_9113,N_8713,N_8721);
or U9114 (N_9114,N_8765,N_8777);
nor U9115 (N_9115,N_8457,N_8590);
nand U9116 (N_9116,N_8422,N_8583);
nand U9117 (N_9117,N_8578,N_8719);
xnor U9118 (N_9118,N_8540,N_8787);
xor U9119 (N_9119,N_8617,N_8536);
nand U9120 (N_9120,N_8557,N_8750);
nand U9121 (N_9121,N_8527,N_8420);
nand U9122 (N_9122,N_8620,N_8582);
nor U9123 (N_9123,N_8549,N_8472);
nor U9124 (N_9124,N_8706,N_8760);
and U9125 (N_9125,N_8647,N_8721);
nand U9126 (N_9126,N_8463,N_8596);
xor U9127 (N_9127,N_8497,N_8406);
or U9128 (N_9128,N_8443,N_8454);
nand U9129 (N_9129,N_8517,N_8611);
nand U9130 (N_9130,N_8470,N_8702);
and U9131 (N_9131,N_8647,N_8412);
and U9132 (N_9132,N_8647,N_8629);
and U9133 (N_9133,N_8504,N_8480);
or U9134 (N_9134,N_8437,N_8670);
or U9135 (N_9135,N_8589,N_8527);
or U9136 (N_9136,N_8684,N_8589);
nor U9137 (N_9137,N_8532,N_8477);
nor U9138 (N_9138,N_8497,N_8555);
and U9139 (N_9139,N_8747,N_8401);
or U9140 (N_9140,N_8586,N_8537);
xor U9141 (N_9141,N_8480,N_8584);
and U9142 (N_9142,N_8723,N_8777);
nor U9143 (N_9143,N_8571,N_8427);
and U9144 (N_9144,N_8573,N_8443);
or U9145 (N_9145,N_8409,N_8422);
or U9146 (N_9146,N_8765,N_8475);
and U9147 (N_9147,N_8607,N_8584);
xnor U9148 (N_9148,N_8465,N_8446);
nor U9149 (N_9149,N_8616,N_8754);
xnor U9150 (N_9150,N_8652,N_8600);
nand U9151 (N_9151,N_8672,N_8680);
nand U9152 (N_9152,N_8671,N_8471);
nor U9153 (N_9153,N_8527,N_8767);
xor U9154 (N_9154,N_8482,N_8605);
or U9155 (N_9155,N_8425,N_8627);
nand U9156 (N_9156,N_8750,N_8690);
or U9157 (N_9157,N_8665,N_8624);
or U9158 (N_9158,N_8664,N_8701);
nor U9159 (N_9159,N_8612,N_8593);
nand U9160 (N_9160,N_8409,N_8792);
xnor U9161 (N_9161,N_8764,N_8457);
and U9162 (N_9162,N_8517,N_8465);
or U9163 (N_9163,N_8632,N_8747);
nor U9164 (N_9164,N_8611,N_8493);
and U9165 (N_9165,N_8431,N_8563);
or U9166 (N_9166,N_8531,N_8505);
nand U9167 (N_9167,N_8488,N_8472);
xor U9168 (N_9168,N_8621,N_8741);
nand U9169 (N_9169,N_8551,N_8574);
xor U9170 (N_9170,N_8690,N_8685);
nor U9171 (N_9171,N_8721,N_8518);
or U9172 (N_9172,N_8584,N_8707);
nor U9173 (N_9173,N_8633,N_8473);
or U9174 (N_9174,N_8681,N_8504);
nor U9175 (N_9175,N_8641,N_8608);
and U9176 (N_9176,N_8429,N_8547);
or U9177 (N_9177,N_8678,N_8461);
nand U9178 (N_9178,N_8715,N_8565);
xor U9179 (N_9179,N_8529,N_8616);
xor U9180 (N_9180,N_8759,N_8747);
nand U9181 (N_9181,N_8691,N_8692);
or U9182 (N_9182,N_8779,N_8729);
nor U9183 (N_9183,N_8772,N_8774);
xor U9184 (N_9184,N_8694,N_8747);
nand U9185 (N_9185,N_8580,N_8693);
or U9186 (N_9186,N_8667,N_8775);
and U9187 (N_9187,N_8589,N_8760);
nand U9188 (N_9188,N_8794,N_8543);
nor U9189 (N_9189,N_8651,N_8699);
nor U9190 (N_9190,N_8753,N_8430);
and U9191 (N_9191,N_8613,N_8724);
nor U9192 (N_9192,N_8575,N_8731);
xor U9193 (N_9193,N_8437,N_8683);
xor U9194 (N_9194,N_8759,N_8537);
or U9195 (N_9195,N_8799,N_8678);
or U9196 (N_9196,N_8444,N_8585);
nor U9197 (N_9197,N_8431,N_8496);
and U9198 (N_9198,N_8594,N_8624);
xor U9199 (N_9199,N_8517,N_8557);
nor U9200 (N_9200,N_8953,N_9189);
nor U9201 (N_9201,N_9027,N_8910);
nor U9202 (N_9202,N_8954,N_9157);
or U9203 (N_9203,N_8919,N_9191);
nand U9204 (N_9204,N_9033,N_8957);
or U9205 (N_9205,N_9041,N_8909);
xor U9206 (N_9206,N_9054,N_9156);
and U9207 (N_9207,N_9133,N_9056);
nor U9208 (N_9208,N_9097,N_9000);
xor U9209 (N_9209,N_8906,N_9175);
or U9210 (N_9210,N_8849,N_9153);
nand U9211 (N_9211,N_9063,N_8986);
or U9212 (N_9212,N_9155,N_8877);
and U9213 (N_9213,N_8895,N_8948);
and U9214 (N_9214,N_8868,N_9198);
xor U9215 (N_9215,N_8829,N_8854);
xnor U9216 (N_9216,N_9137,N_8968);
nor U9217 (N_9217,N_9001,N_9092);
or U9218 (N_9218,N_9106,N_8813);
and U9219 (N_9219,N_9003,N_8977);
and U9220 (N_9220,N_8822,N_9023);
and U9221 (N_9221,N_8860,N_8988);
and U9222 (N_9222,N_9008,N_8894);
nand U9223 (N_9223,N_8924,N_8866);
or U9224 (N_9224,N_9125,N_8956);
xnor U9225 (N_9225,N_8883,N_8819);
xnor U9226 (N_9226,N_9029,N_8992);
or U9227 (N_9227,N_8801,N_9192);
or U9228 (N_9228,N_9166,N_9094);
xnor U9229 (N_9229,N_8980,N_9121);
or U9230 (N_9230,N_8820,N_9176);
or U9231 (N_9231,N_9120,N_9140);
nand U9232 (N_9232,N_8961,N_9050);
nand U9233 (N_9233,N_9026,N_8929);
nor U9234 (N_9234,N_9044,N_9193);
nand U9235 (N_9235,N_8971,N_9061);
or U9236 (N_9236,N_8902,N_9078);
nand U9237 (N_9237,N_9196,N_8856);
xor U9238 (N_9238,N_8917,N_8925);
xnor U9239 (N_9239,N_9145,N_8888);
xor U9240 (N_9240,N_9055,N_9177);
and U9241 (N_9241,N_8940,N_9126);
or U9242 (N_9242,N_8809,N_8916);
and U9243 (N_9243,N_9197,N_9031);
and U9244 (N_9244,N_8846,N_9181);
nand U9245 (N_9245,N_8978,N_8833);
or U9246 (N_9246,N_9080,N_9010);
or U9247 (N_9247,N_8999,N_8848);
nand U9248 (N_9248,N_8914,N_8807);
nand U9249 (N_9249,N_8941,N_9062);
or U9250 (N_9250,N_8885,N_8896);
and U9251 (N_9251,N_9169,N_9134);
or U9252 (N_9252,N_8943,N_8951);
and U9253 (N_9253,N_9194,N_8959);
nor U9254 (N_9254,N_8963,N_9038);
and U9255 (N_9255,N_9084,N_9128);
nor U9256 (N_9256,N_8931,N_8964);
and U9257 (N_9257,N_8975,N_8950);
and U9258 (N_9258,N_9099,N_8826);
nand U9259 (N_9259,N_8926,N_9188);
xor U9260 (N_9260,N_9164,N_9087);
and U9261 (N_9261,N_8874,N_9129);
xnor U9262 (N_9262,N_9086,N_8840);
nand U9263 (N_9263,N_9187,N_9180);
and U9264 (N_9264,N_8811,N_8928);
and U9265 (N_9265,N_9105,N_9146);
nor U9266 (N_9266,N_9014,N_9048);
and U9267 (N_9267,N_8852,N_8962);
and U9268 (N_9268,N_8845,N_8984);
and U9269 (N_9269,N_9082,N_9045);
and U9270 (N_9270,N_9047,N_8979);
nor U9271 (N_9271,N_9163,N_8861);
nor U9272 (N_9272,N_8990,N_9037);
or U9273 (N_9273,N_8881,N_9046);
nor U9274 (N_9274,N_8805,N_8998);
or U9275 (N_9275,N_8933,N_9117);
and U9276 (N_9276,N_9182,N_9111);
nand U9277 (N_9277,N_9081,N_9042);
or U9278 (N_9278,N_9132,N_8994);
nor U9279 (N_9279,N_8955,N_8882);
or U9280 (N_9280,N_9100,N_8976);
and U9281 (N_9281,N_9183,N_8974);
nor U9282 (N_9282,N_9002,N_8891);
nor U9283 (N_9283,N_8949,N_9085);
nand U9284 (N_9284,N_8808,N_9112);
nor U9285 (N_9285,N_9013,N_9067);
nor U9286 (N_9286,N_8923,N_9124);
or U9287 (N_9287,N_8960,N_8837);
and U9288 (N_9288,N_9165,N_8899);
nor U9289 (N_9289,N_9119,N_9095);
xor U9290 (N_9290,N_8875,N_8841);
nor U9291 (N_9291,N_8814,N_9077);
and U9292 (N_9292,N_9016,N_9186);
and U9293 (N_9293,N_9007,N_9104);
or U9294 (N_9294,N_9174,N_8871);
xor U9295 (N_9295,N_9028,N_9079);
or U9296 (N_9296,N_9072,N_9139);
or U9297 (N_9297,N_9185,N_9049);
and U9298 (N_9298,N_8907,N_8869);
xor U9299 (N_9299,N_8802,N_8810);
and U9300 (N_9300,N_8939,N_9110);
nor U9301 (N_9301,N_9096,N_8985);
and U9302 (N_9302,N_9162,N_9093);
and U9303 (N_9303,N_8942,N_8884);
and U9304 (N_9304,N_8927,N_8838);
or U9305 (N_9305,N_9123,N_8993);
xor U9306 (N_9306,N_8872,N_9158);
and U9307 (N_9307,N_8911,N_9030);
xor U9308 (N_9308,N_8946,N_9136);
and U9309 (N_9309,N_8890,N_8969);
or U9310 (N_9310,N_8855,N_8997);
or U9311 (N_9311,N_9076,N_9089);
xnor U9312 (N_9312,N_8835,N_8870);
or U9313 (N_9313,N_8967,N_8815);
or U9314 (N_9314,N_8828,N_9103);
nor U9315 (N_9315,N_9160,N_9102);
nand U9316 (N_9316,N_9011,N_8818);
nor U9317 (N_9317,N_8966,N_9058);
nor U9318 (N_9318,N_8834,N_8862);
xnor U9319 (N_9319,N_8920,N_8832);
and U9320 (N_9320,N_9015,N_8867);
nand U9321 (N_9321,N_8847,N_8844);
xnor U9322 (N_9322,N_8842,N_9098);
or U9323 (N_9323,N_9149,N_8938);
or U9324 (N_9324,N_8937,N_8913);
xnor U9325 (N_9325,N_9069,N_9017);
or U9326 (N_9326,N_9118,N_8898);
xnor U9327 (N_9327,N_9195,N_8886);
nand U9328 (N_9328,N_9004,N_8887);
nor U9329 (N_9329,N_9068,N_9184);
and U9330 (N_9330,N_8851,N_9148);
or U9331 (N_9331,N_8973,N_9152);
nand U9332 (N_9332,N_8823,N_8982);
nor U9333 (N_9333,N_9108,N_8893);
xor U9334 (N_9334,N_9060,N_8857);
xor U9335 (N_9335,N_8825,N_8836);
and U9336 (N_9336,N_9170,N_9154);
or U9337 (N_9337,N_8880,N_8915);
nor U9338 (N_9338,N_9144,N_9130);
nand U9339 (N_9339,N_9053,N_9088);
and U9340 (N_9340,N_9059,N_9024);
nand U9341 (N_9341,N_8865,N_8903);
nand U9342 (N_9342,N_8981,N_9022);
and U9343 (N_9343,N_9074,N_9025);
and U9344 (N_9344,N_8863,N_9116);
xor U9345 (N_9345,N_8816,N_8876);
nand U9346 (N_9346,N_8804,N_9035);
xor U9347 (N_9347,N_8904,N_8803);
and U9348 (N_9348,N_8878,N_8912);
or U9349 (N_9349,N_9115,N_8864);
xnor U9350 (N_9350,N_9135,N_9173);
nand U9351 (N_9351,N_9159,N_9161);
or U9352 (N_9352,N_8905,N_9178);
xnor U9353 (N_9353,N_9065,N_8987);
nand U9354 (N_9354,N_8995,N_9199);
nor U9355 (N_9355,N_8947,N_9032);
or U9356 (N_9356,N_9009,N_8853);
or U9357 (N_9357,N_9142,N_9131);
xor U9358 (N_9358,N_9114,N_9127);
and U9359 (N_9359,N_9066,N_9113);
and U9360 (N_9360,N_9147,N_8945);
and U9361 (N_9361,N_9107,N_8934);
nor U9362 (N_9362,N_8989,N_8839);
nor U9363 (N_9363,N_9019,N_8996);
nor U9364 (N_9364,N_9083,N_8827);
or U9365 (N_9365,N_8983,N_9075);
xor U9366 (N_9366,N_9021,N_8830);
nand U9367 (N_9367,N_9143,N_9090);
nand U9368 (N_9368,N_8817,N_9150);
nor U9369 (N_9369,N_8944,N_8935);
nor U9370 (N_9370,N_8824,N_8873);
nor U9371 (N_9371,N_9109,N_9167);
nor U9372 (N_9372,N_9091,N_8858);
nand U9373 (N_9373,N_8831,N_9073);
or U9374 (N_9374,N_9071,N_8821);
nor U9375 (N_9375,N_8921,N_9043);
nand U9376 (N_9376,N_8850,N_9171);
nor U9377 (N_9377,N_8879,N_8901);
and U9378 (N_9378,N_8859,N_9057);
or U9379 (N_9379,N_8812,N_9006);
nand U9380 (N_9380,N_9020,N_8958);
xor U9381 (N_9381,N_9151,N_8908);
nor U9382 (N_9382,N_8952,N_9168);
nor U9383 (N_9383,N_8892,N_8932);
or U9384 (N_9384,N_8918,N_9101);
nand U9385 (N_9385,N_9122,N_9012);
xnor U9386 (N_9386,N_8843,N_9005);
or U9387 (N_9387,N_8930,N_9172);
nor U9388 (N_9388,N_8965,N_9141);
or U9389 (N_9389,N_9034,N_8936);
and U9390 (N_9390,N_9052,N_8806);
xor U9391 (N_9391,N_9064,N_9190);
xnor U9392 (N_9392,N_8800,N_8889);
nand U9393 (N_9393,N_8897,N_9051);
nor U9394 (N_9394,N_8972,N_9039);
nor U9395 (N_9395,N_8991,N_9070);
nor U9396 (N_9396,N_9018,N_9040);
or U9397 (N_9397,N_9138,N_8970);
nor U9398 (N_9398,N_8922,N_8900);
xnor U9399 (N_9399,N_9179,N_9036);
nand U9400 (N_9400,N_8828,N_8882);
and U9401 (N_9401,N_8811,N_8834);
xor U9402 (N_9402,N_8832,N_8994);
xnor U9403 (N_9403,N_9140,N_8927);
nand U9404 (N_9404,N_8843,N_9027);
xnor U9405 (N_9405,N_9052,N_8928);
and U9406 (N_9406,N_8972,N_8929);
or U9407 (N_9407,N_8829,N_8916);
or U9408 (N_9408,N_8908,N_8899);
xor U9409 (N_9409,N_8942,N_8839);
and U9410 (N_9410,N_9043,N_8806);
or U9411 (N_9411,N_8827,N_8973);
or U9412 (N_9412,N_9010,N_9009);
nand U9413 (N_9413,N_8997,N_8913);
nor U9414 (N_9414,N_8860,N_9028);
nand U9415 (N_9415,N_8898,N_8883);
and U9416 (N_9416,N_8821,N_9087);
or U9417 (N_9417,N_9022,N_9170);
and U9418 (N_9418,N_9000,N_8840);
and U9419 (N_9419,N_9002,N_9181);
nand U9420 (N_9420,N_8970,N_8931);
nand U9421 (N_9421,N_9190,N_8945);
or U9422 (N_9422,N_9096,N_8897);
nor U9423 (N_9423,N_8805,N_8936);
and U9424 (N_9424,N_9055,N_8910);
and U9425 (N_9425,N_9149,N_8861);
and U9426 (N_9426,N_8943,N_8904);
nand U9427 (N_9427,N_8851,N_9038);
xnor U9428 (N_9428,N_9142,N_8838);
nand U9429 (N_9429,N_9058,N_9162);
xor U9430 (N_9430,N_8920,N_9195);
xor U9431 (N_9431,N_8862,N_9055);
and U9432 (N_9432,N_9110,N_8867);
nor U9433 (N_9433,N_8924,N_9061);
xnor U9434 (N_9434,N_8808,N_8922);
nand U9435 (N_9435,N_8873,N_9156);
and U9436 (N_9436,N_9047,N_8866);
nand U9437 (N_9437,N_8886,N_8812);
xnor U9438 (N_9438,N_8958,N_8844);
nor U9439 (N_9439,N_9037,N_8975);
xor U9440 (N_9440,N_9053,N_8808);
nand U9441 (N_9441,N_9181,N_9075);
xor U9442 (N_9442,N_9112,N_9062);
xnor U9443 (N_9443,N_9012,N_8865);
nand U9444 (N_9444,N_9072,N_9000);
xnor U9445 (N_9445,N_8857,N_9184);
xnor U9446 (N_9446,N_8944,N_9160);
and U9447 (N_9447,N_8884,N_8883);
and U9448 (N_9448,N_8845,N_8969);
or U9449 (N_9449,N_9131,N_8909);
and U9450 (N_9450,N_9047,N_9042);
xor U9451 (N_9451,N_9112,N_9109);
xnor U9452 (N_9452,N_8807,N_9016);
nor U9453 (N_9453,N_8884,N_9162);
xor U9454 (N_9454,N_8940,N_9183);
xnor U9455 (N_9455,N_8924,N_9161);
xor U9456 (N_9456,N_8879,N_9184);
nand U9457 (N_9457,N_9138,N_8826);
and U9458 (N_9458,N_9005,N_9157);
and U9459 (N_9459,N_9046,N_8937);
and U9460 (N_9460,N_8938,N_9137);
or U9461 (N_9461,N_9191,N_9131);
xnor U9462 (N_9462,N_8871,N_8966);
or U9463 (N_9463,N_9115,N_9071);
xnor U9464 (N_9464,N_8864,N_9151);
nand U9465 (N_9465,N_8969,N_8979);
and U9466 (N_9466,N_9164,N_8934);
and U9467 (N_9467,N_9138,N_8899);
nand U9468 (N_9468,N_8895,N_9170);
and U9469 (N_9469,N_8914,N_8866);
and U9470 (N_9470,N_8807,N_9130);
or U9471 (N_9471,N_8978,N_8913);
and U9472 (N_9472,N_8910,N_8879);
nand U9473 (N_9473,N_8899,N_8866);
and U9474 (N_9474,N_8971,N_8994);
or U9475 (N_9475,N_9117,N_9107);
nor U9476 (N_9476,N_9173,N_9058);
or U9477 (N_9477,N_9016,N_9023);
nor U9478 (N_9478,N_8987,N_9113);
or U9479 (N_9479,N_8951,N_9154);
nand U9480 (N_9480,N_9102,N_8907);
nand U9481 (N_9481,N_9125,N_9085);
nand U9482 (N_9482,N_9035,N_9044);
nor U9483 (N_9483,N_8961,N_8950);
and U9484 (N_9484,N_8957,N_9183);
nor U9485 (N_9485,N_9123,N_9156);
and U9486 (N_9486,N_9008,N_9147);
nor U9487 (N_9487,N_9153,N_8882);
or U9488 (N_9488,N_9000,N_8825);
nor U9489 (N_9489,N_9004,N_8926);
nor U9490 (N_9490,N_9075,N_9048);
or U9491 (N_9491,N_9143,N_8875);
nand U9492 (N_9492,N_9102,N_8910);
and U9493 (N_9493,N_9036,N_8812);
xor U9494 (N_9494,N_8936,N_8818);
and U9495 (N_9495,N_9109,N_9023);
and U9496 (N_9496,N_9063,N_8889);
and U9497 (N_9497,N_8873,N_8858);
nor U9498 (N_9498,N_8817,N_8822);
xnor U9499 (N_9499,N_8837,N_9033);
nand U9500 (N_9500,N_9139,N_8971);
or U9501 (N_9501,N_8981,N_9040);
and U9502 (N_9502,N_9134,N_9088);
xor U9503 (N_9503,N_9033,N_9024);
nor U9504 (N_9504,N_8904,N_8908);
and U9505 (N_9505,N_9007,N_8923);
xor U9506 (N_9506,N_8909,N_9026);
nor U9507 (N_9507,N_8958,N_9058);
nand U9508 (N_9508,N_8881,N_9195);
xor U9509 (N_9509,N_8817,N_8939);
nand U9510 (N_9510,N_9093,N_9058);
and U9511 (N_9511,N_9119,N_9109);
or U9512 (N_9512,N_9054,N_9150);
nand U9513 (N_9513,N_9135,N_8875);
nor U9514 (N_9514,N_9087,N_8841);
nor U9515 (N_9515,N_9086,N_9064);
or U9516 (N_9516,N_9056,N_9017);
nor U9517 (N_9517,N_8935,N_8950);
nand U9518 (N_9518,N_9070,N_8996);
or U9519 (N_9519,N_9197,N_9026);
nor U9520 (N_9520,N_8856,N_9197);
xor U9521 (N_9521,N_9161,N_9082);
and U9522 (N_9522,N_8867,N_9090);
nor U9523 (N_9523,N_8888,N_9127);
nand U9524 (N_9524,N_9134,N_8928);
xor U9525 (N_9525,N_9134,N_8938);
or U9526 (N_9526,N_9174,N_9198);
and U9527 (N_9527,N_9033,N_8841);
nor U9528 (N_9528,N_9197,N_8834);
and U9529 (N_9529,N_8924,N_8912);
or U9530 (N_9530,N_9129,N_8901);
nand U9531 (N_9531,N_9057,N_8942);
nand U9532 (N_9532,N_8993,N_8919);
nor U9533 (N_9533,N_8878,N_8868);
and U9534 (N_9534,N_8878,N_8948);
and U9535 (N_9535,N_9117,N_9036);
and U9536 (N_9536,N_8977,N_9113);
and U9537 (N_9537,N_9035,N_9116);
xor U9538 (N_9538,N_8836,N_9079);
nand U9539 (N_9539,N_8938,N_8912);
and U9540 (N_9540,N_8846,N_9161);
nor U9541 (N_9541,N_8820,N_9198);
or U9542 (N_9542,N_8979,N_9120);
xor U9543 (N_9543,N_8993,N_8964);
xnor U9544 (N_9544,N_8812,N_8933);
and U9545 (N_9545,N_9049,N_9128);
nor U9546 (N_9546,N_9060,N_9073);
or U9547 (N_9547,N_9002,N_9193);
and U9548 (N_9548,N_9072,N_8831);
nand U9549 (N_9549,N_8854,N_8935);
xnor U9550 (N_9550,N_9133,N_9165);
nor U9551 (N_9551,N_8994,N_8987);
nor U9552 (N_9552,N_9017,N_8908);
nor U9553 (N_9553,N_8944,N_8858);
nand U9554 (N_9554,N_8819,N_9021);
nor U9555 (N_9555,N_8870,N_8836);
xor U9556 (N_9556,N_8897,N_8804);
nand U9557 (N_9557,N_8987,N_9198);
nor U9558 (N_9558,N_9061,N_9146);
nand U9559 (N_9559,N_8802,N_9083);
or U9560 (N_9560,N_9094,N_9040);
nand U9561 (N_9561,N_8857,N_8921);
and U9562 (N_9562,N_8972,N_8953);
nor U9563 (N_9563,N_8930,N_8810);
or U9564 (N_9564,N_8901,N_9137);
nand U9565 (N_9565,N_8895,N_8962);
nand U9566 (N_9566,N_9018,N_8860);
and U9567 (N_9567,N_9004,N_8849);
xor U9568 (N_9568,N_8908,N_9188);
or U9569 (N_9569,N_8895,N_9162);
or U9570 (N_9570,N_8971,N_9182);
nand U9571 (N_9571,N_9105,N_8856);
nand U9572 (N_9572,N_9128,N_8984);
nand U9573 (N_9573,N_8835,N_9171);
and U9574 (N_9574,N_9192,N_9181);
xor U9575 (N_9575,N_9149,N_9005);
and U9576 (N_9576,N_9146,N_9079);
nor U9577 (N_9577,N_8964,N_9185);
nor U9578 (N_9578,N_8932,N_9116);
and U9579 (N_9579,N_9164,N_9061);
nand U9580 (N_9580,N_9088,N_9004);
nand U9581 (N_9581,N_8892,N_9101);
nand U9582 (N_9582,N_8900,N_9003);
xor U9583 (N_9583,N_9146,N_9164);
or U9584 (N_9584,N_9037,N_9005);
xor U9585 (N_9585,N_9138,N_8971);
or U9586 (N_9586,N_8943,N_8881);
or U9587 (N_9587,N_9199,N_8967);
xor U9588 (N_9588,N_9090,N_9129);
nand U9589 (N_9589,N_9140,N_9090);
nand U9590 (N_9590,N_8890,N_9039);
and U9591 (N_9591,N_9181,N_8942);
and U9592 (N_9592,N_8845,N_9188);
or U9593 (N_9593,N_9139,N_9128);
nand U9594 (N_9594,N_9036,N_8933);
xnor U9595 (N_9595,N_9093,N_9020);
and U9596 (N_9596,N_8958,N_9097);
nor U9597 (N_9597,N_8968,N_9075);
or U9598 (N_9598,N_9006,N_9087);
and U9599 (N_9599,N_9178,N_8966);
or U9600 (N_9600,N_9541,N_9333);
xor U9601 (N_9601,N_9203,N_9436);
or U9602 (N_9602,N_9201,N_9451);
nand U9603 (N_9603,N_9434,N_9459);
nand U9604 (N_9604,N_9221,N_9574);
nand U9605 (N_9605,N_9249,N_9314);
nand U9606 (N_9606,N_9253,N_9258);
or U9607 (N_9607,N_9468,N_9293);
nand U9608 (N_9608,N_9353,N_9594);
and U9609 (N_9609,N_9402,N_9396);
nor U9610 (N_9610,N_9472,N_9483);
or U9611 (N_9611,N_9467,N_9323);
and U9612 (N_9612,N_9565,N_9235);
xnor U9613 (N_9613,N_9330,N_9456);
nand U9614 (N_9614,N_9567,N_9208);
or U9615 (N_9615,N_9283,N_9465);
and U9616 (N_9616,N_9386,N_9507);
nor U9617 (N_9617,N_9417,N_9497);
nor U9618 (N_9618,N_9534,N_9561);
xor U9619 (N_9619,N_9485,N_9550);
and U9620 (N_9620,N_9492,N_9343);
xor U9621 (N_9621,N_9202,N_9505);
nand U9622 (N_9622,N_9575,N_9345);
and U9623 (N_9623,N_9357,N_9511);
and U9624 (N_9624,N_9557,N_9289);
and U9625 (N_9625,N_9597,N_9522);
xor U9626 (N_9626,N_9301,N_9421);
or U9627 (N_9627,N_9475,N_9388);
nor U9628 (N_9628,N_9391,N_9564);
nor U9629 (N_9629,N_9205,N_9338);
nor U9630 (N_9630,N_9471,N_9241);
and U9631 (N_9631,N_9570,N_9577);
nor U9632 (N_9632,N_9429,N_9490);
nor U9633 (N_9633,N_9339,N_9347);
xnor U9634 (N_9634,N_9369,N_9584);
or U9635 (N_9635,N_9406,N_9445);
xor U9636 (N_9636,N_9237,N_9446);
nor U9637 (N_9637,N_9212,N_9447);
nor U9638 (N_9638,N_9498,N_9276);
or U9639 (N_9639,N_9502,N_9555);
nor U9640 (N_9640,N_9273,N_9458);
xor U9641 (N_9641,N_9440,N_9544);
and U9642 (N_9642,N_9482,N_9287);
nor U9643 (N_9643,N_9401,N_9332);
or U9644 (N_9644,N_9397,N_9556);
or U9645 (N_9645,N_9248,N_9500);
or U9646 (N_9646,N_9523,N_9364);
nand U9647 (N_9647,N_9243,N_9344);
xor U9648 (N_9648,N_9239,N_9449);
or U9649 (N_9649,N_9506,N_9317);
xor U9650 (N_9650,N_9328,N_9381);
nand U9651 (N_9651,N_9515,N_9372);
and U9652 (N_9652,N_9257,N_9540);
xnor U9653 (N_9653,N_9495,N_9304);
or U9654 (N_9654,N_9348,N_9591);
nand U9655 (N_9655,N_9399,N_9480);
or U9656 (N_9656,N_9285,N_9268);
nor U9657 (N_9657,N_9366,N_9494);
xor U9658 (N_9658,N_9501,N_9275);
nand U9659 (N_9659,N_9546,N_9443);
or U9660 (N_9660,N_9300,N_9519);
nor U9661 (N_9661,N_9595,N_9576);
and U9662 (N_9662,N_9588,N_9251);
nor U9663 (N_9663,N_9566,N_9309);
xor U9664 (N_9664,N_9466,N_9389);
and U9665 (N_9665,N_9259,N_9234);
or U9666 (N_9666,N_9213,N_9313);
nor U9667 (N_9667,N_9463,N_9418);
nor U9668 (N_9668,N_9263,N_9581);
and U9669 (N_9669,N_9315,N_9378);
nand U9670 (N_9670,N_9363,N_9413);
or U9671 (N_9671,N_9382,N_9593);
or U9672 (N_9672,N_9598,N_9295);
nand U9673 (N_9673,N_9512,N_9530);
nor U9674 (N_9674,N_9592,N_9298);
xnor U9675 (N_9675,N_9403,N_9392);
xor U9676 (N_9676,N_9587,N_9228);
or U9677 (N_9677,N_9279,N_9262);
and U9678 (N_9678,N_9528,N_9361);
nand U9679 (N_9679,N_9284,N_9321);
nand U9680 (N_9680,N_9337,N_9573);
nor U9681 (N_9681,N_9291,N_9329);
and U9682 (N_9682,N_9335,N_9322);
nand U9683 (N_9683,N_9521,N_9422);
nand U9684 (N_9684,N_9416,N_9297);
nor U9685 (N_9685,N_9231,N_9487);
nor U9686 (N_9686,N_9400,N_9367);
nor U9687 (N_9687,N_9374,N_9513);
xor U9688 (N_9688,N_9387,N_9486);
nor U9689 (N_9689,N_9217,N_9572);
and U9690 (N_9690,N_9256,N_9390);
nor U9691 (N_9691,N_9375,N_9219);
xnor U9692 (N_9692,N_9368,N_9305);
xor U9693 (N_9693,N_9408,N_9341);
or U9694 (N_9694,N_9517,N_9254);
nor U9695 (N_9695,N_9537,N_9438);
nand U9696 (N_9696,N_9450,N_9462);
xor U9697 (N_9697,N_9525,N_9342);
or U9698 (N_9698,N_9288,N_9373);
and U9699 (N_9699,N_9596,N_9479);
or U9700 (N_9700,N_9245,N_9589);
and U9701 (N_9701,N_9407,N_9412);
xor U9702 (N_9702,N_9457,N_9398);
and U9703 (N_9703,N_9559,N_9599);
nand U9704 (N_9704,N_9553,N_9433);
xnor U9705 (N_9705,N_9299,N_9265);
and U9706 (N_9706,N_9376,N_9370);
or U9707 (N_9707,N_9394,N_9281);
or U9708 (N_9708,N_9496,N_9210);
xor U9709 (N_9709,N_9377,N_9385);
nor U9710 (N_9710,N_9223,N_9358);
and U9711 (N_9711,N_9325,N_9215);
nor U9712 (N_9712,N_9426,N_9430);
nor U9713 (N_9713,N_9324,N_9542);
xnor U9714 (N_9714,N_9218,N_9545);
nor U9715 (N_9715,N_9539,N_9543);
xnor U9716 (N_9716,N_9508,N_9527);
or U9717 (N_9717,N_9535,N_9340);
xor U9718 (N_9718,N_9439,N_9504);
or U9719 (N_9719,N_9516,N_9461);
xor U9720 (N_9720,N_9225,N_9308);
xor U9721 (N_9721,N_9585,N_9319);
and U9722 (N_9722,N_9380,N_9520);
nor U9723 (N_9723,N_9247,N_9562);
and U9724 (N_9724,N_9278,N_9282);
xnor U9725 (N_9725,N_9242,N_9538);
xnor U9726 (N_9726,N_9514,N_9404);
and U9727 (N_9727,N_9209,N_9227);
nand U9728 (N_9728,N_9365,N_9302);
nand U9729 (N_9729,N_9316,N_9229);
nand U9730 (N_9730,N_9267,N_9427);
and U9731 (N_9731,N_9260,N_9336);
xor U9732 (N_9732,N_9533,N_9464);
xnor U9733 (N_9733,N_9435,N_9224);
or U9734 (N_9734,N_9294,N_9454);
and U9735 (N_9735,N_9264,N_9424);
and U9736 (N_9736,N_9230,N_9211);
xnor U9737 (N_9737,N_9232,N_9405);
xor U9738 (N_9738,N_9478,N_9437);
nand U9739 (N_9739,N_9200,N_9214);
and U9740 (N_9740,N_9549,N_9310);
nor U9741 (N_9741,N_9226,N_9583);
nor U9742 (N_9742,N_9448,N_9460);
or U9743 (N_9743,N_9477,N_9469);
nand U9744 (N_9744,N_9547,N_9306);
or U9745 (N_9745,N_9334,N_9356);
nor U9746 (N_9746,N_9270,N_9240);
nand U9747 (N_9747,N_9428,N_9238);
xor U9748 (N_9748,N_9255,N_9509);
or U9749 (N_9749,N_9425,N_9346);
or U9750 (N_9750,N_9423,N_9586);
nand U9751 (N_9751,N_9216,N_9488);
nor U9752 (N_9752,N_9371,N_9491);
or U9753 (N_9753,N_9307,N_9415);
nor U9754 (N_9754,N_9327,N_9420);
xor U9755 (N_9755,N_9350,N_9384);
xor U9756 (N_9756,N_9532,N_9452);
xor U9757 (N_9757,N_9571,N_9431);
or U9758 (N_9758,N_9455,N_9272);
nor U9759 (N_9759,N_9579,N_9551);
nand U9760 (N_9760,N_9531,N_9410);
nand U9761 (N_9761,N_9296,N_9362);
or U9762 (N_9762,N_9442,N_9470);
or U9763 (N_9763,N_9526,N_9548);
xor U9764 (N_9764,N_9578,N_9580);
and U9765 (N_9765,N_9499,N_9590);
xnor U9766 (N_9766,N_9252,N_9563);
nand U9767 (N_9767,N_9236,N_9354);
xnor U9768 (N_9768,N_9393,N_9569);
and U9769 (N_9769,N_9360,N_9441);
and U9770 (N_9770,N_9277,N_9331);
nor U9771 (N_9771,N_9453,N_9474);
xnor U9772 (N_9772,N_9473,N_9395);
and U9773 (N_9773,N_9383,N_9582);
and U9774 (N_9774,N_9286,N_9220);
xor U9775 (N_9775,N_9552,N_9529);
and U9776 (N_9776,N_9558,N_9351);
nand U9777 (N_9777,N_9419,N_9355);
xor U9778 (N_9778,N_9489,N_9311);
and U9779 (N_9779,N_9503,N_9484);
xor U9780 (N_9780,N_9444,N_9292);
or U9781 (N_9781,N_9414,N_9244);
or U9782 (N_9782,N_9207,N_9554);
xor U9783 (N_9783,N_9352,N_9280);
xor U9784 (N_9784,N_9560,N_9518);
xnor U9785 (N_9785,N_9326,N_9379);
and U9786 (N_9786,N_9432,N_9269);
xor U9787 (N_9787,N_9204,N_9303);
and U9788 (N_9788,N_9411,N_9409);
nor U9789 (N_9789,N_9493,N_9318);
and U9790 (N_9790,N_9320,N_9261);
nor U9791 (N_9791,N_9274,N_9266);
nand U9792 (N_9792,N_9206,N_9476);
and U9793 (N_9793,N_9271,N_9233);
and U9794 (N_9794,N_9510,N_9568);
nand U9795 (N_9795,N_9481,N_9359);
or U9796 (N_9796,N_9536,N_9349);
nor U9797 (N_9797,N_9290,N_9222);
and U9798 (N_9798,N_9524,N_9250);
nand U9799 (N_9799,N_9246,N_9312);
xor U9800 (N_9800,N_9354,N_9214);
nand U9801 (N_9801,N_9216,N_9568);
nand U9802 (N_9802,N_9397,N_9525);
nand U9803 (N_9803,N_9536,N_9270);
nand U9804 (N_9804,N_9507,N_9235);
xnor U9805 (N_9805,N_9255,N_9448);
nor U9806 (N_9806,N_9282,N_9489);
xnor U9807 (N_9807,N_9398,N_9502);
xnor U9808 (N_9808,N_9275,N_9420);
nand U9809 (N_9809,N_9475,N_9505);
xor U9810 (N_9810,N_9561,N_9518);
or U9811 (N_9811,N_9288,N_9509);
nand U9812 (N_9812,N_9288,N_9272);
nand U9813 (N_9813,N_9410,N_9465);
and U9814 (N_9814,N_9587,N_9461);
nand U9815 (N_9815,N_9533,N_9333);
and U9816 (N_9816,N_9460,N_9598);
and U9817 (N_9817,N_9476,N_9301);
nand U9818 (N_9818,N_9588,N_9396);
nor U9819 (N_9819,N_9351,N_9422);
nand U9820 (N_9820,N_9349,N_9422);
nand U9821 (N_9821,N_9376,N_9314);
or U9822 (N_9822,N_9291,N_9296);
xor U9823 (N_9823,N_9433,N_9465);
nor U9824 (N_9824,N_9452,N_9384);
nand U9825 (N_9825,N_9506,N_9397);
and U9826 (N_9826,N_9322,N_9455);
xnor U9827 (N_9827,N_9437,N_9315);
xnor U9828 (N_9828,N_9344,N_9284);
nor U9829 (N_9829,N_9357,N_9411);
or U9830 (N_9830,N_9580,N_9457);
xor U9831 (N_9831,N_9210,N_9545);
and U9832 (N_9832,N_9284,N_9526);
xnor U9833 (N_9833,N_9272,N_9319);
nand U9834 (N_9834,N_9505,N_9559);
or U9835 (N_9835,N_9322,N_9479);
or U9836 (N_9836,N_9407,N_9488);
nor U9837 (N_9837,N_9253,N_9537);
and U9838 (N_9838,N_9530,N_9485);
nor U9839 (N_9839,N_9201,N_9228);
or U9840 (N_9840,N_9599,N_9363);
nand U9841 (N_9841,N_9223,N_9301);
xnor U9842 (N_9842,N_9265,N_9264);
nand U9843 (N_9843,N_9423,N_9302);
xor U9844 (N_9844,N_9479,N_9348);
nor U9845 (N_9845,N_9240,N_9530);
and U9846 (N_9846,N_9436,N_9272);
nor U9847 (N_9847,N_9266,N_9359);
nor U9848 (N_9848,N_9499,N_9553);
nand U9849 (N_9849,N_9589,N_9581);
or U9850 (N_9850,N_9308,N_9266);
nand U9851 (N_9851,N_9440,N_9558);
and U9852 (N_9852,N_9247,N_9335);
xnor U9853 (N_9853,N_9296,N_9300);
and U9854 (N_9854,N_9551,N_9404);
nand U9855 (N_9855,N_9448,N_9459);
and U9856 (N_9856,N_9475,N_9301);
and U9857 (N_9857,N_9542,N_9411);
nor U9858 (N_9858,N_9551,N_9329);
and U9859 (N_9859,N_9551,N_9469);
nor U9860 (N_9860,N_9345,N_9305);
nor U9861 (N_9861,N_9507,N_9412);
nor U9862 (N_9862,N_9517,N_9392);
or U9863 (N_9863,N_9546,N_9241);
nor U9864 (N_9864,N_9348,N_9512);
nand U9865 (N_9865,N_9567,N_9280);
or U9866 (N_9866,N_9560,N_9212);
nor U9867 (N_9867,N_9468,N_9344);
and U9868 (N_9868,N_9222,N_9403);
nor U9869 (N_9869,N_9340,N_9577);
xnor U9870 (N_9870,N_9588,N_9534);
xor U9871 (N_9871,N_9213,N_9399);
or U9872 (N_9872,N_9389,N_9476);
nand U9873 (N_9873,N_9565,N_9339);
nand U9874 (N_9874,N_9219,N_9334);
or U9875 (N_9875,N_9398,N_9395);
nand U9876 (N_9876,N_9521,N_9450);
or U9877 (N_9877,N_9203,N_9480);
nand U9878 (N_9878,N_9368,N_9271);
xnor U9879 (N_9879,N_9468,N_9560);
or U9880 (N_9880,N_9500,N_9382);
or U9881 (N_9881,N_9498,N_9492);
xnor U9882 (N_9882,N_9330,N_9468);
and U9883 (N_9883,N_9451,N_9575);
xor U9884 (N_9884,N_9421,N_9308);
or U9885 (N_9885,N_9201,N_9492);
and U9886 (N_9886,N_9404,N_9343);
xnor U9887 (N_9887,N_9498,N_9456);
and U9888 (N_9888,N_9383,N_9406);
or U9889 (N_9889,N_9418,N_9385);
nor U9890 (N_9890,N_9559,N_9314);
xnor U9891 (N_9891,N_9450,N_9380);
and U9892 (N_9892,N_9573,N_9369);
or U9893 (N_9893,N_9596,N_9211);
xnor U9894 (N_9894,N_9402,N_9537);
nand U9895 (N_9895,N_9399,N_9243);
xor U9896 (N_9896,N_9389,N_9577);
or U9897 (N_9897,N_9567,N_9209);
nand U9898 (N_9898,N_9458,N_9397);
nor U9899 (N_9899,N_9519,N_9266);
nor U9900 (N_9900,N_9266,N_9279);
nand U9901 (N_9901,N_9547,N_9340);
and U9902 (N_9902,N_9491,N_9370);
xnor U9903 (N_9903,N_9449,N_9317);
and U9904 (N_9904,N_9241,N_9331);
nand U9905 (N_9905,N_9306,N_9471);
xor U9906 (N_9906,N_9282,N_9360);
or U9907 (N_9907,N_9216,N_9439);
nand U9908 (N_9908,N_9523,N_9317);
xnor U9909 (N_9909,N_9303,N_9502);
and U9910 (N_9910,N_9484,N_9585);
nor U9911 (N_9911,N_9330,N_9475);
and U9912 (N_9912,N_9520,N_9495);
nor U9913 (N_9913,N_9272,N_9507);
and U9914 (N_9914,N_9316,N_9586);
nand U9915 (N_9915,N_9570,N_9586);
or U9916 (N_9916,N_9464,N_9361);
nand U9917 (N_9917,N_9291,N_9230);
or U9918 (N_9918,N_9588,N_9567);
xor U9919 (N_9919,N_9504,N_9456);
or U9920 (N_9920,N_9372,N_9370);
xnor U9921 (N_9921,N_9324,N_9258);
nand U9922 (N_9922,N_9540,N_9492);
nor U9923 (N_9923,N_9226,N_9237);
xnor U9924 (N_9924,N_9247,N_9280);
nand U9925 (N_9925,N_9571,N_9403);
nand U9926 (N_9926,N_9289,N_9264);
nor U9927 (N_9927,N_9520,N_9234);
xnor U9928 (N_9928,N_9440,N_9406);
or U9929 (N_9929,N_9206,N_9201);
nor U9930 (N_9930,N_9216,N_9596);
xnor U9931 (N_9931,N_9564,N_9555);
nand U9932 (N_9932,N_9453,N_9331);
xor U9933 (N_9933,N_9399,N_9573);
xnor U9934 (N_9934,N_9202,N_9393);
or U9935 (N_9935,N_9468,N_9596);
and U9936 (N_9936,N_9415,N_9208);
nor U9937 (N_9937,N_9406,N_9253);
or U9938 (N_9938,N_9427,N_9442);
or U9939 (N_9939,N_9400,N_9350);
and U9940 (N_9940,N_9289,N_9597);
nor U9941 (N_9941,N_9282,N_9425);
nor U9942 (N_9942,N_9553,N_9267);
nand U9943 (N_9943,N_9325,N_9582);
nor U9944 (N_9944,N_9287,N_9338);
nor U9945 (N_9945,N_9491,N_9437);
or U9946 (N_9946,N_9547,N_9526);
and U9947 (N_9947,N_9575,N_9515);
nand U9948 (N_9948,N_9231,N_9558);
nor U9949 (N_9949,N_9287,N_9518);
or U9950 (N_9950,N_9346,N_9511);
and U9951 (N_9951,N_9345,N_9213);
xor U9952 (N_9952,N_9482,N_9242);
nor U9953 (N_9953,N_9428,N_9204);
nand U9954 (N_9954,N_9563,N_9569);
and U9955 (N_9955,N_9217,N_9230);
xor U9956 (N_9956,N_9375,N_9247);
xnor U9957 (N_9957,N_9378,N_9527);
nor U9958 (N_9958,N_9228,N_9317);
xor U9959 (N_9959,N_9553,N_9464);
nor U9960 (N_9960,N_9467,N_9443);
xnor U9961 (N_9961,N_9582,N_9464);
nor U9962 (N_9962,N_9350,N_9518);
or U9963 (N_9963,N_9257,N_9414);
or U9964 (N_9964,N_9326,N_9470);
xnor U9965 (N_9965,N_9556,N_9313);
or U9966 (N_9966,N_9335,N_9591);
nor U9967 (N_9967,N_9217,N_9529);
and U9968 (N_9968,N_9330,N_9409);
nand U9969 (N_9969,N_9319,N_9414);
nor U9970 (N_9970,N_9241,N_9446);
xnor U9971 (N_9971,N_9334,N_9247);
nor U9972 (N_9972,N_9576,N_9265);
nand U9973 (N_9973,N_9392,N_9336);
nor U9974 (N_9974,N_9369,N_9292);
and U9975 (N_9975,N_9587,N_9415);
and U9976 (N_9976,N_9393,N_9329);
xnor U9977 (N_9977,N_9440,N_9300);
nor U9978 (N_9978,N_9408,N_9224);
nor U9979 (N_9979,N_9496,N_9229);
or U9980 (N_9980,N_9451,N_9204);
and U9981 (N_9981,N_9335,N_9243);
nand U9982 (N_9982,N_9249,N_9349);
xor U9983 (N_9983,N_9220,N_9422);
and U9984 (N_9984,N_9295,N_9584);
nand U9985 (N_9985,N_9219,N_9566);
xor U9986 (N_9986,N_9260,N_9215);
nand U9987 (N_9987,N_9487,N_9287);
nand U9988 (N_9988,N_9271,N_9584);
or U9989 (N_9989,N_9378,N_9221);
or U9990 (N_9990,N_9282,N_9598);
nor U9991 (N_9991,N_9469,N_9369);
and U9992 (N_9992,N_9411,N_9235);
nor U9993 (N_9993,N_9380,N_9325);
or U9994 (N_9994,N_9563,N_9452);
and U9995 (N_9995,N_9434,N_9299);
xnor U9996 (N_9996,N_9200,N_9201);
nand U9997 (N_9997,N_9432,N_9510);
nand U9998 (N_9998,N_9553,N_9373);
nand U9999 (N_9999,N_9355,N_9225);
nor U10000 (N_10000,N_9650,N_9767);
nand U10001 (N_10001,N_9955,N_9969);
nand U10002 (N_10002,N_9823,N_9795);
nand U10003 (N_10003,N_9663,N_9886);
xor U10004 (N_10004,N_9732,N_9911);
nand U10005 (N_10005,N_9759,N_9742);
and U10006 (N_10006,N_9706,N_9646);
nor U10007 (N_10007,N_9756,N_9999);
and U10008 (N_10008,N_9679,N_9947);
and U10009 (N_10009,N_9612,N_9837);
or U10010 (N_10010,N_9858,N_9889);
or U10011 (N_10011,N_9676,N_9764);
xor U10012 (N_10012,N_9816,N_9623);
xnor U10013 (N_10013,N_9888,N_9794);
xnor U10014 (N_10014,N_9840,N_9920);
and U10015 (N_10015,N_9956,N_9899);
and U10016 (N_10016,N_9791,N_9687);
xnor U10017 (N_10017,N_9939,N_9748);
or U10018 (N_10018,N_9806,N_9730);
nand U10019 (N_10019,N_9965,N_9785);
and U10020 (N_10020,N_9616,N_9815);
or U10021 (N_10021,N_9707,N_9984);
nor U10022 (N_10022,N_9617,N_9949);
or U10023 (N_10023,N_9698,N_9752);
nand U10024 (N_10024,N_9803,N_9941);
or U10025 (N_10025,N_9692,N_9711);
xnor U10026 (N_10026,N_9709,N_9611);
nor U10027 (N_10027,N_9885,N_9626);
or U10028 (N_10028,N_9662,N_9808);
or U10029 (N_10029,N_9643,N_9772);
or U10030 (N_10030,N_9813,N_9876);
or U10031 (N_10031,N_9856,N_9935);
nand U10032 (N_10032,N_9980,N_9873);
xor U10033 (N_10033,N_9774,N_9710);
nand U10034 (N_10034,N_9838,N_9700);
nor U10035 (N_10035,N_9930,N_9918);
or U10036 (N_10036,N_9660,N_9685);
or U10037 (N_10037,N_9995,N_9655);
xnor U10038 (N_10038,N_9725,N_9983);
nor U10039 (N_10039,N_9945,N_9981);
nand U10040 (N_10040,N_9914,N_9847);
nor U10041 (N_10041,N_9619,N_9821);
nor U10042 (N_10042,N_9990,N_9627);
nor U10043 (N_10043,N_9780,N_9827);
xor U10044 (N_10044,N_9799,N_9971);
or U10045 (N_10045,N_9950,N_9943);
or U10046 (N_10046,N_9738,N_9970);
nor U10047 (N_10047,N_9861,N_9757);
or U10048 (N_10048,N_9686,N_9665);
xor U10049 (N_10049,N_9713,N_9677);
and U10050 (N_10050,N_9865,N_9620);
and U10051 (N_10051,N_9834,N_9849);
or U10052 (N_10052,N_9652,N_9664);
nor U10053 (N_10053,N_9609,N_9807);
xor U10054 (N_10054,N_9960,N_9697);
or U10055 (N_10055,N_9951,N_9605);
nor U10056 (N_10056,N_9681,N_9860);
xor U10057 (N_10057,N_9841,N_9831);
nand U10058 (N_10058,N_9937,N_9726);
or U10059 (N_10059,N_9670,N_9962);
nand U10060 (N_10060,N_9653,N_9910);
nand U10061 (N_10061,N_9703,N_9731);
nand U10062 (N_10062,N_9810,N_9695);
and U10063 (N_10063,N_9781,N_9933);
nand U10064 (N_10064,N_9690,N_9651);
and U10065 (N_10065,N_9875,N_9779);
nand U10066 (N_10066,N_9790,N_9606);
nand U10067 (N_10067,N_9744,N_9890);
or U10068 (N_10068,N_9870,N_9735);
and U10069 (N_10069,N_9901,N_9978);
nand U10070 (N_10070,N_9678,N_9832);
nor U10071 (N_10071,N_9966,N_9874);
nand U10072 (N_10072,N_9919,N_9629);
nand U10073 (N_10073,N_9701,N_9814);
or U10074 (N_10074,N_9603,N_9642);
nand U10075 (N_10075,N_9625,N_9777);
and U10076 (N_10076,N_9801,N_9867);
xnor U10077 (N_10077,N_9699,N_9908);
nor U10078 (N_10078,N_9974,N_9968);
nor U10079 (N_10079,N_9773,N_9887);
or U10080 (N_10080,N_9638,N_9724);
or U10081 (N_10081,N_9762,N_9877);
xnor U10082 (N_10082,N_9957,N_9891);
nand U10083 (N_10083,N_9739,N_9654);
nand U10084 (N_10084,N_9833,N_9944);
and U10085 (N_10085,N_9977,N_9909);
or U10086 (N_10086,N_9749,N_9880);
or U10087 (N_10087,N_9723,N_9936);
and U10088 (N_10088,N_9976,N_9751);
nand U10089 (N_10089,N_9859,N_9758);
xor U10090 (N_10090,N_9761,N_9649);
nand U10091 (N_10091,N_9932,N_9967);
or U10092 (N_10092,N_9869,N_9636);
or U10093 (N_10093,N_9826,N_9693);
and U10094 (N_10094,N_9668,N_9618);
xor U10095 (N_10095,N_9648,N_9997);
nor U10096 (N_10096,N_9953,N_9682);
and U10097 (N_10097,N_9848,N_9916);
or U10098 (N_10098,N_9793,N_9783);
nand U10099 (N_10099,N_9672,N_9963);
xor U10100 (N_10100,N_9893,N_9923);
or U10101 (N_10101,N_9716,N_9985);
and U10102 (N_10102,N_9982,N_9640);
and U10103 (N_10103,N_9647,N_9631);
nand U10104 (N_10104,N_9776,N_9720);
xor U10105 (N_10105,N_9610,N_9796);
xor U10106 (N_10106,N_9778,N_9879);
and U10107 (N_10107,N_9804,N_9721);
nand U10108 (N_10108,N_9775,N_9769);
nor U10109 (N_10109,N_9922,N_9798);
nor U10110 (N_10110,N_9819,N_9747);
nor U10111 (N_10111,N_9658,N_9750);
nor U10112 (N_10112,N_9714,N_9902);
nand U10113 (N_10113,N_9844,N_9717);
or U10114 (N_10114,N_9727,N_9866);
or U10115 (N_10115,N_9613,N_9883);
and U10116 (N_10116,N_9639,N_9702);
and U10117 (N_10117,N_9868,N_9818);
or U10118 (N_10118,N_9994,N_9782);
nor U10119 (N_10119,N_9946,N_9755);
and U10120 (N_10120,N_9928,N_9737);
nand U10121 (N_10121,N_9600,N_9952);
nor U10122 (N_10122,N_9975,N_9900);
xnor U10123 (N_10123,N_9671,N_9872);
and U10124 (N_10124,N_9661,N_9854);
nand U10125 (N_10125,N_9830,N_9674);
nor U10126 (N_10126,N_9934,N_9789);
or U10127 (N_10127,N_9787,N_9688);
nand U10128 (N_10128,N_9924,N_9903);
nor U10129 (N_10129,N_9728,N_9921);
xnor U10130 (N_10130,N_9917,N_9666);
and U10131 (N_10131,N_9855,N_9958);
nand U10132 (N_10132,N_9637,N_9753);
or U10133 (N_10133,N_9857,N_9766);
xor U10134 (N_10134,N_9635,N_9797);
or U10135 (N_10135,N_9771,N_9973);
and U10136 (N_10136,N_9878,N_9992);
or U10137 (N_10137,N_9770,N_9954);
nor U10138 (N_10138,N_9864,N_9927);
nor U10139 (N_10139,N_9843,N_9835);
and U10140 (N_10140,N_9667,N_9656);
nand U10141 (N_10141,N_9708,N_9897);
nand U10142 (N_10142,N_9628,N_9839);
nand U10143 (N_10143,N_9754,N_9904);
xor U10144 (N_10144,N_9733,N_9938);
xnor U10145 (N_10145,N_9895,N_9959);
nand U10146 (N_10146,N_9915,N_9632);
and U10147 (N_10147,N_9608,N_9786);
and U10148 (N_10148,N_9745,N_9998);
xor U10149 (N_10149,N_9669,N_9729);
nor U10150 (N_10150,N_9659,N_9817);
nand U10151 (N_10151,N_9683,N_9913);
or U10152 (N_10152,N_9705,N_9604);
xor U10153 (N_10153,N_9675,N_9800);
and U10154 (N_10154,N_9828,N_9940);
xor U10155 (N_10155,N_9722,N_9630);
xnor U10156 (N_10156,N_9906,N_9882);
xor U10157 (N_10157,N_9846,N_9602);
xor U10158 (N_10158,N_9607,N_9614);
xnor U10159 (N_10159,N_9948,N_9684);
nand U10160 (N_10160,N_9929,N_9993);
and U10161 (N_10161,N_9622,N_9746);
and U10162 (N_10162,N_9601,N_9760);
or U10163 (N_10163,N_9768,N_9712);
nand U10164 (N_10164,N_9972,N_9853);
nor U10165 (N_10165,N_9898,N_9740);
nor U10166 (N_10166,N_9905,N_9788);
and U10167 (N_10167,N_9765,N_9991);
or U10168 (N_10168,N_9633,N_9986);
nand U10169 (N_10169,N_9641,N_9734);
or U10170 (N_10170,N_9979,N_9704);
and U10171 (N_10171,N_9802,N_9812);
xor U10172 (N_10172,N_9996,N_9715);
nand U10173 (N_10173,N_9621,N_9842);
xor U10174 (N_10174,N_9926,N_9907);
and U10175 (N_10175,N_9634,N_9863);
and U10176 (N_10176,N_9894,N_9743);
xor U10177 (N_10177,N_9852,N_9696);
xnor U10178 (N_10178,N_9896,N_9942);
and U10179 (N_10179,N_9763,N_9884);
xnor U10180 (N_10180,N_9871,N_9736);
or U10181 (N_10181,N_9719,N_9836);
or U10182 (N_10182,N_9931,N_9673);
nor U10183 (N_10183,N_9718,N_9811);
xor U10184 (N_10184,N_9680,N_9689);
nor U10185 (N_10185,N_9912,N_9987);
or U10186 (N_10186,N_9694,N_9784);
xor U10187 (N_10187,N_9845,N_9851);
and U10188 (N_10188,N_9644,N_9615);
nand U10189 (N_10189,N_9824,N_9961);
nand U10190 (N_10190,N_9850,N_9829);
nor U10191 (N_10191,N_9881,N_9691);
nor U10192 (N_10192,N_9792,N_9741);
xor U10193 (N_10193,N_9820,N_9925);
or U10194 (N_10194,N_9989,N_9657);
and U10195 (N_10195,N_9825,N_9805);
nand U10196 (N_10196,N_9964,N_9645);
xnor U10197 (N_10197,N_9988,N_9892);
or U10198 (N_10198,N_9624,N_9862);
nand U10199 (N_10199,N_9822,N_9809);
and U10200 (N_10200,N_9656,N_9952);
nand U10201 (N_10201,N_9857,N_9649);
or U10202 (N_10202,N_9907,N_9815);
or U10203 (N_10203,N_9878,N_9932);
nor U10204 (N_10204,N_9974,N_9984);
and U10205 (N_10205,N_9747,N_9635);
nor U10206 (N_10206,N_9827,N_9752);
xor U10207 (N_10207,N_9860,N_9863);
nand U10208 (N_10208,N_9782,N_9917);
nand U10209 (N_10209,N_9817,N_9737);
nand U10210 (N_10210,N_9897,N_9603);
or U10211 (N_10211,N_9885,N_9989);
and U10212 (N_10212,N_9669,N_9998);
or U10213 (N_10213,N_9828,N_9992);
or U10214 (N_10214,N_9910,N_9603);
xnor U10215 (N_10215,N_9757,N_9838);
nor U10216 (N_10216,N_9655,N_9687);
or U10217 (N_10217,N_9721,N_9717);
and U10218 (N_10218,N_9925,N_9669);
or U10219 (N_10219,N_9640,N_9812);
xnor U10220 (N_10220,N_9926,N_9807);
or U10221 (N_10221,N_9688,N_9714);
xnor U10222 (N_10222,N_9839,N_9980);
and U10223 (N_10223,N_9634,N_9893);
or U10224 (N_10224,N_9967,N_9952);
or U10225 (N_10225,N_9900,N_9913);
or U10226 (N_10226,N_9698,N_9955);
nand U10227 (N_10227,N_9877,N_9741);
xnor U10228 (N_10228,N_9963,N_9983);
xor U10229 (N_10229,N_9881,N_9904);
xor U10230 (N_10230,N_9676,N_9987);
nor U10231 (N_10231,N_9703,N_9729);
xnor U10232 (N_10232,N_9681,N_9958);
nor U10233 (N_10233,N_9819,N_9949);
and U10234 (N_10234,N_9962,N_9920);
nand U10235 (N_10235,N_9950,N_9645);
or U10236 (N_10236,N_9940,N_9991);
nand U10237 (N_10237,N_9661,N_9626);
xor U10238 (N_10238,N_9631,N_9929);
nand U10239 (N_10239,N_9857,N_9675);
nor U10240 (N_10240,N_9621,N_9869);
or U10241 (N_10241,N_9821,N_9661);
xor U10242 (N_10242,N_9821,N_9642);
nand U10243 (N_10243,N_9869,N_9967);
nand U10244 (N_10244,N_9647,N_9704);
nand U10245 (N_10245,N_9929,N_9889);
and U10246 (N_10246,N_9887,N_9855);
xor U10247 (N_10247,N_9825,N_9640);
nor U10248 (N_10248,N_9910,N_9973);
or U10249 (N_10249,N_9856,N_9885);
xnor U10250 (N_10250,N_9758,N_9918);
and U10251 (N_10251,N_9901,N_9777);
xnor U10252 (N_10252,N_9722,N_9993);
or U10253 (N_10253,N_9713,N_9692);
xnor U10254 (N_10254,N_9940,N_9984);
or U10255 (N_10255,N_9882,N_9886);
nor U10256 (N_10256,N_9778,N_9979);
and U10257 (N_10257,N_9610,N_9674);
xnor U10258 (N_10258,N_9645,N_9916);
or U10259 (N_10259,N_9906,N_9744);
xnor U10260 (N_10260,N_9735,N_9813);
nor U10261 (N_10261,N_9939,N_9723);
nor U10262 (N_10262,N_9994,N_9907);
nor U10263 (N_10263,N_9872,N_9758);
or U10264 (N_10264,N_9646,N_9833);
xor U10265 (N_10265,N_9952,N_9729);
nor U10266 (N_10266,N_9732,N_9946);
or U10267 (N_10267,N_9945,N_9879);
xor U10268 (N_10268,N_9653,N_9793);
and U10269 (N_10269,N_9753,N_9977);
nor U10270 (N_10270,N_9941,N_9894);
nand U10271 (N_10271,N_9829,N_9981);
and U10272 (N_10272,N_9735,N_9885);
and U10273 (N_10273,N_9966,N_9885);
nand U10274 (N_10274,N_9903,N_9714);
or U10275 (N_10275,N_9871,N_9884);
xor U10276 (N_10276,N_9790,N_9827);
nor U10277 (N_10277,N_9806,N_9835);
xor U10278 (N_10278,N_9640,N_9976);
nand U10279 (N_10279,N_9697,N_9638);
xor U10280 (N_10280,N_9619,N_9891);
xnor U10281 (N_10281,N_9638,N_9937);
xor U10282 (N_10282,N_9838,N_9969);
nor U10283 (N_10283,N_9998,N_9816);
xor U10284 (N_10284,N_9737,N_9921);
and U10285 (N_10285,N_9698,N_9879);
xor U10286 (N_10286,N_9872,N_9621);
nor U10287 (N_10287,N_9834,N_9764);
xor U10288 (N_10288,N_9912,N_9913);
nor U10289 (N_10289,N_9825,N_9860);
xnor U10290 (N_10290,N_9609,N_9815);
or U10291 (N_10291,N_9999,N_9924);
or U10292 (N_10292,N_9640,N_9738);
or U10293 (N_10293,N_9993,N_9631);
and U10294 (N_10294,N_9996,N_9755);
or U10295 (N_10295,N_9742,N_9695);
nor U10296 (N_10296,N_9619,N_9657);
xor U10297 (N_10297,N_9667,N_9626);
nand U10298 (N_10298,N_9789,N_9871);
or U10299 (N_10299,N_9886,N_9613);
nand U10300 (N_10300,N_9708,N_9644);
nand U10301 (N_10301,N_9805,N_9863);
and U10302 (N_10302,N_9872,N_9980);
or U10303 (N_10303,N_9863,N_9735);
nor U10304 (N_10304,N_9826,N_9713);
nand U10305 (N_10305,N_9904,N_9840);
nor U10306 (N_10306,N_9706,N_9687);
and U10307 (N_10307,N_9944,N_9972);
and U10308 (N_10308,N_9636,N_9916);
or U10309 (N_10309,N_9941,N_9823);
and U10310 (N_10310,N_9610,N_9688);
nor U10311 (N_10311,N_9639,N_9632);
nor U10312 (N_10312,N_9671,N_9907);
and U10313 (N_10313,N_9887,N_9673);
or U10314 (N_10314,N_9807,N_9956);
xnor U10315 (N_10315,N_9662,N_9696);
or U10316 (N_10316,N_9899,N_9948);
or U10317 (N_10317,N_9963,N_9954);
and U10318 (N_10318,N_9888,N_9746);
and U10319 (N_10319,N_9876,N_9864);
xnor U10320 (N_10320,N_9934,N_9778);
nand U10321 (N_10321,N_9689,N_9932);
nor U10322 (N_10322,N_9822,N_9718);
or U10323 (N_10323,N_9921,N_9824);
and U10324 (N_10324,N_9685,N_9788);
nor U10325 (N_10325,N_9825,N_9866);
nand U10326 (N_10326,N_9706,N_9665);
and U10327 (N_10327,N_9751,N_9942);
and U10328 (N_10328,N_9668,N_9647);
nand U10329 (N_10329,N_9974,N_9737);
nor U10330 (N_10330,N_9784,N_9842);
and U10331 (N_10331,N_9638,N_9765);
nor U10332 (N_10332,N_9820,N_9662);
xor U10333 (N_10333,N_9786,N_9975);
nand U10334 (N_10334,N_9839,N_9651);
nand U10335 (N_10335,N_9631,N_9686);
and U10336 (N_10336,N_9819,N_9742);
and U10337 (N_10337,N_9925,N_9751);
nand U10338 (N_10338,N_9673,N_9624);
or U10339 (N_10339,N_9982,N_9979);
and U10340 (N_10340,N_9946,N_9777);
nor U10341 (N_10341,N_9616,N_9945);
nand U10342 (N_10342,N_9985,N_9932);
xnor U10343 (N_10343,N_9600,N_9617);
xnor U10344 (N_10344,N_9654,N_9626);
and U10345 (N_10345,N_9898,N_9678);
nor U10346 (N_10346,N_9864,N_9659);
xor U10347 (N_10347,N_9841,N_9696);
and U10348 (N_10348,N_9674,N_9700);
or U10349 (N_10349,N_9678,N_9619);
and U10350 (N_10350,N_9896,N_9673);
or U10351 (N_10351,N_9982,N_9903);
xnor U10352 (N_10352,N_9862,N_9977);
xnor U10353 (N_10353,N_9929,N_9770);
or U10354 (N_10354,N_9607,N_9613);
and U10355 (N_10355,N_9758,N_9894);
and U10356 (N_10356,N_9877,N_9756);
nor U10357 (N_10357,N_9746,N_9615);
xor U10358 (N_10358,N_9794,N_9626);
and U10359 (N_10359,N_9778,N_9637);
and U10360 (N_10360,N_9643,N_9704);
or U10361 (N_10361,N_9609,N_9635);
nand U10362 (N_10362,N_9655,N_9660);
nor U10363 (N_10363,N_9660,N_9859);
nor U10364 (N_10364,N_9912,N_9629);
xnor U10365 (N_10365,N_9776,N_9840);
nand U10366 (N_10366,N_9751,N_9957);
nand U10367 (N_10367,N_9602,N_9954);
nand U10368 (N_10368,N_9804,N_9966);
and U10369 (N_10369,N_9939,N_9729);
or U10370 (N_10370,N_9703,N_9759);
nand U10371 (N_10371,N_9663,N_9836);
nand U10372 (N_10372,N_9766,N_9719);
nand U10373 (N_10373,N_9900,N_9982);
xnor U10374 (N_10374,N_9617,N_9847);
nor U10375 (N_10375,N_9771,N_9876);
nor U10376 (N_10376,N_9777,N_9642);
or U10377 (N_10377,N_9788,N_9613);
nor U10378 (N_10378,N_9701,N_9789);
xor U10379 (N_10379,N_9623,N_9823);
or U10380 (N_10380,N_9951,N_9647);
nor U10381 (N_10381,N_9606,N_9973);
xor U10382 (N_10382,N_9981,N_9838);
nor U10383 (N_10383,N_9673,N_9895);
and U10384 (N_10384,N_9915,N_9985);
xnor U10385 (N_10385,N_9668,N_9868);
nor U10386 (N_10386,N_9736,N_9974);
nor U10387 (N_10387,N_9929,N_9998);
nor U10388 (N_10388,N_9976,N_9679);
or U10389 (N_10389,N_9647,N_9766);
xor U10390 (N_10390,N_9977,N_9641);
or U10391 (N_10391,N_9638,N_9979);
or U10392 (N_10392,N_9750,N_9996);
nand U10393 (N_10393,N_9776,N_9662);
and U10394 (N_10394,N_9938,N_9878);
nor U10395 (N_10395,N_9699,N_9973);
or U10396 (N_10396,N_9682,N_9817);
nand U10397 (N_10397,N_9600,N_9886);
nor U10398 (N_10398,N_9825,N_9725);
or U10399 (N_10399,N_9614,N_9932);
and U10400 (N_10400,N_10014,N_10217);
nand U10401 (N_10401,N_10054,N_10147);
and U10402 (N_10402,N_10202,N_10394);
xor U10403 (N_10403,N_10062,N_10192);
nand U10404 (N_10404,N_10281,N_10084);
nor U10405 (N_10405,N_10249,N_10396);
and U10406 (N_10406,N_10016,N_10384);
xor U10407 (N_10407,N_10068,N_10223);
xnor U10408 (N_10408,N_10166,N_10365);
nor U10409 (N_10409,N_10096,N_10033);
and U10410 (N_10410,N_10375,N_10034);
nor U10411 (N_10411,N_10133,N_10279);
and U10412 (N_10412,N_10051,N_10292);
nor U10413 (N_10413,N_10218,N_10081);
and U10414 (N_10414,N_10216,N_10162);
or U10415 (N_10415,N_10350,N_10304);
xnor U10416 (N_10416,N_10267,N_10328);
or U10417 (N_10417,N_10209,N_10040);
nand U10418 (N_10418,N_10399,N_10242);
and U10419 (N_10419,N_10335,N_10229);
nor U10420 (N_10420,N_10352,N_10036);
or U10421 (N_10421,N_10358,N_10385);
xor U10422 (N_10422,N_10230,N_10269);
xor U10423 (N_10423,N_10026,N_10342);
or U10424 (N_10424,N_10330,N_10397);
nand U10425 (N_10425,N_10232,N_10079);
xnor U10426 (N_10426,N_10088,N_10067);
nor U10427 (N_10427,N_10072,N_10241);
nor U10428 (N_10428,N_10271,N_10136);
xor U10429 (N_10429,N_10163,N_10322);
xnor U10430 (N_10430,N_10323,N_10295);
xnor U10431 (N_10431,N_10265,N_10102);
nor U10432 (N_10432,N_10076,N_10256);
or U10433 (N_10433,N_10336,N_10203);
nor U10434 (N_10434,N_10078,N_10128);
xnor U10435 (N_10435,N_10190,N_10169);
nor U10436 (N_10436,N_10387,N_10125);
xor U10437 (N_10437,N_10134,N_10297);
and U10438 (N_10438,N_10367,N_10383);
or U10439 (N_10439,N_10178,N_10082);
xnor U10440 (N_10440,N_10266,N_10346);
nor U10441 (N_10441,N_10332,N_10362);
and U10442 (N_10442,N_10161,N_10174);
nor U10443 (N_10443,N_10086,N_10364);
xnor U10444 (N_10444,N_10069,N_10188);
or U10445 (N_10445,N_10182,N_10318);
and U10446 (N_10446,N_10368,N_10061);
xnor U10447 (N_10447,N_10000,N_10184);
xor U10448 (N_10448,N_10371,N_10064);
and U10449 (N_10449,N_10018,N_10046);
and U10450 (N_10450,N_10165,N_10058);
nand U10451 (N_10451,N_10246,N_10329);
nand U10452 (N_10452,N_10037,N_10354);
and U10453 (N_10453,N_10199,N_10243);
or U10454 (N_10454,N_10347,N_10284);
and U10455 (N_10455,N_10282,N_10127);
nor U10456 (N_10456,N_10052,N_10020);
nor U10457 (N_10457,N_10010,N_10154);
nor U10458 (N_10458,N_10280,N_10025);
and U10459 (N_10459,N_10003,N_10255);
nand U10460 (N_10460,N_10183,N_10380);
and U10461 (N_10461,N_10213,N_10240);
or U10462 (N_10462,N_10310,N_10179);
and U10463 (N_10463,N_10032,N_10160);
nand U10464 (N_10464,N_10103,N_10348);
xor U10465 (N_10465,N_10234,N_10198);
nor U10466 (N_10466,N_10315,N_10378);
xor U10467 (N_10467,N_10044,N_10035);
nor U10468 (N_10468,N_10113,N_10248);
and U10469 (N_10469,N_10108,N_10028);
xnor U10470 (N_10470,N_10222,N_10070);
or U10471 (N_10471,N_10366,N_10355);
or U10472 (N_10472,N_10264,N_10293);
nand U10473 (N_10473,N_10090,N_10320);
nand U10474 (N_10474,N_10135,N_10272);
xnor U10475 (N_10475,N_10359,N_10050);
and U10476 (N_10476,N_10283,N_10080);
nor U10477 (N_10477,N_10122,N_10205);
nor U10478 (N_10478,N_10087,N_10031);
nor U10479 (N_10479,N_10057,N_10262);
and U10480 (N_10480,N_10009,N_10100);
nor U10481 (N_10481,N_10126,N_10194);
nor U10482 (N_10482,N_10305,N_10245);
nand U10483 (N_10483,N_10120,N_10116);
nor U10484 (N_10484,N_10024,N_10237);
or U10485 (N_10485,N_10388,N_10021);
and U10486 (N_10486,N_10075,N_10381);
nor U10487 (N_10487,N_10150,N_10290);
xnor U10488 (N_10488,N_10337,N_10309);
nand U10489 (N_10489,N_10112,N_10321);
nor U10490 (N_10490,N_10228,N_10386);
xnor U10491 (N_10491,N_10208,N_10093);
xor U10492 (N_10492,N_10236,N_10285);
or U10493 (N_10493,N_10200,N_10224);
xnor U10494 (N_10494,N_10171,N_10053);
nand U10495 (N_10495,N_10130,N_10042);
and U10496 (N_10496,N_10197,N_10370);
nand U10497 (N_10497,N_10164,N_10319);
and U10498 (N_10498,N_10141,N_10007);
xor U10499 (N_10499,N_10157,N_10047);
nor U10500 (N_10500,N_10176,N_10143);
and U10501 (N_10501,N_10220,N_10379);
or U10502 (N_10502,N_10107,N_10244);
xor U10503 (N_10503,N_10211,N_10065);
and U10504 (N_10504,N_10300,N_10251);
nor U10505 (N_10505,N_10250,N_10258);
nor U10506 (N_10506,N_10340,N_10351);
or U10507 (N_10507,N_10288,N_10104);
nand U10508 (N_10508,N_10095,N_10390);
or U10509 (N_10509,N_10312,N_10227);
xnor U10510 (N_10510,N_10252,N_10142);
or U10511 (N_10511,N_10226,N_10094);
and U10512 (N_10512,N_10274,N_10311);
and U10513 (N_10513,N_10123,N_10008);
nor U10514 (N_10514,N_10105,N_10317);
nand U10515 (N_10515,N_10187,N_10038);
and U10516 (N_10516,N_10303,N_10231);
nand U10517 (N_10517,N_10361,N_10324);
nand U10518 (N_10518,N_10151,N_10060);
xor U10519 (N_10519,N_10114,N_10132);
or U10520 (N_10520,N_10389,N_10089);
or U10521 (N_10521,N_10349,N_10006);
xnor U10522 (N_10522,N_10148,N_10149);
nand U10523 (N_10523,N_10158,N_10015);
nor U10524 (N_10524,N_10377,N_10259);
nor U10525 (N_10525,N_10019,N_10353);
nor U10526 (N_10526,N_10001,N_10212);
xnor U10527 (N_10527,N_10181,N_10291);
nand U10528 (N_10528,N_10398,N_10278);
and U10529 (N_10529,N_10005,N_10153);
or U10530 (N_10530,N_10055,N_10144);
or U10531 (N_10531,N_10030,N_10041);
nand U10532 (N_10532,N_10185,N_10201);
or U10533 (N_10533,N_10382,N_10193);
nor U10534 (N_10534,N_10085,N_10017);
or U10535 (N_10535,N_10146,N_10296);
or U10536 (N_10536,N_10239,N_10048);
nor U10537 (N_10537,N_10273,N_10191);
nand U10538 (N_10538,N_10339,N_10173);
and U10539 (N_10539,N_10257,N_10097);
and U10540 (N_10540,N_10119,N_10121);
xnor U10541 (N_10541,N_10345,N_10207);
or U10542 (N_10542,N_10083,N_10356);
xor U10543 (N_10543,N_10287,N_10045);
xor U10544 (N_10544,N_10253,N_10277);
nor U10545 (N_10545,N_10155,N_10013);
nor U10546 (N_10546,N_10314,N_10374);
and U10547 (N_10547,N_10391,N_10056);
xor U10548 (N_10548,N_10022,N_10106);
and U10549 (N_10549,N_10170,N_10063);
and U10550 (N_10550,N_10074,N_10325);
or U10551 (N_10551,N_10066,N_10189);
nor U10552 (N_10552,N_10306,N_10168);
nand U10553 (N_10553,N_10115,N_10118);
xor U10554 (N_10554,N_10326,N_10221);
or U10555 (N_10555,N_10011,N_10331);
nor U10556 (N_10556,N_10139,N_10393);
nor U10557 (N_10557,N_10073,N_10175);
nand U10558 (N_10558,N_10333,N_10111);
nand U10559 (N_10559,N_10233,N_10302);
xnor U10560 (N_10560,N_10254,N_10219);
nor U10561 (N_10561,N_10145,N_10204);
nor U10562 (N_10562,N_10180,N_10156);
and U10563 (N_10563,N_10289,N_10210);
and U10564 (N_10564,N_10343,N_10195);
and U10565 (N_10565,N_10196,N_10334);
xnor U10566 (N_10566,N_10294,N_10110);
nand U10567 (N_10567,N_10215,N_10131);
or U10568 (N_10568,N_10101,N_10327);
and U10569 (N_10569,N_10360,N_10307);
nor U10570 (N_10570,N_10099,N_10071);
nor U10571 (N_10571,N_10276,N_10167);
and U10572 (N_10572,N_10238,N_10338);
or U10573 (N_10573,N_10124,N_10138);
nor U10574 (N_10574,N_10263,N_10369);
and U10575 (N_10575,N_10376,N_10027);
nand U10576 (N_10576,N_10395,N_10392);
nor U10577 (N_10577,N_10373,N_10129);
nor U10578 (N_10578,N_10039,N_10247);
or U10579 (N_10579,N_10268,N_10137);
and U10580 (N_10580,N_10172,N_10159);
xor U10581 (N_10581,N_10043,N_10117);
nand U10582 (N_10582,N_10270,N_10225);
nor U10583 (N_10583,N_10301,N_10077);
or U10584 (N_10584,N_10140,N_10177);
nor U10585 (N_10585,N_10316,N_10357);
nand U10586 (N_10586,N_10235,N_10186);
or U10587 (N_10587,N_10260,N_10152);
xor U10588 (N_10588,N_10261,N_10091);
nand U10589 (N_10589,N_10098,N_10092);
nor U10590 (N_10590,N_10059,N_10004);
xor U10591 (N_10591,N_10299,N_10372);
nor U10592 (N_10592,N_10214,N_10313);
and U10593 (N_10593,N_10308,N_10109);
or U10594 (N_10594,N_10275,N_10206);
nor U10595 (N_10595,N_10298,N_10344);
nand U10596 (N_10596,N_10002,N_10023);
or U10597 (N_10597,N_10012,N_10341);
nand U10598 (N_10598,N_10363,N_10029);
xnor U10599 (N_10599,N_10286,N_10049);
nor U10600 (N_10600,N_10357,N_10394);
xnor U10601 (N_10601,N_10229,N_10074);
xor U10602 (N_10602,N_10292,N_10327);
xor U10603 (N_10603,N_10008,N_10137);
xnor U10604 (N_10604,N_10195,N_10140);
or U10605 (N_10605,N_10384,N_10116);
or U10606 (N_10606,N_10146,N_10241);
xnor U10607 (N_10607,N_10358,N_10345);
or U10608 (N_10608,N_10051,N_10387);
nand U10609 (N_10609,N_10250,N_10081);
nand U10610 (N_10610,N_10249,N_10309);
nor U10611 (N_10611,N_10054,N_10110);
nor U10612 (N_10612,N_10101,N_10347);
xor U10613 (N_10613,N_10054,N_10047);
xor U10614 (N_10614,N_10168,N_10153);
nand U10615 (N_10615,N_10060,N_10180);
nor U10616 (N_10616,N_10355,N_10243);
and U10617 (N_10617,N_10080,N_10148);
nor U10618 (N_10618,N_10107,N_10077);
xor U10619 (N_10619,N_10003,N_10289);
nand U10620 (N_10620,N_10277,N_10039);
and U10621 (N_10621,N_10166,N_10338);
xor U10622 (N_10622,N_10346,N_10137);
nand U10623 (N_10623,N_10039,N_10368);
and U10624 (N_10624,N_10252,N_10175);
or U10625 (N_10625,N_10192,N_10366);
or U10626 (N_10626,N_10153,N_10054);
nand U10627 (N_10627,N_10013,N_10141);
nand U10628 (N_10628,N_10353,N_10257);
xor U10629 (N_10629,N_10173,N_10159);
or U10630 (N_10630,N_10125,N_10051);
nand U10631 (N_10631,N_10223,N_10188);
nor U10632 (N_10632,N_10251,N_10157);
xnor U10633 (N_10633,N_10117,N_10061);
nor U10634 (N_10634,N_10312,N_10298);
nor U10635 (N_10635,N_10142,N_10300);
and U10636 (N_10636,N_10172,N_10239);
xor U10637 (N_10637,N_10250,N_10027);
xnor U10638 (N_10638,N_10068,N_10080);
xor U10639 (N_10639,N_10182,N_10372);
or U10640 (N_10640,N_10158,N_10336);
xor U10641 (N_10641,N_10228,N_10383);
and U10642 (N_10642,N_10133,N_10381);
and U10643 (N_10643,N_10326,N_10299);
nand U10644 (N_10644,N_10186,N_10159);
or U10645 (N_10645,N_10076,N_10224);
or U10646 (N_10646,N_10096,N_10388);
and U10647 (N_10647,N_10203,N_10110);
nor U10648 (N_10648,N_10096,N_10276);
and U10649 (N_10649,N_10162,N_10035);
xnor U10650 (N_10650,N_10002,N_10234);
or U10651 (N_10651,N_10236,N_10391);
or U10652 (N_10652,N_10113,N_10318);
nor U10653 (N_10653,N_10092,N_10248);
or U10654 (N_10654,N_10037,N_10393);
nor U10655 (N_10655,N_10244,N_10366);
nand U10656 (N_10656,N_10099,N_10335);
or U10657 (N_10657,N_10033,N_10038);
nor U10658 (N_10658,N_10262,N_10170);
and U10659 (N_10659,N_10120,N_10156);
nand U10660 (N_10660,N_10071,N_10166);
nand U10661 (N_10661,N_10014,N_10205);
or U10662 (N_10662,N_10073,N_10118);
and U10663 (N_10663,N_10330,N_10347);
nor U10664 (N_10664,N_10389,N_10150);
xnor U10665 (N_10665,N_10082,N_10294);
xor U10666 (N_10666,N_10226,N_10016);
nand U10667 (N_10667,N_10054,N_10007);
and U10668 (N_10668,N_10134,N_10037);
nor U10669 (N_10669,N_10020,N_10322);
and U10670 (N_10670,N_10287,N_10254);
and U10671 (N_10671,N_10207,N_10295);
nand U10672 (N_10672,N_10389,N_10119);
nand U10673 (N_10673,N_10245,N_10276);
xnor U10674 (N_10674,N_10105,N_10389);
xor U10675 (N_10675,N_10028,N_10013);
nor U10676 (N_10676,N_10339,N_10069);
xnor U10677 (N_10677,N_10212,N_10264);
or U10678 (N_10678,N_10285,N_10175);
or U10679 (N_10679,N_10190,N_10348);
nand U10680 (N_10680,N_10267,N_10059);
nand U10681 (N_10681,N_10071,N_10186);
nor U10682 (N_10682,N_10055,N_10291);
nor U10683 (N_10683,N_10138,N_10154);
and U10684 (N_10684,N_10024,N_10298);
or U10685 (N_10685,N_10173,N_10251);
xor U10686 (N_10686,N_10318,N_10256);
nor U10687 (N_10687,N_10220,N_10076);
and U10688 (N_10688,N_10390,N_10347);
nor U10689 (N_10689,N_10246,N_10166);
or U10690 (N_10690,N_10273,N_10288);
xnor U10691 (N_10691,N_10007,N_10000);
xnor U10692 (N_10692,N_10002,N_10190);
nand U10693 (N_10693,N_10226,N_10388);
and U10694 (N_10694,N_10190,N_10295);
nor U10695 (N_10695,N_10189,N_10138);
nor U10696 (N_10696,N_10240,N_10229);
xor U10697 (N_10697,N_10111,N_10211);
and U10698 (N_10698,N_10290,N_10101);
nor U10699 (N_10699,N_10158,N_10137);
nor U10700 (N_10700,N_10007,N_10061);
xnor U10701 (N_10701,N_10084,N_10231);
and U10702 (N_10702,N_10335,N_10118);
xor U10703 (N_10703,N_10021,N_10378);
xnor U10704 (N_10704,N_10391,N_10135);
nor U10705 (N_10705,N_10135,N_10388);
and U10706 (N_10706,N_10219,N_10107);
xnor U10707 (N_10707,N_10151,N_10067);
xor U10708 (N_10708,N_10180,N_10389);
nand U10709 (N_10709,N_10338,N_10210);
nor U10710 (N_10710,N_10029,N_10156);
and U10711 (N_10711,N_10311,N_10227);
or U10712 (N_10712,N_10053,N_10147);
and U10713 (N_10713,N_10044,N_10279);
or U10714 (N_10714,N_10303,N_10234);
or U10715 (N_10715,N_10313,N_10087);
or U10716 (N_10716,N_10391,N_10251);
nand U10717 (N_10717,N_10244,N_10352);
and U10718 (N_10718,N_10019,N_10048);
xor U10719 (N_10719,N_10077,N_10320);
and U10720 (N_10720,N_10167,N_10064);
and U10721 (N_10721,N_10302,N_10207);
xor U10722 (N_10722,N_10214,N_10018);
and U10723 (N_10723,N_10074,N_10047);
or U10724 (N_10724,N_10074,N_10298);
nor U10725 (N_10725,N_10219,N_10215);
nor U10726 (N_10726,N_10166,N_10184);
nor U10727 (N_10727,N_10039,N_10376);
and U10728 (N_10728,N_10019,N_10010);
xor U10729 (N_10729,N_10379,N_10030);
nand U10730 (N_10730,N_10288,N_10317);
and U10731 (N_10731,N_10076,N_10157);
xnor U10732 (N_10732,N_10165,N_10100);
or U10733 (N_10733,N_10323,N_10130);
nor U10734 (N_10734,N_10068,N_10107);
and U10735 (N_10735,N_10116,N_10392);
and U10736 (N_10736,N_10057,N_10152);
nor U10737 (N_10737,N_10113,N_10374);
nor U10738 (N_10738,N_10333,N_10227);
nor U10739 (N_10739,N_10149,N_10268);
nor U10740 (N_10740,N_10211,N_10069);
nand U10741 (N_10741,N_10217,N_10243);
and U10742 (N_10742,N_10382,N_10223);
or U10743 (N_10743,N_10020,N_10194);
or U10744 (N_10744,N_10354,N_10225);
nor U10745 (N_10745,N_10127,N_10261);
nor U10746 (N_10746,N_10125,N_10363);
nor U10747 (N_10747,N_10176,N_10133);
xnor U10748 (N_10748,N_10001,N_10346);
or U10749 (N_10749,N_10086,N_10063);
nand U10750 (N_10750,N_10076,N_10059);
or U10751 (N_10751,N_10145,N_10002);
nand U10752 (N_10752,N_10229,N_10081);
nand U10753 (N_10753,N_10028,N_10242);
and U10754 (N_10754,N_10222,N_10226);
xor U10755 (N_10755,N_10119,N_10269);
nand U10756 (N_10756,N_10339,N_10044);
and U10757 (N_10757,N_10020,N_10132);
xnor U10758 (N_10758,N_10235,N_10381);
or U10759 (N_10759,N_10017,N_10027);
or U10760 (N_10760,N_10322,N_10398);
nor U10761 (N_10761,N_10365,N_10225);
and U10762 (N_10762,N_10345,N_10070);
nor U10763 (N_10763,N_10396,N_10047);
nor U10764 (N_10764,N_10015,N_10026);
nand U10765 (N_10765,N_10173,N_10385);
or U10766 (N_10766,N_10240,N_10123);
xnor U10767 (N_10767,N_10059,N_10175);
nand U10768 (N_10768,N_10045,N_10047);
or U10769 (N_10769,N_10023,N_10339);
or U10770 (N_10770,N_10126,N_10064);
and U10771 (N_10771,N_10076,N_10249);
nor U10772 (N_10772,N_10152,N_10282);
or U10773 (N_10773,N_10258,N_10126);
nand U10774 (N_10774,N_10273,N_10393);
and U10775 (N_10775,N_10038,N_10073);
and U10776 (N_10776,N_10160,N_10147);
and U10777 (N_10777,N_10286,N_10269);
and U10778 (N_10778,N_10292,N_10346);
or U10779 (N_10779,N_10142,N_10085);
nor U10780 (N_10780,N_10126,N_10375);
xnor U10781 (N_10781,N_10346,N_10149);
or U10782 (N_10782,N_10238,N_10178);
nand U10783 (N_10783,N_10149,N_10270);
xor U10784 (N_10784,N_10202,N_10059);
or U10785 (N_10785,N_10243,N_10333);
and U10786 (N_10786,N_10286,N_10356);
or U10787 (N_10787,N_10374,N_10129);
nor U10788 (N_10788,N_10128,N_10037);
and U10789 (N_10789,N_10381,N_10270);
or U10790 (N_10790,N_10372,N_10373);
nor U10791 (N_10791,N_10263,N_10141);
nand U10792 (N_10792,N_10388,N_10272);
nor U10793 (N_10793,N_10112,N_10397);
xor U10794 (N_10794,N_10203,N_10318);
nand U10795 (N_10795,N_10100,N_10060);
and U10796 (N_10796,N_10381,N_10105);
nand U10797 (N_10797,N_10198,N_10277);
and U10798 (N_10798,N_10027,N_10117);
nor U10799 (N_10799,N_10233,N_10243);
or U10800 (N_10800,N_10432,N_10546);
xnor U10801 (N_10801,N_10655,N_10714);
nor U10802 (N_10802,N_10532,N_10765);
or U10803 (N_10803,N_10507,N_10550);
nor U10804 (N_10804,N_10686,N_10680);
and U10805 (N_10805,N_10509,N_10695);
or U10806 (N_10806,N_10707,N_10616);
and U10807 (N_10807,N_10403,N_10434);
xnor U10808 (N_10808,N_10768,N_10510);
nand U10809 (N_10809,N_10548,N_10437);
and U10810 (N_10810,N_10682,N_10769);
nand U10811 (N_10811,N_10776,N_10461);
or U10812 (N_10812,N_10749,N_10486);
and U10813 (N_10813,N_10475,N_10780);
and U10814 (N_10814,N_10577,N_10662);
nor U10815 (N_10815,N_10628,N_10429);
nand U10816 (N_10816,N_10585,N_10715);
nand U10817 (N_10817,N_10406,N_10445);
nor U10818 (N_10818,N_10524,N_10479);
or U10819 (N_10819,N_10702,N_10743);
nand U10820 (N_10820,N_10565,N_10551);
nor U10821 (N_10821,N_10725,N_10783);
or U10822 (N_10822,N_10692,N_10549);
and U10823 (N_10823,N_10449,N_10764);
nor U10824 (N_10824,N_10665,N_10763);
nand U10825 (N_10825,N_10790,N_10558);
or U10826 (N_10826,N_10610,N_10463);
nand U10827 (N_10827,N_10469,N_10466);
xnor U10828 (N_10828,N_10418,N_10739);
nand U10829 (N_10829,N_10428,N_10408);
xnor U10830 (N_10830,N_10552,N_10646);
or U10831 (N_10831,N_10709,N_10414);
xor U10832 (N_10832,N_10774,N_10799);
nor U10833 (N_10833,N_10599,N_10643);
xor U10834 (N_10834,N_10751,N_10529);
or U10835 (N_10835,N_10520,N_10781);
nor U10836 (N_10836,N_10736,N_10566);
nand U10837 (N_10837,N_10436,N_10630);
nor U10838 (N_10838,N_10402,N_10731);
nand U10839 (N_10839,N_10416,N_10409);
and U10840 (N_10840,N_10775,N_10490);
nand U10841 (N_10841,N_10626,N_10487);
xor U10842 (N_10842,N_10459,N_10443);
xor U10843 (N_10843,N_10600,N_10735);
and U10844 (N_10844,N_10627,N_10573);
or U10845 (N_10845,N_10439,N_10491);
nor U10846 (N_10846,N_10644,N_10420);
or U10847 (N_10847,N_10571,N_10531);
xor U10848 (N_10848,N_10767,N_10415);
nand U10849 (N_10849,N_10779,N_10794);
nor U10850 (N_10850,N_10563,N_10688);
xnor U10851 (N_10851,N_10467,N_10586);
nand U10852 (N_10852,N_10498,N_10511);
nand U10853 (N_10853,N_10504,N_10535);
or U10854 (N_10854,N_10710,N_10441);
and U10855 (N_10855,N_10724,N_10588);
xnor U10856 (N_10856,N_10587,N_10796);
and U10857 (N_10857,N_10537,N_10401);
nand U10858 (N_10858,N_10668,N_10419);
and U10859 (N_10859,N_10632,N_10508);
nor U10860 (N_10860,N_10618,N_10698);
nand U10861 (N_10861,N_10620,N_10578);
nor U10862 (N_10862,N_10638,N_10525);
or U10863 (N_10863,N_10417,N_10575);
or U10864 (N_10864,N_10499,N_10497);
nor U10865 (N_10865,N_10758,N_10798);
nand U10866 (N_10866,N_10601,N_10517);
nor U10867 (N_10867,N_10773,N_10460);
xnor U10868 (N_10868,N_10755,N_10592);
and U10869 (N_10869,N_10683,N_10591);
and U10870 (N_10870,N_10624,N_10659);
and U10871 (N_10871,N_10666,N_10580);
xnor U10872 (N_10872,N_10635,N_10621);
nand U10873 (N_10873,N_10738,N_10533);
or U10874 (N_10874,N_10421,N_10720);
or U10875 (N_10875,N_10742,N_10413);
nand U10876 (N_10876,N_10450,N_10653);
nand U10877 (N_10877,N_10583,N_10716);
and U10878 (N_10878,N_10703,N_10663);
xor U10879 (N_10879,N_10718,N_10759);
and U10880 (N_10880,N_10660,N_10641);
or U10881 (N_10881,N_10501,N_10762);
nand U10882 (N_10882,N_10785,N_10699);
xor U10883 (N_10883,N_10502,N_10664);
or U10884 (N_10884,N_10771,N_10602);
and U10885 (N_10885,N_10748,N_10730);
xor U10886 (N_10886,N_10723,N_10564);
and U10887 (N_10887,N_10608,N_10582);
xnor U10888 (N_10888,N_10435,N_10741);
nor U10889 (N_10889,N_10757,N_10713);
or U10890 (N_10890,N_10470,N_10426);
and U10891 (N_10891,N_10649,N_10687);
nor U10892 (N_10892,N_10677,N_10539);
nand U10893 (N_10893,N_10651,N_10792);
nand U10894 (N_10894,N_10481,N_10473);
or U10895 (N_10895,N_10747,N_10642);
nand U10896 (N_10896,N_10574,N_10777);
and U10897 (N_10897,N_10672,N_10744);
xnor U10898 (N_10898,N_10711,N_10633);
xor U10899 (N_10899,N_10440,N_10772);
xnor U10900 (N_10900,N_10614,N_10400);
nor U10901 (N_10901,N_10536,N_10685);
xnor U10902 (N_10902,N_10562,N_10619);
nand U10903 (N_10903,N_10729,N_10447);
nand U10904 (N_10904,N_10732,N_10615);
nand U10905 (N_10905,N_10705,N_10407);
or U10906 (N_10906,N_10760,N_10594);
nor U10907 (N_10907,N_10750,N_10468);
or U10908 (N_10908,N_10639,N_10595);
xor U10909 (N_10909,N_10589,N_10488);
nand U10910 (N_10910,N_10675,N_10493);
or U10911 (N_10911,N_10778,N_10523);
or U10912 (N_10912,N_10625,N_10700);
xnor U10913 (N_10913,N_10694,N_10598);
nand U10914 (N_10914,N_10512,N_10706);
or U10915 (N_10915,N_10726,N_10431);
nand U10916 (N_10916,N_10503,N_10788);
or U10917 (N_10917,N_10697,N_10527);
and U10918 (N_10918,N_10622,N_10456);
xnor U10919 (N_10919,N_10753,N_10451);
and U10920 (N_10920,N_10422,N_10679);
xor U10921 (N_10921,N_10654,N_10495);
nor U10922 (N_10922,N_10534,N_10477);
xor U10923 (N_10923,N_10482,N_10541);
and U10924 (N_10924,N_10737,N_10793);
or U10925 (N_10925,N_10430,N_10690);
or U10926 (N_10926,N_10542,N_10500);
or U10927 (N_10927,N_10433,N_10656);
nand U10928 (N_10928,N_10717,N_10727);
or U10929 (N_10929,N_10648,N_10719);
and U10930 (N_10930,N_10576,N_10458);
nor U10931 (N_10931,N_10448,N_10636);
and U10932 (N_10932,N_10721,N_10661);
xnor U10933 (N_10933,N_10645,N_10561);
nand U10934 (N_10934,N_10609,N_10530);
or U10935 (N_10935,N_10631,N_10789);
nand U10936 (N_10936,N_10667,N_10637);
nor U10937 (N_10937,N_10514,N_10590);
and U10938 (N_10938,N_10634,N_10733);
xor U10939 (N_10939,N_10681,N_10745);
nor U10940 (N_10940,N_10712,N_10693);
xor U10941 (N_10941,N_10555,N_10569);
xnor U10942 (N_10942,N_10612,N_10770);
and U10943 (N_10943,N_10607,N_10684);
nand U10944 (N_10944,N_10480,N_10472);
or U10945 (N_10945,N_10557,N_10674);
or U10946 (N_10946,N_10673,N_10584);
xnor U10947 (N_10947,N_10545,N_10476);
or U10948 (N_10948,N_10411,N_10567);
nand U10949 (N_10949,N_10784,N_10526);
nand U10950 (N_10950,N_10521,N_10404);
nor U10951 (N_10951,N_10427,N_10658);
xor U10952 (N_10952,N_10579,N_10442);
nor U10953 (N_10953,N_10424,N_10671);
nand U10954 (N_10954,N_10797,N_10761);
xnor U10955 (N_10955,N_10701,N_10756);
nand U10956 (N_10956,N_10528,N_10540);
or U10957 (N_10957,N_10494,N_10740);
nand U10958 (N_10958,N_10652,N_10556);
or U10959 (N_10959,N_10474,N_10568);
xor U10960 (N_10960,N_10596,N_10543);
nand U10961 (N_10961,N_10734,N_10787);
or U10962 (N_10962,N_10611,N_10453);
nand U10963 (N_10963,N_10412,N_10465);
nand U10964 (N_10964,N_10471,N_10650);
nor U10965 (N_10965,N_10462,N_10613);
or U10966 (N_10966,N_10452,N_10559);
or U10967 (N_10967,N_10505,N_10519);
nand U10968 (N_10968,N_10678,N_10605);
nor U10969 (N_10969,N_10405,N_10766);
or U10970 (N_10970,N_10464,N_10676);
nor U10971 (N_10971,N_10593,N_10786);
and U10972 (N_10972,N_10506,N_10604);
nand U10973 (N_10973,N_10444,N_10489);
nor U10974 (N_10974,N_10544,N_10513);
nor U10975 (N_10975,N_10425,N_10455);
or U10976 (N_10976,N_10554,N_10617);
xnor U10977 (N_10977,N_10485,N_10722);
nor U10978 (N_10978,N_10696,N_10581);
xor U10979 (N_10979,N_10446,N_10478);
nand U10980 (N_10980,N_10657,N_10484);
and U10981 (N_10981,N_10728,N_10518);
nand U10982 (N_10982,N_10522,N_10640);
nand U10983 (N_10983,N_10538,N_10629);
xnor U10984 (N_10984,N_10496,N_10410);
xnor U10985 (N_10985,N_10560,N_10457);
nor U10986 (N_10986,N_10689,N_10572);
xnor U10987 (N_10987,N_10454,N_10603);
nand U10988 (N_10988,N_10669,N_10483);
or U10989 (N_10989,N_10547,N_10746);
nand U10990 (N_10990,N_10795,N_10791);
xnor U10991 (N_10991,N_10623,N_10553);
nand U10992 (N_10992,N_10782,N_10492);
nand U10993 (N_10993,N_10704,N_10516);
and U10994 (N_10994,N_10752,N_10515);
or U10995 (N_10995,N_10754,N_10670);
or U10996 (N_10996,N_10423,N_10691);
xnor U10997 (N_10997,N_10708,N_10606);
xnor U10998 (N_10998,N_10647,N_10570);
nand U10999 (N_10999,N_10438,N_10597);
or U11000 (N_11000,N_10600,N_10782);
or U11001 (N_11001,N_10623,N_10683);
or U11002 (N_11002,N_10407,N_10710);
nor U11003 (N_11003,N_10542,N_10510);
and U11004 (N_11004,N_10634,N_10500);
and U11005 (N_11005,N_10654,N_10582);
nor U11006 (N_11006,N_10580,N_10535);
or U11007 (N_11007,N_10682,N_10529);
or U11008 (N_11008,N_10471,N_10473);
nand U11009 (N_11009,N_10776,N_10777);
and U11010 (N_11010,N_10512,N_10709);
nor U11011 (N_11011,N_10543,N_10518);
nor U11012 (N_11012,N_10580,N_10449);
nor U11013 (N_11013,N_10728,N_10624);
or U11014 (N_11014,N_10708,N_10705);
xnor U11015 (N_11015,N_10700,N_10683);
nand U11016 (N_11016,N_10478,N_10613);
xor U11017 (N_11017,N_10632,N_10552);
xnor U11018 (N_11018,N_10655,N_10780);
and U11019 (N_11019,N_10539,N_10706);
nor U11020 (N_11020,N_10659,N_10603);
nor U11021 (N_11021,N_10622,N_10771);
xor U11022 (N_11022,N_10666,N_10648);
and U11023 (N_11023,N_10401,N_10571);
or U11024 (N_11024,N_10697,N_10410);
and U11025 (N_11025,N_10461,N_10525);
or U11026 (N_11026,N_10678,N_10488);
or U11027 (N_11027,N_10479,N_10689);
or U11028 (N_11028,N_10769,N_10519);
or U11029 (N_11029,N_10487,N_10736);
nor U11030 (N_11030,N_10475,N_10734);
or U11031 (N_11031,N_10501,N_10408);
or U11032 (N_11032,N_10745,N_10546);
and U11033 (N_11033,N_10416,N_10566);
nor U11034 (N_11034,N_10692,N_10402);
and U11035 (N_11035,N_10755,N_10756);
nand U11036 (N_11036,N_10505,N_10406);
nor U11037 (N_11037,N_10715,N_10411);
and U11038 (N_11038,N_10794,N_10511);
nand U11039 (N_11039,N_10716,N_10625);
nand U11040 (N_11040,N_10572,N_10432);
xnor U11041 (N_11041,N_10517,N_10735);
nand U11042 (N_11042,N_10740,N_10688);
and U11043 (N_11043,N_10518,N_10519);
nand U11044 (N_11044,N_10798,N_10649);
nor U11045 (N_11045,N_10788,N_10502);
xor U11046 (N_11046,N_10629,N_10487);
and U11047 (N_11047,N_10444,N_10716);
and U11048 (N_11048,N_10540,N_10711);
nand U11049 (N_11049,N_10547,N_10440);
and U11050 (N_11050,N_10470,N_10446);
xnor U11051 (N_11051,N_10601,N_10674);
and U11052 (N_11052,N_10634,N_10714);
and U11053 (N_11053,N_10404,N_10774);
or U11054 (N_11054,N_10515,N_10775);
nor U11055 (N_11055,N_10732,N_10691);
and U11056 (N_11056,N_10792,N_10527);
and U11057 (N_11057,N_10777,N_10542);
or U11058 (N_11058,N_10710,N_10640);
or U11059 (N_11059,N_10514,N_10456);
nor U11060 (N_11060,N_10682,N_10413);
nor U11061 (N_11061,N_10517,N_10700);
nor U11062 (N_11062,N_10755,N_10723);
and U11063 (N_11063,N_10638,N_10569);
or U11064 (N_11064,N_10756,N_10730);
and U11065 (N_11065,N_10465,N_10573);
or U11066 (N_11066,N_10558,N_10539);
nand U11067 (N_11067,N_10700,N_10706);
xnor U11068 (N_11068,N_10558,N_10497);
nor U11069 (N_11069,N_10526,N_10437);
nor U11070 (N_11070,N_10677,N_10514);
nor U11071 (N_11071,N_10437,N_10639);
xnor U11072 (N_11072,N_10679,N_10555);
and U11073 (N_11073,N_10508,N_10729);
nand U11074 (N_11074,N_10674,N_10661);
nand U11075 (N_11075,N_10754,N_10529);
nor U11076 (N_11076,N_10641,N_10419);
or U11077 (N_11077,N_10414,N_10707);
and U11078 (N_11078,N_10537,N_10405);
nor U11079 (N_11079,N_10591,N_10725);
nand U11080 (N_11080,N_10400,N_10763);
xor U11081 (N_11081,N_10530,N_10543);
or U11082 (N_11082,N_10533,N_10605);
xnor U11083 (N_11083,N_10565,N_10409);
nand U11084 (N_11084,N_10564,N_10567);
or U11085 (N_11085,N_10711,N_10425);
or U11086 (N_11086,N_10738,N_10583);
and U11087 (N_11087,N_10709,N_10738);
or U11088 (N_11088,N_10719,N_10526);
nand U11089 (N_11089,N_10735,N_10611);
nand U11090 (N_11090,N_10560,N_10569);
nor U11091 (N_11091,N_10676,N_10644);
or U11092 (N_11092,N_10577,N_10568);
xor U11093 (N_11093,N_10740,N_10588);
and U11094 (N_11094,N_10721,N_10644);
and U11095 (N_11095,N_10662,N_10686);
and U11096 (N_11096,N_10415,N_10722);
xnor U11097 (N_11097,N_10473,N_10554);
nand U11098 (N_11098,N_10514,N_10756);
and U11099 (N_11099,N_10569,N_10529);
xnor U11100 (N_11100,N_10505,N_10462);
and U11101 (N_11101,N_10610,N_10558);
xor U11102 (N_11102,N_10548,N_10540);
and U11103 (N_11103,N_10585,N_10741);
nor U11104 (N_11104,N_10541,N_10534);
or U11105 (N_11105,N_10734,N_10701);
and U11106 (N_11106,N_10450,N_10691);
or U11107 (N_11107,N_10678,N_10618);
or U11108 (N_11108,N_10403,N_10712);
xnor U11109 (N_11109,N_10540,N_10674);
or U11110 (N_11110,N_10610,N_10742);
or U11111 (N_11111,N_10445,N_10591);
and U11112 (N_11112,N_10688,N_10593);
or U11113 (N_11113,N_10691,N_10506);
xor U11114 (N_11114,N_10523,N_10625);
or U11115 (N_11115,N_10475,N_10456);
or U11116 (N_11116,N_10517,N_10557);
nor U11117 (N_11117,N_10427,N_10440);
nor U11118 (N_11118,N_10550,N_10530);
or U11119 (N_11119,N_10734,N_10710);
nand U11120 (N_11120,N_10635,N_10563);
xor U11121 (N_11121,N_10668,N_10654);
nor U11122 (N_11122,N_10476,N_10540);
nor U11123 (N_11123,N_10608,N_10513);
xor U11124 (N_11124,N_10607,N_10770);
nor U11125 (N_11125,N_10572,N_10404);
xor U11126 (N_11126,N_10434,N_10479);
xor U11127 (N_11127,N_10694,N_10466);
or U11128 (N_11128,N_10627,N_10424);
or U11129 (N_11129,N_10623,N_10724);
or U11130 (N_11130,N_10676,N_10536);
nor U11131 (N_11131,N_10401,N_10666);
nand U11132 (N_11132,N_10795,N_10751);
xor U11133 (N_11133,N_10728,N_10683);
and U11134 (N_11134,N_10473,N_10655);
xor U11135 (N_11135,N_10544,N_10460);
nor U11136 (N_11136,N_10735,N_10463);
nor U11137 (N_11137,N_10653,N_10414);
xor U11138 (N_11138,N_10404,N_10742);
nand U11139 (N_11139,N_10525,N_10604);
and U11140 (N_11140,N_10655,N_10777);
and U11141 (N_11141,N_10765,N_10769);
or U11142 (N_11142,N_10574,N_10784);
nor U11143 (N_11143,N_10738,N_10726);
or U11144 (N_11144,N_10711,N_10770);
nor U11145 (N_11145,N_10616,N_10770);
or U11146 (N_11146,N_10556,N_10502);
nand U11147 (N_11147,N_10766,N_10782);
nand U11148 (N_11148,N_10689,N_10427);
and U11149 (N_11149,N_10679,N_10606);
and U11150 (N_11150,N_10469,N_10738);
nand U11151 (N_11151,N_10591,N_10692);
nor U11152 (N_11152,N_10610,N_10691);
and U11153 (N_11153,N_10673,N_10533);
or U11154 (N_11154,N_10590,N_10739);
or U11155 (N_11155,N_10549,N_10783);
nand U11156 (N_11156,N_10634,N_10771);
or U11157 (N_11157,N_10417,N_10783);
or U11158 (N_11158,N_10697,N_10493);
nand U11159 (N_11159,N_10577,N_10770);
or U11160 (N_11160,N_10437,N_10773);
xnor U11161 (N_11161,N_10452,N_10501);
or U11162 (N_11162,N_10405,N_10779);
xnor U11163 (N_11163,N_10728,N_10798);
nand U11164 (N_11164,N_10538,N_10698);
or U11165 (N_11165,N_10581,N_10761);
or U11166 (N_11166,N_10770,N_10663);
nand U11167 (N_11167,N_10480,N_10483);
and U11168 (N_11168,N_10426,N_10659);
and U11169 (N_11169,N_10530,N_10754);
xnor U11170 (N_11170,N_10475,N_10718);
xor U11171 (N_11171,N_10461,N_10550);
xor U11172 (N_11172,N_10780,N_10726);
nand U11173 (N_11173,N_10444,N_10771);
xor U11174 (N_11174,N_10635,N_10795);
or U11175 (N_11175,N_10464,N_10501);
nand U11176 (N_11176,N_10671,N_10561);
and U11177 (N_11177,N_10786,N_10476);
nand U11178 (N_11178,N_10627,N_10773);
and U11179 (N_11179,N_10544,N_10764);
or U11180 (N_11180,N_10670,N_10588);
xnor U11181 (N_11181,N_10755,N_10598);
or U11182 (N_11182,N_10566,N_10556);
nor U11183 (N_11183,N_10546,N_10592);
xnor U11184 (N_11184,N_10577,N_10485);
nand U11185 (N_11185,N_10406,N_10504);
nand U11186 (N_11186,N_10729,N_10528);
nand U11187 (N_11187,N_10542,N_10560);
and U11188 (N_11188,N_10491,N_10733);
xnor U11189 (N_11189,N_10593,N_10625);
or U11190 (N_11190,N_10491,N_10598);
nor U11191 (N_11191,N_10445,N_10754);
and U11192 (N_11192,N_10552,N_10713);
and U11193 (N_11193,N_10696,N_10599);
nor U11194 (N_11194,N_10617,N_10433);
nor U11195 (N_11195,N_10547,N_10764);
nand U11196 (N_11196,N_10489,N_10539);
or U11197 (N_11197,N_10630,N_10560);
nand U11198 (N_11198,N_10482,N_10444);
xnor U11199 (N_11199,N_10633,N_10571);
and U11200 (N_11200,N_10986,N_10991);
nand U11201 (N_11201,N_11048,N_11194);
or U11202 (N_11202,N_10908,N_11055);
and U11203 (N_11203,N_10947,N_11119);
nor U11204 (N_11204,N_10969,N_11143);
nor U11205 (N_11205,N_10904,N_10811);
or U11206 (N_11206,N_11156,N_11164);
and U11207 (N_11207,N_10882,N_11124);
nor U11208 (N_11208,N_10897,N_10815);
or U11209 (N_11209,N_10981,N_10930);
or U11210 (N_11210,N_11199,N_10984);
nand U11211 (N_11211,N_10824,N_11182);
nand U11212 (N_11212,N_10855,N_10940);
nand U11213 (N_11213,N_10982,N_10818);
and U11214 (N_11214,N_10819,N_11073);
nand U11215 (N_11215,N_10888,N_11008);
xnor U11216 (N_11216,N_11168,N_10836);
nor U11217 (N_11217,N_11062,N_10929);
and U11218 (N_11218,N_10808,N_10825);
xnor U11219 (N_11219,N_11079,N_10881);
nor U11220 (N_11220,N_11170,N_10883);
or U11221 (N_11221,N_11053,N_11031);
nor U11222 (N_11222,N_11067,N_10804);
xnor U11223 (N_11223,N_10886,N_10922);
and U11224 (N_11224,N_10920,N_11126);
nor U11225 (N_11225,N_11049,N_10857);
or U11226 (N_11226,N_11037,N_10895);
nand U11227 (N_11227,N_11021,N_11063);
nor U11228 (N_11228,N_10803,N_11129);
nand U11229 (N_11229,N_10887,N_10959);
and U11230 (N_11230,N_10851,N_10975);
nor U11231 (N_11231,N_11198,N_11189);
xnor U11232 (N_11232,N_11030,N_10946);
or U11233 (N_11233,N_10977,N_10864);
nor U11234 (N_11234,N_10802,N_10954);
and U11235 (N_11235,N_11099,N_11057);
nand U11236 (N_11236,N_11191,N_11052);
xor U11237 (N_11237,N_10944,N_10898);
nor U11238 (N_11238,N_11101,N_10834);
nand U11239 (N_11239,N_11065,N_11023);
nor U11240 (N_11240,N_11097,N_10958);
nor U11241 (N_11241,N_10970,N_10837);
xnor U11242 (N_11242,N_10863,N_10997);
nand U11243 (N_11243,N_10848,N_11142);
or U11244 (N_11244,N_10994,N_10880);
xnor U11245 (N_11245,N_10905,N_10936);
and U11246 (N_11246,N_11035,N_10906);
nand U11247 (N_11247,N_11153,N_10916);
and U11248 (N_11248,N_10890,N_11110);
xnor U11249 (N_11249,N_10843,N_10853);
xor U11250 (N_11250,N_11162,N_10974);
xnor U11251 (N_11251,N_11032,N_10980);
or U11252 (N_11252,N_10865,N_11090);
and U11253 (N_11253,N_10813,N_10907);
nor U11254 (N_11254,N_10827,N_11084);
nand U11255 (N_11255,N_11135,N_11093);
nor U11256 (N_11256,N_11076,N_10987);
or U11257 (N_11257,N_11096,N_11165);
xor U11258 (N_11258,N_11196,N_11034);
nor U11259 (N_11259,N_10933,N_11138);
or U11260 (N_11260,N_10938,N_10823);
or U11261 (N_11261,N_11010,N_10932);
nand U11262 (N_11262,N_10927,N_11100);
nand U11263 (N_11263,N_11178,N_11108);
nor U11264 (N_11264,N_11074,N_10893);
or U11265 (N_11265,N_10846,N_11072);
or U11266 (N_11266,N_10874,N_11116);
nor U11267 (N_11267,N_10894,N_11060);
nor U11268 (N_11268,N_10948,N_11029);
xor U11269 (N_11269,N_11145,N_10988);
nand U11270 (N_11270,N_10999,N_11175);
xnor U11271 (N_11271,N_11033,N_11174);
and U11272 (N_11272,N_11131,N_10939);
xor U11273 (N_11273,N_11095,N_10963);
or U11274 (N_11274,N_10915,N_10909);
nand U11275 (N_11275,N_11140,N_10800);
xnor U11276 (N_11276,N_11000,N_11181);
nor U11277 (N_11277,N_10891,N_11085);
and U11278 (N_11278,N_10919,N_10901);
and U11279 (N_11279,N_11128,N_10910);
and U11280 (N_11280,N_11011,N_11184);
xor U11281 (N_11281,N_10877,N_11167);
and U11282 (N_11282,N_11121,N_10951);
nor U11283 (N_11283,N_10868,N_11027);
and U11284 (N_11284,N_11009,N_10928);
xor U11285 (N_11285,N_11115,N_10816);
nand U11286 (N_11286,N_10976,N_11046);
xnor U11287 (N_11287,N_11080,N_11088);
xor U11288 (N_11288,N_10860,N_10810);
xor U11289 (N_11289,N_11012,N_10854);
and U11290 (N_11290,N_11177,N_11120);
nor U11291 (N_11291,N_11082,N_11105);
nor U11292 (N_11292,N_10858,N_10992);
nand U11293 (N_11293,N_11154,N_10964);
nor U11294 (N_11294,N_10990,N_11061);
nor U11295 (N_11295,N_11050,N_10937);
nor U11296 (N_11296,N_11019,N_10934);
nor U11297 (N_11297,N_10978,N_10801);
or U11298 (N_11298,N_10950,N_11045);
nand U11299 (N_11299,N_11089,N_10844);
or U11300 (N_11300,N_10966,N_10838);
xor U11301 (N_11301,N_11109,N_10955);
nand U11302 (N_11302,N_10989,N_10983);
or U11303 (N_11303,N_11051,N_11146);
nand U11304 (N_11304,N_11007,N_11077);
and U11305 (N_11305,N_11058,N_10931);
xor U11306 (N_11306,N_11002,N_11180);
nand U11307 (N_11307,N_11188,N_10971);
nor U11308 (N_11308,N_10847,N_10878);
and U11309 (N_11309,N_10949,N_10841);
xor U11310 (N_11310,N_11043,N_10822);
xnor U11311 (N_11311,N_11147,N_11044);
or U11312 (N_11312,N_10856,N_10842);
or U11313 (N_11313,N_10852,N_11195);
or U11314 (N_11314,N_10965,N_10945);
nor U11315 (N_11315,N_11103,N_10879);
nor U11316 (N_11316,N_10889,N_10960);
and U11317 (N_11317,N_10876,N_10941);
nor U11318 (N_11318,N_11070,N_11091);
nand U11319 (N_11319,N_10961,N_10830);
nand U11320 (N_11320,N_10872,N_10985);
nor U11321 (N_11321,N_11104,N_11183);
nand U11322 (N_11322,N_11106,N_10885);
nor U11323 (N_11323,N_11102,N_10814);
nand U11324 (N_11324,N_10917,N_11150);
nand U11325 (N_11325,N_11132,N_10918);
nand U11326 (N_11326,N_10820,N_10921);
nand U11327 (N_11327,N_11185,N_10925);
xnor U11328 (N_11328,N_11197,N_11173);
and U11329 (N_11329,N_11172,N_10926);
and U11330 (N_11330,N_10866,N_11159);
or U11331 (N_11331,N_11098,N_10845);
nor U11332 (N_11332,N_11014,N_10867);
or U11333 (N_11333,N_11040,N_11148);
or U11334 (N_11334,N_10972,N_11176);
or U11335 (N_11335,N_11190,N_10826);
or U11336 (N_11336,N_11169,N_10979);
xnor U11337 (N_11337,N_11114,N_10862);
or U11338 (N_11338,N_11094,N_11078);
and U11339 (N_11339,N_10903,N_11160);
xor U11340 (N_11340,N_11004,N_11163);
xor U11341 (N_11341,N_11017,N_10833);
or U11342 (N_11342,N_10896,N_11054);
or U11343 (N_11343,N_11001,N_11113);
or U11344 (N_11344,N_10993,N_10806);
nor U11345 (N_11345,N_11028,N_11186);
nor U11346 (N_11346,N_10849,N_11015);
or U11347 (N_11347,N_10821,N_11179);
nor U11348 (N_11348,N_11018,N_10817);
or U11349 (N_11349,N_11161,N_11069);
xor U11350 (N_11350,N_10840,N_10807);
and U11351 (N_11351,N_10943,N_11059);
or U11352 (N_11352,N_10952,N_10924);
or U11353 (N_11353,N_10870,N_10899);
or U11354 (N_11354,N_11149,N_10996);
nor U11355 (N_11355,N_11112,N_11118);
or U11356 (N_11356,N_11130,N_11122);
and U11357 (N_11357,N_10859,N_10832);
xor U11358 (N_11358,N_10902,N_11144);
xnor U11359 (N_11359,N_11064,N_10869);
xor U11360 (N_11360,N_11157,N_11134);
or U11361 (N_11361,N_11056,N_11125);
and U11362 (N_11362,N_11042,N_10911);
and U11363 (N_11363,N_11016,N_10967);
nor U11364 (N_11364,N_11193,N_10884);
nor U11365 (N_11365,N_11107,N_10839);
xor U11366 (N_11366,N_10812,N_10850);
xor U11367 (N_11367,N_11075,N_11155);
or U11368 (N_11368,N_11003,N_10809);
or U11369 (N_11369,N_11083,N_11039);
or U11370 (N_11370,N_10923,N_10831);
nor U11371 (N_11371,N_11166,N_11136);
nor U11372 (N_11372,N_10935,N_11127);
xnor U11373 (N_11373,N_11066,N_11139);
nand U11374 (N_11374,N_11086,N_11036);
and U11375 (N_11375,N_11068,N_11020);
xnor U11376 (N_11376,N_11081,N_11092);
and U11377 (N_11377,N_11187,N_11141);
and U11378 (N_11378,N_11013,N_10953);
xor U11379 (N_11379,N_11151,N_10892);
and U11380 (N_11380,N_10871,N_11171);
xor U11381 (N_11381,N_11038,N_11087);
and U11382 (N_11382,N_11071,N_11152);
and U11383 (N_11383,N_11006,N_11047);
or U11384 (N_11384,N_10962,N_11022);
and U11385 (N_11385,N_11111,N_10942);
and U11386 (N_11386,N_11123,N_10829);
and U11387 (N_11387,N_10914,N_11005);
nand U11388 (N_11388,N_10995,N_10968);
nor U11389 (N_11389,N_10873,N_11026);
or U11390 (N_11390,N_10805,N_11041);
or U11391 (N_11391,N_11137,N_10998);
nor U11392 (N_11392,N_10912,N_10861);
or U11393 (N_11393,N_10973,N_11117);
nor U11394 (N_11394,N_11158,N_10828);
and U11395 (N_11395,N_10900,N_10875);
or U11396 (N_11396,N_10913,N_11192);
xor U11397 (N_11397,N_11025,N_11024);
nor U11398 (N_11398,N_10957,N_10956);
nand U11399 (N_11399,N_10835,N_11133);
xnor U11400 (N_11400,N_11138,N_11120);
or U11401 (N_11401,N_10892,N_10844);
nand U11402 (N_11402,N_11121,N_11171);
xnor U11403 (N_11403,N_10940,N_11157);
or U11404 (N_11404,N_11072,N_11124);
or U11405 (N_11405,N_11151,N_10909);
xnor U11406 (N_11406,N_10836,N_10827);
nor U11407 (N_11407,N_10920,N_10911);
nand U11408 (N_11408,N_11181,N_11052);
nand U11409 (N_11409,N_11157,N_11136);
xor U11410 (N_11410,N_10898,N_11147);
and U11411 (N_11411,N_10920,N_10843);
or U11412 (N_11412,N_10828,N_11159);
xor U11413 (N_11413,N_10835,N_11193);
or U11414 (N_11414,N_11133,N_10967);
nor U11415 (N_11415,N_10938,N_10854);
nor U11416 (N_11416,N_10853,N_11179);
or U11417 (N_11417,N_11044,N_11155);
xnor U11418 (N_11418,N_11019,N_11184);
xor U11419 (N_11419,N_11090,N_10896);
and U11420 (N_11420,N_11140,N_10896);
nor U11421 (N_11421,N_10947,N_11151);
nand U11422 (N_11422,N_10853,N_11021);
or U11423 (N_11423,N_11065,N_11054);
or U11424 (N_11424,N_10881,N_10891);
xnor U11425 (N_11425,N_11046,N_11086);
or U11426 (N_11426,N_10858,N_10987);
nor U11427 (N_11427,N_10842,N_11108);
nor U11428 (N_11428,N_11081,N_10907);
and U11429 (N_11429,N_11133,N_10857);
nor U11430 (N_11430,N_10872,N_11059);
or U11431 (N_11431,N_10917,N_10872);
nor U11432 (N_11432,N_11181,N_11135);
nor U11433 (N_11433,N_11048,N_11151);
xnor U11434 (N_11434,N_11028,N_11049);
nand U11435 (N_11435,N_11182,N_11147);
nor U11436 (N_11436,N_10985,N_11197);
xor U11437 (N_11437,N_11007,N_11198);
nor U11438 (N_11438,N_11074,N_10941);
nand U11439 (N_11439,N_11059,N_10927);
xnor U11440 (N_11440,N_10954,N_11075);
or U11441 (N_11441,N_11101,N_11138);
nor U11442 (N_11442,N_11164,N_11140);
and U11443 (N_11443,N_11198,N_11079);
xnor U11444 (N_11444,N_10978,N_11087);
or U11445 (N_11445,N_11154,N_11132);
and U11446 (N_11446,N_11085,N_11187);
nand U11447 (N_11447,N_10856,N_10911);
nand U11448 (N_11448,N_10855,N_10857);
nor U11449 (N_11449,N_10818,N_11087);
nor U11450 (N_11450,N_11021,N_11191);
or U11451 (N_11451,N_11063,N_11083);
and U11452 (N_11452,N_11074,N_10884);
nor U11453 (N_11453,N_10996,N_11133);
and U11454 (N_11454,N_10915,N_10968);
nand U11455 (N_11455,N_11169,N_11189);
and U11456 (N_11456,N_10869,N_10903);
xor U11457 (N_11457,N_10810,N_10973);
xor U11458 (N_11458,N_11029,N_11186);
and U11459 (N_11459,N_11050,N_11081);
xnor U11460 (N_11460,N_11015,N_11008);
or U11461 (N_11461,N_10894,N_10919);
nand U11462 (N_11462,N_10980,N_10861);
nor U11463 (N_11463,N_11051,N_10925);
or U11464 (N_11464,N_11182,N_11190);
nor U11465 (N_11465,N_10901,N_10881);
nor U11466 (N_11466,N_10959,N_10968);
nor U11467 (N_11467,N_11112,N_11150);
xor U11468 (N_11468,N_11099,N_11167);
or U11469 (N_11469,N_10879,N_10929);
or U11470 (N_11470,N_11086,N_11191);
or U11471 (N_11471,N_11110,N_11196);
nand U11472 (N_11472,N_10944,N_10961);
nor U11473 (N_11473,N_10991,N_10882);
or U11474 (N_11474,N_10943,N_11021);
nand U11475 (N_11475,N_10928,N_11037);
nor U11476 (N_11476,N_11144,N_11007);
xor U11477 (N_11477,N_10919,N_11077);
or U11478 (N_11478,N_11043,N_10935);
or U11479 (N_11479,N_11084,N_11179);
nand U11480 (N_11480,N_11060,N_10953);
xor U11481 (N_11481,N_10851,N_11054);
nor U11482 (N_11482,N_11087,N_11138);
and U11483 (N_11483,N_10958,N_10855);
nand U11484 (N_11484,N_11008,N_11147);
xnor U11485 (N_11485,N_11077,N_11037);
and U11486 (N_11486,N_11175,N_10868);
or U11487 (N_11487,N_10811,N_10943);
and U11488 (N_11488,N_10925,N_10875);
and U11489 (N_11489,N_11165,N_10862);
nor U11490 (N_11490,N_10921,N_11091);
or U11491 (N_11491,N_11198,N_10861);
nand U11492 (N_11492,N_10816,N_10808);
or U11493 (N_11493,N_10877,N_11104);
nand U11494 (N_11494,N_10988,N_10984);
xor U11495 (N_11495,N_11149,N_10974);
or U11496 (N_11496,N_10888,N_11103);
and U11497 (N_11497,N_10861,N_10867);
xor U11498 (N_11498,N_10915,N_10977);
xor U11499 (N_11499,N_11040,N_11182);
nand U11500 (N_11500,N_10828,N_11064);
and U11501 (N_11501,N_10988,N_11128);
xnor U11502 (N_11502,N_10921,N_11186);
xnor U11503 (N_11503,N_10803,N_11047);
xor U11504 (N_11504,N_10943,N_10915);
or U11505 (N_11505,N_10850,N_10878);
nor U11506 (N_11506,N_11155,N_10983);
and U11507 (N_11507,N_10882,N_11196);
xnor U11508 (N_11508,N_10819,N_11111);
nand U11509 (N_11509,N_11178,N_10932);
xnor U11510 (N_11510,N_10868,N_11052);
nor U11511 (N_11511,N_10934,N_11132);
xnor U11512 (N_11512,N_11093,N_11067);
nand U11513 (N_11513,N_10987,N_11167);
xor U11514 (N_11514,N_11176,N_10862);
xor U11515 (N_11515,N_11177,N_11135);
nand U11516 (N_11516,N_11038,N_10996);
or U11517 (N_11517,N_11051,N_11136);
nor U11518 (N_11518,N_11072,N_11008);
nand U11519 (N_11519,N_11116,N_10963);
xnor U11520 (N_11520,N_10819,N_11046);
or U11521 (N_11521,N_10954,N_10952);
and U11522 (N_11522,N_11120,N_11180);
and U11523 (N_11523,N_10913,N_11120);
nor U11524 (N_11524,N_11194,N_11145);
nand U11525 (N_11525,N_11083,N_10835);
nand U11526 (N_11526,N_10974,N_11129);
and U11527 (N_11527,N_11001,N_11132);
nand U11528 (N_11528,N_11067,N_10951);
nand U11529 (N_11529,N_11093,N_10802);
nand U11530 (N_11530,N_10820,N_10937);
and U11531 (N_11531,N_10977,N_11151);
nand U11532 (N_11532,N_11142,N_11145);
xnor U11533 (N_11533,N_10887,N_10802);
or U11534 (N_11534,N_11115,N_10824);
xor U11535 (N_11535,N_10998,N_10941);
nand U11536 (N_11536,N_11067,N_10866);
xnor U11537 (N_11537,N_10888,N_10893);
or U11538 (N_11538,N_11181,N_10854);
and U11539 (N_11539,N_11199,N_11123);
nand U11540 (N_11540,N_11010,N_10975);
nor U11541 (N_11541,N_10900,N_11075);
and U11542 (N_11542,N_11037,N_10891);
nand U11543 (N_11543,N_11096,N_10892);
nand U11544 (N_11544,N_10915,N_10934);
nor U11545 (N_11545,N_11156,N_10889);
xnor U11546 (N_11546,N_11140,N_10883);
and U11547 (N_11547,N_11115,N_10938);
xnor U11548 (N_11548,N_10982,N_11176);
nand U11549 (N_11549,N_11002,N_10922);
nand U11550 (N_11550,N_10884,N_11060);
nor U11551 (N_11551,N_11132,N_10923);
nor U11552 (N_11552,N_11012,N_11075);
nand U11553 (N_11553,N_10870,N_11118);
or U11554 (N_11554,N_11170,N_11127);
xnor U11555 (N_11555,N_10859,N_11060);
nand U11556 (N_11556,N_11110,N_11192);
nand U11557 (N_11557,N_11105,N_11012);
xor U11558 (N_11558,N_10978,N_11121);
nor U11559 (N_11559,N_11090,N_10803);
nor U11560 (N_11560,N_11030,N_11140);
nand U11561 (N_11561,N_11095,N_11136);
xor U11562 (N_11562,N_11175,N_11119);
and U11563 (N_11563,N_11160,N_10830);
nor U11564 (N_11564,N_10962,N_11031);
and U11565 (N_11565,N_10840,N_11197);
nand U11566 (N_11566,N_10981,N_11121);
or U11567 (N_11567,N_10960,N_10827);
and U11568 (N_11568,N_11137,N_11156);
and U11569 (N_11569,N_11107,N_11045);
or U11570 (N_11570,N_11004,N_10941);
and U11571 (N_11571,N_10809,N_10812);
and U11572 (N_11572,N_10913,N_11052);
nand U11573 (N_11573,N_10825,N_11149);
or U11574 (N_11574,N_11071,N_10884);
and U11575 (N_11575,N_11106,N_10904);
nand U11576 (N_11576,N_11136,N_10922);
nor U11577 (N_11577,N_11074,N_10811);
nor U11578 (N_11578,N_10822,N_11133);
xnor U11579 (N_11579,N_11195,N_11007);
or U11580 (N_11580,N_10890,N_11141);
and U11581 (N_11581,N_10851,N_10816);
nand U11582 (N_11582,N_11145,N_11111);
nor U11583 (N_11583,N_10957,N_10823);
nor U11584 (N_11584,N_11134,N_11155);
nand U11585 (N_11585,N_10888,N_10845);
xnor U11586 (N_11586,N_11144,N_10841);
nand U11587 (N_11587,N_11076,N_11013);
nand U11588 (N_11588,N_11180,N_11130);
xor U11589 (N_11589,N_11077,N_10972);
nor U11590 (N_11590,N_11163,N_11152);
or U11591 (N_11591,N_11185,N_11019);
xor U11592 (N_11592,N_11026,N_11163);
nand U11593 (N_11593,N_10809,N_10802);
xor U11594 (N_11594,N_11076,N_11109);
and U11595 (N_11595,N_10809,N_11001);
and U11596 (N_11596,N_10951,N_11175);
nand U11597 (N_11597,N_10998,N_10999);
and U11598 (N_11598,N_10900,N_11167);
or U11599 (N_11599,N_10907,N_11164);
nor U11600 (N_11600,N_11366,N_11288);
and U11601 (N_11601,N_11582,N_11447);
or U11602 (N_11602,N_11528,N_11579);
nand U11603 (N_11603,N_11502,N_11598);
nor U11604 (N_11604,N_11309,N_11355);
and U11605 (N_11605,N_11445,N_11406);
xnor U11606 (N_11606,N_11563,N_11398);
nor U11607 (N_11607,N_11274,N_11360);
nor U11608 (N_11608,N_11488,N_11489);
nor U11609 (N_11609,N_11555,N_11464);
and U11610 (N_11610,N_11408,N_11432);
and U11611 (N_11611,N_11479,N_11420);
and U11612 (N_11612,N_11258,N_11379);
nor U11613 (N_11613,N_11315,N_11374);
nand U11614 (N_11614,N_11252,N_11293);
and U11615 (N_11615,N_11317,N_11525);
nor U11616 (N_11616,N_11536,N_11373);
nand U11617 (N_11617,N_11491,N_11433);
nor U11618 (N_11618,N_11565,N_11456);
and U11619 (N_11619,N_11364,N_11338);
xor U11620 (N_11620,N_11519,N_11537);
xor U11621 (N_11621,N_11508,N_11544);
nand U11622 (N_11622,N_11229,N_11271);
and U11623 (N_11623,N_11291,N_11477);
and U11624 (N_11624,N_11560,N_11367);
nor U11625 (N_11625,N_11214,N_11391);
or U11626 (N_11626,N_11388,N_11351);
xnor U11627 (N_11627,N_11213,N_11302);
xor U11628 (N_11628,N_11549,N_11590);
or U11629 (N_11629,N_11381,N_11311);
nor U11630 (N_11630,N_11266,N_11558);
or U11631 (N_11631,N_11574,N_11468);
nor U11632 (N_11632,N_11368,N_11486);
xor U11633 (N_11633,N_11513,N_11298);
nand U11634 (N_11634,N_11474,N_11324);
or U11635 (N_11635,N_11539,N_11262);
and U11636 (N_11636,N_11542,N_11418);
nor U11637 (N_11637,N_11578,N_11591);
and U11638 (N_11638,N_11310,N_11500);
or U11639 (N_11639,N_11340,N_11399);
nand U11640 (N_11640,N_11201,N_11583);
nand U11641 (N_11641,N_11575,N_11530);
xor U11642 (N_11642,N_11345,N_11236);
nor U11643 (N_11643,N_11208,N_11339);
xnor U11644 (N_11644,N_11596,N_11313);
nand U11645 (N_11645,N_11454,N_11270);
xnor U11646 (N_11646,N_11304,N_11209);
nand U11647 (N_11647,N_11292,N_11365);
and U11648 (N_11648,N_11487,N_11325);
or U11649 (N_11649,N_11511,N_11218);
nand U11650 (N_11650,N_11535,N_11248);
nand U11651 (N_11651,N_11279,N_11257);
or U11652 (N_11652,N_11427,N_11382);
and U11653 (N_11653,N_11561,N_11587);
nand U11654 (N_11654,N_11435,N_11370);
and U11655 (N_11655,N_11282,N_11543);
and U11656 (N_11656,N_11241,N_11392);
nand U11657 (N_11657,N_11532,N_11523);
nand U11658 (N_11658,N_11425,N_11553);
xnor U11659 (N_11659,N_11520,N_11571);
nor U11660 (N_11660,N_11592,N_11232);
or U11661 (N_11661,N_11349,N_11299);
nand U11662 (N_11662,N_11417,N_11450);
nand U11663 (N_11663,N_11243,N_11323);
and U11664 (N_11664,N_11576,N_11550);
xor U11665 (N_11665,N_11333,N_11397);
nand U11666 (N_11666,N_11480,N_11261);
or U11667 (N_11667,N_11372,N_11551);
nand U11668 (N_11668,N_11371,N_11342);
xnor U11669 (N_11669,N_11572,N_11348);
nand U11670 (N_11670,N_11205,N_11586);
xnor U11671 (N_11671,N_11496,N_11581);
xor U11672 (N_11672,N_11303,N_11395);
nor U11673 (N_11673,N_11457,N_11356);
nand U11674 (N_11674,N_11440,N_11529);
or U11675 (N_11675,N_11259,N_11231);
and U11676 (N_11676,N_11444,N_11273);
and U11677 (N_11677,N_11240,N_11285);
nor U11678 (N_11678,N_11396,N_11272);
and U11679 (N_11679,N_11443,N_11305);
xnor U11680 (N_11680,N_11300,N_11376);
nand U11681 (N_11681,N_11416,N_11483);
and U11682 (N_11682,N_11434,N_11386);
and U11683 (N_11683,N_11552,N_11531);
xnor U11684 (N_11684,N_11517,N_11385);
and U11685 (N_11685,N_11541,N_11234);
nor U11686 (N_11686,N_11383,N_11283);
nand U11687 (N_11687,N_11327,N_11225);
xor U11688 (N_11688,N_11343,N_11286);
and U11689 (N_11689,N_11211,N_11393);
xnor U11690 (N_11690,N_11405,N_11465);
nor U11691 (N_11691,N_11331,N_11238);
xnor U11692 (N_11692,N_11458,N_11490);
and U11693 (N_11693,N_11577,N_11202);
nand U11694 (N_11694,N_11461,N_11492);
nor U11695 (N_11695,N_11438,N_11384);
and U11696 (N_11696,N_11481,N_11516);
xnor U11697 (N_11697,N_11413,N_11320);
or U11698 (N_11698,N_11495,N_11589);
xor U11699 (N_11699,N_11219,N_11290);
and U11700 (N_11700,N_11295,N_11599);
nor U11701 (N_11701,N_11221,N_11540);
nor U11702 (N_11702,N_11280,N_11319);
nor U11703 (N_11703,N_11498,N_11350);
xnor U11704 (N_11704,N_11469,N_11436);
nand U11705 (N_11705,N_11570,N_11449);
or U11706 (N_11706,N_11321,N_11501);
xor U11707 (N_11707,N_11462,N_11220);
nor U11708 (N_11708,N_11289,N_11448);
or U11709 (N_11709,N_11245,N_11346);
nor U11710 (N_11710,N_11242,N_11287);
or U11711 (N_11711,N_11318,N_11276);
or U11712 (N_11712,N_11470,N_11564);
nor U11713 (N_11713,N_11494,N_11200);
nor U11714 (N_11714,N_11375,N_11472);
nand U11715 (N_11715,N_11277,N_11475);
and U11716 (N_11716,N_11250,N_11446);
and U11717 (N_11717,N_11352,N_11460);
nand U11718 (N_11718,N_11204,N_11344);
and U11719 (N_11719,N_11584,N_11510);
nor U11720 (N_11720,N_11554,N_11562);
nor U11721 (N_11721,N_11267,N_11216);
or U11722 (N_11722,N_11301,N_11453);
xor U11723 (N_11723,N_11473,N_11235);
nand U11724 (N_11724,N_11329,N_11451);
nor U11725 (N_11725,N_11484,N_11422);
or U11726 (N_11726,N_11297,N_11357);
nand U11727 (N_11727,N_11330,N_11559);
or U11728 (N_11728,N_11233,N_11354);
or U11729 (N_11729,N_11217,N_11478);
and U11730 (N_11730,N_11253,N_11585);
nand U11731 (N_11731,N_11332,N_11249);
xor U11732 (N_11732,N_11380,N_11254);
nor U11733 (N_11733,N_11482,N_11230);
nand U11734 (N_11734,N_11509,N_11215);
or U11735 (N_11735,N_11410,N_11275);
nand U11736 (N_11736,N_11402,N_11506);
xnor U11737 (N_11737,N_11505,N_11244);
nor U11738 (N_11738,N_11308,N_11573);
or U11739 (N_11739,N_11264,N_11538);
nor U11740 (N_11740,N_11207,N_11423);
nand U11741 (N_11741,N_11296,N_11314);
nor U11742 (N_11742,N_11306,N_11463);
and U11743 (N_11743,N_11265,N_11206);
nand U11744 (N_11744,N_11476,N_11222);
nand U11745 (N_11745,N_11493,N_11336);
nor U11746 (N_11746,N_11358,N_11515);
nand U11747 (N_11747,N_11322,N_11326);
and U11748 (N_11748,N_11534,N_11504);
or U11749 (N_11749,N_11518,N_11566);
xor U11750 (N_11750,N_11316,N_11369);
or U11751 (N_11751,N_11588,N_11414);
or U11752 (N_11752,N_11228,N_11394);
and U11753 (N_11753,N_11593,N_11419);
xnor U11754 (N_11754,N_11328,N_11260);
nor U11755 (N_11755,N_11203,N_11455);
and U11756 (N_11756,N_11441,N_11268);
nor U11757 (N_11757,N_11431,N_11485);
xnor U11758 (N_11758,N_11467,N_11421);
nor U11759 (N_11759,N_11557,N_11514);
and U11760 (N_11760,N_11497,N_11212);
nand U11761 (N_11761,N_11246,N_11353);
nand U11762 (N_11762,N_11237,N_11503);
and U11763 (N_11763,N_11341,N_11407);
xnor U11764 (N_11764,N_11442,N_11580);
or U11765 (N_11765,N_11400,N_11334);
nor U11766 (N_11766,N_11512,N_11378);
nor U11767 (N_11767,N_11526,N_11404);
or U11768 (N_11768,N_11430,N_11223);
or U11769 (N_11769,N_11426,N_11361);
xnor U11770 (N_11770,N_11412,N_11227);
nor U11771 (N_11771,N_11210,N_11567);
xnor U11772 (N_11772,N_11337,N_11389);
nor U11773 (N_11773,N_11499,N_11347);
xor U11774 (N_11774,N_11521,N_11439);
and U11775 (N_11775,N_11522,N_11507);
nand U11776 (N_11776,N_11403,N_11556);
nor U11777 (N_11777,N_11401,N_11466);
and U11778 (N_11778,N_11459,N_11411);
xor U11779 (N_11779,N_11545,N_11597);
or U11780 (N_11780,N_11256,N_11224);
nor U11781 (N_11781,N_11278,N_11527);
nor U11782 (N_11782,N_11359,N_11546);
or U11783 (N_11783,N_11595,N_11428);
nand U11784 (N_11784,N_11387,N_11377);
xnor U11785 (N_11785,N_11363,N_11362);
and U11786 (N_11786,N_11548,N_11239);
nor U11787 (N_11787,N_11437,N_11452);
or U11788 (N_11788,N_11284,N_11424);
nand U11789 (N_11789,N_11263,N_11307);
or U11790 (N_11790,N_11226,N_11594);
xor U11791 (N_11791,N_11415,N_11524);
nand U11792 (N_11792,N_11390,N_11533);
or U11793 (N_11793,N_11251,N_11471);
nand U11794 (N_11794,N_11269,N_11568);
nand U11795 (N_11795,N_11281,N_11547);
nand U11796 (N_11796,N_11247,N_11312);
xnor U11797 (N_11797,N_11409,N_11429);
xnor U11798 (N_11798,N_11335,N_11294);
and U11799 (N_11799,N_11569,N_11255);
or U11800 (N_11800,N_11495,N_11278);
or U11801 (N_11801,N_11265,N_11251);
or U11802 (N_11802,N_11581,N_11264);
xor U11803 (N_11803,N_11337,N_11243);
nand U11804 (N_11804,N_11563,N_11327);
nand U11805 (N_11805,N_11450,N_11571);
nor U11806 (N_11806,N_11233,N_11546);
nor U11807 (N_11807,N_11217,N_11364);
or U11808 (N_11808,N_11484,N_11310);
xor U11809 (N_11809,N_11240,N_11309);
and U11810 (N_11810,N_11207,N_11282);
or U11811 (N_11811,N_11456,N_11205);
and U11812 (N_11812,N_11524,N_11430);
nor U11813 (N_11813,N_11344,N_11294);
and U11814 (N_11814,N_11569,N_11261);
nor U11815 (N_11815,N_11233,N_11400);
xnor U11816 (N_11816,N_11212,N_11244);
nand U11817 (N_11817,N_11222,N_11424);
xnor U11818 (N_11818,N_11256,N_11210);
xnor U11819 (N_11819,N_11301,N_11278);
nand U11820 (N_11820,N_11433,N_11287);
or U11821 (N_11821,N_11312,N_11228);
xnor U11822 (N_11822,N_11369,N_11562);
and U11823 (N_11823,N_11461,N_11345);
or U11824 (N_11824,N_11268,N_11569);
or U11825 (N_11825,N_11300,N_11234);
or U11826 (N_11826,N_11323,N_11560);
xor U11827 (N_11827,N_11344,N_11290);
xnor U11828 (N_11828,N_11550,N_11453);
nand U11829 (N_11829,N_11565,N_11462);
xnor U11830 (N_11830,N_11387,N_11228);
and U11831 (N_11831,N_11283,N_11206);
or U11832 (N_11832,N_11300,N_11593);
xor U11833 (N_11833,N_11296,N_11461);
and U11834 (N_11834,N_11216,N_11277);
nand U11835 (N_11835,N_11399,N_11372);
or U11836 (N_11836,N_11432,N_11599);
or U11837 (N_11837,N_11338,N_11211);
and U11838 (N_11838,N_11329,N_11519);
or U11839 (N_11839,N_11268,N_11278);
and U11840 (N_11840,N_11589,N_11466);
or U11841 (N_11841,N_11244,N_11421);
or U11842 (N_11842,N_11551,N_11504);
nor U11843 (N_11843,N_11438,N_11265);
nand U11844 (N_11844,N_11509,N_11500);
nand U11845 (N_11845,N_11221,N_11265);
nor U11846 (N_11846,N_11251,N_11304);
nor U11847 (N_11847,N_11400,N_11227);
xnor U11848 (N_11848,N_11542,N_11513);
nor U11849 (N_11849,N_11338,N_11554);
xnor U11850 (N_11850,N_11587,N_11498);
or U11851 (N_11851,N_11438,N_11519);
xor U11852 (N_11852,N_11467,N_11309);
nand U11853 (N_11853,N_11579,N_11285);
nand U11854 (N_11854,N_11458,N_11497);
xnor U11855 (N_11855,N_11213,N_11554);
xor U11856 (N_11856,N_11512,N_11527);
and U11857 (N_11857,N_11399,N_11524);
or U11858 (N_11858,N_11384,N_11410);
xor U11859 (N_11859,N_11459,N_11516);
and U11860 (N_11860,N_11502,N_11406);
xor U11861 (N_11861,N_11288,N_11279);
nor U11862 (N_11862,N_11507,N_11390);
or U11863 (N_11863,N_11212,N_11565);
xnor U11864 (N_11864,N_11469,N_11349);
xnor U11865 (N_11865,N_11290,N_11376);
and U11866 (N_11866,N_11445,N_11238);
xnor U11867 (N_11867,N_11475,N_11263);
nor U11868 (N_11868,N_11585,N_11383);
nand U11869 (N_11869,N_11555,N_11225);
nand U11870 (N_11870,N_11332,N_11269);
or U11871 (N_11871,N_11206,N_11325);
xnor U11872 (N_11872,N_11401,N_11439);
or U11873 (N_11873,N_11325,N_11511);
or U11874 (N_11874,N_11299,N_11325);
and U11875 (N_11875,N_11459,N_11433);
and U11876 (N_11876,N_11289,N_11414);
or U11877 (N_11877,N_11507,N_11297);
and U11878 (N_11878,N_11495,N_11517);
and U11879 (N_11879,N_11304,N_11533);
xor U11880 (N_11880,N_11463,N_11324);
nand U11881 (N_11881,N_11440,N_11332);
nand U11882 (N_11882,N_11301,N_11445);
and U11883 (N_11883,N_11305,N_11348);
and U11884 (N_11884,N_11547,N_11524);
nor U11885 (N_11885,N_11577,N_11483);
or U11886 (N_11886,N_11443,N_11263);
nor U11887 (N_11887,N_11562,N_11318);
xor U11888 (N_11888,N_11359,N_11267);
nor U11889 (N_11889,N_11329,N_11238);
nor U11890 (N_11890,N_11284,N_11339);
or U11891 (N_11891,N_11425,N_11345);
and U11892 (N_11892,N_11393,N_11337);
and U11893 (N_11893,N_11312,N_11525);
and U11894 (N_11894,N_11462,N_11311);
nor U11895 (N_11895,N_11217,N_11329);
or U11896 (N_11896,N_11321,N_11326);
nand U11897 (N_11897,N_11221,N_11433);
and U11898 (N_11898,N_11513,N_11311);
xnor U11899 (N_11899,N_11525,N_11205);
or U11900 (N_11900,N_11440,N_11385);
or U11901 (N_11901,N_11262,N_11532);
and U11902 (N_11902,N_11414,N_11432);
xor U11903 (N_11903,N_11202,N_11534);
nand U11904 (N_11904,N_11598,N_11217);
and U11905 (N_11905,N_11386,N_11521);
nand U11906 (N_11906,N_11214,N_11527);
or U11907 (N_11907,N_11487,N_11538);
or U11908 (N_11908,N_11292,N_11316);
nand U11909 (N_11909,N_11367,N_11211);
nor U11910 (N_11910,N_11382,N_11275);
and U11911 (N_11911,N_11354,N_11411);
or U11912 (N_11912,N_11596,N_11285);
and U11913 (N_11913,N_11559,N_11550);
and U11914 (N_11914,N_11384,N_11416);
nand U11915 (N_11915,N_11276,N_11451);
xnor U11916 (N_11916,N_11519,N_11343);
or U11917 (N_11917,N_11323,N_11491);
nand U11918 (N_11918,N_11560,N_11341);
nor U11919 (N_11919,N_11283,N_11241);
or U11920 (N_11920,N_11502,N_11573);
nor U11921 (N_11921,N_11328,N_11460);
nor U11922 (N_11922,N_11592,N_11207);
and U11923 (N_11923,N_11457,N_11367);
or U11924 (N_11924,N_11325,N_11252);
and U11925 (N_11925,N_11497,N_11328);
nand U11926 (N_11926,N_11389,N_11572);
or U11927 (N_11927,N_11402,N_11494);
nand U11928 (N_11928,N_11396,N_11531);
xor U11929 (N_11929,N_11474,N_11370);
and U11930 (N_11930,N_11464,N_11301);
xnor U11931 (N_11931,N_11521,N_11345);
xnor U11932 (N_11932,N_11522,N_11465);
xnor U11933 (N_11933,N_11285,N_11482);
xnor U11934 (N_11934,N_11296,N_11445);
nor U11935 (N_11935,N_11262,N_11234);
or U11936 (N_11936,N_11442,N_11534);
nand U11937 (N_11937,N_11590,N_11205);
xor U11938 (N_11938,N_11522,N_11594);
nand U11939 (N_11939,N_11531,N_11451);
and U11940 (N_11940,N_11377,N_11201);
or U11941 (N_11941,N_11357,N_11400);
xnor U11942 (N_11942,N_11305,N_11337);
nand U11943 (N_11943,N_11397,N_11591);
and U11944 (N_11944,N_11297,N_11489);
nand U11945 (N_11945,N_11220,N_11459);
or U11946 (N_11946,N_11423,N_11377);
and U11947 (N_11947,N_11338,N_11580);
nor U11948 (N_11948,N_11556,N_11497);
nor U11949 (N_11949,N_11287,N_11223);
and U11950 (N_11950,N_11335,N_11233);
nand U11951 (N_11951,N_11233,N_11415);
nor U11952 (N_11952,N_11317,N_11240);
or U11953 (N_11953,N_11393,N_11322);
or U11954 (N_11954,N_11246,N_11418);
nor U11955 (N_11955,N_11203,N_11516);
or U11956 (N_11956,N_11207,N_11407);
nand U11957 (N_11957,N_11257,N_11553);
nand U11958 (N_11958,N_11407,N_11423);
xnor U11959 (N_11959,N_11376,N_11260);
nand U11960 (N_11960,N_11461,N_11554);
xnor U11961 (N_11961,N_11291,N_11374);
nand U11962 (N_11962,N_11332,N_11212);
nor U11963 (N_11963,N_11269,N_11397);
and U11964 (N_11964,N_11368,N_11592);
or U11965 (N_11965,N_11213,N_11372);
xnor U11966 (N_11966,N_11493,N_11520);
nand U11967 (N_11967,N_11559,N_11487);
nor U11968 (N_11968,N_11410,N_11568);
xnor U11969 (N_11969,N_11443,N_11325);
nor U11970 (N_11970,N_11570,N_11320);
or U11971 (N_11971,N_11357,N_11380);
nor U11972 (N_11972,N_11533,N_11542);
nor U11973 (N_11973,N_11498,N_11308);
nor U11974 (N_11974,N_11248,N_11319);
and U11975 (N_11975,N_11436,N_11400);
and U11976 (N_11976,N_11506,N_11269);
xor U11977 (N_11977,N_11277,N_11421);
nand U11978 (N_11978,N_11253,N_11349);
nor U11979 (N_11979,N_11385,N_11451);
xnor U11980 (N_11980,N_11228,N_11471);
xnor U11981 (N_11981,N_11251,N_11400);
nand U11982 (N_11982,N_11373,N_11443);
xor U11983 (N_11983,N_11290,N_11364);
nand U11984 (N_11984,N_11312,N_11519);
xnor U11985 (N_11985,N_11301,N_11437);
or U11986 (N_11986,N_11401,N_11463);
and U11987 (N_11987,N_11558,N_11225);
nor U11988 (N_11988,N_11566,N_11588);
nor U11989 (N_11989,N_11213,N_11379);
or U11990 (N_11990,N_11349,N_11301);
and U11991 (N_11991,N_11305,N_11550);
nand U11992 (N_11992,N_11385,N_11311);
or U11993 (N_11993,N_11471,N_11516);
nor U11994 (N_11994,N_11380,N_11477);
or U11995 (N_11995,N_11246,N_11565);
nor U11996 (N_11996,N_11452,N_11465);
and U11997 (N_11997,N_11572,N_11424);
xor U11998 (N_11998,N_11529,N_11499);
nor U11999 (N_11999,N_11581,N_11273);
xor U12000 (N_12000,N_11747,N_11764);
nand U12001 (N_12001,N_11840,N_11816);
xor U12002 (N_12002,N_11895,N_11633);
xor U12003 (N_12003,N_11653,N_11805);
and U12004 (N_12004,N_11953,N_11920);
xor U12005 (N_12005,N_11841,N_11718);
nand U12006 (N_12006,N_11916,N_11806);
nor U12007 (N_12007,N_11776,N_11898);
xnor U12008 (N_12008,N_11715,N_11921);
nand U12009 (N_12009,N_11643,N_11970);
xor U12010 (N_12010,N_11654,N_11629);
nor U12011 (N_12011,N_11964,N_11761);
or U12012 (N_12012,N_11635,N_11780);
nand U12013 (N_12013,N_11742,N_11914);
nor U12014 (N_12014,N_11675,N_11753);
nor U12015 (N_12015,N_11620,N_11913);
xor U12016 (N_12016,N_11927,N_11652);
and U12017 (N_12017,N_11834,N_11951);
xor U12018 (N_12018,N_11986,N_11711);
nor U12019 (N_12019,N_11932,N_11706);
xnor U12020 (N_12020,N_11952,N_11782);
xnor U12021 (N_12021,N_11878,N_11601);
nor U12022 (N_12022,N_11904,N_11939);
or U12023 (N_12023,N_11682,N_11650);
and U12024 (N_12024,N_11809,N_11801);
or U12025 (N_12025,N_11857,N_11720);
and U12026 (N_12026,N_11619,N_11866);
nand U12027 (N_12027,N_11680,N_11681);
or U12028 (N_12028,N_11657,N_11956);
xnor U12029 (N_12029,N_11838,N_11661);
nor U12030 (N_12030,N_11665,N_11976);
or U12031 (N_12031,N_11797,N_11911);
or U12032 (N_12032,N_11645,N_11971);
xor U12033 (N_12033,N_11957,N_11900);
and U12034 (N_12034,N_11905,N_11626);
or U12035 (N_12035,N_11859,N_11979);
nor U12036 (N_12036,N_11658,N_11663);
nand U12037 (N_12037,N_11723,N_11978);
nor U12038 (N_12038,N_11694,N_11656);
or U12039 (N_12039,N_11984,N_11710);
and U12040 (N_12040,N_11707,N_11977);
and U12041 (N_12041,N_11798,N_11766);
and U12042 (N_12042,N_11883,N_11750);
and U12043 (N_12043,N_11667,N_11774);
xnor U12044 (N_12044,N_11703,N_11642);
and U12045 (N_12045,N_11655,N_11755);
or U12046 (N_12046,N_11649,N_11947);
xor U12047 (N_12047,N_11968,N_11807);
nor U12048 (N_12048,N_11851,N_11901);
xor U12049 (N_12049,N_11749,N_11818);
and U12050 (N_12050,N_11686,N_11634);
nand U12051 (N_12051,N_11950,N_11821);
or U12052 (N_12052,N_11909,N_11882);
nor U12053 (N_12053,N_11941,N_11704);
or U12054 (N_12054,N_11796,N_11881);
or U12055 (N_12055,N_11611,N_11980);
or U12056 (N_12056,N_11985,N_11736);
nand U12057 (N_12057,N_11922,N_11770);
nor U12058 (N_12058,N_11690,N_11842);
and U12059 (N_12059,N_11726,N_11773);
or U12060 (N_12060,N_11728,N_11600);
nand U12061 (N_12061,N_11676,N_11779);
xnor U12062 (N_12062,N_11751,N_11948);
or U12063 (N_12063,N_11765,N_11693);
and U12064 (N_12064,N_11739,N_11999);
nand U12065 (N_12065,N_11981,N_11908);
nor U12066 (N_12066,N_11931,N_11785);
nand U12067 (N_12067,N_11732,N_11758);
xor U12068 (N_12068,N_11887,N_11983);
nor U12069 (N_12069,N_11695,N_11727);
or U12070 (N_12070,N_11722,N_11616);
nor U12071 (N_12071,N_11832,N_11926);
nor U12072 (N_12072,N_11700,N_11713);
nor U12073 (N_12073,N_11987,N_11836);
or U12074 (N_12074,N_11996,N_11954);
or U12075 (N_12075,N_11698,N_11928);
and U12076 (N_12076,N_11647,N_11624);
xor U12077 (N_12077,N_11648,N_11712);
or U12078 (N_12078,N_11990,N_11828);
xnor U12079 (N_12079,N_11746,N_11991);
nand U12080 (N_12080,N_11839,N_11897);
and U12081 (N_12081,N_11888,N_11877);
xnor U12082 (N_12082,N_11741,N_11691);
and U12083 (N_12083,N_11812,N_11795);
nor U12084 (N_12084,N_11673,N_11874);
xor U12085 (N_12085,N_11783,N_11856);
and U12086 (N_12086,N_11730,N_11872);
xnor U12087 (N_12087,N_11625,N_11992);
nor U12088 (N_12088,N_11603,N_11793);
nand U12089 (N_12089,N_11903,N_11825);
xnor U12090 (N_12090,N_11724,N_11640);
or U12091 (N_12091,N_11889,N_11679);
nand U12092 (N_12092,N_11860,N_11771);
nand U12093 (N_12093,N_11702,N_11989);
xnor U12094 (N_12094,N_11855,N_11631);
xor U12095 (N_12095,N_11623,N_11830);
and U12096 (N_12096,N_11848,N_11811);
nor U12097 (N_12097,N_11775,N_11674);
nand U12098 (N_12098,N_11787,N_11884);
and U12099 (N_12099,N_11791,N_11618);
xnor U12100 (N_12100,N_11824,N_11886);
or U12101 (N_12101,N_11870,N_11973);
and U12102 (N_12102,N_11819,N_11890);
nand U12103 (N_12103,N_11871,N_11891);
and U12104 (N_12104,N_11684,N_11937);
xnor U12105 (N_12105,N_11678,N_11759);
or U12106 (N_12106,N_11935,N_11827);
xor U12107 (N_12107,N_11810,N_11745);
xnor U12108 (N_12108,N_11837,N_11615);
nor U12109 (N_12109,N_11705,N_11716);
nand U12110 (N_12110,N_11627,N_11664);
and U12111 (N_12111,N_11958,N_11781);
or U12112 (N_12112,N_11847,N_11923);
and U12113 (N_12113,N_11636,N_11995);
or U12114 (N_12114,N_11942,N_11902);
and U12115 (N_12115,N_11709,N_11917);
or U12116 (N_12116,N_11862,N_11630);
nand U12117 (N_12117,N_11943,N_11945);
or U12118 (N_12118,N_11814,N_11788);
or U12119 (N_12119,N_11833,N_11609);
or U12120 (N_12120,N_11641,N_11784);
nor U12121 (N_12121,N_11843,N_11602);
or U12122 (N_12122,N_11893,N_11934);
nand U12123 (N_12123,N_11972,N_11734);
nor U12124 (N_12124,N_11683,N_11622);
nor U12125 (N_12125,N_11869,N_11868);
nand U12126 (N_12126,N_11865,N_11974);
nor U12127 (N_12127,N_11685,N_11769);
nand U12128 (N_12128,N_11689,N_11763);
nor U12129 (N_12129,N_11670,N_11799);
nor U12130 (N_12130,N_11725,N_11846);
nor U12131 (N_12131,N_11800,N_11610);
and U12132 (N_12132,N_11899,N_11961);
nand U12133 (N_12133,N_11697,N_11997);
xnor U12134 (N_12134,N_11994,N_11644);
nor U12135 (N_12135,N_11731,N_11614);
or U12136 (N_12136,N_11613,N_11998);
xnor U12137 (N_12137,N_11864,N_11938);
and U12138 (N_12138,N_11925,N_11852);
or U12139 (N_12139,N_11936,N_11786);
or U12140 (N_12140,N_11850,N_11982);
nor U12141 (N_12141,N_11835,N_11919);
or U12142 (N_12142,N_11820,N_11699);
nor U12143 (N_12143,N_11826,N_11965);
and U12144 (N_12144,N_11677,N_11778);
nand U12145 (N_12145,N_11858,N_11912);
nor U12146 (N_12146,N_11845,N_11894);
nor U12147 (N_12147,N_11907,N_11748);
or U12148 (N_12148,N_11831,N_11967);
or U12149 (N_12149,N_11606,N_11687);
or U12150 (N_12150,N_11933,N_11651);
or U12151 (N_12151,N_11662,N_11632);
nand U12152 (N_12152,N_11671,N_11607);
or U12153 (N_12153,N_11815,N_11754);
and U12154 (N_12154,N_11804,N_11849);
nor U12155 (N_12155,N_11744,N_11993);
nand U12156 (N_12156,N_11608,N_11962);
nand U12157 (N_12157,N_11760,N_11692);
or U12158 (N_12158,N_11672,N_11817);
xnor U12159 (N_12159,N_11915,N_11743);
and U12160 (N_12160,N_11949,N_11863);
nand U12161 (N_12161,N_11910,N_11719);
nand U12162 (N_12162,N_11659,N_11930);
xnor U12163 (N_12163,N_11756,N_11975);
nor U12164 (N_12164,N_11861,N_11808);
or U12165 (N_12165,N_11717,N_11792);
nor U12166 (N_12166,N_11822,N_11823);
nand U12167 (N_12167,N_11639,N_11637);
and U12168 (N_12168,N_11892,N_11772);
nand U12169 (N_12169,N_11646,N_11789);
nor U12170 (N_12170,N_11794,N_11621);
xnor U12171 (N_12171,N_11873,N_11735);
xor U12172 (N_12172,N_11924,N_11963);
and U12173 (N_12173,N_11777,N_11737);
nand U12174 (N_12174,N_11701,N_11729);
and U12175 (N_12175,N_11969,N_11966);
nand U12176 (N_12176,N_11929,N_11605);
and U12177 (N_12177,N_11628,N_11733);
xnor U12178 (N_12178,N_11853,N_11767);
nor U12179 (N_12179,N_11802,N_11867);
xor U12180 (N_12180,N_11612,N_11960);
and U12181 (N_12181,N_11803,N_11876);
nor U12182 (N_12182,N_11940,N_11955);
nand U12183 (N_12183,N_11854,N_11813);
and U12184 (N_12184,N_11669,N_11875);
or U12185 (N_12185,N_11738,N_11708);
xnor U12186 (N_12186,N_11638,N_11757);
nor U12187 (N_12187,N_11959,N_11829);
xnor U12188 (N_12188,N_11768,N_11906);
xor U12189 (N_12189,N_11885,N_11988);
and U12190 (N_12190,N_11879,N_11790);
nand U12191 (N_12191,N_11688,N_11668);
or U12192 (N_12192,N_11944,N_11946);
xor U12193 (N_12193,N_11696,N_11762);
nand U12194 (N_12194,N_11660,N_11918);
xor U12195 (N_12195,N_11740,N_11880);
xor U12196 (N_12196,N_11721,N_11666);
nor U12197 (N_12197,N_11617,N_11604);
and U12198 (N_12198,N_11896,N_11714);
nor U12199 (N_12199,N_11844,N_11752);
and U12200 (N_12200,N_11645,N_11761);
nand U12201 (N_12201,N_11686,N_11621);
and U12202 (N_12202,N_11664,N_11992);
nor U12203 (N_12203,N_11637,N_11803);
nand U12204 (N_12204,N_11620,N_11965);
nand U12205 (N_12205,N_11910,N_11611);
xor U12206 (N_12206,N_11857,N_11682);
nor U12207 (N_12207,N_11944,N_11872);
nand U12208 (N_12208,N_11843,N_11778);
nor U12209 (N_12209,N_11708,N_11624);
nand U12210 (N_12210,N_11977,N_11971);
or U12211 (N_12211,N_11743,N_11987);
or U12212 (N_12212,N_11988,N_11896);
nor U12213 (N_12213,N_11654,N_11906);
and U12214 (N_12214,N_11908,N_11652);
nor U12215 (N_12215,N_11859,N_11720);
nand U12216 (N_12216,N_11607,N_11753);
or U12217 (N_12217,N_11671,N_11862);
nand U12218 (N_12218,N_11983,N_11969);
nand U12219 (N_12219,N_11836,N_11891);
and U12220 (N_12220,N_11889,N_11914);
and U12221 (N_12221,N_11678,N_11963);
or U12222 (N_12222,N_11969,N_11622);
xnor U12223 (N_12223,N_11943,N_11743);
nor U12224 (N_12224,N_11823,N_11880);
or U12225 (N_12225,N_11775,N_11824);
or U12226 (N_12226,N_11823,N_11837);
or U12227 (N_12227,N_11662,N_11746);
nor U12228 (N_12228,N_11674,N_11779);
or U12229 (N_12229,N_11977,N_11884);
xor U12230 (N_12230,N_11750,N_11636);
or U12231 (N_12231,N_11805,N_11771);
nor U12232 (N_12232,N_11606,N_11814);
nand U12233 (N_12233,N_11629,N_11655);
xor U12234 (N_12234,N_11909,N_11625);
xor U12235 (N_12235,N_11974,N_11620);
nor U12236 (N_12236,N_11980,N_11623);
or U12237 (N_12237,N_11677,N_11868);
nand U12238 (N_12238,N_11744,N_11642);
nand U12239 (N_12239,N_11684,N_11650);
nor U12240 (N_12240,N_11801,N_11777);
or U12241 (N_12241,N_11670,N_11899);
nor U12242 (N_12242,N_11931,N_11858);
xnor U12243 (N_12243,N_11949,N_11604);
nand U12244 (N_12244,N_11719,N_11972);
nor U12245 (N_12245,N_11852,N_11928);
nor U12246 (N_12246,N_11823,N_11899);
xnor U12247 (N_12247,N_11647,N_11757);
or U12248 (N_12248,N_11727,N_11650);
nor U12249 (N_12249,N_11862,N_11993);
and U12250 (N_12250,N_11609,N_11626);
nor U12251 (N_12251,N_11704,N_11912);
nor U12252 (N_12252,N_11807,N_11735);
or U12253 (N_12253,N_11970,N_11727);
nand U12254 (N_12254,N_11671,N_11832);
nand U12255 (N_12255,N_11976,N_11878);
nand U12256 (N_12256,N_11803,N_11775);
and U12257 (N_12257,N_11796,N_11842);
nand U12258 (N_12258,N_11687,N_11706);
or U12259 (N_12259,N_11843,N_11669);
nor U12260 (N_12260,N_11612,N_11820);
nand U12261 (N_12261,N_11941,N_11987);
nor U12262 (N_12262,N_11772,N_11941);
or U12263 (N_12263,N_11978,N_11767);
nand U12264 (N_12264,N_11794,N_11957);
or U12265 (N_12265,N_11932,N_11658);
xnor U12266 (N_12266,N_11809,N_11663);
and U12267 (N_12267,N_11950,N_11683);
nand U12268 (N_12268,N_11771,N_11994);
and U12269 (N_12269,N_11735,N_11695);
nand U12270 (N_12270,N_11958,N_11725);
nor U12271 (N_12271,N_11648,N_11717);
nand U12272 (N_12272,N_11977,N_11857);
xnor U12273 (N_12273,N_11953,N_11730);
nand U12274 (N_12274,N_11779,N_11788);
and U12275 (N_12275,N_11835,N_11615);
or U12276 (N_12276,N_11699,N_11940);
nor U12277 (N_12277,N_11807,N_11912);
xnor U12278 (N_12278,N_11852,N_11806);
nor U12279 (N_12279,N_11810,N_11684);
nand U12280 (N_12280,N_11691,N_11783);
or U12281 (N_12281,N_11746,N_11797);
xnor U12282 (N_12282,N_11888,N_11683);
nand U12283 (N_12283,N_11657,N_11871);
and U12284 (N_12284,N_11754,N_11919);
or U12285 (N_12285,N_11696,N_11767);
nor U12286 (N_12286,N_11927,N_11930);
and U12287 (N_12287,N_11785,N_11704);
nand U12288 (N_12288,N_11976,N_11620);
or U12289 (N_12289,N_11963,N_11786);
nand U12290 (N_12290,N_11802,N_11614);
nor U12291 (N_12291,N_11792,N_11738);
nand U12292 (N_12292,N_11852,N_11912);
xor U12293 (N_12293,N_11740,N_11778);
and U12294 (N_12294,N_11855,N_11798);
nand U12295 (N_12295,N_11713,N_11910);
or U12296 (N_12296,N_11885,N_11947);
nand U12297 (N_12297,N_11857,N_11784);
and U12298 (N_12298,N_11902,N_11739);
nand U12299 (N_12299,N_11981,N_11821);
xnor U12300 (N_12300,N_11770,N_11670);
and U12301 (N_12301,N_11804,N_11953);
nand U12302 (N_12302,N_11739,N_11670);
and U12303 (N_12303,N_11618,N_11950);
or U12304 (N_12304,N_11679,N_11663);
or U12305 (N_12305,N_11616,N_11764);
nor U12306 (N_12306,N_11628,N_11603);
or U12307 (N_12307,N_11869,N_11881);
xnor U12308 (N_12308,N_11793,N_11837);
xor U12309 (N_12309,N_11636,N_11753);
xor U12310 (N_12310,N_11798,N_11918);
or U12311 (N_12311,N_11741,N_11730);
nand U12312 (N_12312,N_11754,N_11934);
xnor U12313 (N_12313,N_11891,N_11672);
nand U12314 (N_12314,N_11679,N_11953);
nor U12315 (N_12315,N_11651,N_11629);
xor U12316 (N_12316,N_11699,N_11990);
nand U12317 (N_12317,N_11804,N_11887);
xor U12318 (N_12318,N_11920,N_11917);
and U12319 (N_12319,N_11705,N_11725);
and U12320 (N_12320,N_11914,N_11604);
nand U12321 (N_12321,N_11989,N_11843);
xnor U12322 (N_12322,N_11601,N_11986);
nand U12323 (N_12323,N_11857,N_11769);
nor U12324 (N_12324,N_11773,N_11883);
nand U12325 (N_12325,N_11647,N_11772);
nand U12326 (N_12326,N_11665,N_11969);
and U12327 (N_12327,N_11996,N_11697);
nor U12328 (N_12328,N_11824,N_11637);
nand U12329 (N_12329,N_11624,N_11786);
nor U12330 (N_12330,N_11956,N_11730);
nand U12331 (N_12331,N_11681,N_11987);
or U12332 (N_12332,N_11816,N_11652);
nand U12333 (N_12333,N_11780,N_11787);
nand U12334 (N_12334,N_11749,N_11973);
xnor U12335 (N_12335,N_11947,N_11618);
xor U12336 (N_12336,N_11959,N_11686);
nor U12337 (N_12337,N_11753,N_11618);
or U12338 (N_12338,N_11710,N_11645);
or U12339 (N_12339,N_11897,N_11681);
nor U12340 (N_12340,N_11703,N_11984);
and U12341 (N_12341,N_11770,N_11812);
and U12342 (N_12342,N_11641,N_11971);
xor U12343 (N_12343,N_11680,N_11776);
and U12344 (N_12344,N_11840,N_11766);
and U12345 (N_12345,N_11930,N_11753);
nand U12346 (N_12346,N_11969,N_11787);
nor U12347 (N_12347,N_11781,N_11957);
nor U12348 (N_12348,N_11640,N_11766);
and U12349 (N_12349,N_11768,N_11600);
nand U12350 (N_12350,N_11746,N_11891);
nand U12351 (N_12351,N_11685,N_11789);
and U12352 (N_12352,N_11778,N_11605);
xor U12353 (N_12353,N_11904,N_11712);
xor U12354 (N_12354,N_11775,N_11891);
xnor U12355 (N_12355,N_11601,N_11800);
xor U12356 (N_12356,N_11724,N_11836);
and U12357 (N_12357,N_11911,N_11619);
or U12358 (N_12358,N_11900,N_11973);
xnor U12359 (N_12359,N_11750,N_11993);
nor U12360 (N_12360,N_11821,N_11854);
and U12361 (N_12361,N_11624,N_11669);
or U12362 (N_12362,N_11622,N_11777);
or U12363 (N_12363,N_11788,N_11678);
nand U12364 (N_12364,N_11678,N_11973);
nor U12365 (N_12365,N_11911,N_11999);
and U12366 (N_12366,N_11760,N_11770);
nand U12367 (N_12367,N_11630,N_11874);
or U12368 (N_12368,N_11838,N_11691);
and U12369 (N_12369,N_11887,N_11779);
and U12370 (N_12370,N_11685,N_11884);
and U12371 (N_12371,N_11701,N_11992);
xor U12372 (N_12372,N_11775,N_11847);
xnor U12373 (N_12373,N_11904,N_11611);
nor U12374 (N_12374,N_11984,N_11944);
and U12375 (N_12375,N_11639,N_11973);
nand U12376 (N_12376,N_11603,N_11709);
or U12377 (N_12377,N_11749,N_11635);
nand U12378 (N_12378,N_11629,N_11803);
or U12379 (N_12379,N_11757,N_11633);
xnor U12380 (N_12380,N_11823,N_11986);
or U12381 (N_12381,N_11631,N_11986);
nand U12382 (N_12382,N_11906,N_11816);
nor U12383 (N_12383,N_11954,N_11681);
xnor U12384 (N_12384,N_11639,N_11645);
xnor U12385 (N_12385,N_11815,N_11641);
nor U12386 (N_12386,N_11698,N_11689);
nand U12387 (N_12387,N_11795,N_11944);
and U12388 (N_12388,N_11714,N_11917);
nand U12389 (N_12389,N_11817,N_11910);
nand U12390 (N_12390,N_11664,N_11828);
and U12391 (N_12391,N_11924,N_11897);
and U12392 (N_12392,N_11775,N_11703);
nand U12393 (N_12393,N_11964,N_11901);
xor U12394 (N_12394,N_11752,N_11902);
xor U12395 (N_12395,N_11883,N_11943);
nor U12396 (N_12396,N_11965,N_11730);
nand U12397 (N_12397,N_11750,N_11791);
nor U12398 (N_12398,N_11759,N_11877);
nor U12399 (N_12399,N_11932,N_11652);
xor U12400 (N_12400,N_12071,N_12006);
or U12401 (N_12401,N_12285,N_12094);
nand U12402 (N_12402,N_12267,N_12025);
nor U12403 (N_12403,N_12233,N_12398);
xnor U12404 (N_12404,N_12184,N_12309);
nor U12405 (N_12405,N_12042,N_12275);
or U12406 (N_12406,N_12041,N_12258);
nor U12407 (N_12407,N_12347,N_12009);
xnor U12408 (N_12408,N_12290,N_12052);
nor U12409 (N_12409,N_12159,N_12167);
or U12410 (N_12410,N_12246,N_12277);
and U12411 (N_12411,N_12260,N_12352);
or U12412 (N_12412,N_12008,N_12075);
xor U12413 (N_12413,N_12093,N_12118);
and U12414 (N_12414,N_12336,N_12179);
and U12415 (N_12415,N_12023,N_12280);
nor U12416 (N_12416,N_12324,N_12395);
xor U12417 (N_12417,N_12091,N_12252);
or U12418 (N_12418,N_12058,N_12357);
xnor U12419 (N_12419,N_12278,N_12100);
and U12420 (N_12420,N_12232,N_12081);
nand U12421 (N_12421,N_12027,N_12107);
nand U12422 (N_12422,N_12211,N_12222);
nand U12423 (N_12423,N_12339,N_12004);
nand U12424 (N_12424,N_12351,N_12151);
and U12425 (N_12425,N_12036,N_12143);
xnor U12426 (N_12426,N_12349,N_12360);
xor U12427 (N_12427,N_12015,N_12029);
nand U12428 (N_12428,N_12030,N_12354);
nor U12429 (N_12429,N_12127,N_12343);
or U12430 (N_12430,N_12097,N_12202);
or U12431 (N_12431,N_12087,N_12072);
or U12432 (N_12432,N_12055,N_12155);
and U12433 (N_12433,N_12163,N_12134);
nand U12434 (N_12434,N_12189,N_12158);
nand U12435 (N_12435,N_12390,N_12310);
and U12436 (N_12436,N_12197,N_12065);
and U12437 (N_12437,N_12335,N_12371);
nand U12438 (N_12438,N_12079,N_12243);
or U12439 (N_12439,N_12121,N_12085);
xnor U12440 (N_12440,N_12053,N_12021);
xor U12441 (N_12441,N_12133,N_12294);
or U12442 (N_12442,N_12177,N_12399);
nand U12443 (N_12443,N_12005,N_12368);
or U12444 (N_12444,N_12288,N_12261);
or U12445 (N_12445,N_12296,N_12378);
xor U12446 (N_12446,N_12328,N_12176);
nor U12447 (N_12447,N_12314,N_12255);
or U12448 (N_12448,N_12321,N_12325);
nand U12449 (N_12449,N_12376,N_12069);
and U12450 (N_12450,N_12039,N_12082);
or U12451 (N_12451,N_12326,N_12056);
nand U12452 (N_12452,N_12122,N_12073);
nor U12453 (N_12453,N_12161,N_12224);
nand U12454 (N_12454,N_12305,N_12103);
nor U12455 (N_12455,N_12312,N_12283);
xor U12456 (N_12456,N_12044,N_12385);
and U12457 (N_12457,N_12175,N_12026);
nand U12458 (N_12458,N_12210,N_12120);
and U12459 (N_12459,N_12198,N_12199);
xor U12460 (N_12460,N_12397,N_12236);
xnor U12461 (N_12461,N_12353,N_12102);
nand U12462 (N_12462,N_12392,N_12219);
or U12463 (N_12463,N_12089,N_12051);
nor U12464 (N_12464,N_12387,N_12215);
or U12465 (N_12465,N_12111,N_12286);
or U12466 (N_12466,N_12345,N_12342);
nand U12467 (N_12467,N_12311,N_12186);
nor U12468 (N_12468,N_12194,N_12284);
or U12469 (N_12469,N_12396,N_12003);
xor U12470 (N_12470,N_12138,N_12374);
nor U12471 (N_12471,N_12046,N_12054);
or U12472 (N_12472,N_12274,N_12217);
xor U12473 (N_12473,N_12037,N_12237);
nand U12474 (N_12474,N_12361,N_12332);
or U12475 (N_12475,N_12185,N_12156);
nor U12476 (N_12476,N_12050,N_12307);
xnor U12477 (N_12477,N_12128,N_12016);
nor U12478 (N_12478,N_12316,N_12337);
xor U12479 (N_12479,N_12173,N_12221);
and U12480 (N_12480,N_12112,N_12209);
and U12481 (N_12481,N_12295,N_12126);
or U12482 (N_12482,N_12125,N_12287);
nand U12483 (N_12483,N_12379,N_12329);
nand U12484 (N_12484,N_12077,N_12256);
or U12485 (N_12485,N_12187,N_12250);
xor U12486 (N_12486,N_12317,N_12205);
and U12487 (N_12487,N_12190,N_12164);
and U12488 (N_12488,N_12124,N_12377);
nand U12489 (N_12489,N_12137,N_12235);
xnor U12490 (N_12490,N_12240,N_12251);
xnor U12491 (N_12491,N_12109,N_12359);
nor U12492 (N_12492,N_12154,N_12034);
or U12493 (N_12493,N_12262,N_12289);
nand U12494 (N_12494,N_12062,N_12273);
nor U12495 (N_12495,N_12135,N_12007);
xnor U12496 (N_12496,N_12099,N_12270);
nand U12497 (N_12497,N_12227,N_12017);
and U12498 (N_12498,N_12153,N_12279);
or U12499 (N_12499,N_12024,N_12370);
or U12500 (N_12500,N_12226,N_12152);
xor U12501 (N_12501,N_12178,N_12063);
nor U12502 (N_12502,N_12001,N_12191);
nand U12503 (N_12503,N_12031,N_12132);
nand U12504 (N_12504,N_12308,N_12149);
xor U12505 (N_12505,N_12231,N_12192);
nor U12506 (N_12506,N_12047,N_12358);
and U12507 (N_12507,N_12291,N_12384);
nor U12508 (N_12508,N_12220,N_12101);
or U12509 (N_12509,N_12306,N_12105);
xnor U12510 (N_12510,N_12259,N_12180);
nor U12511 (N_12511,N_12011,N_12320);
nand U12512 (N_12512,N_12067,N_12060);
nand U12513 (N_12513,N_12012,N_12083);
nand U12514 (N_12514,N_12264,N_12282);
and U12515 (N_12515,N_12172,N_12193);
nand U12516 (N_12516,N_12207,N_12212);
nor U12517 (N_12517,N_12281,N_12057);
or U12518 (N_12518,N_12302,N_12117);
nor U12519 (N_12519,N_12228,N_12114);
nor U12520 (N_12520,N_12182,N_12223);
and U12521 (N_12521,N_12363,N_12171);
nor U12522 (N_12522,N_12214,N_12014);
and U12523 (N_12523,N_12315,N_12200);
or U12524 (N_12524,N_12070,N_12365);
or U12525 (N_12525,N_12327,N_12375);
or U12526 (N_12526,N_12206,N_12218);
xnor U12527 (N_12527,N_12096,N_12247);
nor U12528 (N_12528,N_12268,N_12033);
nand U12529 (N_12529,N_12139,N_12254);
or U12530 (N_12530,N_12131,N_12130);
nor U12531 (N_12531,N_12391,N_12263);
nor U12532 (N_12532,N_12393,N_12145);
and U12533 (N_12533,N_12098,N_12108);
and U12534 (N_12534,N_12350,N_12043);
nand U12535 (N_12535,N_12230,N_12066);
nand U12536 (N_12536,N_12330,N_12338);
nor U12537 (N_12537,N_12297,N_12257);
nor U12538 (N_12538,N_12367,N_12394);
nand U12539 (N_12539,N_12382,N_12276);
nor U12540 (N_12540,N_12319,N_12340);
nor U12541 (N_12541,N_12389,N_12115);
nand U12542 (N_12542,N_12271,N_12265);
xnor U12543 (N_12543,N_12157,N_12344);
xor U12544 (N_12544,N_12076,N_12068);
nand U12545 (N_12545,N_12322,N_12346);
or U12546 (N_12546,N_12301,N_12086);
and U12547 (N_12547,N_12242,N_12110);
nor U12548 (N_12548,N_12123,N_12196);
or U12549 (N_12549,N_12292,N_12141);
and U12550 (N_12550,N_12356,N_12388);
xor U12551 (N_12551,N_12298,N_12341);
and U12552 (N_12552,N_12165,N_12216);
nand U12553 (N_12553,N_12059,N_12383);
or U12554 (N_12554,N_12244,N_12362);
nand U12555 (N_12555,N_12084,N_12048);
xor U12556 (N_12556,N_12020,N_12148);
or U12557 (N_12557,N_12300,N_12095);
xor U12558 (N_12558,N_12304,N_12239);
nand U12559 (N_12559,N_12106,N_12090);
nand U12560 (N_12560,N_12355,N_12266);
or U12561 (N_12561,N_12245,N_12174);
nand U12562 (N_12562,N_12299,N_12144);
and U12563 (N_12563,N_12038,N_12116);
and U12564 (N_12564,N_12147,N_12334);
nand U12565 (N_12565,N_12045,N_12201);
xor U12566 (N_12566,N_12035,N_12160);
and U12567 (N_12567,N_12204,N_12104);
nand U12568 (N_12568,N_12373,N_12170);
xor U12569 (N_12569,N_12019,N_12140);
nand U12570 (N_12570,N_12195,N_12129);
and U12571 (N_12571,N_12188,N_12022);
and U12572 (N_12572,N_12119,N_12241);
nor U12573 (N_12573,N_12078,N_12168);
nor U12574 (N_12574,N_12313,N_12028);
or U12575 (N_12575,N_12213,N_12293);
xor U12576 (N_12576,N_12162,N_12272);
and U12577 (N_12577,N_12253,N_12183);
or U12578 (N_12578,N_12136,N_12366);
nand U12579 (N_12579,N_12203,N_12364);
or U12580 (N_12580,N_12269,N_12323);
nand U12581 (N_12581,N_12331,N_12372);
nor U12582 (N_12582,N_12169,N_12208);
nand U12583 (N_12583,N_12234,N_12088);
nor U12584 (N_12584,N_12040,N_12381);
or U12585 (N_12585,N_12013,N_12049);
xor U12586 (N_12586,N_12303,N_12064);
nor U12587 (N_12587,N_12181,N_12074);
nand U12588 (N_12588,N_12225,N_12142);
nor U12589 (N_12589,N_12032,N_12080);
nor U12590 (N_12590,N_12318,N_12348);
or U12591 (N_12591,N_12369,N_12386);
and U12592 (N_12592,N_12150,N_12238);
nor U12593 (N_12593,N_12380,N_12113);
or U12594 (N_12594,N_12146,N_12010);
nand U12595 (N_12595,N_12061,N_12248);
nor U12596 (N_12596,N_12092,N_12018);
or U12597 (N_12597,N_12166,N_12249);
nor U12598 (N_12598,N_12002,N_12333);
nor U12599 (N_12599,N_12000,N_12229);
or U12600 (N_12600,N_12087,N_12196);
or U12601 (N_12601,N_12373,N_12263);
xor U12602 (N_12602,N_12352,N_12198);
or U12603 (N_12603,N_12368,N_12371);
xnor U12604 (N_12604,N_12165,N_12010);
or U12605 (N_12605,N_12368,N_12056);
nand U12606 (N_12606,N_12048,N_12054);
nand U12607 (N_12607,N_12252,N_12191);
nor U12608 (N_12608,N_12229,N_12361);
and U12609 (N_12609,N_12373,N_12293);
or U12610 (N_12610,N_12346,N_12264);
nor U12611 (N_12611,N_12366,N_12030);
and U12612 (N_12612,N_12273,N_12346);
xor U12613 (N_12613,N_12233,N_12376);
or U12614 (N_12614,N_12152,N_12102);
nor U12615 (N_12615,N_12046,N_12372);
nor U12616 (N_12616,N_12107,N_12176);
and U12617 (N_12617,N_12344,N_12353);
or U12618 (N_12618,N_12326,N_12138);
and U12619 (N_12619,N_12121,N_12277);
nor U12620 (N_12620,N_12071,N_12195);
nor U12621 (N_12621,N_12220,N_12086);
and U12622 (N_12622,N_12169,N_12109);
and U12623 (N_12623,N_12070,N_12333);
or U12624 (N_12624,N_12100,N_12363);
nand U12625 (N_12625,N_12081,N_12316);
nor U12626 (N_12626,N_12145,N_12108);
nand U12627 (N_12627,N_12218,N_12137);
nor U12628 (N_12628,N_12189,N_12314);
nor U12629 (N_12629,N_12080,N_12367);
xnor U12630 (N_12630,N_12184,N_12393);
and U12631 (N_12631,N_12124,N_12197);
nor U12632 (N_12632,N_12187,N_12228);
and U12633 (N_12633,N_12396,N_12339);
nor U12634 (N_12634,N_12203,N_12158);
xor U12635 (N_12635,N_12074,N_12342);
nand U12636 (N_12636,N_12326,N_12382);
and U12637 (N_12637,N_12094,N_12280);
nand U12638 (N_12638,N_12066,N_12170);
xnor U12639 (N_12639,N_12099,N_12151);
xnor U12640 (N_12640,N_12269,N_12142);
and U12641 (N_12641,N_12338,N_12005);
and U12642 (N_12642,N_12162,N_12176);
or U12643 (N_12643,N_12082,N_12348);
nand U12644 (N_12644,N_12246,N_12148);
or U12645 (N_12645,N_12260,N_12177);
nand U12646 (N_12646,N_12100,N_12398);
nand U12647 (N_12647,N_12053,N_12302);
nor U12648 (N_12648,N_12234,N_12061);
nand U12649 (N_12649,N_12182,N_12103);
xor U12650 (N_12650,N_12111,N_12132);
or U12651 (N_12651,N_12073,N_12255);
xnor U12652 (N_12652,N_12028,N_12078);
or U12653 (N_12653,N_12133,N_12128);
nor U12654 (N_12654,N_12368,N_12298);
xor U12655 (N_12655,N_12139,N_12122);
or U12656 (N_12656,N_12179,N_12341);
and U12657 (N_12657,N_12003,N_12318);
nor U12658 (N_12658,N_12089,N_12006);
nor U12659 (N_12659,N_12268,N_12170);
nor U12660 (N_12660,N_12348,N_12156);
xnor U12661 (N_12661,N_12071,N_12106);
nand U12662 (N_12662,N_12294,N_12103);
nand U12663 (N_12663,N_12308,N_12304);
and U12664 (N_12664,N_12391,N_12163);
or U12665 (N_12665,N_12044,N_12094);
xnor U12666 (N_12666,N_12048,N_12304);
nor U12667 (N_12667,N_12295,N_12276);
and U12668 (N_12668,N_12183,N_12206);
and U12669 (N_12669,N_12294,N_12168);
or U12670 (N_12670,N_12105,N_12191);
or U12671 (N_12671,N_12246,N_12132);
or U12672 (N_12672,N_12241,N_12100);
or U12673 (N_12673,N_12098,N_12021);
and U12674 (N_12674,N_12213,N_12167);
nand U12675 (N_12675,N_12354,N_12277);
nand U12676 (N_12676,N_12342,N_12286);
or U12677 (N_12677,N_12362,N_12105);
nand U12678 (N_12678,N_12321,N_12085);
nor U12679 (N_12679,N_12059,N_12374);
nor U12680 (N_12680,N_12147,N_12276);
and U12681 (N_12681,N_12156,N_12138);
xnor U12682 (N_12682,N_12208,N_12078);
nand U12683 (N_12683,N_12180,N_12262);
xnor U12684 (N_12684,N_12348,N_12281);
xor U12685 (N_12685,N_12377,N_12208);
or U12686 (N_12686,N_12372,N_12303);
nor U12687 (N_12687,N_12022,N_12257);
xor U12688 (N_12688,N_12370,N_12251);
or U12689 (N_12689,N_12387,N_12228);
nor U12690 (N_12690,N_12213,N_12246);
xor U12691 (N_12691,N_12004,N_12284);
and U12692 (N_12692,N_12352,N_12358);
or U12693 (N_12693,N_12111,N_12163);
or U12694 (N_12694,N_12348,N_12387);
and U12695 (N_12695,N_12298,N_12103);
nor U12696 (N_12696,N_12181,N_12323);
or U12697 (N_12697,N_12111,N_12004);
nor U12698 (N_12698,N_12263,N_12181);
or U12699 (N_12699,N_12105,N_12177);
nand U12700 (N_12700,N_12174,N_12172);
and U12701 (N_12701,N_12285,N_12082);
nand U12702 (N_12702,N_12182,N_12203);
or U12703 (N_12703,N_12217,N_12242);
and U12704 (N_12704,N_12371,N_12362);
and U12705 (N_12705,N_12175,N_12394);
xnor U12706 (N_12706,N_12366,N_12198);
and U12707 (N_12707,N_12244,N_12054);
xor U12708 (N_12708,N_12326,N_12074);
nor U12709 (N_12709,N_12293,N_12066);
xnor U12710 (N_12710,N_12013,N_12232);
nand U12711 (N_12711,N_12014,N_12330);
nor U12712 (N_12712,N_12386,N_12058);
nand U12713 (N_12713,N_12338,N_12344);
xor U12714 (N_12714,N_12125,N_12306);
nor U12715 (N_12715,N_12338,N_12346);
nand U12716 (N_12716,N_12235,N_12001);
or U12717 (N_12717,N_12189,N_12166);
xor U12718 (N_12718,N_12370,N_12189);
nor U12719 (N_12719,N_12138,N_12388);
and U12720 (N_12720,N_12128,N_12222);
nand U12721 (N_12721,N_12276,N_12041);
or U12722 (N_12722,N_12288,N_12065);
or U12723 (N_12723,N_12346,N_12189);
nand U12724 (N_12724,N_12363,N_12039);
and U12725 (N_12725,N_12101,N_12050);
and U12726 (N_12726,N_12353,N_12183);
nand U12727 (N_12727,N_12254,N_12197);
nor U12728 (N_12728,N_12098,N_12384);
and U12729 (N_12729,N_12388,N_12363);
xor U12730 (N_12730,N_12241,N_12062);
or U12731 (N_12731,N_12329,N_12248);
nor U12732 (N_12732,N_12180,N_12041);
nor U12733 (N_12733,N_12295,N_12083);
xor U12734 (N_12734,N_12376,N_12078);
or U12735 (N_12735,N_12178,N_12168);
nor U12736 (N_12736,N_12095,N_12161);
nor U12737 (N_12737,N_12032,N_12356);
nor U12738 (N_12738,N_12397,N_12132);
nor U12739 (N_12739,N_12229,N_12311);
nand U12740 (N_12740,N_12042,N_12045);
nand U12741 (N_12741,N_12155,N_12323);
nand U12742 (N_12742,N_12359,N_12300);
nand U12743 (N_12743,N_12340,N_12361);
nor U12744 (N_12744,N_12387,N_12379);
nand U12745 (N_12745,N_12141,N_12101);
and U12746 (N_12746,N_12263,N_12247);
xnor U12747 (N_12747,N_12375,N_12070);
or U12748 (N_12748,N_12159,N_12382);
xnor U12749 (N_12749,N_12034,N_12145);
xnor U12750 (N_12750,N_12392,N_12063);
or U12751 (N_12751,N_12253,N_12120);
and U12752 (N_12752,N_12322,N_12139);
xnor U12753 (N_12753,N_12248,N_12153);
or U12754 (N_12754,N_12311,N_12335);
xor U12755 (N_12755,N_12278,N_12019);
nor U12756 (N_12756,N_12066,N_12135);
or U12757 (N_12757,N_12060,N_12138);
xnor U12758 (N_12758,N_12278,N_12176);
xnor U12759 (N_12759,N_12208,N_12163);
xnor U12760 (N_12760,N_12384,N_12184);
nand U12761 (N_12761,N_12312,N_12399);
and U12762 (N_12762,N_12046,N_12210);
nor U12763 (N_12763,N_12244,N_12075);
nor U12764 (N_12764,N_12227,N_12366);
nor U12765 (N_12765,N_12392,N_12225);
or U12766 (N_12766,N_12388,N_12212);
nor U12767 (N_12767,N_12241,N_12390);
and U12768 (N_12768,N_12342,N_12108);
xnor U12769 (N_12769,N_12086,N_12382);
nand U12770 (N_12770,N_12323,N_12278);
and U12771 (N_12771,N_12065,N_12250);
nor U12772 (N_12772,N_12313,N_12361);
and U12773 (N_12773,N_12327,N_12220);
nand U12774 (N_12774,N_12252,N_12259);
and U12775 (N_12775,N_12386,N_12063);
nor U12776 (N_12776,N_12117,N_12044);
nor U12777 (N_12777,N_12185,N_12064);
or U12778 (N_12778,N_12323,N_12066);
and U12779 (N_12779,N_12080,N_12168);
nand U12780 (N_12780,N_12202,N_12171);
and U12781 (N_12781,N_12156,N_12095);
nand U12782 (N_12782,N_12092,N_12222);
nor U12783 (N_12783,N_12384,N_12390);
or U12784 (N_12784,N_12150,N_12053);
nor U12785 (N_12785,N_12174,N_12357);
xor U12786 (N_12786,N_12035,N_12371);
xor U12787 (N_12787,N_12202,N_12000);
or U12788 (N_12788,N_12249,N_12344);
and U12789 (N_12789,N_12196,N_12033);
or U12790 (N_12790,N_12351,N_12172);
and U12791 (N_12791,N_12219,N_12338);
nor U12792 (N_12792,N_12022,N_12244);
or U12793 (N_12793,N_12222,N_12125);
nand U12794 (N_12794,N_12333,N_12154);
nand U12795 (N_12795,N_12102,N_12285);
xor U12796 (N_12796,N_12378,N_12370);
and U12797 (N_12797,N_12121,N_12337);
and U12798 (N_12798,N_12313,N_12120);
nor U12799 (N_12799,N_12249,N_12395);
and U12800 (N_12800,N_12694,N_12658);
or U12801 (N_12801,N_12553,N_12732);
nand U12802 (N_12802,N_12442,N_12405);
and U12803 (N_12803,N_12478,N_12521);
nand U12804 (N_12804,N_12655,N_12578);
nand U12805 (N_12805,N_12600,N_12642);
nand U12806 (N_12806,N_12494,N_12515);
nand U12807 (N_12807,N_12487,N_12627);
and U12808 (N_12808,N_12477,N_12464);
and U12809 (N_12809,N_12593,N_12712);
or U12810 (N_12810,N_12581,N_12713);
nor U12811 (N_12811,N_12696,N_12723);
or U12812 (N_12812,N_12577,N_12678);
nand U12813 (N_12813,N_12454,N_12508);
or U12814 (N_12814,N_12741,N_12419);
nor U12815 (N_12815,N_12591,N_12795);
nor U12816 (N_12816,N_12637,N_12674);
or U12817 (N_12817,N_12728,N_12413);
nand U12818 (N_12818,N_12681,N_12597);
xnor U12819 (N_12819,N_12672,N_12606);
xnor U12820 (N_12820,N_12663,N_12539);
or U12821 (N_12821,N_12613,N_12484);
nor U12822 (N_12822,N_12433,N_12463);
and U12823 (N_12823,N_12408,N_12540);
or U12824 (N_12824,N_12565,N_12476);
nor U12825 (N_12825,N_12799,N_12495);
nand U12826 (N_12826,N_12654,N_12435);
nor U12827 (N_12827,N_12756,N_12783);
or U12828 (N_12828,N_12664,N_12760);
nand U12829 (N_12829,N_12559,N_12744);
or U12830 (N_12830,N_12447,N_12411);
and U12831 (N_12831,N_12762,N_12451);
nand U12832 (N_12832,N_12468,N_12499);
xnor U12833 (N_12833,N_12716,N_12482);
and U12834 (N_12834,N_12523,N_12704);
nor U12835 (N_12835,N_12595,N_12432);
xnor U12836 (N_12836,N_12656,N_12511);
nor U12837 (N_12837,N_12603,N_12786);
or U12838 (N_12838,N_12772,N_12736);
and U12839 (N_12839,N_12586,N_12640);
xor U12840 (N_12840,N_12552,N_12737);
and U12841 (N_12841,N_12645,N_12519);
nand U12842 (N_12842,N_12438,N_12702);
or U12843 (N_12843,N_12682,N_12501);
nand U12844 (N_12844,N_12685,N_12714);
or U12845 (N_12845,N_12507,N_12527);
nor U12846 (N_12846,N_12441,N_12695);
nor U12847 (N_12847,N_12444,N_12479);
xnor U12848 (N_12848,N_12779,N_12576);
or U12849 (N_12849,N_12584,N_12406);
nand U12850 (N_12850,N_12749,N_12746);
or U12851 (N_12851,N_12776,N_12763);
nand U12852 (N_12852,N_12687,N_12427);
and U12853 (N_12853,N_12548,N_12498);
nor U12854 (N_12854,N_12415,N_12619);
nor U12855 (N_12855,N_12780,N_12503);
or U12856 (N_12856,N_12446,N_12797);
nor U12857 (N_12857,N_12489,N_12409);
nand U12858 (N_12858,N_12631,N_12570);
nor U12859 (N_12859,N_12452,N_12416);
nand U12860 (N_12860,N_12531,N_12679);
nand U12861 (N_12861,N_12533,N_12676);
or U12862 (N_12862,N_12480,N_12556);
xor U12863 (N_12863,N_12580,N_12575);
nor U12864 (N_12864,N_12668,N_12569);
xor U12865 (N_12865,N_12688,N_12607);
and U12866 (N_12866,N_12598,N_12758);
or U12867 (N_12867,N_12430,N_12529);
or U12868 (N_12868,N_12750,N_12617);
nand U12869 (N_12869,N_12740,N_12757);
nand U12870 (N_12870,N_12618,N_12517);
and U12871 (N_12871,N_12417,N_12693);
nor U12872 (N_12872,N_12789,N_12555);
or U12873 (N_12873,N_12609,N_12530);
nor U12874 (N_12874,N_12491,N_12662);
nor U12875 (N_12875,N_12751,N_12660);
nor U12876 (N_12876,N_12761,N_12557);
nor U12877 (N_12877,N_12493,N_12599);
nor U12878 (N_12878,N_12766,N_12460);
nor U12879 (N_12879,N_12722,N_12458);
and U12880 (N_12880,N_12437,N_12615);
nand U12881 (N_12881,N_12745,N_12686);
or U12882 (N_12882,N_12407,N_12512);
and U12883 (N_12883,N_12453,N_12610);
nand U12884 (N_12884,N_12703,N_12765);
or U12885 (N_12885,N_12455,N_12720);
nand U12886 (N_12886,N_12743,N_12572);
or U12887 (N_12887,N_12735,N_12585);
nor U12888 (N_12888,N_12680,N_12462);
or U12889 (N_12889,N_12418,N_12469);
nand U12890 (N_12890,N_12709,N_12425);
xor U12891 (N_12891,N_12421,N_12629);
and U12892 (N_12892,N_12796,N_12520);
and U12893 (N_12893,N_12510,N_12546);
xnor U12894 (N_12894,N_12788,N_12544);
xor U12895 (N_12895,N_12504,N_12675);
xor U12896 (N_12896,N_12538,N_12592);
xnor U12897 (N_12897,N_12730,N_12422);
nor U12898 (N_12898,N_12719,N_12759);
xor U12899 (N_12899,N_12456,N_12535);
and U12900 (N_12900,N_12781,N_12646);
nand U12901 (N_12901,N_12601,N_12459);
nand U12902 (N_12902,N_12628,N_12566);
xnor U12903 (N_12903,N_12414,N_12708);
nor U12904 (N_12904,N_12647,N_12638);
nand U12905 (N_12905,N_12697,N_12505);
nand U12906 (N_12906,N_12567,N_12784);
or U12907 (N_12907,N_12400,N_12727);
nor U12908 (N_12908,N_12604,N_12428);
or U12909 (N_12909,N_12614,N_12725);
or U12910 (N_12910,N_12733,N_12516);
nor U12911 (N_12911,N_12542,N_12549);
xor U12912 (N_12912,N_12475,N_12653);
or U12913 (N_12913,N_12785,N_12470);
nand U12914 (N_12914,N_12424,N_12777);
nand U12915 (N_12915,N_12648,N_12691);
or U12916 (N_12916,N_12473,N_12547);
xnor U12917 (N_12917,N_12689,N_12624);
and U12918 (N_12918,N_12699,N_12594);
nor U12919 (N_12919,N_12589,N_12650);
xor U12920 (N_12920,N_12449,N_12561);
nor U12921 (N_12921,N_12753,N_12402);
nor U12922 (N_12922,N_12734,N_12706);
nor U12923 (N_12923,N_12790,N_12457);
and U12924 (N_12924,N_12560,N_12673);
xnor U12925 (N_12925,N_12573,N_12621);
xor U12926 (N_12926,N_12775,N_12711);
or U12927 (N_12927,N_12490,N_12543);
xnor U12928 (N_12928,N_12429,N_12792);
nor U12929 (N_12929,N_12541,N_12602);
or U12930 (N_12930,N_12705,N_12724);
or U12931 (N_12931,N_12536,N_12665);
nor U12932 (N_12932,N_12738,N_12562);
and U12933 (N_12933,N_12509,N_12483);
nor U12934 (N_12934,N_12692,N_12485);
nand U12935 (N_12935,N_12563,N_12558);
and U12936 (N_12936,N_12525,N_12568);
xor U12937 (N_12937,N_12742,N_12467);
and U12938 (N_12938,N_12590,N_12574);
and U12939 (N_12939,N_12798,N_12502);
nor U12940 (N_12940,N_12644,N_12439);
nor U12941 (N_12941,N_12683,N_12532);
nor U12942 (N_12942,N_12634,N_12731);
or U12943 (N_12943,N_12528,N_12434);
and U12944 (N_12944,N_12793,N_12671);
and U12945 (N_12945,N_12461,N_12641);
nor U12946 (N_12946,N_12710,N_12666);
or U12947 (N_12947,N_12623,N_12774);
nor U12948 (N_12948,N_12534,N_12769);
and U12949 (N_12949,N_12481,N_12657);
and U12950 (N_12950,N_12471,N_12684);
and U12951 (N_12951,N_12496,N_12729);
and U12952 (N_12952,N_12787,N_12423);
or U12953 (N_12953,N_12707,N_12773);
xor U12954 (N_12954,N_12669,N_12583);
and U12955 (N_12955,N_12667,N_12513);
or U12956 (N_12956,N_12582,N_12690);
nor U12957 (N_12957,N_12497,N_12551);
nand U12958 (N_12958,N_12721,N_12401);
nand U12959 (N_12959,N_12472,N_12649);
nor U12960 (N_12960,N_12625,N_12782);
nor U12961 (N_12961,N_12550,N_12701);
xor U12962 (N_12962,N_12518,N_12404);
or U12963 (N_12963,N_12545,N_12770);
and U12964 (N_12964,N_12571,N_12436);
and U12965 (N_12965,N_12755,N_12426);
and U12966 (N_12966,N_12611,N_12474);
nor U12967 (N_12967,N_12537,N_12431);
nand U12968 (N_12968,N_12588,N_12514);
or U12969 (N_12969,N_12651,N_12596);
and U12970 (N_12970,N_12486,N_12506);
and U12971 (N_12971,N_12605,N_12739);
xor U12972 (N_12972,N_12522,N_12492);
xor U12973 (N_12973,N_12791,N_12677);
and U12974 (N_12974,N_12587,N_12718);
xnor U12975 (N_12975,N_12659,N_12630);
and U12976 (N_12976,N_12620,N_12639);
xor U12977 (N_12977,N_12445,N_12440);
nor U12978 (N_12978,N_12700,N_12715);
or U12979 (N_12979,N_12554,N_12579);
and U12980 (N_12980,N_12420,N_12726);
nor U12981 (N_12981,N_12500,N_12643);
nor U12982 (N_12982,N_12717,N_12448);
xnor U12983 (N_12983,N_12636,N_12626);
xor U12984 (N_12984,N_12403,N_12564);
nor U12985 (N_12985,N_12764,N_12635);
xor U12986 (N_12986,N_12612,N_12661);
xnor U12987 (N_12987,N_12632,N_12652);
and U12988 (N_12988,N_12771,N_12616);
nor U12989 (N_12989,N_12443,N_12768);
or U12990 (N_12990,N_12752,N_12488);
xor U12991 (N_12991,N_12670,N_12767);
nor U12992 (N_12992,N_12450,N_12633);
xor U12993 (N_12993,N_12622,N_12410);
or U12994 (N_12994,N_12466,N_12748);
or U12995 (N_12995,N_12698,N_12794);
or U12996 (N_12996,N_12747,N_12524);
nand U12997 (N_12997,N_12608,N_12778);
or U12998 (N_12998,N_12754,N_12526);
or U12999 (N_12999,N_12412,N_12465);
or U13000 (N_13000,N_12522,N_12771);
xor U13001 (N_13001,N_12408,N_12786);
and U13002 (N_13002,N_12469,N_12690);
nor U13003 (N_13003,N_12672,N_12500);
nand U13004 (N_13004,N_12761,N_12462);
nand U13005 (N_13005,N_12732,N_12686);
xor U13006 (N_13006,N_12658,N_12705);
or U13007 (N_13007,N_12662,N_12472);
xnor U13008 (N_13008,N_12509,N_12697);
or U13009 (N_13009,N_12622,N_12453);
xor U13010 (N_13010,N_12761,N_12570);
nor U13011 (N_13011,N_12781,N_12569);
nor U13012 (N_13012,N_12445,N_12751);
xor U13013 (N_13013,N_12487,N_12546);
nand U13014 (N_13014,N_12450,N_12512);
xor U13015 (N_13015,N_12731,N_12482);
nor U13016 (N_13016,N_12613,N_12727);
xnor U13017 (N_13017,N_12783,N_12550);
xor U13018 (N_13018,N_12769,N_12512);
xor U13019 (N_13019,N_12421,N_12734);
or U13020 (N_13020,N_12591,N_12517);
and U13021 (N_13021,N_12596,N_12465);
xnor U13022 (N_13022,N_12625,N_12513);
xor U13023 (N_13023,N_12689,N_12782);
and U13024 (N_13024,N_12606,N_12499);
nor U13025 (N_13025,N_12556,N_12509);
xnor U13026 (N_13026,N_12733,N_12671);
nor U13027 (N_13027,N_12622,N_12598);
xor U13028 (N_13028,N_12439,N_12700);
nor U13029 (N_13029,N_12552,N_12545);
xnor U13030 (N_13030,N_12470,N_12565);
or U13031 (N_13031,N_12579,N_12725);
nand U13032 (N_13032,N_12624,N_12505);
nor U13033 (N_13033,N_12592,N_12470);
nor U13034 (N_13034,N_12553,N_12525);
nand U13035 (N_13035,N_12480,N_12765);
nor U13036 (N_13036,N_12788,N_12467);
and U13037 (N_13037,N_12519,N_12457);
or U13038 (N_13038,N_12702,N_12452);
nand U13039 (N_13039,N_12544,N_12754);
nor U13040 (N_13040,N_12720,N_12514);
nand U13041 (N_13041,N_12640,N_12731);
or U13042 (N_13042,N_12627,N_12471);
or U13043 (N_13043,N_12777,N_12513);
nand U13044 (N_13044,N_12574,N_12566);
nand U13045 (N_13045,N_12439,N_12494);
and U13046 (N_13046,N_12707,N_12765);
nand U13047 (N_13047,N_12758,N_12455);
xor U13048 (N_13048,N_12596,N_12688);
and U13049 (N_13049,N_12559,N_12441);
nand U13050 (N_13050,N_12554,N_12434);
nand U13051 (N_13051,N_12404,N_12478);
xor U13052 (N_13052,N_12490,N_12788);
xor U13053 (N_13053,N_12692,N_12741);
nor U13054 (N_13054,N_12474,N_12432);
nor U13055 (N_13055,N_12747,N_12456);
or U13056 (N_13056,N_12773,N_12579);
or U13057 (N_13057,N_12551,N_12523);
and U13058 (N_13058,N_12672,N_12456);
nand U13059 (N_13059,N_12616,N_12456);
xor U13060 (N_13060,N_12569,N_12550);
and U13061 (N_13061,N_12624,N_12411);
nand U13062 (N_13062,N_12609,N_12523);
and U13063 (N_13063,N_12713,N_12434);
xor U13064 (N_13064,N_12648,N_12713);
or U13065 (N_13065,N_12634,N_12494);
or U13066 (N_13066,N_12504,N_12497);
nor U13067 (N_13067,N_12768,N_12451);
nand U13068 (N_13068,N_12668,N_12498);
and U13069 (N_13069,N_12408,N_12720);
nor U13070 (N_13070,N_12487,N_12619);
nand U13071 (N_13071,N_12412,N_12686);
xor U13072 (N_13072,N_12666,N_12692);
xnor U13073 (N_13073,N_12552,N_12773);
nor U13074 (N_13074,N_12681,N_12622);
xnor U13075 (N_13075,N_12499,N_12485);
nor U13076 (N_13076,N_12491,N_12708);
and U13077 (N_13077,N_12603,N_12479);
nand U13078 (N_13078,N_12446,N_12698);
xor U13079 (N_13079,N_12613,N_12442);
nor U13080 (N_13080,N_12571,N_12424);
and U13081 (N_13081,N_12645,N_12638);
xor U13082 (N_13082,N_12647,N_12745);
nand U13083 (N_13083,N_12715,N_12629);
and U13084 (N_13084,N_12673,N_12457);
nand U13085 (N_13085,N_12551,N_12621);
nor U13086 (N_13086,N_12434,N_12674);
and U13087 (N_13087,N_12487,N_12622);
nor U13088 (N_13088,N_12458,N_12409);
or U13089 (N_13089,N_12522,N_12442);
nand U13090 (N_13090,N_12669,N_12688);
or U13091 (N_13091,N_12401,N_12652);
nor U13092 (N_13092,N_12404,N_12603);
xor U13093 (N_13093,N_12613,N_12642);
nor U13094 (N_13094,N_12664,N_12598);
nand U13095 (N_13095,N_12653,N_12594);
and U13096 (N_13096,N_12539,N_12774);
nand U13097 (N_13097,N_12601,N_12587);
nor U13098 (N_13098,N_12714,N_12678);
nor U13099 (N_13099,N_12439,N_12707);
nand U13100 (N_13100,N_12458,N_12612);
xnor U13101 (N_13101,N_12743,N_12697);
or U13102 (N_13102,N_12596,N_12627);
xor U13103 (N_13103,N_12797,N_12576);
or U13104 (N_13104,N_12625,N_12778);
or U13105 (N_13105,N_12509,N_12637);
nor U13106 (N_13106,N_12672,N_12571);
nor U13107 (N_13107,N_12702,N_12433);
nor U13108 (N_13108,N_12564,N_12531);
and U13109 (N_13109,N_12443,N_12618);
nor U13110 (N_13110,N_12453,N_12515);
or U13111 (N_13111,N_12692,N_12634);
and U13112 (N_13112,N_12679,N_12532);
nor U13113 (N_13113,N_12629,N_12720);
or U13114 (N_13114,N_12794,N_12549);
xnor U13115 (N_13115,N_12749,N_12687);
nor U13116 (N_13116,N_12418,N_12617);
or U13117 (N_13117,N_12793,N_12609);
nand U13118 (N_13118,N_12757,N_12466);
or U13119 (N_13119,N_12579,N_12494);
or U13120 (N_13120,N_12572,N_12506);
and U13121 (N_13121,N_12530,N_12535);
nor U13122 (N_13122,N_12718,N_12776);
or U13123 (N_13123,N_12402,N_12648);
or U13124 (N_13124,N_12618,N_12600);
and U13125 (N_13125,N_12458,N_12637);
and U13126 (N_13126,N_12674,N_12528);
nor U13127 (N_13127,N_12727,N_12770);
or U13128 (N_13128,N_12779,N_12750);
xnor U13129 (N_13129,N_12418,N_12526);
and U13130 (N_13130,N_12427,N_12495);
or U13131 (N_13131,N_12738,N_12707);
nor U13132 (N_13132,N_12459,N_12761);
and U13133 (N_13133,N_12555,N_12712);
nand U13134 (N_13134,N_12789,N_12477);
nand U13135 (N_13135,N_12614,N_12667);
xor U13136 (N_13136,N_12593,N_12702);
xnor U13137 (N_13137,N_12475,N_12644);
xor U13138 (N_13138,N_12662,N_12407);
nor U13139 (N_13139,N_12717,N_12439);
xnor U13140 (N_13140,N_12475,N_12547);
nand U13141 (N_13141,N_12539,N_12451);
xor U13142 (N_13142,N_12730,N_12779);
and U13143 (N_13143,N_12614,N_12592);
and U13144 (N_13144,N_12545,N_12430);
xnor U13145 (N_13145,N_12469,N_12734);
or U13146 (N_13146,N_12580,N_12520);
nand U13147 (N_13147,N_12684,N_12740);
xor U13148 (N_13148,N_12497,N_12565);
and U13149 (N_13149,N_12511,N_12514);
and U13150 (N_13150,N_12453,N_12731);
nand U13151 (N_13151,N_12614,N_12768);
nor U13152 (N_13152,N_12636,N_12432);
nor U13153 (N_13153,N_12792,N_12461);
and U13154 (N_13154,N_12658,N_12781);
xor U13155 (N_13155,N_12611,N_12428);
and U13156 (N_13156,N_12766,N_12527);
nor U13157 (N_13157,N_12692,N_12578);
nor U13158 (N_13158,N_12470,N_12451);
nor U13159 (N_13159,N_12762,N_12405);
or U13160 (N_13160,N_12780,N_12445);
and U13161 (N_13161,N_12433,N_12559);
nor U13162 (N_13162,N_12606,N_12644);
nor U13163 (N_13163,N_12587,N_12460);
xnor U13164 (N_13164,N_12461,N_12529);
or U13165 (N_13165,N_12740,N_12512);
or U13166 (N_13166,N_12530,N_12718);
or U13167 (N_13167,N_12538,N_12674);
nor U13168 (N_13168,N_12720,N_12667);
and U13169 (N_13169,N_12494,N_12703);
and U13170 (N_13170,N_12526,N_12417);
xnor U13171 (N_13171,N_12739,N_12612);
or U13172 (N_13172,N_12716,N_12417);
nor U13173 (N_13173,N_12646,N_12423);
xor U13174 (N_13174,N_12604,N_12704);
nand U13175 (N_13175,N_12543,N_12593);
nor U13176 (N_13176,N_12534,N_12758);
nor U13177 (N_13177,N_12607,N_12611);
xnor U13178 (N_13178,N_12784,N_12492);
nand U13179 (N_13179,N_12491,N_12593);
xnor U13180 (N_13180,N_12535,N_12450);
or U13181 (N_13181,N_12639,N_12703);
and U13182 (N_13182,N_12659,N_12663);
nand U13183 (N_13183,N_12707,N_12762);
nor U13184 (N_13184,N_12578,N_12671);
xnor U13185 (N_13185,N_12469,N_12521);
xor U13186 (N_13186,N_12796,N_12408);
or U13187 (N_13187,N_12569,N_12646);
and U13188 (N_13188,N_12789,N_12558);
xor U13189 (N_13189,N_12427,N_12675);
and U13190 (N_13190,N_12453,N_12774);
and U13191 (N_13191,N_12789,N_12740);
nand U13192 (N_13192,N_12619,N_12759);
xor U13193 (N_13193,N_12619,N_12723);
nor U13194 (N_13194,N_12636,N_12585);
nand U13195 (N_13195,N_12594,N_12752);
or U13196 (N_13196,N_12657,N_12736);
and U13197 (N_13197,N_12448,N_12635);
or U13198 (N_13198,N_12774,N_12504);
or U13199 (N_13199,N_12663,N_12749);
and U13200 (N_13200,N_12828,N_13090);
nand U13201 (N_13201,N_12946,N_12903);
nor U13202 (N_13202,N_13089,N_12809);
xnor U13203 (N_13203,N_13142,N_12922);
and U13204 (N_13204,N_12837,N_13026);
or U13205 (N_13205,N_13047,N_13073);
nor U13206 (N_13206,N_12917,N_12910);
and U13207 (N_13207,N_12921,N_13196);
and U13208 (N_13208,N_13034,N_13116);
nor U13209 (N_13209,N_13160,N_12934);
nand U13210 (N_13210,N_12938,N_12931);
nor U13211 (N_13211,N_12945,N_12930);
and U13212 (N_13212,N_12865,N_12973);
nor U13213 (N_13213,N_13003,N_12836);
and U13214 (N_13214,N_12825,N_12804);
xor U13215 (N_13215,N_13053,N_13050);
nand U13216 (N_13216,N_12982,N_13017);
and U13217 (N_13217,N_12887,N_13146);
nor U13218 (N_13218,N_13183,N_13173);
nor U13219 (N_13219,N_12966,N_13113);
xnor U13220 (N_13220,N_12877,N_13145);
xor U13221 (N_13221,N_12901,N_13054);
xor U13222 (N_13222,N_12944,N_13038);
and U13223 (N_13223,N_12974,N_12801);
and U13224 (N_13224,N_13152,N_13141);
nor U13225 (N_13225,N_12972,N_13168);
xnor U13226 (N_13226,N_13013,N_13198);
nand U13227 (N_13227,N_13129,N_12895);
and U13228 (N_13228,N_13051,N_12948);
nor U13229 (N_13229,N_12950,N_13179);
nor U13230 (N_13230,N_13134,N_13072);
xnor U13231 (N_13231,N_12955,N_12826);
nor U13232 (N_13232,N_13043,N_13192);
or U13233 (N_13233,N_13078,N_12847);
nor U13234 (N_13234,N_12981,N_13062);
nand U13235 (N_13235,N_12858,N_13005);
and U13236 (N_13236,N_13185,N_13060);
or U13237 (N_13237,N_12889,N_12928);
nor U13238 (N_13238,N_12841,N_12811);
or U13239 (N_13239,N_13040,N_12983);
nor U13240 (N_13240,N_13092,N_13166);
nand U13241 (N_13241,N_12853,N_12833);
nor U13242 (N_13242,N_12961,N_13197);
nand U13243 (N_13243,N_12845,N_12834);
xnor U13244 (N_13244,N_13044,N_12846);
and U13245 (N_13245,N_12879,N_12906);
and U13246 (N_13246,N_12997,N_13079);
and U13247 (N_13247,N_13021,N_13112);
and U13248 (N_13248,N_12940,N_12912);
nor U13249 (N_13249,N_12868,N_12867);
nor U13250 (N_13250,N_12820,N_12898);
and U13251 (N_13251,N_13107,N_13023);
or U13252 (N_13252,N_13057,N_13189);
or U13253 (N_13253,N_13187,N_12990);
xnor U13254 (N_13254,N_13071,N_12883);
xnor U13255 (N_13255,N_13042,N_13161);
xnor U13256 (N_13256,N_13188,N_13110);
xor U13257 (N_13257,N_13065,N_13132);
nor U13258 (N_13258,N_12861,N_12908);
nand U13259 (N_13259,N_13122,N_12829);
nor U13260 (N_13260,N_13037,N_12823);
xnor U13261 (N_13261,N_13104,N_12992);
nand U13262 (N_13262,N_12943,N_12999);
xor U13263 (N_13263,N_12806,N_13182);
or U13264 (N_13264,N_12919,N_12905);
xor U13265 (N_13265,N_13033,N_12953);
or U13266 (N_13266,N_13036,N_13027);
and U13267 (N_13267,N_13158,N_13138);
or U13268 (N_13268,N_13130,N_12960);
nor U13269 (N_13269,N_13151,N_13119);
xnor U13270 (N_13270,N_12862,N_12936);
nand U13271 (N_13271,N_13140,N_13084);
nor U13272 (N_13272,N_12863,N_12860);
or U13273 (N_13273,N_12838,N_13105);
nand U13274 (N_13274,N_12880,N_12888);
nand U13275 (N_13275,N_12967,N_12812);
nor U13276 (N_13276,N_13020,N_13157);
and U13277 (N_13277,N_13070,N_12968);
or U13278 (N_13278,N_13127,N_13147);
and U13279 (N_13279,N_13063,N_12926);
xor U13280 (N_13280,N_13099,N_13039);
nand U13281 (N_13281,N_13135,N_13010);
nand U13282 (N_13282,N_13056,N_13093);
nand U13283 (N_13283,N_13159,N_12832);
and U13284 (N_13284,N_13153,N_13199);
or U13285 (N_13285,N_13114,N_12890);
and U13286 (N_13286,N_12991,N_13004);
nand U13287 (N_13287,N_13195,N_12927);
xor U13288 (N_13288,N_13048,N_12881);
nand U13289 (N_13289,N_12870,N_12979);
and U13290 (N_13290,N_13067,N_13006);
nand U13291 (N_13291,N_13111,N_13095);
xnor U13292 (N_13292,N_13131,N_13186);
nand U13293 (N_13293,N_12929,N_12909);
xnor U13294 (N_13294,N_12850,N_12977);
nand U13295 (N_13295,N_12987,N_12876);
xor U13296 (N_13296,N_12873,N_12884);
nor U13297 (N_13297,N_12859,N_12819);
nand U13298 (N_13298,N_12869,N_13069);
xnor U13299 (N_13299,N_12989,N_13046);
xor U13300 (N_13300,N_12904,N_12965);
nand U13301 (N_13301,N_13167,N_12937);
xor U13302 (N_13302,N_13088,N_13029);
or U13303 (N_13303,N_13103,N_13101);
nor U13304 (N_13304,N_13156,N_12822);
nand U13305 (N_13305,N_12815,N_12800);
nor U13306 (N_13306,N_13175,N_13143);
and U13307 (N_13307,N_12896,N_13125);
xor U13308 (N_13308,N_13117,N_13162);
nor U13309 (N_13309,N_13180,N_13155);
and U13310 (N_13310,N_13016,N_13066);
nand U13311 (N_13311,N_12963,N_12954);
nor U13312 (N_13312,N_13087,N_12856);
nand U13313 (N_13313,N_13121,N_13124);
and U13314 (N_13314,N_13106,N_12851);
or U13315 (N_13315,N_12939,N_13091);
nand U13316 (N_13316,N_13030,N_13190);
or U13317 (N_13317,N_13120,N_12996);
nor U13318 (N_13318,N_13058,N_13194);
and U13319 (N_13319,N_13149,N_12818);
or U13320 (N_13320,N_12994,N_13181);
or U13321 (N_13321,N_12803,N_13144);
nor U13322 (N_13322,N_12897,N_13000);
nand U13323 (N_13323,N_13012,N_13059);
xnor U13324 (N_13324,N_13028,N_12843);
or U13325 (N_13325,N_12902,N_13064);
nand U13326 (N_13326,N_12915,N_12805);
nor U13327 (N_13327,N_13068,N_12933);
or U13328 (N_13328,N_13024,N_12857);
nand U13329 (N_13329,N_13025,N_13137);
or U13330 (N_13330,N_13102,N_13018);
nand U13331 (N_13331,N_12891,N_12894);
xor U13332 (N_13332,N_13154,N_12925);
nand U13333 (N_13333,N_12947,N_13108);
nand U13334 (N_13334,N_12932,N_13061);
xnor U13335 (N_13335,N_12866,N_13126);
and U13336 (N_13336,N_12882,N_12830);
nor U13337 (N_13337,N_13001,N_12924);
xnor U13338 (N_13338,N_12913,N_13193);
and U13339 (N_13339,N_12802,N_12985);
and U13340 (N_13340,N_13019,N_12864);
nor U13341 (N_13341,N_12824,N_12813);
or U13342 (N_13342,N_12885,N_13080);
and U13343 (N_13343,N_13177,N_12918);
and U13344 (N_13344,N_12831,N_12976);
or U13345 (N_13345,N_13032,N_13164);
or U13346 (N_13346,N_13052,N_12911);
or U13347 (N_13347,N_13083,N_13074);
xor U13348 (N_13348,N_12808,N_13165);
and U13349 (N_13349,N_12842,N_12920);
nor U13350 (N_13350,N_13148,N_12923);
nand U13351 (N_13351,N_12814,N_12949);
or U13352 (N_13352,N_12935,N_12962);
nor U13353 (N_13353,N_12986,N_13076);
or U13354 (N_13354,N_12871,N_13171);
and U13355 (N_13355,N_12874,N_13176);
or U13356 (N_13356,N_13085,N_12964);
nor U13357 (N_13357,N_12956,N_12951);
nand U13358 (N_13358,N_13008,N_12816);
nor U13359 (N_13359,N_12899,N_12839);
nand U13360 (N_13360,N_13100,N_13150);
xor U13361 (N_13361,N_12840,N_12852);
or U13362 (N_13362,N_13115,N_13049);
or U13363 (N_13363,N_12907,N_13077);
and U13364 (N_13364,N_12886,N_13174);
and U13365 (N_13365,N_12978,N_13045);
nor U13366 (N_13366,N_13022,N_12941);
nand U13367 (N_13367,N_13097,N_12952);
and U13368 (N_13368,N_12854,N_13094);
and U13369 (N_13369,N_12959,N_13014);
and U13370 (N_13370,N_13082,N_12892);
nor U13371 (N_13371,N_13031,N_13002);
xnor U13372 (N_13372,N_13011,N_13139);
xnor U13373 (N_13373,N_13184,N_12875);
nor U13374 (N_13374,N_13118,N_13086);
and U13375 (N_13375,N_12835,N_13191);
xor U13376 (N_13376,N_12984,N_13172);
or U13377 (N_13377,N_12998,N_13055);
nand U13378 (N_13378,N_12980,N_12995);
nor U13379 (N_13379,N_12942,N_12810);
nand U13380 (N_13380,N_12807,N_12821);
or U13381 (N_13381,N_12849,N_12916);
nand U13382 (N_13382,N_13009,N_13015);
xor U13383 (N_13383,N_12817,N_13081);
and U13384 (N_13384,N_13136,N_12878);
nor U13385 (N_13385,N_12975,N_13123);
or U13386 (N_13386,N_12844,N_12914);
and U13387 (N_13387,N_13128,N_13178);
and U13388 (N_13388,N_12971,N_12957);
nor U13389 (N_13389,N_12855,N_13109);
xor U13390 (N_13390,N_13075,N_13133);
or U13391 (N_13391,N_12970,N_13007);
nand U13392 (N_13392,N_12993,N_13169);
or U13393 (N_13393,N_13163,N_12893);
nor U13394 (N_13394,N_13170,N_12827);
nand U13395 (N_13395,N_13098,N_12988);
xnor U13396 (N_13396,N_13041,N_13096);
nand U13397 (N_13397,N_13035,N_12848);
or U13398 (N_13398,N_12958,N_12900);
xor U13399 (N_13399,N_12969,N_12872);
xnor U13400 (N_13400,N_13034,N_13062);
xnor U13401 (N_13401,N_12944,N_13004);
nor U13402 (N_13402,N_13046,N_12906);
nand U13403 (N_13403,N_12925,N_13027);
or U13404 (N_13404,N_12951,N_13181);
and U13405 (N_13405,N_12824,N_12847);
nor U13406 (N_13406,N_12852,N_13056);
and U13407 (N_13407,N_12850,N_12980);
and U13408 (N_13408,N_13179,N_12916);
xor U13409 (N_13409,N_13142,N_12854);
or U13410 (N_13410,N_12978,N_13055);
nand U13411 (N_13411,N_13129,N_12880);
nand U13412 (N_13412,N_12885,N_12966);
and U13413 (N_13413,N_13075,N_13172);
and U13414 (N_13414,N_12875,N_13146);
nand U13415 (N_13415,N_13008,N_13059);
nand U13416 (N_13416,N_13119,N_13106);
and U13417 (N_13417,N_13099,N_12991);
nand U13418 (N_13418,N_13143,N_12969);
xnor U13419 (N_13419,N_13110,N_13105);
and U13420 (N_13420,N_12976,N_13108);
and U13421 (N_13421,N_12875,N_13106);
nand U13422 (N_13422,N_13163,N_13143);
and U13423 (N_13423,N_13180,N_12912);
nand U13424 (N_13424,N_13169,N_12864);
or U13425 (N_13425,N_12808,N_12878);
or U13426 (N_13426,N_13125,N_13073);
xnor U13427 (N_13427,N_12908,N_12870);
and U13428 (N_13428,N_13035,N_12983);
and U13429 (N_13429,N_13163,N_13022);
xnor U13430 (N_13430,N_13065,N_12927);
or U13431 (N_13431,N_13187,N_12912);
and U13432 (N_13432,N_12857,N_13129);
nor U13433 (N_13433,N_12800,N_13095);
or U13434 (N_13434,N_13144,N_13044);
and U13435 (N_13435,N_12808,N_12912);
nor U13436 (N_13436,N_13123,N_13006);
nor U13437 (N_13437,N_13154,N_13020);
or U13438 (N_13438,N_13086,N_12863);
xor U13439 (N_13439,N_12910,N_12982);
or U13440 (N_13440,N_12995,N_12937);
nand U13441 (N_13441,N_12987,N_13061);
and U13442 (N_13442,N_13052,N_12879);
nand U13443 (N_13443,N_12945,N_12995);
xnor U13444 (N_13444,N_12975,N_13167);
or U13445 (N_13445,N_13148,N_12893);
xnor U13446 (N_13446,N_13004,N_12934);
and U13447 (N_13447,N_12993,N_12991);
xnor U13448 (N_13448,N_12980,N_12883);
nor U13449 (N_13449,N_13071,N_13188);
xnor U13450 (N_13450,N_12933,N_13187);
nand U13451 (N_13451,N_12857,N_12942);
or U13452 (N_13452,N_13190,N_13090);
and U13453 (N_13453,N_12929,N_12932);
nand U13454 (N_13454,N_12975,N_12888);
and U13455 (N_13455,N_12988,N_13018);
xnor U13456 (N_13456,N_13071,N_13148);
nor U13457 (N_13457,N_12868,N_12971);
nor U13458 (N_13458,N_13119,N_13080);
nor U13459 (N_13459,N_13011,N_12923);
nor U13460 (N_13460,N_12919,N_12877);
nand U13461 (N_13461,N_12884,N_13100);
nor U13462 (N_13462,N_13141,N_12860);
xnor U13463 (N_13463,N_12847,N_13010);
nand U13464 (N_13464,N_12984,N_13035);
nand U13465 (N_13465,N_13024,N_12897);
or U13466 (N_13466,N_13087,N_12984);
or U13467 (N_13467,N_12825,N_12990);
xor U13468 (N_13468,N_12850,N_12928);
xnor U13469 (N_13469,N_12919,N_12939);
xor U13470 (N_13470,N_13069,N_13035);
and U13471 (N_13471,N_13156,N_12848);
or U13472 (N_13472,N_12939,N_12955);
nor U13473 (N_13473,N_13054,N_13138);
nor U13474 (N_13474,N_12984,N_12853);
nand U13475 (N_13475,N_12956,N_12918);
nor U13476 (N_13476,N_13113,N_13124);
nand U13477 (N_13477,N_12879,N_12856);
xor U13478 (N_13478,N_13121,N_13166);
nor U13479 (N_13479,N_12887,N_13132);
nor U13480 (N_13480,N_13168,N_12934);
nand U13481 (N_13481,N_13105,N_13102);
nand U13482 (N_13482,N_12902,N_13198);
nor U13483 (N_13483,N_13127,N_13068);
and U13484 (N_13484,N_13120,N_13083);
nand U13485 (N_13485,N_12836,N_13124);
nor U13486 (N_13486,N_12920,N_13097);
nand U13487 (N_13487,N_12915,N_12862);
nand U13488 (N_13488,N_12889,N_12971);
nand U13489 (N_13489,N_13096,N_13135);
xnor U13490 (N_13490,N_13054,N_12879);
or U13491 (N_13491,N_12863,N_13096);
xnor U13492 (N_13492,N_12847,N_13138);
or U13493 (N_13493,N_12851,N_12859);
nand U13494 (N_13494,N_13029,N_12886);
or U13495 (N_13495,N_12993,N_12807);
or U13496 (N_13496,N_12976,N_12911);
nor U13497 (N_13497,N_13111,N_13015);
xor U13498 (N_13498,N_13031,N_13185);
nand U13499 (N_13499,N_12896,N_12894);
nor U13500 (N_13500,N_13179,N_12993);
xnor U13501 (N_13501,N_13114,N_13177);
nand U13502 (N_13502,N_12949,N_13047);
and U13503 (N_13503,N_12805,N_13019);
and U13504 (N_13504,N_12821,N_12866);
or U13505 (N_13505,N_12908,N_13012);
or U13506 (N_13506,N_12948,N_13071);
nand U13507 (N_13507,N_12974,N_12868);
or U13508 (N_13508,N_12908,N_12845);
and U13509 (N_13509,N_13027,N_12908);
nand U13510 (N_13510,N_13000,N_12987);
xnor U13511 (N_13511,N_13143,N_12960);
or U13512 (N_13512,N_13037,N_13079);
nor U13513 (N_13513,N_12962,N_13122);
nor U13514 (N_13514,N_13048,N_12827);
and U13515 (N_13515,N_12996,N_12964);
nor U13516 (N_13516,N_13009,N_13024);
nor U13517 (N_13517,N_13175,N_13026);
or U13518 (N_13518,N_12884,N_12889);
xor U13519 (N_13519,N_13112,N_13014);
or U13520 (N_13520,N_12897,N_13156);
or U13521 (N_13521,N_13125,N_12830);
xnor U13522 (N_13522,N_12952,N_12964);
and U13523 (N_13523,N_13128,N_12933);
nor U13524 (N_13524,N_13133,N_13115);
or U13525 (N_13525,N_13032,N_12977);
or U13526 (N_13526,N_13141,N_13083);
nor U13527 (N_13527,N_12831,N_13141);
nor U13528 (N_13528,N_12970,N_13135);
or U13529 (N_13529,N_13169,N_12963);
xor U13530 (N_13530,N_13121,N_13030);
xnor U13531 (N_13531,N_12991,N_13038);
nand U13532 (N_13532,N_13076,N_13165);
or U13533 (N_13533,N_12843,N_13034);
nor U13534 (N_13534,N_12831,N_12844);
nor U13535 (N_13535,N_13021,N_13152);
or U13536 (N_13536,N_13085,N_12925);
xor U13537 (N_13537,N_13135,N_13015);
or U13538 (N_13538,N_12962,N_12910);
nor U13539 (N_13539,N_13024,N_12834);
xor U13540 (N_13540,N_13139,N_13095);
or U13541 (N_13541,N_12829,N_12897);
nand U13542 (N_13542,N_12858,N_12965);
xnor U13543 (N_13543,N_13075,N_12882);
nand U13544 (N_13544,N_12964,N_13027);
nand U13545 (N_13545,N_12953,N_12956);
xor U13546 (N_13546,N_13012,N_12997);
nor U13547 (N_13547,N_12823,N_12923);
or U13548 (N_13548,N_13111,N_12886);
nor U13549 (N_13549,N_12939,N_12935);
nor U13550 (N_13550,N_13003,N_12983);
xor U13551 (N_13551,N_12853,N_12930);
nor U13552 (N_13552,N_12846,N_12855);
nor U13553 (N_13553,N_13175,N_12925);
or U13554 (N_13554,N_12883,N_12852);
xnor U13555 (N_13555,N_13003,N_12843);
or U13556 (N_13556,N_12842,N_13144);
and U13557 (N_13557,N_13107,N_12854);
or U13558 (N_13558,N_13141,N_12937);
nor U13559 (N_13559,N_13069,N_12957);
xnor U13560 (N_13560,N_13132,N_13098);
nor U13561 (N_13561,N_13013,N_13126);
xor U13562 (N_13562,N_12826,N_13171);
xnor U13563 (N_13563,N_12850,N_12983);
and U13564 (N_13564,N_12855,N_13086);
nor U13565 (N_13565,N_13053,N_13006);
xnor U13566 (N_13566,N_13007,N_13072);
or U13567 (N_13567,N_13050,N_13095);
or U13568 (N_13568,N_13121,N_12871);
and U13569 (N_13569,N_12999,N_12985);
nand U13570 (N_13570,N_13091,N_12857);
nor U13571 (N_13571,N_13187,N_12817);
or U13572 (N_13572,N_12837,N_12931);
nand U13573 (N_13573,N_12883,N_13035);
nand U13574 (N_13574,N_13047,N_13042);
xnor U13575 (N_13575,N_13091,N_13086);
and U13576 (N_13576,N_12861,N_13049);
and U13577 (N_13577,N_12923,N_13193);
or U13578 (N_13578,N_13105,N_12835);
nand U13579 (N_13579,N_12855,N_12838);
xor U13580 (N_13580,N_12812,N_13097);
and U13581 (N_13581,N_13011,N_13167);
and U13582 (N_13582,N_13055,N_13069);
nor U13583 (N_13583,N_12883,N_13025);
or U13584 (N_13584,N_13055,N_12916);
xor U13585 (N_13585,N_13136,N_13189);
nand U13586 (N_13586,N_12875,N_13162);
nor U13587 (N_13587,N_13187,N_13000);
nand U13588 (N_13588,N_12975,N_13126);
and U13589 (N_13589,N_12877,N_13065);
nand U13590 (N_13590,N_13118,N_12818);
nor U13591 (N_13591,N_13154,N_12876);
nor U13592 (N_13592,N_12871,N_13127);
nor U13593 (N_13593,N_13053,N_13103);
nand U13594 (N_13594,N_13130,N_13190);
or U13595 (N_13595,N_12988,N_12956);
and U13596 (N_13596,N_12817,N_12883);
xor U13597 (N_13597,N_12846,N_12946);
nand U13598 (N_13598,N_12813,N_12815);
and U13599 (N_13599,N_12910,N_13025);
nor U13600 (N_13600,N_13413,N_13339);
nand U13601 (N_13601,N_13430,N_13565);
and U13602 (N_13602,N_13563,N_13543);
or U13603 (N_13603,N_13441,N_13364);
nand U13604 (N_13604,N_13418,N_13366);
nand U13605 (N_13605,N_13511,N_13204);
nor U13606 (N_13606,N_13229,N_13479);
nor U13607 (N_13607,N_13362,N_13289);
nand U13608 (N_13608,N_13460,N_13560);
or U13609 (N_13609,N_13461,N_13412);
or U13610 (N_13610,N_13395,N_13286);
nor U13611 (N_13611,N_13564,N_13228);
and U13612 (N_13612,N_13530,N_13219);
and U13613 (N_13613,N_13213,N_13275);
nand U13614 (N_13614,N_13284,N_13436);
xnor U13615 (N_13615,N_13209,N_13405);
or U13616 (N_13616,N_13313,N_13583);
nor U13617 (N_13617,N_13484,N_13205);
xor U13618 (N_13618,N_13216,N_13473);
nand U13619 (N_13619,N_13534,N_13510);
and U13620 (N_13620,N_13292,N_13337);
nor U13621 (N_13621,N_13212,N_13300);
nor U13622 (N_13622,N_13513,N_13307);
xnor U13623 (N_13623,N_13450,N_13537);
xor U13624 (N_13624,N_13231,N_13222);
and U13625 (N_13625,N_13414,N_13569);
xnor U13626 (N_13626,N_13294,N_13252);
or U13627 (N_13627,N_13211,N_13482);
nand U13628 (N_13628,N_13454,N_13278);
and U13629 (N_13629,N_13262,N_13535);
xor U13630 (N_13630,N_13524,N_13580);
nor U13631 (N_13631,N_13378,N_13576);
and U13632 (N_13632,N_13380,N_13253);
xnor U13633 (N_13633,N_13235,N_13372);
nor U13634 (N_13634,N_13499,N_13221);
xnor U13635 (N_13635,N_13588,N_13434);
nor U13636 (N_13636,N_13207,N_13467);
or U13637 (N_13637,N_13203,N_13483);
and U13638 (N_13638,N_13308,N_13587);
and U13639 (N_13639,N_13383,N_13266);
or U13640 (N_13640,N_13363,N_13554);
nand U13641 (N_13641,N_13239,N_13352);
nor U13642 (N_13642,N_13310,N_13287);
nor U13643 (N_13643,N_13448,N_13476);
xor U13644 (N_13644,N_13485,N_13265);
or U13645 (N_13645,N_13516,N_13474);
nor U13646 (N_13646,N_13403,N_13542);
nor U13647 (N_13647,N_13517,N_13399);
xnor U13648 (N_13648,N_13246,N_13504);
xnor U13649 (N_13649,N_13404,N_13206);
nor U13650 (N_13650,N_13311,N_13387);
nand U13651 (N_13651,N_13316,N_13407);
or U13652 (N_13652,N_13477,N_13301);
xor U13653 (N_13653,N_13263,N_13274);
xor U13654 (N_13654,N_13438,N_13507);
xnor U13655 (N_13655,N_13324,N_13547);
nor U13656 (N_13656,N_13200,N_13243);
or U13657 (N_13657,N_13329,N_13567);
and U13658 (N_13658,N_13515,N_13536);
xor U13659 (N_13659,N_13401,N_13549);
nor U13660 (N_13660,N_13502,N_13561);
and U13661 (N_13661,N_13323,N_13346);
nand U13662 (N_13662,N_13505,N_13487);
xor U13663 (N_13663,N_13533,N_13402);
or U13664 (N_13664,N_13259,N_13334);
and U13665 (N_13665,N_13356,N_13280);
nor U13666 (N_13666,N_13371,N_13432);
or U13667 (N_13667,N_13489,N_13447);
or U13668 (N_13668,N_13330,N_13331);
nor U13669 (N_13669,N_13336,N_13443);
and U13670 (N_13670,N_13445,N_13390);
and U13671 (N_13671,N_13251,N_13288);
and U13672 (N_13672,N_13540,N_13321);
nand U13673 (N_13673,N_13410,N_13349);
or U13674 (N_13674,N_13492,N_13462);
nor U13675 (N_13675,N_13315,N_13271);
nand U13676 (N_13676,N_13224,N_13250);
nor U13677 (N_13677,N_13532,N_13437);
nor U13678 (N_13678,N_13365,N_13320);
or U13679 (N_13679,N_13539,N_13545);
xnor U13680 (N_13680,N_13225,N_13348);
or U13681 (N_13681,N_13506,N_13431);
nor U13682 (N_13682,N_13248,N_13258);
or U13683 (N_13683,N_13455,N_13202);
and U13684 (N_13684,N_13305,N_13503);
xor U13685 (N_13685,N_13464,N_13465);
xor U13686 (N_13686,N_13242,N_13245);
or U13687 (N_13687,N_13234,N_13261);
nor U13688 (N_13688,N_13572,N_13354);
and U13689 (N_13689,N_13327,N_13550);
and U13690 (N_13690,N_13574,N_13217);
or U13691 (N_13691,N_13514,N_13367);
nand U13692 (N_13692,N_13230,N_13398);
xnor U13693 (N_13693,N_13531,N_13306);
nand U13694 (N_13694,N_13433,N_13406);
and U13695 (N_13695,N_13598,N_13309);
or U13696 (N_13696,N_13451,N_13472);
nor U13697 (N_13697,N_13596,N_13281);
and U13698 (N_13698,N_13589,N_13595);
xnor U13699 (N_13699,N_13557,N_13385);
or U13700 (N_13700,N_13422,N_13298);
xnor U13701 (N_13701,N_13525,N_13397);
and U13702 (N_13702,N_13335,N_13201);
xor U13703 (N_13703,N_13495,N_13396);
nand U13704 (N_13704,N_13421,N_13297);
nor U13705 (N_13705,N_13386,N_13457);
xor U13706 (N_13706,N_13355,N_13254);
or U13707 (N_13707,N_13586,N_13490);
and U13708 (N_13708,N_13359,N_13255);
and U13709 (N_13709,N_13351,N_13446);
xor U13710 (N_13710,N_13344,N_13326);
or U13711 (N_13711,N_13444,N_13353);
or U13712 (N_13712,N_13293,N_13568);
and U13713 (N_13713,N_13374,N_13345);
or U13714 (N_13714,N_13585,N_13541);
nand U13715 (N_13715,N_13481,N_13459);
xor U13716 (N_13716,N_13578,N_13361);
and U13717 (N_13717,N_13456,N_13290);
nor U13718 (N_13718,N_13343,N_13424);
xnor U13719 (N_13719,N_13478,N_13594);
nand U13720 (N_13720,N_13333,N_13220);
xor U13721 (N_13721,N_13597,N_13392);
xor U13722 (N_13722,N_13579,N_13419);
nor U13723 (N_13723,N_13295,N_13526);
xor U13724 (N_13724,N_13332,N_13268);
nand U13725 (N_13725,N_13318,N_13591);
and U13726 (N_13726,N_13282,N_13210);
nor U13727 (N_13727,N_13599,N_13249);
and U13728 (N_13728,N_13475,N_13411);
or U13729 (N_13729,N_13256,N_13304);
nor U13730 (N_13730,N_13529,N_13555);
or U13731 (N_13731,N_13581,N_13575);
xnor U13732 (N_13732,N_13237,N_13215);
nand U13733 (N_13733,N_13512,N_13496);
or U13734 (N_13734,N_13379,N_13571);
xor U13735 (N_13735,N_13466,N_13494);
nand U13736 (N_13736,N_13223,N_13238);
xor U13737 (N_13737,N_13538,N_13415);
and U13738 (N_13738,N_13241,N_13573);
xnor U13739 (N_13739,N_13393,N_13470);
and U13740 (N_13740,N_13592,N_13435);
nand U13741 (N_13741,N_13214,N_13528);
xnor U13742 (N_13742,N_13527,N_13376);
nand U13743 (N_13743,N_13232,N_13391);
and U13744 (N_13744,N_13508,N_13291);
and U13745 (N_13745,N_13553,N_13208);
and U13746 (N_13746,N_13244,N_13226);
nor U13747 (N_13747,N_13381,N_13570);
and U13748 (N_13748,N_13400,N_13509);
or U13749 (N_13749,N_13272,N_13270);
nor U13750 (N_13750,N_13340,N_13522);
nand U13751 (N_13751,N_13427,N_13236);
or U13752 (N_13752,N_13350,N_13521);
xor U13753 (N_13753,N_13471,N_13314);
nand U13754 (N_13754,N_13590,N_13468);
xor U13755 (N_13755,N_13518,N_13267);
nand U13756 (N_13756,N_13500,N_13369);
or U13757 (N_13757,N_13269,N_13317);
nand U13758 (N_13758,N_13375,N_13382);
xnor U13759 (N_13759,N_13544,N_13368);
and U13760 (N_13760,N_13417,N_13370);
and U13761 (N_13761,N_13491,N_13312);
or U13762 (N_13762,N_13338,N_13260);
or U13763 (N_13763,N_13240,N_13373);
xnor U13764 (N_13764,N_13322,N_13426);
xor U13765 (N_13765,N_13452,N_13389);
and U13766 (N_13766,N_13501,N_13552);
nand U13767 (N_13767,N_13388,N_13342);
and U13768 (N_13768,N_13486,N_13546);
or U13769 (N_13769,N_13299,N_13227);
nand U13770 (N_13770,N_13562,N_13384);
xnor U13771 (N_13771,N_13328,N_13325);
xnor U13772 (N_13772,N_13360,N_13439);
nand U13773 (N_13773,N_13264,N_13520);
nand U13774 (N_13774,N_13469,N_13449);
nand U13775 (N_13775,N_13218,N_13303);
xnor U13776 (N_13776,N_13302,N_13558);
nand U13777 (N_13777,N_13493,N_13556);
or U13778 (N_13778,N_13425,N_13285);
or U13779 (N_13779,N_13488,N_13428);
and U13780 (N_13780,N_13551,N_13423);
nor U13781 (N_13781,N_13440,N_13420);
or U13782 (N_13782,N_13408,N_13416);
nor U13783 (N_13783,N_13283,N_13233);
xor U13784 (N_13784,N_13442,N_13347);
and U13785 (N_13785,N_13519,N_13341);
nor U13786 (N_13786,N_13394,N_13498);
and U13787 (N_13787,N_13276,N_13577);
and U13788 (N_13788,N_13463,N_13480);
nor U13789 (N_13789,N_13593,N_13458);
nand U13790 (N_13790,N_13257,N_13357);
or U13791 (N_13791,N_13279,N_13319);
or U13792 (N_13792,N_13559,N_13277);
or U13793 (N_13793,N_13566,N_13296);
and U13794 (N_13794,N_13523,N_13582);
xor U13795 (N_13795,N_13247,N_13377);
nor U13796 (N_13796,N_13358,N_13584);
and U13797 (N_13797,N_13497,N_13273);
nand U13798 (N_13798,N_13409,N_13429);
nand U13799 (N_13799,N_13548,N_13453);
or U13800 (N_13800,N_13258,N_13582);
nand U13801 (N_13801,N_13288,N_13212);
nand U13802 (N_13802,N_13335,N_13326);
xnor U13803 (N_13803,N_13550,N_13383);
xnor U13804 (N_13804,N_13245,N_13459);
xnor U13805 (N_13805,N_13356,N_13586);
and U13806 (N_13806,N_13201,N_13472);
and U13807 (N_13807,N_13351,N_13584);
and U13808 (N_13808,N_13387,N_13358);
nand U13809 (N_13809,N_13346,N_13514);
xnor U13810 (N_13810,N_13404,N_13454);
or U13811 (N_13811,N_13501,N_13491);
nor U13812 (N_13812,N_13311,N_13505);
and U13813 (N_13813,N_13229,N_13316);
and U13814 (N_13814,N_13294,N_13505);
xnor U13815 (N_13815,N_13465,N_13302);
xnor U13816 (N_13816,N_13318,N_13352);
nor U13817 (N_13817,N_13414,N_13206);
nor U13818 (N_13818,N_13571,N_13499);
nor U13819 (N_13819,N_13452,N_13481);
nand U13820 (N_13820,N_13269,N_13508);
and U13821 (N_13821,N_13528,N_13304);
nand U13822 (N_13822,N_13363,N_13525);
and U13823 (N_13823,N_13385,N_13575);
xor U13824 (N_13824,N_13323,N_13529);
xor U13825 (N_13825,N_13242,N_13539);
nand U13826 (N_13826,N_13433,N_13329);
or U13827 (N_13827,N_13564,N_13408);
nand U13828 (N_13828,N_13442,N_13252);
nor U13829 (N_13829,N_13395,N_13536);
nor U13830 (N_13830,N_13503,N_13378);
xnor U13831 (N_13831,N_13218,N_13296);
or U13832 (N_13832,N_13578,N_13287);
nor U13833 (N_13833,N_13248,N_13505);
nand U13834 (N_13834,N_13406,N_13252);
nand U13835 (N_13835,N_13485,N_13501);
or U13836 (N_13836,N_13473,N_13434);
nor U13837 (N_13837,N_13331,N_13254);
nand U13838 (N_13838,N_13482,N_13479);
and U13839 (N_13839,N_13347,N_13395);
or U13840 (N_13840,N_13221,N_13470);
xnor U13841 (N_13841,N_13238,N_13443);
nor U13842 (N_13842,N_13202,N_13237);
and U13843 (N_13843,N_13369,N_13537);
nand U13844 (N_13844,N_13527,N_13334);
nand U13845 (N_13845,N_13304,N_13290);
xnor U13846 (N_13846,N_13333,N_13247);
nor U13847 (N_13847,N_13344,N_13590);
or U13848 (N_13848,N_13325,N_13413);
nor U13849 (N_13849,N_13507,N_13574);
xnor U13850 (N_13850,N_13309,N_13483);
nand U13851 (N_13851,N_13422,N_13567);
xor U13852 (N_13852,N_13487,N_13545);
nor U13853 (N_13853,N_13455,N_13569);
or U13854 (N_13854,N_13584,N_13308);
xnor U13855 (N_13855,N_13584,N_13480);
or U13856 (N_13856,N_13534,N_13348);
or U13857 (N_13857,N_13384,N_13396);
and U13858 (N_13858,N_13389,N_13400);
xnor U13859 (N_13859,N_13533,N_13365);
nand U13860 (N_13860,N_13217,N_13483);
or U13861 (N_13861,N_13296,N_13282);
xnor U13862 (N_13862,N_13305,N_13526);
nor U13863 (N_13863,N_13587,N_13494);
nor U13864 (N_13864,N_13230,N_13314);
nand U13865 (N_13865,N_13263,N_13277);
and U13866 (N_13866,N_13520,N_13476);
xor U13867 (N_13867,N_13388,N_13482);
xnor U13868 (N_13868,N_13274,N_13214);
or U13869 (N_13869,N_13369,N_13259);
xor U13870 (N_13870,N_13484,N_13327);
nand U13871 (N_13871,N_13512,N_13281);
nand U13872 (N_13872,N_13424,N_13403);
and U13873 (N_13873,N_13213,N_13423);
or U13874 (N_13874,N_13578,N_13509);
xnor U13875 (N_13875,N_13460,N_13405);
and U13876 (N_13876,N_13248,N_13217);
or U13877 (N_13877,N_13227,N_13582);
nand U13878 (N_13878,N_13547,N_13349);
nor U13879 (N_13879,N_13296,N_13490);
or U13880 (N_13880,N_13215,N_13515);
and U13881 (N_13881,N_13445,N_13353);
nor U13882 (N_13882,N_13470,N_13369);
xnor U13883 (N_13883,N_13277,N_13518);
nand U13884 (N_13884,N_13276,N_13489);
and U13885 (N_13885,N_13530,N_13239);
xor U13886 (N_13886,N_13426,N_13290);
xor U13887 (N_13887,N_13312,N_13371);
and U13888 (N_13888,N_13361,N_13522);
nor U13889 (N_13889,N_13493,N_13225);
nand U13890 (N_13890,N_13493,N_13234);
nand U13891 (N_13891,N_13273,N_13520);
xor U13892 (N_13892,N_13270,N_13221);
nor U13893 (N_13893,N_13301,N_13273);
and U13894 (N_13894,N_13389,N_13243);
nand U13895 (N_13895,N_13280,N_13373);
nor U13896 (N_13896,N_13403,N_13209);
xnor U13897 (N_13897,N_13464,N_13295);
or U13898 (N_13898,N_13282,N_13351);
or U13899 (N_13899,N_13282,N_13592);
xnor U13900 (N_13900,N_13552,N_13229);
nand U13901 (N_13901,N_13515,N_13475);
nand U13902 (N_13902,N_13469,N_13453);
and U13903 (N_13903,N_13427,N_13320);
nand U13904 (N_13904,N_13291,N_13545);
nand U13905 (N_13905,N_13484,N_13292);
nor U13906 (N_13906,N_13313,N_13212);
nor U13907 (N_13907,N_13497,N_13462);
nor U13908 (N_13908,N_13466,N_13292);
xnor U13909 (N_13909,N_13367,N_13349);
or U13910 (N_13910,N_13364,N_13428);
and U13911 (N_13911,N_13339,N_13539);
or U13912 (N_13912,N_13441,N_13481);
xnor U13913 (N_13913,N_13317,N_13278);
and U13914 (N_13914,N_13569,N_13222);
and U13915 (N_13915,N_13444,N_13340);
and U13916 (N_13916,N_13599,N_13202);
xnor U13917 (N_13917,N_13250,N_13261);
and U13918 (N_13918,N_13317,N_13581);
xnor U13919 (N_13919,N_13213,N_13508);
nor U13920 (N_13920,N_13256,N_13346);
nor U13921 (N_13921,N_13411,N_13356);
nand U13922 (N_13922,N_13251,N_13349);
or U13923 (N_13923,N_13472,N_13541);
nand U13924 (N_13924,N_13298,N_13439);
nor U13925 (N_13925,N_13313,N_13332);
xor U13926 (N_13926,N_13444,N_13524);
or U13927 (N_13927,N_13566,N_13504);
nor U13928 (N_13928,N_13414,N_13285);
and U13929 (N_13929,N_13250,N_13431);
xnor U13930 (N_13930,N_13217,N_13204);
xnor U13931 (N_13931,N_13299,N_13242);
xnor U13932 (N_13932,N_13263,N_13365);
nor U13933 (N_13933,N_13571,N_13432);
nand U13934 (N_13934,N_13248,N_13559);
or U13935 (N_13935,N_13366,N_13273);
and U13936 (N_13936,N_13553,N_13449);
and U13937 (N_13937,N_13319,N_13533);
and U13938 (N_13938,N_13336,N_13420);
and U13939 (N_13939,N_13348,N_13240);
or U13940 (N_13940,N_13224,N_13346);
xnor U13941 (N_13941,N_13286,N_13326);
nor U13942 (N_13942,N_13410,N_13266);
and U13943 (N_13943,N_13232,N_13507);
or U13944 (N_13944,N_13482,N_13462);
nand U13945 (N_13945,N_13479,N_13469);
and U13946 (N_13946,N_13271,N_13354);
or U13947 (N_13947,N_13411,N_13534);
nor U13948 (N_13948,N_13558,N_13207);
xnor U13949 (N_13949,N_13514,N_13572);
and U13950 (N_13950,N_13424,N_13565);
or U13951 (N_13951,N_13506,N_13429);
nand U13952 (N_13952,N_13571,N_13262);
or U13953 (N_13953,N_13559,N_13430);
or U13954 (N_13954,N_13438,N_13280);
nor U13955 (N_13955,N_13554,N_13427);
xnor U13956 (N_13956,N_13426,N_13267);
nor U13957 (N_13957,N_13383,N_13212);
nand U13958 (N_13958,N_13480,N_13520);
nand U13959 (N_13959,N_13453,N_13528);
nor U13960 (N_13960,N_13579,N_13275);
xnor U13961 (N_13961,N_13279,N_13498);
nand U13962 (N_13962,N_13548,N_13269);
nand U13963 (N_13963,N_13518,N_13589);
nor U13964 (N_13964,N_13423,N_13238);
nor U13965 (N_13965,N_13417,N_13279);
xor U13966 (N_13966,N_13504,N_13253);
or U13967 (N_13967,N_13508,N_13312);
nand U13968 (N_13968,N_13415,N_13541);
and U13969 (N_13969,N_13256,N_13310);
nor U13970 (N_13970,N_13445,N_13342);
xnor U13971 (N_13971,N_13544,N_13209);
or U13972 (N_13972,N_13216,N_13306);
nor U13973 (N_13973,N_13308,N_13249);
or U13974 (N_13974,N_13574,N_13288);
xor U13975 (N_13975,N_13516,N_13579);
and U13976 (N_13976,N_13200,N_13216);
or U13977 (N_13977,N_13543,N_13282);
and U13978 (N_13978,N_13319,N_13259);
nand U13979 (N_13979,N_13586,N_13300);
xor U13980 (N_13980,N_13241,N_13397);
or U13981 (N_13981,N_13556,N_13509);
nor U13982 (N_13982,N_13419,N_13329);
nand U13983 (N_13983,N_13257,N_13441);
xor U13984 (N_13984,N_13214,N_13388);
or U13985 (N_13985,N_13403,N_13318);
or U13986 (N_13986,N_13322,N_13443);
nor U13987 (N_13987,N_13223,N_13485);
nor U13988 (N_13988,N_13531,N_13420);
and U13989 (N_13989,N_13350,N_13301);
nand U13990 (N_13990,N_13338,N_13440);
nor U13991 (N_13991,N_13387,N_13235);
and U13992 (N_13992,N_13534,N_13305);
nand U13993 (N_13993,N_13278,N_13555);
xnor U13994 (N_13994,N_13513,N_13564);
xor U13995 (N_13995,N_13580,N_13488);
and U13996 (N_13996,N_13339,N_13552);
or U13997 (N_13997,N_13359,N_13535);
nor U13998 (N_13998,N_13229,N_13329);
nor U13999 (N_13999,N_13541,N_13495);
or U14000 (N_14000,N_13639,N_13699);
nor U14001 (N_14001,N_13831,N_13744);
or U14002 (N_14002,N_13771,N_13824);
or U14003 (N_14003,N_13983,N_13890);
and U14004 (N_14004,N_13974,N_13614);
nand U14005 (N_14005,N_13713,N_13768);
and U14006 (N_14006,N_13737,N_13620);
or U14007 (N_14007,N_13663,N_13843);
and U14008 (N_14008,N_13923,N_13984);
nor U14009 (N_14009,N_13792,N_13960);
nor U14010 (N_14010,N_13731,N_13864);
nand U14011 (N_14011,N_13697,N_13658);
nor U14012 (N_14012,N_13806,N_13956);
xor U14013 (N_14013,N_13778,N_13851);
and U14014 (N_14014,N_13701,N_13797);
nor U14015 (N_14015,N_13998,N_13964);
and U14016 (N_14016,N_13705,N_13607);
nor U14017 (N_14017,N_13674,N_13861);
or U14018 (N_14018,N_13911,N_13606);
nor U14019 (N_14019,N_13858,N_13753);
and U14020 (N_14020,N_13800,N_13885);
xnor U14021 (N_14021,N_13736,N_13835);
xor U14022 (N_14022,N_13640,N_13622);
nand U14023 (N_14023,N_13632,N_13905);
xor U14024 (N_14024,N_13869,N_13857);
and U14025 (N_14025,N_13810,N_13794);
or U14026 (N_14026,N_13747,N_13822);
nor U14027 (N_14027,N_13657,N_13793);
nor U14028 (N_14028,N_13827,N_13939);
or U14029 (N_14029,N_13791,N_13689);
xnor U14030 (N_14030,N_13881,N_13787);
nand U14031 (N_14031,N_13758,N_13702);
and U14032 (N_14032,N_13766,N_13803);
xor U14033 (N_14033,N_13669,N_13917);
and U14034 (N_14034,N_13954,N_13722);
nand U14035 (N_14035,N_13946,N_13756);
and U14036 (N_14036,N_13783,N_13664);
nor U14037 (N_14037,N_13764,N_13666);
nor U14038 (N_14038,N_13932,N_13748);
nand U14039 (N_14039,N_13973,N_13780);
and U14040 (N_14040,N_13818,N_13690);
and U14041 (N_14041,N_13661,N_13995);
or U14042 (N_14042,N_13990,N_13601);
nand U14043 (N_14043,N_13903,N_13681);
xor U14044 (N_14044,N_13976,N_13865);
xor U14045 (N_14045,N_13838,N_13720);
and U14046 (N_14046,N_13776,N_13817);
nor U14047 (N_14047,N_13910,N_13668);
nor U14048 (N_14048,N_13618,N_13804);
nand U14049 (N_14049,N_13936,N_13915);
nor U14050 (N_14050,N_13683,N_13892);
xor U14051 (N_14051,N_13934,N_13698);
nor U14052 (N_14052,N_13878,N_13845);
xor U14053 (N_14053,N_13708,N_13906);
and U14054 (N_14054,N_13985,N_13965);
or U14055 (N_14055,N_13949,N_13650);
nand U14056 (N_14056,N_13888,N_13959);
and U14057 (N_14057,N_13920,N_13757);
and U14058 (N_14058,N_13922,N_13833);
nor U14059 (N_14059,N_13740,N_13945);
nor U14060 (N_14060,N_13978,N_13755);
nand U14061 (N_14061,N_13672,N_13953);
nor U14062 (N_14062,N_13642,N_13608);
and U14063 (N_14063,N_13777,N_13633);
or U14064 (N_14064,N_13981,N_13918);
or U14065 (N_14065,N_13723,N_13805);
nand U14066 (N_14066,N_13788,N_13763);
xor U14067 (N_14067,N_13996,N_13929);
nor U14068 (N_14068,N_13704,N_13972);
and U14069 (N_14069,N_13914,N_13616);
or U14070 (N_14070,N_13840,N_13726);
or U14071 (N_14071,N_13774,N_13979);
and U14072 (N_14072,N_13844,N_13826);
nor U14073 (N_14073,N_13629,N_13625);
and U14074 (N_14074,N_13935,N_13814);
xor U14075 (N_14075,N_13837,N_13925);
and U14076 (N_14076,N_13604,N_13971);
nor U14077 (N_14077,N_13801,N_13717);
and U14078 (N_14078,N_13679,N_13928);
xor U14079 (N_14079,N_13933,N_13796);
xnor U14080 (N_14080,N_13786,N_13635);
nand U14081 (N_14081,N_13694,N_13961);
and U14082 (N_14082,N_13887,N_13942);
xor U14083 (N_14083,N_13916,N_13733);
nor U14084 (N_14084,N_13807,N_13876);
xor U14085 (N_14085,N_13686,N_13921);
xor U14086 (N_14086,N_13955,N_13931);
or U14087 (N_14087,N_13641,N_13856);
nand U14088 (N_14088,N_13852,N_13693);
nand U14089 (N_14089,N_13685,N_13868);
xnor U14090 (N_14090,N_13902,N_13623);
xnor U14091 (N_14091,N_13741,N_13784);
xor U14092 (N_14092,N_13710,N_13779);
and U14093 (N_14093,N_13675,N_13926);
or U14094 (N_14094,N_13765,N_13912);
and U14095 (N_14095,N_13671,N_13654);
xor U14096 (N_14096,N_13612,N_13636);
or U14097 (N_14097,N_13884,N_13759);
or U14098 (N_14098,N_13621,N_13725);
xnor U14099 (N_14099,N_13941,N_13651);
nand U14100 (N_14100,N_13615,N_13820);
or U14101 (N_14101,N_13982,N_13893);
nand U14102 (N_14102,N_13677,N_13882);
and U14103 (N_14103,N_13706,N_13847);
xor U14104 (N_14104,N_13825,N_13696);
and U14105 (N_14105,N_13957,N_13752);
and U14106 (N_14106,N_13966,N_13785);
nand U14107 (N_14107,N_13832,N_13962);
or U14108 (N_14108,N_13927,N_13754);
nor U14109 (N_14109,N_13815,N_13789);
xor U14110 (N_14110,N_13695,N_13691);
xor U14111 (N_14111,N_13734,N_13943);
xnor U14112 (N_14112,N_13970,N_13709);
nor U14113 (N_14113,N_13812,N_13853);
nor U14114 (N_14114,N_13711,N_13782);
nand U14115 (N_14115,N_13829,N_13952);
xnor U14116 (N_14116,N_13721,N_13848);
or U14117 (N_14117,N_13714,N_13886);
or U14118 (N_14118,N_13940,N_13988);
or U14119 (N_14119,N_13999,N_13638);
nand U14120 (N_14120,N_13863,N_13894);
nand U14121 (N_14121,N_13617,N_13670);
nor U14122 (N_14122,N_13900,N_13652);
or U14123 (N_14123,N_13680,N_13889);
nor U14124 (N_14124,N_13781,N_13951);
and U14125 (N_14125,N_13687,N_13898);
and U14126 (N_14126,N_13839,N_13950);
or U14127 (N_14127,N_13676,N_13854);
nand U14128 (N_14128,N_13655,N_13647);
xnor U14129 (N_14129,N_13603,N_13909);
nor U14130 (N_14130,N_13877,N_13611);
or U14131 (N_14131,N_13682,N_13773);
nand U14132 (N_14132,N_13767,N_13891);
xor U14133 (N_14133,N_13867,N_13850);
nor U14134 (N_14134,N_13937,N_13707);
or U14135 (N_14135,N_13862,N_13866);
or U14136 (N_14136,N_13762,N_13645);
xor U14137 (N_14137,N_13948,N_13649);
and U14138 (N_14138,N_13798,N_13630);
nand U14139 (N_14139,N_13997,N_13975);
nand U14140 (N_14140,N_13930,N_13944);
and U14141 (N_14141,N_13828,N_13727);
and U14142 (N_14142,N_13846,N_13730);
xnor U14143 (N_14143,N_13684,N_13994);
nor U14144 (N_14144,N_13991,N_13875);
and U14145 (N_14145,N_13656,N_13624);
and U14146 (N_14146,N_13977,N_13712);
nor U14147 (N_14147,N_13986,N_13855);
xor U14148 (N_14148,N_13790,N_13989);
and U14149 (N_14149,N_13770,N_13969);
nor U14150 (N_14150,N_13749,N_13883);
xnor U14151 (N_14151,N_13746,N_13963);
or U14152 (N_14152,N_13735,N_13819);
nand U14153 (N_14153,N_13769,N_13841);
and U14154 (N_14154,N_13719,N_13751);
and U14155 (N_14155,N_13742,N_13688);
xnor U14156 (N_14156,N_13610,N_13924);
xnor U14157 (N_14157,N_13772,N_13662);
or U14158 (N_14158,N_13795,N_13646);
xnor U14159 (N_14159,N_13860,N_13987);
and U14160 (N_14160,N_13874,N_13821);
and U14161 (N_14161,N_13605,N_13830);
nor U14162 (N_14162,N_13648,N_13897);
xor U14163 (N_14163,N_13834,N_13958);
xnor U14164 (N_14164,N_13813,N_13745);
xor U14165 (N_14165,N_13724,N_13667);
xor U14166 (N_14166,N_13967,N_13859);
xnor U14167 (N_14167,N_13993,N_13643);
nand U14168 (N_14168,N_13901,N_13842);
xnor U14169 (N_14169,N_13673,N_13904);
xor U14170 (N_14170,N_13718,N_13872);
nor U14171 (N_14171,N_13716,N_13634);
and U14172 (N_14172,N_13613,N_13913);
and U14173 (N_14173,N_13644,N_13637);
nand U14174 (N_14174,N_13700,N_13760);
and U14175 (N_14175,N_13619,N_13678);
or U14176 (N_14176,N_13665,N_13715);
xor U14177 (N_14177,N_13811,N_13609);
and U14178 (N_14178,N_13750,N_13732);
nor U14179 (N_14179,N_13908,N_13879);
nor U14180 (N_14180,N_13602,N_13880);
nor U14181 (N_14181,N_13775,N_13799);
xnor U14182 (N_14182,N_13692,N_13836);
and U14183 (N_14183,N_13660,N_13600);
nor U14184 (N_14184,N_13627,N_13895);
nand U14185 (N_14185,N_13980,N_13703);
and U14186 (N_14186,N_13899,N_13870);
or U14187 (N_14187,N_13738,N_13628);
or U14188 (N_14188,N_13802,N_13729);
nor U14189 (N_14189,N_13849,N_13743);
nor U14190 (N_14190,N_13907,N_13992);
nor U14191 (N_14191,N_13739,N_13938);
and U14192 (N_14192,N_13816,N_13631);
nand U14193 (N_14193,N_13968,N_13809);
xor U14194 (N_14194,N_13871,N_13896);
nor U14195 (N_14195,N_13761,N_13873);
or U14196 (N_14196,N_13808,N_13728);
nand U14197 (N_14197,N_13823,N_13919);
and U14198 (N_14198,N_13659,N_13947);
xor U14199 (N_14199,N_13653,N_13626);
and U14200 (N_14200,N_13800,N_13982);
and U14201 (N_14201,N_13979,N_13872);
nand U14202 (N_14202,N_13614,N_13938);
and U14203 (N_14203,N_13950,N_13813);
or U14204 (N_14204,N_13894,N_13968);
or U14205 (N_14205,N_13966,N_13830);
nor U14206 (N_14206,N_13893,N_13781);
nor U14207 (N_14207,N_13871,N_13603);
or U14208 (N_14208,N_13719,N_13948);
nor U14209 (N_14209,N_13873,N_13700);
xnor U14210 (N_14210,N_13655,N_13939);
and U14211 (N_14211,N_13673,N_13759);
xor U14212 (N_14212,N_13891,N_13880);
xnor U14213 (N_14213,N_13997,N_13718);
nand U14214 (N_14214,N_13683,N_13609);
nor U14215 (N_14215,N_13680,N_13809);
nor U14216 (N_14216,N_13604,N_13640);
nand U14217 (N_14217,N_13844,N_13706);
or U14218 (N_14218,N_13989,N_13910);
and U14219 (N_14219,N_13818,N_13892);
xor U14220 (N_14220,N_13930,N_13931);
nand U14221 (N_14221,N_13612,N_13703);
xnor U14222 (N_14222,N_13791,N_13755);
or U14223 (N_14223,N_13704,N_13736);
and U14224 (N_14224,N_13721,N_13765);
nand U14225 (N_14225,N_13781,N_13652);
or U14226 (N_14226,N_13894,N_13727);
or U14227 (N_14227,N_13825,N_13877);
xor U14228 (N_14228,N_13741,N_13679);
nor U14229 (N_14229,N_13873,N_13746);
nor U14230 (N_14230,N_13607,N_13638);
nor U14231 (N_14231,N_13699,N_13764);
and U14232 (N_14232,N_13903,N_13969);
nand U14233 (N_14233,N_13899,N_13817);
nand U14234 (N_14234,N_13739,N_13635);
or U14235 (N_14235,N_13748,N_13776);
or U14236 (N_14236,N_13700,N_13655);
or U14237 (N_14237,N_13948,N_13798);
nand U14238 (N_14238,N_13843,N_13910);
or U14239 (N_14239,N_13833,N_13942);
and U14240 (N_14240,N_13888,N_13639);
nor U14241 (N_14241,N_13646,N_13930);
nand U14242 (N_14242,N_13945,N_13817);
and U14243 (N_14243,N_13914,N_13692);
or U14244 (N_14244,N_13979,N_13935);
nor U14245 (N_14245,N_13720,N_13911);
xor U14246 (N_14246,N_13963,N_13660);
or U14247 (N_14247,N_13825,N_13764);
nor U14248 (N_14248,N_13702,N_13705);
or U14249 (N_14249,N_13930,N_13951);
or U14250 (N_14250,N_13770,N_13722);
nor U14251 (N_14251,N_13612,N_13691);
or U14252 (N_14252,N_13666,N_13833);
nand U14253 (N_14253,N_13776,N_13623);
nand U14254 (N_14254,N_13901,N_13659);
nand U14255 (N_14255,N_13686,N_13894);
xor U14256 (N_14256,N_13943,N_13940);
xor U14257 (N_14257,N_13815,N_13976);
xnor U14258 (N_14258,N_13678,N_13921);
or U14259 (N_14259,N_13776,N_13860);
or U14260 (N_14260,N_13890,N_13699);
nor U14261 (N_14261,N_13886,N_13682);
and U14262 (N_14262,N_13836,N_13933);
nand U14263 (N_14263,N_13958,N_13823);
and U14264 (N_14264,N_13704,N_13819);
and U14265 (N_14265,N_13626,N_13680);
and U14266 (N_14266,N_13804,N_13916);
xnor U14267 (N_14267,N_13689,N_13769);
nand U14268 (N_14268,N_13999,N_13692);
or U14269 (N_14269,N_13707,N_13819);
nand U14270 (N_14270,N_13626,N_13904);
nor U14271 (N_14271,N_13903,N_13953);
or U14272 (N_14272,N_13811,N_13689);
or U14273 (N_14273,N_13879,N_13657);
nor U14274 (N_14274,N_13818,N_13710);
xor U14275 (N_14275,N_13734,N_13949);
or U14276 (N_14276,N_13947,N_13876);
nor U14277 (N_14277,N_13898,N_13891);
or U14278 (N_14278,N_13839,N_13623);
nor U14279 (N_14279,N_13728,N_13768);
and U14280 (N_14280,N_13886,N_13810);
xnor U14281 (N_14281,N_13892,N_13705);
nor U14282 (N_14282,N_13996,N_13843);
and U14283 (N_14283,N_13765,N_13684);
nand U14284 (N_14284,N_13756,N_13664);
and U14285 (N_14285,N_13738,N_13973);
or U14286 (N_14286,N_13923,N_13652);
and U14287 (N_14287,N_13608,N_13784);
xnor U14288 (N_14288,N_13612,N_13856);
nor U14289 (N_14289,N_13981,N_13754);
or U14290 (N_14290,N_13889,N_13832);
and U14291 (N_14291,N_13632,N_13928);
or U14292 (N_14292,N_13976,N_13707);
and U14293 (N_14293,N_13895,N_13622);
xnor U14294 (N_14294,N_13709,N_13967);
nor U14295 (N_14295,N_13635,N_13748);
or U14296 (N_14296,N_13775,N_13762);
nor U14297 (N_14297,N_13885,N_13676);
xnor U14298 (N_14298,N_13691,N_13831);
and U14299 (N_14299,N_13834,N_13994);
or U14300 (N_14300,N_13635,N_13939);
or U14301 (N_14301,N_13600,N_13806);
nand U14302 (N_14302,N_13945,N_13994);
or U14303 (N_14303,N_13817,N_13755);
xnor U14304 (N_14304,N_13931,N_13952);
nor U14305 (N_14305,N_13846,N_13934);
and U14306 (N_14306,N_13797,N_13964);
nor U14307 (N_14307,N_13816,N_13616);
and U14308 (N_14308,N_13918,N_13633);
or U14309 (N_14309,N_13606,N_13695);
nor U14310 (N_14310,N_13734,N_13601);
nand U14311 (N_14311,N_13864,N_13757);
or U14312 (N_14312,N_13848,N_13903);
xor U14313 (N_14313,N_13825,N_13671);
nor U14314 (N_14314,N_13728,N_13824);
or U14315 (N_14315,N_13659,N_13785);
and U14316 (N_14316,N_13631,N_13637);
or U14317 (N_14317,N_13791,N_13606);
or U14318 (N_14318,N_13663,N_13785);
or U14319 (N_14319,N_13988,N_13627);
nor U14320 (N_14320,N_13978,N_13775);
nand U14321 (N_14321,N_13935,N_13910);
and U14322 (N_14322,N_13889,N_13749);
xnor U14323 (N_14323,N_13799,N_13900);
nand U14324 (N_14324,N_13995,N_13718);
xor U14325 (N_14325,N_13703,N_13830);
nor U14326 (N_14326,N_13802,N_13739);
xnor U14327 (N_14327,N_13754,N_13624);
or U14328 (N_14328,N_13914,N_13974);
or U14329 (N_14329,N_13972,N_13817);
nor U14330 (N_14330,N_13811,N_13769);
and U14331 (N_14331,N_13853,N_13999);
or U14332 (N_14332,N_13694,N_13897);
and U14333 (N_14333,N_13860,N_13732);
nor U14334 (N_14334,N_13963,N_13998);
or U14335 (N_14335,N_13606,N_13867);
or U14336 (N_14336,N_13788,N_13930);
xor U14337 (N_14337,N_13838,N_13697);
or U14338 (N_14338,N_13958,N_13652);
nand U14339 (N_14339,N_13624,N_13778);
xnor U14340 (N_14340,N_13739,N_13639);
nand U14341 (N_14341,N_13672,N_13889);
nor U14342 (N_14342,N_13709,N_13952);
nand U14343 (N_14343,N_13792,N_13733);
nor U14344 (N_14344,N_13669,N_13660);
nand U14345 (N_14345,N_13894,N_13854);
and U14346 (N_14346,N_13723,N_13605);
nand U14347 (N_14347,N_13652,N_13931);
and U14348 (N_14348,N_13633,N_13698);
or U14349 (N_14349,N_13627,N_13677);
and U14350 (N_14350,N_13892,N_13703);
nand U14351 (N_14351,N_13749,N_13912);
nor U14352 (N_14352,N_13605,N_13688);
nand U14353 (N_14353,N_13742,N_13953);
nor U14354 (N_14354,N_13844,N_13869);
nor U14355 (N_14355,N_13760,N_13978);
or U14356 (N_14356,N_13761,N_13808);
xor U14357 (N_14357,N_13655,N_13806);
nand U14358 (N_14358,N_13928,N_13610);
or U14359 (N_14359,N_13835,N_13646);
nor U14360 (N_14360,N_13918,N_13631);
or U14361 (N_14361,N_13680,N_13678);
xnor U14362 (N_14362,N_13966,N_13687);
or U14363 (N_14363,N_13846,N_13784);
nor U14364 (N_14364,N_13968,N_13815);
nand U14365 (N_14365,N_13790,N_13777);
xnor U14366 (N_14366,N_13803,N_13687);
xor U14367 (N_14367,N_13885,N_13964);
or U14368 (N_14368,N_13984,N_13667);
nor U14369 (N_14369,N_13600,N_13798);
or U14370 (N_14370,N_13704,N_13853);
or U14371 (N_14371,N_13922,N_13747);
or U14372 (N_14372,N_13605,N_13894);
nand U14373 (N_14373,N_13877,N_13780);
nor U14374 (N_14374,N_13689,N_13744);
and U14375 (N_14375,N_13684,N_13704);
and U14376 (N_14376,N_13674,N_13825);
xor U14377 (N_14377,N_13890,N_13870);
xor U14378 (N_14378,N_13690,N_13832);
or U14379 (N_14379,N_13911,N_13956);
or U14380 (N_14380,N_13861,N_13866);
and U14381 (N_14381,N_13903,N_13950);
or U14382 (N_14382,N_13783,N_13828);
nor U14383 (N_14383,N_13701,N_13991);
nor U14384 (N_14384,N_13602,N_13992);
nor U14385 (N_14385,N_13751,N_13718);
or U14386 (N_14386,N_13763,N_13923);
nand U14387 (N_14387,N_13732,N_13751);
and U14388 (N_14388,N_13946,N_13769);
nand U14389 (N_14389,N_13797,N_13866);
xnor U14390 (N_14390,N_13603,N_13845);
xnor U14391 (N_14391,N_13805,N_13956);
xor U14392 (N_14392,N_13911,N_13631);
or U14393 (N_14393,N_13974,N_13933);
nor U14394 (N_14394,N_13761,N_13712);
nor U14395 (N_14395,N_13869,N_13605);
or U14396 (N_14396,N_13611,N_13962);
nand U14397 (N_14397,N_13685,N_13764);
nand U14398 (N_14398,N_13992,N_13669);
xor U14399 (N_14399,N_13842,N_13726);
nand U14400 (N_14400,N_14219,N_14158);
and U14401 (N_14401,N_14231,N_14322);
xnor U14402 (N_14402,N_14034,N_14311);
xnor U14403 (N_14403,N_14205,N_14126);
and U14404 (N_14404,N_14188,N_14167);
nor U14405 (N_14405,N_14261,N_14294);
nor U14406 (N_14406,N_14060,N_14170);
xor U14407 (N_14407,N_14397,N_14276);
nor U14408 (N_14408,N_14324,N_14341);
or U14409 (N_14409,N_14332,N_14108);
nand U14410 (N_14410,N_14070,N_14107);
and U14411 (N_14411,N_14307,N_14267);
xor U14412 (N_14412,N_14043,N_14373);
xor U14413 (N_14413,N_14003,N_14216);
and U14414 (N_14414,N_14147,N_14016);
nand U14415 (N_14415,N_14377,N_14193);
or U14416 (N_14416,N_14222,N_14114);
nand U14417 (N_14417,N_14177,N_14235);
nor U14418 (N_14418,N_14331,N_14249);
or U14419 (N_14419,N_14385,N_14381);
and U14420 (N_14420,N_14323,N_14066);
nand U14421 (N_14421,N_14176,N_14252);
and U14422 (N_14422,N_14269,N_14358);
nand U14423 (N_14423,N_14181,N_14037);
nand U14424 (N_14424,N_14364,N_14325);
xor U14425 (N_14425,N_14163,N_14334);
nor U14426 (N_14426,N_14336,N_14308);
and U14427 (N_14427,N_14251,N_14208);
or U14428 (N_14428,N_14053,N_14335);
nor U14429 (N_14429,N_14321,N_14085);
nand U14430 (N_14430,N_14094,N_14215);
and U14431 (N_14431,N_14286,N_14345);
and U14432 (N_14432,N_14206,N_14309);
nor U14433 (N_14433,N_14050,N_14125);
and U14434 (N_14434,N_14081,N_14116);
xnor U14435 (N_14435,N_14368,N_14120);
xnor U14436 (N_14436,N_14029,N_14390);
and U14437 (N_14437,N_14351,N_14207);
nand U14438 (N_14438,N_14357,N_14100);
xnor U14439 (N_14439,N_14056,N_14164);
xor U14440 (N_14440,N_14315,N_14020);
and U14441 (N_14441,N_14233,N_14004);
nor U14442 (N_14442,N_14068,N_14184);
xnor U14443 (N_14443,N_14212,N_14393);
nor U14444 (N_14444,N_14001,N_14186);
and U14445 (N_14445,N_14041,N_14312);
and U14446 (N_14446,N_14237,N_14096);
nand U14447 (N_14447,N_14040,N_14217);
and U14448 (N_14448,N_14011,N_14305);
xnor U14449 (N_14449,N_14282,N_14145);
nand U14450 (N_14450,N_14287,N_14022);
or U14451 (N_14451,N_14062,N_14234);
nor U14452 (N_14452,N_14326,N_14248);
and U14453 (N_14453,N_14297,N_14241);
and U14454 (N_14454,N_14365,N_14306);
and U14455 (N_14455,N_14013,N_14347);
nor U14456 (N_14456,N_14372,N_14106);
nand U14457 (N_14457,N_14002,N_14187);
nor U14458 (N_14458,N_14348,N_14105);
xnor U14459 (N_14459,N_14151,N_14396);
nor U14460 (N_14460,N_14032,N_14366);
nand U14461 (N_14461,N_14354,N_14242);
nor U14462 (N_14462,N_14224,N_14098);
nor U14463 (N_14463,N_14239,N_14376);
or U14464 (N_14464,N_14179,N_14300);
nor U14465 (N_14465,N_14229,N_14007);
nand U14466 (N_14466,N_14015,N_14012);
xnor U14467 (N_14467,N_14061,N_14127);
xor U14468 (N_14468,N_14389,N_14173);
xnor U14469 (N_14469,N_14175,N_14008);
or U14470 (N_14470,N_14257,N_14262);
nor U14471 (N_14471,N_14316,N_14327);
nor U14472 (N_14472,N_14250,N_14374);
or U14473 (N_14473,N_14087,N_14018);
and U14474 (N_14474,N_14292,N_14386);
or U14475 (N_14475,N_14046,N_14117);
xor U14476 (N_14476,N_14048,N_14161);
and U14477 (N_14477,N_14255,N_14076);
nand U14478 (N_14478,N_14168,N_14112);
xnor U14479 (N_14479,N_14165,N_14099);
nor U14480 (N_14480,N_14221,N_14140);
and U14481 (N_14481,N_14042,N_14333);
or U14482 (N_14482,N_14135,N_14329);
nor U14483 (N_14483,N_14047,N_14361);
nand U14484 (N_14484,N_14088,N_14392);
or U14485 (N_14485,N_14367,N_14128);
and U14486 (N_14486,N_14166,N_14134);
or U14487 (N_14487,N_14356,N_14330);
nand U14488 (N_14488,N_14343,N_14119);
nor U14489 (N_14489,N_14057,N_14203);
and U14490 (N_14490,N_14084,N_14279);
xor U14491 (N_14491,N_14038,N_14264);
and U14492 (N_14492,N_14129,N_14228);
nand U14493 (N_14493,N_14246,N_14194);
nand U14494 (N_14494,N_14073,N_14245);
nand U14495 (N_14495,N_14148,N_14236);
and U14496 (N_14496,N_14258,N_14254);
nor U14497 (N_14497,N_14318,N_14154);
nor U14498 (N_14498,N_14362,N_14072);
nand U14499 (N_14499,N_14266,N_14380);
nor U14500 (N_14500,N_14124,N_14394);
nor U14501 (N_14501,N_14150,N_14025);
nor U14502 (N_14502,N_14083,N_14023);
nor U14503 (N_14503,N_14388,N_14133);
nand U14504 (N_14504,N_14328,N_14155);
or U14505 (N_14505,N_14178,N_14378);
and U14506 (N_14506,N_14058,N_14280);
and U14507 (N_14507,N_14283,N_14277);
nor U14508 (N_14508,N_14055,N_14353);
nand U14509 (N_14509,N_14370,N_14159);
and U14510 (N_14510,N_14162,N_14244);
nor U14511 (N_14511,N_14202,N_14174);
and U14512 (N_14512,N_14026,N_14115);
and U14513 (N_14513,N_14340,N_14288);
xnor U14514 (N_14514,N_14144,N_14247);
xor U14515 (N_14515,N_14319,N_14296);
and U14516 (N_14516,N_14395,N_14320);
and U14517 (N_14517,N_14180,N_14338);
nor U14518 (N_14518,N_14349,N_14101);
and U14519 (N_14519,N_14227,N_14028);
nand U14520 (N_14520,N_14146,N_14149);
nand U14521 (N_14521,N_14211,N_14295);
and U14522 (N_14522,N_14086,N_14171);
xor U14523 (N_14523,N_14104,N_14342);
and U14524 (N_14524,N_14110,N_14103);
or U14525 (N_14525,N_14024,N_14063);
nor U14526 (N_14526,N_14090,N_14059);
nor U14527 (N_14527,N_14152,N_14278);
nand U14528 (N_14528,N_14274,N_14226);
nor U14529 (N_14529,N_14078,N_14095);
xor U14530 (N_14530,N_14010,N_14253);
nor U14531 (N_14531,N_14017,N_14139);
or U14532 (N_14532,N_14359,N_14137);
xnor U14533 (N_14533,N_14067,N_14153);
xnor U14534 (N_14534,N_14021,N_14214);
and U14535 (N_14535,N_14379,N_14054);
or U14536 (N_14536,N_14169,N_14191);
or U14537 (N_14537,N_14138,N_14293);
nand U14538 (N_14538,N_14006,N_14369);
nand U14539 (N_14539,N_14384,N_14000);
nor U14540 (N_14540,N_14044,N_14182);
or U14541 (N_14541,N_14121,N_14387);
nand U14542 (N_14542,N_14156,N_14232);
and U14543 (N_14543,N_14118,N_14383);
and U14544 (N_14544,N_14009,N_14271);
or U14545 (N_14545,N_14074,N_14375);
nand U14546 (N_14546,N_14035,N_14299);
or U14547 (N_14547,N_14298,N_14049);
or U14548 (N_14548,N_14355,N_14260);
and U14549 (N_14549,N_14122,N_14192);
or U14550 (N_14550,N_14069,N_14132);
or U14551 (N_14551,N_14382,N_14142);
or U14552 (N_14552,N_14268,N_14172);
or U14553 (N_14553,N_14077,N_14230);
nand U14554 (N_14554,N_14102,N_14225);
nand U14555 (N_14555,N_14398,N_14079);
or U14556 (N_14556,N_14189,N_14065);
nor U14557 (N_14557,N_14064,N_14344);
or U14558 (N_14558,N_14310,N_14285);
or U14559 (N_14559,N_14019,N_14196);
or U14560 (N_14560,N_14289,N_14143);
nand U14561 (N_14561,N_14093,N_14201);
or U14562 (N_14562,N_14130,N_14123);
nand U14563 (N_14563,N_14111,N_14045);
and U14564 (N_14564,N_14185,N_14075);
or U14565 (N_14565,N_14238,N_14092);
xnor U14566 (N_14566,N_14314,N_14290);
and U14567 (N_14567,N_14141,N_14030);
xor U14568 (N_14568,N_14218,N_14036);
and U14569 (N_14569,N_14363,N_14273);
or U14570 (N_14570,N_14371,N_14399);
nor U14571 (N_14571,N_14240,N_14303);
and U14572 (N_14572,N_14097,N_14190);
nor U14573 (N_14573,N_14005,N_14339);
xnor U14574 (N_14574,N_14014,N_14027);
and U14575 (N_14575,N_14136,N_14265);
or U14576 (N_14576,N_14197,N_14082);
and U14577 (N_14577,N_14346,N_14033);
nand U14578 (N_14578,N_14272,N_14071);
or U14579 (N_14579,N_14284,N_14223);
nor U14580 (N_14580,N_14113,N_14313);
xnor U14581 (N_14581,N_14256,N_14213);
and U14582 (N_14582,N_14183,N_14352);
or U14583 (N_14583,N_14198,N_14259);
and U14584 (N_14584,N_14391,N_14204);
nand U14585 (N_14585,N_14360,N_14220);
nor U14586 (N_14586,N_14089,N_14209);
or U14587 (N_14587,N_14051,N_14263);
or U14588 (N_14588,N_14131,N_14031);
or U14589 (N_14589,N_14275,N_14052);
or U14590 (N_14590,N_14302,N_14200);
xnor U14591 (N_14591,N_14080,N_14157);
nand U14592 (N_14592,N_14195,N_14304);
nor U14593 (N_14593,N_14270,N_14350);
nand U14594 (N_14594,N_14039,N_14291);
xor U14595 (N_14595,N_14160,N_14281);
and U14596 (N_14596,N_14210,N_14301);
nand U14597 (N_14597,N_14337,N_14317);
nand U14598 (N_14598,N_14109,N_14091);
or U14599 (N_14599,N_14243,N_14199);
xnor U14600 (N_14600,N_14341,N_14217);
nand U14601 (N_14601,N_14390,N_14176);
xnor U14602 (N_14602,N_14082,N_14350);
nand U14603 (N_14603,N_14078,N_14204);
xor U14604 (N_14604,N_14322,N_14224);
nand U14605 (N_14605,N_14243,N_14074);
nor U14606 (N_14606,N_14071,N_14248);
or U14607 (N_14607,N_14113,N_14283);
xnor U14608 (N_14608,N_14115,N_14164);
nand U14609 (N_14609,N_14130,N_14100);
nor U14610 (N_14610,N_14102,N_14314);
or U14611 (N_14611,N_14034,N_14243);
and U14612 (N_14612,N_14272,N_14205);
xnor U14613 (N_14613,N_14010,N_14324);
nor U14614 (N_14614,N_14225,N_14112);
xor U14615 (N_14615,N_14192,N_14377);
nor U14616 (N_14616,N_14286,N_14039);
nand U14617 (N_14617,N_14158,N_14358);
xor U14618 (N_14618,N_14336,N_14340);
nor U14619 (N_14619,N_14024,N_14328);
xnor U14620 (N_14620,N_14317,N_14271);
or U14621 (N_14621,N_14085,N_14223);
and U14622 (N_14622,N_14264,N_14255);
xnor U14623 (N_14623,N_14340,N_14016);
nand U14624 (N_14624,N_14155,N_14353);
or U14625 (N_14625,N_14173,N_14371);
nand U14626 (N_14626,N_14127,N_14134);
or U14627 (N_14627,N_14364,N_14348);
or U14628 (N_14628,N_14182,N_14067);
or U14629 (N_14629,N_14003,N_14035);
nand U14630 (N_14630,N_14156,N_14285);
nand U14631 (N_14631,N_14050,N_14075);
nand U14632 (N_14632,N_14316,N_14396);
or U14633 (N_14633,N_14095,N_14145);
xnor U14634 (N_14634,N_14192,N_14143);
xor U14635 (N_14635,N_14144,N_14242);
xor U14636 (N_14636,N_14158,N_14046);
or U14637 (N_14637,N_14235,N_14061);
nand U14638 (N_14638,N_14358,N_14328);
xnor U14639 (N_14639,N_14213,N_14200);
nor U14640 (N_14640,N_14251,N_14253);
and U14641 (N_14641,N_14061,N_14011);
nand U14642 (N_14642,N_14215,N_14169);
nand U14643 (N_14643,N_14257,N_14178);
xnor U14644 (N_14644,N_14092,N_14124);
nor U14645 (N_14645,N_14225,N_14174);
nor U14646 (N_14646,N_14273,N_14350);
nand U14647 (N_14647,N_14184,N_14008);
nand U14648 (N_14648,N_14027,N_14384);
xnor U14649 (N_14649,N_14064,N_14168);
and U14650 (N_14650,N_14056,N_14346);
and U14651 (N_14651,N_14266,N_14250);
or U14652 (N_14652,N_14264,N_14379);
nor U14653 (N_14653,N_14128,N_14390);
or U14654 (N_14654,N_14353,N_14025);
and U14655 (N_14655,N_14375,N_14217);
and U14656 (N_14656,N_14219,N_14252);
xnor U14657 (N_14657,N_14005,N_14097);
xnor U14658 (N_14658,N_14062,N_14380);
nand U14659 (N_14659,N_14386,N_14128);
and U14660 (N_14660,N_14256,N_14216);
and U14661 (N_14661,N_14064,N_14083);
xnor U14662 (N_14662,N_14396,N_14290);
xor U14663 (N_14663,N_14151,N_14302);
xnor U14664 (N_14664,N_14148,N_14094);
nor U14665 (N_14665,N_14153,N_14314);
nor U14666 (N_14666,N_14244,N_14253);
xor U14667 (N_14667,N_14226,N_14136);
nor U14668 (N_14668,N_14054,N_14293);
or U14669 (N_14669,N_14303,N_14322);
nand U14670 (N_14670,N_14129,N_14125);
or U14671 (N_14671,N_14366,N_14339);
and U14672 (N_14672,N_14392,N_14364);
and U14673 (N_14673,N_14346,N_14083);
xor U14674 (N_14674,N_14059,N_14114);
or U14675 (N_14675,N_14397,N_14224);
nand U14676 (N_14676,N_14174,N_14158);
nand U14677 (N_14677,N_14312,N_14200);
and U14678 (N_14678,N_14158,N_14225);
nand U14679 (N_14679,N_14360,N_14129);
nand U14680 (N_14680,N_14316,N_14137);
nor U14681 (N_14681,N_14239,N_14305);
or U14682 (N_14682,N_14106,N_14073);
or U14683 (N_14683,N_14179,N_14007);
xnor U14684 (N_14684,N_14342,N_14004);
nor U14685 (N_14685,N_14336,N_14234);
nand U14686 (N_14686,N_14298,N_14033);
nor U14687 (N_14687,N_14066,N_14092);
nor U14688 (N_14688,N_14328,N_14350);
nor U14689 (N_14689,N_14091,N_14354);
and U14690 (N_14690,N_14161,N_14204);
or U14691 (N_14691,N_14227,N_14030);
nor U14692 (N_14692,N_14134,N_14111);
and U14693 (N_14693,N_14176,N_14076);
or U14694 (N_14694,N_14334,N_14117);
nand U14695 (N_14695,N_14125,N_14182);
and U14696 (N_14696,N_14101,N_14100);
nand U14697 (N_14697,N_14020,N_14102);
xor U14698 (N_14698,N_14383,N_14190);
nand U14699 (N_14699,N_14236,N_14171);
and U14700 (N_14700,N_14197,N_14232);
xor U14701 (N_14701,N_14132,N_14062);
and U14702 (N_14702,N_14071,N_14396);
nand U14703 (N_14703,N_14132,N_14105);
or U14704 (N_14704,N_14336,N_14191);
and U14705 (N_14705,N_14347,N_14214);
nor U14706 (N_14706,N_14081,N_14066);
and U14707 (N_14707,N_14187,N_14100);
nor U14708 (N_14708,N_14029,N_14039);
xor U14709 (N_14709,N_14196,N_14138);
nand U14710 (N_14710,N_14346,N_14266);
and U14711 (N_14711,N_14057,N_14218);
nor U14712 (N_14712,N_14395,N_14226);
xor U14713 (N_14713,N_14206,N_14024);
xnor U14714 (N_14714,N_14335,N_14249);
nand U14715 (N_14715,N_14088,N_14348);
or U14716 (N_14716,N_14285,N_14349);
nand U14717 (N_14717,N_14211,N_14190);
or U14718 (N_14718,N_14031,N_14080);
xor U14719 (N_14719,N_14031,N_14189);
nand U14720 (N_14720,N_14306,N_14325);
nor U14721 (N_14721,N_14178,N_14151);
or U14722 (N_14722,N_14251,N_14258);
nor U14723 (N_14723,N_14152,N_14393);
nor U14724 (N_14724,N_14229,N_14003);
xnor U14725 (N_14725,N_14360,N_14108);
xnor U14726 (N_14726,N_14234,N_14244);
xnor U14727 (N_14727,N_14316,N_14154);
xnor U14728 (N_14728,N_14390,N_14023);
nand U14729 (N_14729,N_14035,N_14205);
and U14730 (N_14730,N_14146,N_14148);
nor U14731 (N_14731,N_14242,N_14103);
xor U14732 (N_14732,N_14011,N_14007);
nand U14733 (N_14733,N_14273,N_14357);
or U14734 (N_14734,N_14133,N_14315);
nor U14735 (N_14735,N_14001,N_14239);
nor U14736 (N_14736,N_14248,N_14052);
nand U14737 (N_14737,N_14147,N_14199);
nor U14738 (N_14738,N_14070,N_14069);
or U14739 (N_14739,N_14068,N_14145);
nand U14740 (N_14740,N_14067,N_14156);
xor U14741 (N_14741,N_14178,N_14220);
or U14742 (N_14742,N_14083,N_14208);
or U14743 (N_14743,N_14390,N_14245);
or U14744 (N_14744,N_14317,N_14157);
and U14745 (N_14745,N_14307,N_14049);
nand U14746 (N_14746,N_14387,N_14209);
xnor U14747 (N_14747,N_14316,N_14002);
nand U14748 (N_14748,N_14137,N_14257);
or U14749 (N_14749,N_14150,N_14340);
nor U14750 (N_14750,N_14092,N_14244);
xor U14751 (N_14751,N_14082,N_14018);
or U14752 (N_14752,N_14217,N_14054);
and U14753 (N_14753,N_14244,N_14013);
and U14754 (N_14754,N_14008,N_14102);
and U14755 (N_14755,N_14192,N_14298);
nor U14756 (N_14756,N_14035,N_14375);
and U14757 (N_14757,N_14093,N_14344);
xor U14758 (N_14758,N_14088,N_14150);
or U14759 (N_14759,N_14328,N_14009);
xnor U14760 (N_14760,N_14138,N_14137);
nand U14761 (N_14761,N_14191,N_14343);
and U14762 (N_14762,N_14291,N_14367);
or U14763 (N_14763,N_14271,N_14152);
or U14764 (N_14764,N_14259,N_14208);
and U14765 (N_14765,N_14373,N_14125);
and U14766 (N_14766,N_14084,N_14258);
or U14767 (N_14767,N_14058,N_14328);
nor U14768 (N_14768,N_14250,N_14163);
nor U14769 (N_14769,N_14140,N_14162);
nand U14770 (N_14770,N_14089,N_14215);
nor U14771 (N_14771,N_14004,N_14263);
nor U14772 (N_14772,N_14247,N_14191);
or U14773 (N_14773,N_14000,N_14113);
nand U14774 (N_14774,N_14257,N_14383);
nand U14775 (N_14775,N_14257,N_14141);
nor U14776 (N_14776,N_14397,N_14098);
nand U14777 (N_14777,N_14126,N_14022);
and U14778 (N_14778,N_14207,N_14033);
or U14779 (N_14779,N_14254,N_14389);
nand U14780 (N_14780,N_14307,N_14052);
nor U14781 (N_14781,N_14317,N_14280);
xnor U14782 (N_14782,N_14300,N_14127);
nor U14783 (N_14783,N_14083,N_14110);
or U14784 (N_14784,N_14232,N_14364);
and U14785 (N_14785,N_14324,N_14167);
nand U14786 (N_14786,N_14385,N_14356);
and U14787 (N_14787,N_14259,N_14141);
or U14788 (N_14788,N_14192,N_14309);
or U14789 (N_14789,N_14348,N_14350);
or U14790 (N_14790,N_14047,N_14061);
and U14791 (N_14791,N_14073,N_14220);
xnor U14792 (N_14792,N_14087,N_14033);
and U14793 (N_14793,N_14091,N_14347);
xnor U14794 (N_14794,N_14147,N_14152);
or U14795 (N_14795,N_14100,N_14142);
or U14796 (N_14796,N_14235,N_14112);
nor U14797 (N_14797,N_14227,N_14067);
or U14798 (N_14798,N_14209,N_14193);
nand U14799 (N_14799,N_14107,N_14327);
and U14800 (N_14800,N_14559,N_14786);
nor U14801 (N_14801,N_14770,N_14775);
or U14802 (N_14802,N_14730,N_14594);
xor U14803 (N_14803,N_14563,N_14703);
xnor U14804 (N_14804,N_14527,N_14468);
xnor U14805 (N_14805,N_14607,N_14684);
or U14806 (N_14806,N_14420,N_14790);
nand U14807 (N_14807,N_14489,N_14604);
or U14808 (N_14808,N_14476,N_14475);
nor U14809 (N_14809,N_14745,N_14788);
or U14810 (N_14810,N_14682,N_14766);
nor U14811 (N_14811,N_14485,N_14628);
or U14812 (N_14812,N_14542,N_14456);
and U14813 (N_14813,N_14492,N_14680);
nand U14814 (N_14814,N_14421,N_14716);
nor U14815 (N_14815,N_14447,N_14416);
xnor U14816 (N_14816,N_14494,N_14583);
nand U14817 (N_14817,N_14678,N_14548);
nand U14818 (N_14818,N_14496,N_14409);
xor U14819 (N_14819,N_14528,N_14443);
nor U14820 (N_14820,N_14676,N_14731);
xor U14821 (N_14821,N_14799,N_14545);
and U14822 (N_14822,N_14562,N_14778);
nor U14823 (N_14823,N_14408,N_14639);
nor U14824 (N_14824,N_14437,N_14659);
nand U14825 (N_14825,N_14647,N_14631);
xor U14826 (N_14826,N_14585,N_14617);
nor U14827 (N_14827,N_14723,N_14430);
xnor U14828 (N_14828,N_14523,N_14728);
and U14829 (N_14829,N_14720,N_14455);
nand U14830 (N_14830,N_14495,N_14602);
nand U14831 (N_14831,N_14595,N_14640);
nand U14832 (N_14832,N_14406,N_14516);
nand U14833 (N_14833,N_14660,N_14792);
and U14834 (N_14834,N_14736,N_14760);
nand U14835 (N_14835,N_14795,N_14742);
xor U14836 (N_14836,N_14412,N_14439);
nand U14837 (N_14837,N_14605,N_14624);
and U14838 (N_14838,N_14424,N_14546);
nor U14839 (N_14839,N_14571,N_14756);
and U14840 (N_14840,N_14664,N_14428);
and U14841 (N_14841,N_14400,N_14612);
xnor U14842 (N_14842,N_14620,N_14509);
nor U14843 (N_14843,N_14704,N_14774);
nor U14844 (N_14844,N_14515,N_14547);
and U14845 (N_14845,N_14598,N_14635);
nand U14846 (N_14846,N_14779,N_14487);
xor U14847 (N_14847,N_14590,N_14621);
nand U14848 (N_14848,N_14450,N_14535);
nand U14849 (N_14849,N_14435,N_14751);
or U14850 (N_14850,N_14415,N_14434);
or U14851 (N_14851,N_14449,N_14404);
nor U14852 (N_14852,N_14505,N_14674);
xor U14853 (N_14853,N_14477,N_14499);
or U14854 (N_14854,N_14618,N_14473);
or U14855 (N_14855,N_14762,N_14761);
and U14856 (N_14856,N_14502,N_14681);
xor U14857 (N_14857,N_14606,N_14689);
or U14858 (N_14858,N_14462,N_14708);
and U14859 (N_14859,N_14629,N_14789);
and U14860 (N_14860,N_14432,N_14752);
or U14861 (N_14861,N_14705,N_14675);
xor U14862 (N_14862,N_14507,N_14724);
xnor U14863 (N_14863,N_14725,N_14553);
nor U14864 (N_14864,N_14438,N_14407);
nand U14865 (N_14865,N_14481,N_14419);
nor U14866 (N_14866,N_14459,N_14763);
nand U14867 (N_14867,N_14490,N_14539);
xnor U14868 (N_14868,N_14743,N_14471);
nor U14869 (N_14869,N_14798,N_14694);
xnor U14870 (N_14870,N_14622,N_14410);
or U14871 (N_14871,N_14525,N_14533);
xnor U14872 (N_14872,N_14588,N_14727);
nor U14873 (N_14873,N_14740,N_14500);
xnor U14874 (N_14874,N_14579,N_14772);
nor U14875 (N_14875,N_14698,N_14651);
nand U14876 (N_14876,N_14668,N_14710);
nand U14877 (N_14877,N_14702,N_14469);
and U14878 (N_14878,N_14636,N_14638);
xnor U14879 (N_14879,N_14451,N_14654);
nor U14880 (N_14880,N_14461,N_14474);
nand U14881 (N_14881,N_14706,N_14671);
or U14882 (N_14882,N_14572,N_14729);
nor U14883 (N_14883,N_14738,N_14465);
or U14884 (N_14884,N_14422,N_14677);
nand U14885 (N_14885,N_14609,N_14543);
or U14886 (N_14886,N_14458,N_14483);
xnor U14887 (N_14887,N_14445,N_14735);
nor U14888 (N_14888,N_14442,N_14673);
nand U14889 (N_14889,N_14418,N_14749);
nor U14890 (N_14890,N_14470,N_14576);
or U14891 (N_14891,N_14425,N_14567);
and U14892 (N_14892,N_14552,N_14764);
or U14893 (N_14893,N_14557,N_14614);
xor U14894 (N_14894,N_14596,N_14644);
and U14895 (N_14895,N_14601,N_14575);
xnor U14896 (N_14896,N_14611,N_14732);
nor U14897 (N_14897,N_14707,N_14791);
and U14898 (N_14898,N_14454,N_14427);
nor U14899 (N_14899,N_14670,N_14608);
or U14900 (N_14900,N_14769,N_14541);
or U14901 (N_14901,N_14613,N_14662);
and U14902 (N_14902,N_14581,N_14615);
nor U14903 (N_14903,N_14522,N_14561);
xor U14904 (N_14904,N_14593,N_14755);
xor U14905 (N_14905,N_14587,N_14582);
xor U14906 (N_14906,N_14619,N_14460);
xor U14907 (N_14907,N_14782,N_14632);
nor U14908 (N_14908,N_14696,N_14642);
or U14909 (N_14909,N_14544,N_14472);
xor U14910 (N_14910,N_14411,N_14785);
nand U14911 (N_14911,N_14665,N_14506);
xor U14912 (N_14912,N_14580,N_14537);
nor U14913 (N_14913,N_14715,N_14565);
nor U14914 (N_14914,N_14771,N_14610);
xnor U14915 (N_14915,N_14759,N_14777);
nand U14916 (N_14916,N_14574,N_14417);
nor U14917 (N_14917,N_14726,N_14683);
or U14918 (N_14918,N_14555,N_14661);
nor U14919 (N_14919,N_14700,N_14633);
nor U14920 (N_14920,N_14479,N_14637);
and U14921 (N_14921,N_14486,N_14649);
and U14922 (N_14922,N_14484,N_14655);
or U14923 (N_14923,N_14688,N_14734);
nor U14924 (N_14924,N_14603,N_14478);
nor U14925 (N_14925,N_14627,N_14692);
nor U14926 (N_14926,N_14796,N_14467);
nand U14927 (N_14927,N_14737,N_14739);
or U14928 (N_14928,N_14616,N_14656);
and U14929 (N_14929,N_14510,N_14713);
or U14930 (N_14930,N_14672,N_14754);
or U14931 (N_14931,N_14741,N_14488);
or U14932 (N_14932,N_14540,N_14402);
or U14933 (N_14933,N_14657,N_14482);
xor U14934 (N_14934,N_14578,N_14586);
nor U14935 (N_14935,N_14599,N_14685);
and U14936 (N_14936,N_14498,N_14401);
xor U14937 (N_14937,N_14717,N_14570);
xor U14938 (N_14938,N_14667,N_14626);
nand U14939 (N_14939,N_14773,N_14591);
nor U14940 (N_14940,N_14709,N_14554);
or U14941 (N_14941,N_14480,N_14429);
or U14942 (N_14942,N_14560,N_14414);
or U14943 (N_14943,N_14780,N_14767);
xnor U14944 (N_14944,N_14513,N_14690);
nand U14945 (N_14945,N_14797,N_14457);
xor U14946 (N_14946,N_14520,N_14524);
xnor U14947 (N_14947,N_14733,N_14529);
nor U14948 (N_14948,N_14521,N_14503);
nor U14949 (N_14949,N_14758,N_14566);
xnor U14950 (N_14950,N_14719,N_14556);
and U14951 (N_14951,N_14663,N_14508);
nand U14952 (N_14952,N_14721,N_14746);
or U14953 (N_14953,N_14464,N_14514);
nand U14954 (N_14954,N_14491,N_14444);
nor U14955 (N_14955,N_14531,N_14564);
and U14956 (N_14956,N_14433,N_14765);
nor U14957 (N_14957,N_14463,N_14549);
or U14958 (N_14958,N_14781,N_14691);
or U14959 (N_14959,N_14584,N_14568);
or U14960 (N_14960,N_14423,N_14686);
xnor U14961 (N_14961,N_14493,N_14597);
nand U14962 (N_14962,N_14440,N_14592);
nor U14963 (N_14963,N_14431,N_14511);
nor U14964 (N_14964,N_14793,N_14646);
and U14965 (N_14965,N_14641,N_14699);
and U14966 (N_14966,N_14783,N_14526);
nand U14967 (N_14967,N_14446,N_14630);
nand U14968 (N_14968,N_14558,N_14534);
nand U14969 (N_14969,N_14600,N_14530);
or U14970 (N_14970,N_14787,N_14550);
and U14971 (N_14971,N_14711,N_14666);
or U14972 (N_14972,N_14569,N_14744);
and U14973 (N_14973,N_14643,N_14650);
and U14974 (N_14974,N_14448,N_14693);
and U14975 (N_14975,N_14441,N_14536);
and U14976 (N_14976,N_14538,N_14679);
xnor U14977 (N_14977,N_14645,N_14784);
xnor U14978 (N_14978,N_14518,N_14718);
nor U14979 (N_14979,N_14519,N_14747);
xnor U14980 (N_14980,N_14573,N_14697);
xnor U14981 (N_14981,N_14722,N_14517);
nor U14982 (N_14982,N_14625,N_14405);
xor U14983 (N_14983,N_14623,N_14753);
nand U14984 (N_14984,N_14669,N_14634);
nor U14985 (N_14985,N_14653,N_14403);
nand U14986 (N_14986,N_14648,N_14589);
and U14987 (N_14987,N_14512,N_14426);
nor U14988 (N_14988,N_14497,N_14658);
nor U14989 (N_14989,N_14453,N_14413);
nand U14990 (N_14990,N_14466,N_14750);
nor U14991 (N_14991,N_14776,N_14757);
xnor U14992 (N_14992,N_14501,N_14794);
xnor U14993 (N_14993,N_14714,N_14652);
nand U14994 (N_14994,N_14701,N_14687);
or U14995 (N_14995,N_14436,N_14452);
nor U14996 (N_14996,N_14577,N_14551);
nand U14997 (N_14997,N_14712,N_14695);
nor U14998 (N_14998,N_14768,N_14532);
or U14999 (N_14999,N_14504,N_14748);
nand U15000 (N_15000,N_14469,N_14783);
or U15001 (N_15001,N_14520,N_14786);
nor U15002 (N_15002,N_14611,N_14525);
and U15003 (N_15003,N_14745,N_14736);
nor U15004 (N_15004,N_14720,N_14493);
nor U15005 (N_15005,N_14698,N_14705);
nor U15006 (N_15006,N_14705,N_14623);
or U15007 (N_15007,N_14706,N_14732);
or U15008 (N_15008,N_14713,N_14404);
xnor U15009 (N_15009,N_14550,N_14584);
and U15010 (N_15010,N_14569,N_14453);
nor U15011 (N_15011,N_14672,N_14643);
nor U15012 (N_15012,N_14723,N_14605);
or U15013 (N_15013,N_14781,N_14681);
nand U15014 (N_15014,N_14459,N_14766);
xor U15015 (N_15015,N_14424,N_14465);
or U15016 (N_15016,N_14632,N_14630);
nor U15017 (N_15017,N_14628,N_14758);
nor U15018 (N_15018,N_14403,N_14685);
nor U15019 (N_15019,N_14491,N_14588);
xor U15020 (N_15020,N_14736,N_14708);
and U15021 (N_15021,N_14586,N_14734);
xnor U15022 (N_15022,N_14656,N_14717);
nor U15023 (N_15023,N_14544,N_14537);
nor U15024 (N_15024,N_14604,N_14782);
and U15025 (N_15025,N_14571,N_14717);
or U15026 (N_15026,N_14489,N_14402);
xor U15027 (N_15027,N_14488,N_14743);
nor U15028 (N_15028,N_14473,N_14433);
nor U15029 (N_15029,N_14617,N_14444);
nor U15030 (N_15030,N_14592,N_14432);
nor U15031 (N_15031,N_14790,N_14750);
nor U15032 (N_15032,N_14443,N_14798);
and U15033 (N_15033,N_14504,N_14594);
or U15034 (N_15034,N_14673,N_14686);
or U15035 (N_15035,N_14639,N_14571);
nand U15036 (N_15036,N_14591,N_14456);
or U15037 (N_15037,N_14708,N_14509);
or U15038 (N_15038,N_14445,N_14679);
nor U15039 (N_15039,N_14528,N_14650);
and U15040 (N_15040,N_14415,N_14567);
xnor U15041 (N_15041,N_14602,N_14421);
nand U15042 (N_15042,N_14726,N_14490);
nor U15043 (N_15043,N_14524,N_14739);
or U15044 (N_15044,N_14409,N_14567);
nor U15045 (N_15045,N_14706,N_14548);
or U15046 (N_15046,N_14648,N_14556);
nand U15047 (N_15047,N_14435,N_14502);
xnor U15048 (N_15048,N_14448,N_14742);
or U15049 (N_15049,N_14411,N_14782);
nand U15050 (N_15050,N_14466,N_14738);
xor U15051 (N_15051,N_14510,N_14633);
nor U15052 (N_15052,N_14743,N_14594);
xnor U15053 (N_15053,N_14581,N_14662);
and U15054 (N_15054,N_14732,N_14547);
xnor U15055 (N_15055,N_14468,N_14532);
xnor U15056 (N_15056,N_14414,N_14566);
or U15057 (N_15057,N_14580,N_14530);
nor U15058 (N_15058,N_14710,N_14756);
xor U15059 (N_15059,N_14578,N_14475);
xor U15060 (N_15060,N_14694,N_14512);
nand U15061 (N_15061,N_14460,N_14689);
nand U15062 (N_15062,N_14661,N_14750);
nor U15063 (N_15063,N_14566,N_14415);
nand U15064 (N_15064,N_14500,N_14437);
nand U15065 (N_15065,N_14556,N_14486);
and U15066 (N_15066,N_14402,N_14627);
xor U15067 (N_15067,N_14592,N_14643);
or U15068 (N_15068,N_14539,N_14416);
and U15069 (N_15069,N_14632,N_14525);
or U15070 (N_15070,N_14412,N_14755);
xnor U15071 (N_15071,N_14570,N_14709);
and U15072 (N_15072,N_14627,N_14749);
or U15073 (N_15073,N_14637,N_14612);
xor U15074 (N_15074,N_14477,N_14533);
or U15075 (N_15075,N_14508,N_14728);
nor U15076 (N_15076,N_14643,N_14620);
or U15077 (N_15077,N_14645,N_14460);
nor U15078 (N_15078,N_14795,N_14797);
xor U15079 (N_15079,N_14524,N_14478);
and U15080 (N_15080,N_14442,N_14631);
nand U15081 (N_15081,N_14624,N_14650);
nand U15082 (N_15082,N_14758,N_14755);
xor U15083 (N_15083,N_14564,N_14521);
and U15084 (N_15084,N_14632,N_14615);
xor U15085 (N_15085,N_14687,N_14418);
nand U15086 (N_15086,N_14484,N_14688);
nor U15087 (N_15087,N_14510,N_14405);
nand U15088 (N_15088,N_14408,N_14554);
nor U15089 (N_15089,N_14777,N_14790);
xnor U15090 (N_15090,N_14759,N_14580);
nor U15091 (N_15091,N_14788,N_14633);
and U15092 (N_15092,N_14776,N_14501);
xnor U15093 (N_15093,N_14793,N_14487);
or U15094 (N_15094,N_14797,N_14562);
and U15095 (N_15095,N_14758,N_14411);
xor U15096 (N_15096,N_14516,N_14603);
nor U15097 (N_15097,N_14736,N_14722);
xor U15098 (N_15098,N_14467,N_14504);
nor U15099 (N_15099,N_14552,N_14745);
nand U15100 (N_15100,N_14426,N_14659);
nor U15101 (N_15101,N_14699,N_14689);
and U15102 (N_15102,N_14779,N_14410);
nor U15103 (N_15103,N_14723,N_14786);
nor U15104 (N_15104,N_14745,N_14551);
xnor U15105 (N_15105,N_14412,N_14418);
xnor U15106 (N_15106,N_14765,N_14559);
nand U15107 (N_15107,N_14445,N_14582);
nand U15108 (N_15108,N_14603,N_14787);
and U15109 (N_15109,N_14552,N_14780);
xor U15110 (N_15110,N_14632,N_14623);
and U15111 (N_15111,N_14598,N_14449);
and U15112 (N_15112,N_14531,N_14668);
nand U15113 (N_15113,N_14471,N_14472);
or U15114 (N_15114,N_14578,N_14643);
nand U15115 (N_15115,N_14674,N_14754);
nand U15116 (N_15116,N_14736,N_14514);
and U15117 (N_15117,N_14543,N_14547);
nor U15118 (N_15118,N_14742,N_14492);
xor U15119 (N_15119,N_14423,N_14609);
nor U15120 (N_15120,N_14457,N_14425);
nand U15121 (N_15121,N_14799,N_14693);
and U15122 (N_15122,N_14436,N_14666);
nand U15123 (N_15123,N_14764,N_14404);
and U15124 (N_15124,N_14434,N_14621);
or U15125 (N_15125,N_14543,N_14637);
nand U15126 (N_15126,N_14634,N_14575);
nor U15127 (N_15127,N_14562,N_14780);
or U15128 (N_15128,N_14457,N_14592);
xor U15129 (N_15129,N_14639,N_14715);
nand U15130 (N_15130,N_14773,N_14625);
xor U15131 (N_15131,N_14793,N_14555);
or U15132 (N_15132,N_14511,N_14481);
or U15133 (N_15133,N_14573,N_14701);
or U15134 (N_15134,N_14747,N_14729);
nand U15135 (N_15135,N_14561,N_14406);
and U15136 (N_15136,N_14499,N_14700);
and U15137 (N_15137,N_14593,N_14556);
xor U15138 (N_15138,N_14724,N_14407);
nand U15139 (N_15139,N_14737,N_14412);
or U15140 (N_15140,N_14660,N_14451);
xnor U15141 (N_15141,N_14423,N_14567);
nand U15142 (N_15142,N_14737,N_14688);
xor U15143 (N_15143,N_14527,N_14704);
and U15144 (N_15144,N_14739,N_14509);
nor U15145 (N_15145,N_14579,N_14582);
nor U15146 (N_15146,N_14675,N_14550);
or U15147 (N_15147,N_14464,N_14578);
xnor U15148 (N_15148,N_14573,N_14570);
and U15149 (N_15149,N_14454,N_14582);
xor U15150 (N_15150,N_14730,N_14791);
nor U15151 (N_15151,N_14743,N_14714);
nor U15152 (N_15152,N_14569,N_14650);
or U15153 (N_15153,N_14561,N_14481);
xnor U15154 (N_15154,N_14508,N_14526);
or U15155 (N_15155,N_14662,N_14517);
xnor U15156 (N_15156,N_14737,N_14704);
and U15157 (N_15157,N_14773,N_14799);
nor U15158 (N_15158,N_14675,N_14481);
and U15159 (N_15159,N_14567,N_14427);
nand U15160 (N_15160,N_14584,N_14743);
or U15161 (N_15161,N_14587,N_14461);
xor U15162 (N_15162,N_14443,N_14482);
and U15163 (N_15163,N_14566,N_14585);
nor U15164 (N_15164,N_14538,N_14418);
or U15165 (N_15165,N_14768,N_14628);
and U15166 (N_15166,N_14545,N_14762);
and U15167 (N_15167,N_14641,N_14724);
or U15168 (N_15168,N_14724,N_14701);
nand U15169 (N_15169,N_14726,N_14402);
nand U15170 (N_15170,N_14405,N_14733);
nand U15171 (N_15171,N_14791,N_14738);
and U15172 (N_15172,N_14400,N_14696);
nand U15173 (N_15173,N_14744,N_14503);
and U15174 (N_15174,N_14504,N_14508);
nor U15175 (N_15175,N_14701,N_14519);
nor U15176 (N_15176,N_14676,N_14783);
nand U15177 (N_15177,N_14687,N_14634);
or U15178 (N_15178,N_14417,N_14490);
nand U15179 (N_15179,N_14501,N_14563);
nand U15180 (N_15180,N_14562,N_14494);
nor U15181 (N_15181,N_14534,N_14497);
xor U15182 (N_15182,N_14505,N_14409);
or U15183 (N_15183,N_14613,N_14414);
and U15184 (N_15184,N_14698,N_14675);
nor U15185 (N_15185,N_14711,N_14544);
and U15186 (N_15186,N_14431,N_14584);
or U15187 (N_15187,N_14415,N_14728);
and U15188 (N_15188,N_14739,N_14471);
xor U15189 (N_15189,N_14724,N_14784);
and U15190 (N_15190,N_14426,N_14579);
nor U15191 (N_15191,N_14463,N_14575);
or U15192 (N_15192,N_14769,N_14756);
xor U15193 (N_15193,N_14545,N_14478);
and U15194 (N_15194,N_14434,N_14409);
and U15195 (N_15195,N_14552,N_14443);
nand U15196 (N_15196,N_14487,N_14426);
or U15197 (N_15197,N_14686,N_14418);
nand U15198 (N_15198,N_14788,N_14584);
or U15199 (N_15199,N_14618,N_14642);
nand U15200 (N_15200,N_14999,N_15031);
and U15201 (N_15201,N_14987,N_14845);
or U15202 (N_15202,N_15127,N_15091);
and U15203 (N_15203,N_15076,N_14939);
and U15204 (N_15204,N_14921,N_15009);
nor U15205 (N_15205,N_15124,N_15042);
or U15206 (N_15206,N_15101,N_15000);
xor U15207 (N_15207,N_14903,N_14837);
xor U15208 (N_15208,N_15066,N_15104);
xnor U15209 (N_15209,N_14970,N_15097);
xor U15210 (N_15210,N_14800,N_14872);
xnor U15211 (N_15211,N_14883,N_15055);
nor U15212 (N_15212,N_15069,N_14906);
xnor U15213 (N_15213,N_14997,N_14870);
xor U15214 (N_15214,N_15185,N_14828);
nor U15215 (N_15215,N_15022,N_14826);
xor U15216 (N_15216,N_14973,N_14878);
nand U15217 (N_15217,N_14917,N_15155);
xor U15218 (N_15218,N_15165,N_15167);
nand U15219 (N_15219,N_15111,N_15174);
or U15220 (N_15220,N_14927,N_15149);
xor U15221 (N_15221,N_14943,N_15199);
or U15222 (N_15222,N_15032,N_14851);
and U15223 (N_15223,N_15008,N_15057);
nor U15224 (N_15224,N_14983,N_14912);
and U15225 (N_15225,N_14940,N_15035);
or U15226 (N_15226,N_15108,N_14835);
nand U15227 (N_15227,N_14813,N_15193);
xnor U15228 (N_15228,N_14823,N_14991);
nand U15229 (N_15229,N_15078,N_14928);
and U15230 (N_15230,N_14879,N_15045);
xnor U15231 (N_15231,N_15080,N_15190);
and U15232 (N_15232,N_15134,N_14848);
xor U15233 (N_15233,N_14831,N_14911);
nor U15234 (N_15234,N_15038,N_14958);
nand U15235 (N_15235,N_15161,N_15077);
or U15236 (N_15236,N_15178,N_14899);
nor U15237 (N_15237,N_14896,N_14881);
or U15238 (N_15238,N_14989,N_15014);
nand U15239 (N_15239,N_15050,N_14944);
or U15240 (N_15240,N_14996,N_15026);
or U15241 (N_15241,N_15040,N_14971);
or U15242 (N_15242,N_14884,N_15084);
and U15243 (N_15243,N_14876,N_14825);
or U15244 (N_15244,N_15125,N_15043);
xnor U15245 (N_15245,N_14969,N_14956);
nand U15246 (N_15246,N_14961,N_15093);
or U15247 (N_15247,N_15061,N_14886);
or U15248 (N_15248,N_14865,N_14887);
nand U15249 (N_15249,N_15117,N_14807);
and U15250 (N_15250,N_14836,N_14873);
xnor U15251 (N_15251,N_15138,N_15172);
nand U15252 (N_15252,N_15115,N_14804);
nor U15253 (N_15253,N_15012,N_15092);
and U15254 (N_15254,N_14910,N_14947);
or U15255 (N_15255,N_15074,N_14992);
nor U15256 (N_15256,N_15139,N_14888);
and U15257 (N_15257,N_15059,N_14897);
nand U15258 (N_15258,N_14858,N_14880);
and U15259 (N_15259,N_14908,N_14950);
xnor U15260 (N_15260,N_15143,N_15168);
nand U15261 (N_15261,N_15189,N_14859);
nor U15262 (N_15262,N_14934,N_15060);
or U15263 (N_15263,N_14951,N_15196);
or U15264 (N_15264,N_15173,N_14801);
nor U15265 (N_15265,N_15079,N_15192);
nor U15266 (N_15266,N_15051,N_14850);
xnor U15267 (N_15267,N_15015,N_15175);
and U15268 (N_15268,N_15075,N_15004);
or U15269 (N_15269,N_14841,N_15132);
nor U15270 (N_15270,N_14929,N_15123);
and U15271 (N_15271,N_14901,N_14981);
nand U15272 (N_15272,N_15002,N_15072);
and U15273 (N_15273,N_14803,N_15126);
nor U15274 (N_15274,N_14838,N_14984);
or U15275 (N_15275,N_15119,N_15103);
nand U15276 (N_15276,N_14931,N_14864);
xnor U15277 (N_15277,N_14954,N_15120);
nor U15278 (N_15278,N_14948,N_15052);
nand U15279 (N_15279,N_15116,N_14842);
and U15280 (N_15280,N_15156,N_15169);
or U15281 (N_15281,N_14933,N_14898);
or U15282 (N_15282,N_14932,N_15021);
nand U15283 (N_15283,N_14868,N_15157);
nor U15284 (N_15284,N_15023,N_15105);
nand U15285 (N_15285,N_15131,N_14811);
nor U15286 (N_15286,N_15095,N_15140);
and U15287 (N_15287,N_14810,N_14905);
and U15288 (N_15288,N_14855,N_14967);
or U15289 (N_15289,N_14982,N_15086);
xor U15290 (N_15290,N_15028,N_14839);
or U15291 (N_15291,N_14802,N_15017);
and U15292 (N_15292,N_15150,N_14953);
xor U15293 (N_15293,N_15136,N_14893);
nor U15294 (N_15294,N_15144,N_15062);
nor U15295 (N_15295,N_15033,N_15180);
nand U15296 (N_15296,N_14824,N_15016);
and U15297 (N_15297,N_14892,N_14834);
xnor U15298 (N_15298,N_14942,N_15036);
or U15299 (N_15299,N_15037,N_15162);
xor U15300 (N_15300,N_15183,N_14817);
nand U15301 (N_15301,N_15135,N_14985);
xnor U15302 (N_15302,N_15024,N_15058);
nor U15303 (N_15303,N_15068,N_14840);
xnor U15304 (N_15304,N_14874,N_14922);
or U15305 (N_15305,N_15047,N_15018);
nor U15306 (N_15306,N_14949,N_14815);
or U15307 (N_15307,N_14849,N_14854);
nand U15308 (N_15308,N_15194,N_15085);
or U15309 (N_15309,N_15122,N_14968);
nand U15310 (N_15310,N_14833,N_15065);
xor U15311 (N_15311,N_15142,N_14980);
or U15312 (N_15312,N_15109,N_14821);
nand U15313 (N_15313,N_15171,N_14853);
nand U15314 (N_15314,N_15153,N_14889);
and U15315 (N_15315,N_14866,N_15152);
nand U15316 (N_15316,N_15146,N_15130);
or U15317 (N_15317,N_14930,N_14894);
xnor U15318 (N_15318,N_15073,N_15070);
nand U15319 (N_15319,N_14861,N_14990);
nor U15320 (N_15320,N_15044,N_15159);
xnor U15321 (N_15321,N_15141,N_15010);
xnor U15322 (N_15322,N_14946,N_14846);
nand U15323 (N_15323,N_14902,N_15110);
xor U15324 (N_15324,N_14863,N_14805);
xnor U15325 (N_15325,N_14822,N_14925);
nor U15326 (N_15326,N_14945,N_15163);
nand U15327 (N_15327,N_14916,N_15121);
or U15328 (N_15328,N_15160,N_15197);
and U15329 (N_15329,N_15137,N_15013);
xnor U15330 (N_15330,N_14819,N_14900);
nor U15331 (N_15331,N_15071,N_15188);
nor U15332 (N_15332,N_15039,N_14844);
nor U15333 (N_15333,N_14952,N_15081);
nor U15334 (N_15334,N_15102,N_14843);
xor U15335 (N_15335,N_15151,N_14962);
xor U15336 (N_15336,N_14827,N_14808);
or U15337 (N_15337,N_14862,N_14812);
or U15338 (N_15338,N_15182,N_15094);
and U15339 (N_15339,N_14938,N_15096);
or U15340 (N_15340,N_14806,N_15128);
xor U15341 (N_15341,N_14974,N_15030);
and U15342 (N_15342,N_15025,N_14914);
xnor U15343 (N_15343,N_15054,N_15158);
and U15344 (N_15344,N_14993,N_14875);
nor U15345 (N_15345,N_15090,N_14890);
xnor U15346 (N_15346,N_15170,N_14857);
or U15347 (N_15347,N_15053,N_14935);
nand U15348 (N_15348,N_14994,N_14895);
and U15349 (N_15349,N_15087,N_14920);
nand U15350 (N_15350,N_15064,N_15118);
and U15351 (N_15351,N_14869,N_15164);
and U15352 (N_15352,N_14998,N_14814);
and U15353 (N_15353,N_15056,N_14867);
or U15354 (N_15354,N_14904,N_15067);
and U15355 (N_15355,N_15112,N_15154);
nor U15356 (N_15356,N_15186,N_14955);
xor U15357 (N_15357,N_15034,N_14918);
or U15358 (N_15358,N_15083,N_14960);
nand U15359 (N_15359,N_15187,N_14832);
nor U15360 (N_15360,N_15195,N_15198);
nor U15361 (N_15361,N_14877,N_15166);
or U15362 (N_15362,N_15176,N_15027);
nand U15363 (N_15363,N_15191,N_14978);
nor U15364 (N_15364,N_14941,N_14882);
or U15365 (N_15365,N_14976,N_15003);
or U15366 (N_15366,N_14963,N_15001);
xor U15367 (N_15367,N_14926,N_14995);
nand U15368 (N_15368,N_14986,N_15113);
or U15369 (N_15369,N_15046,N_15089);
nor U15370 (N_15370,N_15100,N_14924);
nor U15371 (N_15371,N_15181,N_15147);
nand U15372 (N_15372,N_14988,N_14915);
and U15373 (N_15373,N_14965,N_14964);
or U15374 (N_15374,N_14936,N_15019);
or U15375 (N_15375,N_15184,N_14919);
nor U15376 (N_15376,N_14972,N_15005);
nor U15377 (N_15377,N_15106,N_14830);
and U15378 (N_15378,N_14816,N_15133);
xnor U15379 (N_15379,N_14959,N_14907);
nor U15380 (N_15380,N_14909,N_14891);
xnor U15381 (N_15381,N_14885,N_14923);
xnor U15382 (N_15382,N_15177,N_15041);
or U15383 (N_15383,N_14977,N_15063);
and U15384 (N_15384,N_14957,N_14847);
nor U15385 (N_15385,N_15088,N_15006);
and U15386 (N_15386,N_15029,N_15049);
and U15387 (N_15387,N_15082,N_14975);
nand U15388 (N_15388,N_15099,N_14829);
xnor U15389 (N_15389,N_15148,N_15114);
nand U15390 (N_15390,N_14820,N_14871);
and U15391 (N_15391,N_15129,N_14860);
or U15392 (N_15392,N_14856,N_15145);
or U15393 (N_15393,N_14913,N_15098);
nand U15394 (N_15394,N_15011,N_14979);
or U15395 (N_15395,N_15020,N_14966);
nor U15396 (N_15396,N_14937,N_15048);
xor U15397 (N_15397,N_15179,N_14818);
nor U15398 (N_15398,N_14852,N_15007);
or U15399 (N_15399,N_14809,N_15107);
nor U15400 (N_15400,N_15102,N_14973);
and U15401 (N_15401,N_15151,N_15184);
nand U15402 (N_15402,N_14961,N_15067);
nand U15403 (N_15403,N_15172,N_14819);
xor U15404 (N_15404,N_14897,N_15146);
and U15405 (N_15405,N_14969,N_15064);
nor U15406 (N_15406,N_15138,N_15111);
nand U15407 (N_15407,N_14859,N_15141);
nand U15408 (N_15408,N_15173,N_14875);
nand U15409 (N_15409,N_14849,N_15001);
nand U15410 (N_15410,N_14959,N_14952);
or U15411 (N_15411,N_14835,N_14968);
nor U15412 (N_15412,N_15054,N_15056);
xor U15413 (N_15413,N_14869,N_15154);
and U15414 (N_15414,N_15091,N_14824);
nor U15415 (N_15415,N_15042,N_14846);
or U15416 (N_15416,N_15139,N_14911);
or U15417 (N_15417,N_15027,N_14908);
and U15418 (N_15418,N_15093,N_15132);
nor U15419 (N_15419,N_15044,N_15017);
nand U15420 (N_15420,N_15122,N_14885);
and U15421 (N_15421,N_14873,N_14927);
nor U15422 (N_15422,N_14955,N_15030);
and U15423 (N_15423,N_14811,N_14864);
or U15424 (N_15424,N_15174,N_14882);
and U15425 (N_15425,N_15024,N_15081);
xnor U15426 (N_15426,N_15098,N_15066);
and U15427 (N_15427,N_14889,N_14936);
and U15428 (N_15428,N_14930,N_15011);
and U15429 (N_15429,N_14849,N_15062);
and U15430 (N_15430,N_14811,N_14888);
nand U15431 (N_15431,N_14881,N_14986);
or U15432 (N_15432,N_15043,N_15124);
xnor U15433 (N_15433,N_14851,N_14817);
and U15434 (N_15434,N_14940,N_14898);
or U15435 (N_15435,N_14956,N_15069);
nand U15436 (N_15436,N_14973,N_14862);
xnor U15437 (N_15437,N_14877,N_14819);
nor U15438 (N_15438,N_14914,N_15132);
or U15439 (N_15439,N_15048,N_14835);
or U15440 (N_15440,N_15032,N_14890);
nand U15441 (N_15441,N_14930,N_14917);
or U15442 (N_15442,N_15176,N_14950);
nor U15443 (N_15443,N_15145,N_14968);
nor U15444 (N_15444,N_15058,N_15061);
and U15445 (N_15445,N_14925,N_15117);
xor U15446 (N_15446,N_14948,N_15063);
or U15447 (N_15447,N_14823,N_15184);
and U15448 (N_15448,N_14941,N_14925);
nor U15449 (N_15449,N_15177,N_14856);
xor U15450 (N_15450,N_15079,N_14941);
nand U15451 (N_15451,N_14895,N_14837);
and U15452 (N_15452,N_15093,N_15054);
nor U15453 (N_15453,N_15122,N_15192);
or U15454 (N_15454,N_15141,N_14932);
nor U15455 (N_15455,N_14992,N_14889);
nor U15456 (N_15456,N_14875,N_14862);
nor U15457 (N_15457,N_14971,N_14909);
or U15458 (N_15458,N_15005,N_15136);
and U15459 (N_15459,N_14800,N_14847);
nand U15460 (N_15460,N_15135,N_14880);
and U15461 (N_15461,N_14957,N_15012);
or U15462 (N_15462,N_14981,N_15161);
nor U15463 (N_15463,N_15079,N_14832);
nor U15464 (N_15464,N_15069,N_14944);
nand U15465 (N_15465,N_14813,N_14954);
nand U15466 (N_15466,N_14980,N_14860);
and U15467 (N_15467,N_15188,N_15167);
nand U15468 (N_15468,N_15180,N_14980);
and U15469 (N_15469,N_15180,N_15102);
nand U15470 (N_15470,N_14880,N_14900);
nand U15471 (N_15471,N_15003,N_14809);
or U15472 (N_15472,N_14980,N_14806);
nor U15473 (N_15473,N_14835,N_15034);
nand U15474 (N_15474,N_14819,N_15052);
and U15475 (N_15475,N_15077,N_14877);
and U15476 (N_15476,N_14978,N_15144);
and U15477 (N_15477,N_15101,N_14947);
and U15478 (N_15478,N_15133,N_15135);
and U15479 (N_15479,N_14926,N_15110);
xnor U15480 (N_15480,N_14852,N_15198);
nand U15481 (N_15481,N_14993,N_15161);
nand U15482 (N_15482,N_15085,N_14983);
nor U15483 (N_15483,N_15044,N_14901);
nand U15484 (N_15484,N_15089,N_14951);
or U15485 (N_15485,N_15162,N_14956);
nand U15486 (N_15486,N_15121,N_14845);
and U15487 (N_15487,N_15039,N_15080);
nand U15488 (N_15488,N_14990,N_14881);
and U15489 (N_15489,N_15069,N_14948);
nor U15490 (N_15490,N_14839,N_15045);
xor U15491 (N_15491,N_15038,N_14848);
and U15492 (N_15492,N_15061,N_15177);
or U15493 (N_15493,N_14997,N_14854);
or U15494 (N_15494,N_14818,N_15191);
xnor U15495 (N_15495,N_14956,N_14885);
nor U15496 (N_15496,N_15045,N_14849);
xor U15497 (N_15497,N_14898,N_15183);
or U15498 (N_15498,N_15128,N_14855);
and U15499 (N_15499,N_14972,N_14931);
nand U15500 (N_15500,N_14866,N_15113);
nand U15501 (N_15501,N_14908,N_15167);
and U15502 (N_15502,N_15131,N_14826);
xor U15503 (N_15503,N_15151,N_15109);
nor U15504 (N_15504,N_15095,N_15017);
nor U15505 (N_15505,N_14988,N_15061);
or U15506 (N_15506,N_14898,N_15089);
nand U15507 (N_15507,N_14994,N_14915);
or U15508 (N_15508,N_15085,N_14857);
xnor U15509 (N_15509,N_15105,N_15082);
xnor U15510 (N_15510,N_15093,N_15157);
or U15511 (N_15511,N_14834,N_15143);
nand U15512 (N_15512,N_14890,N_14819);
nand U15513 (N_15513,N_14983,N_15132);
or U15514 (N_15514,N_14923,N_15029);
xnor U15515 (N_15515,N_15090,N_15197);
nand U15516 (N_15516,N_14808,N_14990);
nand U15517 (N_15517,N_14968,N_15099);
nor U15518 (N_15518,N_14974,N_15026);
nor U15519 (N_15519,N_14940,N_15097);
or U15520 (N_15520,N_14992,N_14867);
and U15521 (N_15521,N_14840,N_14864);
xor U15522 (N_15522,N_15098,N_15031);
or U15523 (N_15523,N_14833,N_15189);
nor U15524 (N_15524,N_14891,N_14822);
nand U15525 (N_15525,N_15063,N_14848);
nor U15526 (N_15526,N_14814,N_15191);
xor U15527 (N_15527,N_14882,N_15028);
or U15528 (N_15528,N_15100,N_14809);
and U15529 (N_15529,N_15065,N_14868);
nand U15530 (N_15530,N_15130,N_14914);
or U15531 (N_15531,N_15063,N_14954);
or U15532 (N_15532,N_15134,N_15157);
xor U15533 (N_15533,N_15069,N_15019);
xor U15534 (N_15534,N_14815,N_14946);
xnor U15535 (N_15535,N_14816,N_14948);
and U15536 (N_15536,N_14900,N_15015);
or U15537 (N_15537,N_15095,N_15057);
xor U15538 (N_15538,N_15055,N_14882);
or U15539 (N_15539,N_15122,N_14839);
or U15540 (N_15540,N_14935,N_14827);
nor U15541 (N_15541,N_14964,N_15004);
nand U15542 (N_15542,N_14969,N_14857);
nand U15543 (N_15543,N_14973,N_15106);
nor U15544 (N_15544,N_14885,N_15185);
nor U15545 (N_15545,N_15158,N_15013);
or U15546 (N_15546,N_15040,N_15165);
nor U15547 (N_15547,N_14822,N_14821);
xnor U15548 (N_15548,N_15061,N_15199);
xor U15549 (N_15549,N_15004,N_15112);
nor U15550 (N_15550,N_14851,N_15191);
and U15551 (N_15551,N_15166,N_14990);
xnor U15552 (N_15552,N_15032,N_15072);
or U15553 (N_15553,N_14927,N_15141);
xor U15554 (N_15554,N_15092,N_15015);
xnor U15555 (N_15555,N_15162,N_14948);
or U15556 (N_15556,N_14958,N_14976);
nor U15557 (N_15557,N_15007,N_14809);
nor U15558 (N_15558,N_14904,N_15148);
or U15559 (N_15559,N_15199,N_14814);
or U15560 (N_15560,N_14937,N_15154);
and U15561 (N_15561,N_15059,N_15165);
nand U15562 (N_15562,N_15138,N_14931);
and U15563 (N_15563,N_14996,N_15051);
or U15564 (N_15564,N_15049,N_15004);
nor U15565 (N_15565,N_14843,N_14974);
nor U15566 (N_15566,N_14985,N_15146);
or U15567 (N_15567,N_14892,N_14823);
xor U15568 (N_15568,N_14872,N_14818);
or U15569 (N_15569,N_14820,N_14812);
nor U15570 (N_15570,N_15072,N_15141);
and U15571 (N_15571,N_15095,N_15147);
xnor U15572 (N_15572,N_15162,N_14863);
xor U15573 (N_15573,N_15104,N_14902);
xnor U15574 (N_15574,N_15123,N_15149);
and U15575 (N_15575,N_15010,N_14882);
nand U15576 (N_15576,N_15081,N_15096);
nor U15577 (N_15577,N_14859,N_14973);
and U15578 (N_15578,N_14849,N_14905);
nand U15579 (N_15579,N_14830,N_15064);
nand U15580 (N_15580,N_15005,N_14875);
xor U15581 (N_15581,N_15014,N_14975);
xor U15582 (N_15582,N_15173,N_15143);
nor U15583 (N_15583,N_14947,N_14800);
or U15584 (N_15584,N_15106,N_14801);
nand U15585 (N_15585,N_14905,N_14877);
nor U15586 (N_15586,N_14937,N_15083);
or U15587 (N_15587,N_14851,N_15112);
nand U15588 (N_15588,N_14856,N_14810);
and U15589 (N_15589,N_15081,N_15006);
and U15590 (N_15590,N_14864,N_14966);
and U15591 (N_15591,N_15124,N_14993);
nor U15592 (N_15592,N_15076,N_15184);
xnor U15593 (N_15593,N_14815,N_14806);
xor U15594 (N_15594,N_14872,N_15044);
nand U15595 (N_15595,N_14852,N_14968);
or U15596 (N_15596,N_14824,N_15059);
and U15597 (N_15597,N_14878,N_14951);
and U15598 (N_15598,N_15141,N_15126);
and U15599 (N_15599,N_15184,N_15099);
and U15600 (N_15600,N_15269,N_15336);
nand U15601 (N_15601,N_15585,N_15241);
or U15602 (N_15602,N_15544,N_15338);
nand U15603 (N_15603,N_15281,N_15239);
xor U15604 (N_15604,N_15477,N_15230);
xnor U15605 (N_15605,N_15265,N_15219);
and U15606 (N_15606,N_15541,N_15318);
xor U15607 (N_15607,N_15503,N_15556);
or U15608 (N_15608,N_15533,N_15583);
or U15609 (N_15609,N_15413,N_15314);
xor U15610 (N_15610,N_15291,N_15403);
nand U15611 (N_15611,N_15431,N_15460);
or U15612 (N_15612,N_15342,N_15308);
or U15613 (N_15613,N_15350,N_15211);
nand U15614 (N_15614,N_15236,N_15378);
xnor U15615 (N_15615,N_15373,N_15345);
and U15616 (N_15616,N_15441,N_15598);
and U15617 (N_15617,N_15446,N_15573);
nand U15618 (N_15618,N_15450,N_15509);
xnor U15619 (N_15619,N_15370,N_15325);
nor U15620 (N_15620,N_15531,N_15339);
nand U15621 (N_15621,N_15459,N_15377);
xnor U15622 (N_15622,N_15470,N_15592);
nor U15623 (N_15623,N_15233,N_15250);
xor U15624 (N_15624,N_15232,N_15514);
xor U15625 (N_15625,N_15546,N_15539);
and U15626 (N_15626,N_15499,N_15283);
nand U15627 (N_15627,N_15467,N_15213);
or U15628 (N_15628,N_15466,N_15438);
xnor U15629 (N_15629,N_15374,N_15207);
and U15630 (N_15630,N_15271,N_15449);
and U15631 (N_15631,N_15382,N_15225);
xnor U15632 (N_15632,N_15212,N_15572);
xnor U15633 (N_15633,N_15406,N_15488);
and U15634 (N_15634,N_15465,N_15340);
or U15635 (N_15635,N_15540,N_15506);
xor U15636 (N_15636,N_15589,N_15356);
nand U15637 (N_15637,N_15321,N_15414);
xor U15638 (N_15638,N_15405,N_15278);
xnor U15639 (N_15639,N_15226,N_15423);
and U15640 (N_15640,N_15579,N_15298);
or U15641 (N_15641,N_15381,N_15229);
nand U15642 (N_15642,N_15346,N_15279);
nor U15643 (N_15643,N_15386,N_15555);
nand U15644 (N_15644,N_15272,N_15445);
nor U15645 (N_15645,N_15416,N_15457);
or U15646 (N_15646,N_15549,N_15526);
and U15647 (N_15647,N_15306,N_15483);
nor U15648 (N_15648,N_15428,N_15376);
xor U15649 (N_15649,N_15347,N_15227);
nor U15650 (N_15650,N_15400,N_15390);
xnor U15651 (N_15651,N_15480,N_15288);
nand U15652 (N_15652,N_15204,N_15486);
nand U15653 (N_15653,N_15323,N_15520);
or U15654 (N_15654,N_15551,N_15494);
and U15655 (N_15655,N_15536,N_15261);
nor U15656 (N_15656,N_15537,N_15303);
nand U15657 (N_15657,N_15408,N_15394);
nand U15658 (N_15658,N_15410,N_15440);
and U15659 (N_15659,N_15505,N_15569);
xnor U15660 (N_15660,N_15310,N_15222);
nor U15661 (N_15661,N_15348,N_15472);
nor U15662 (N_15662,N_15392,N_15453);
nand U15663 (N_15663,N_15562,N_15581);
and U15664 (N_15664,N_15240,N_15553);
and U15665 (N_15665,N_15251,N_15586);
nor U15666 (N_15666,N_15424,N_15273);
xnor U15667 (N_15667,N_15257,N_15202);
and U15668 (N_15668,N_15593,N_15471);
nand U15669 (N_15669,N_15341,N_15263);
xnor U15670 (N_15670,N_15497,N_15237);
nor U15671 (N_15671,N_15485,N_15430);
or U15672 (N_15672,N_15206,N_15532);
or U15673 (N_15673,N_15523,N_15482);
nand U15674 (N_15674,N_15337,N_15302);
xor U15675 (N_15675,N_15513,N_15548);
nor U15676 (N_15676,N_15409,N_15436);
nor U15677 (N_15677,N_15312,N_15215);
nand U15678 (N_15678,N_15387,N_15286);
and U15679 (N_15679,N_15481,N_15395);
xor U15680 (N_15680,N_15504,N_15590);
and U15681 (N_15681,N_15254,N_15500);
nand U15682 (N_15682,N_15456,N_15362);
or U15683 (N_15683,N_15412,N_15571);
or U15684 (N_15684,N_15519,N_15260);
xnor U15685 (N_15685,N_15359,N_15476);
or U15686 (N_15686,N_15461,N_15563);
and U15687 (N_15687,N_15311,N_15383);
and U15688 (N_15688,N_15357,N_15448);
nor U15689 (N_15689,N_15420,N_15332);
xor U15690 (N_15690,N_15369,N_15397);
and U15691 (N_15691,N_15524,N_15319);
and U15692 (N_15692,N_15599,N_15309);
nor U15693 (N_15693,N_15530,N_15246);
and U15694 (N_15694,N_15326,N_15554);
or U15695 (N_15695,N_15300,N_15249);
nand U15696 (N_15696,N_15216,N_15401);
nor U15697 (N_15697,N_15452,N_15425);
or U15698 (N_15698,N_15510,N_15349);
xnor U15699 (N_15699,N_15388,N_15508);
xor U15700 (N_15700,N_15447,N_15501);
xor U15701 (N_15701,N_15463,N_15535);
or U15702 (N_15702,N_15360,N_15584);
and U15703 (N_15703,N_15493,N_15258);
nand U15704 (N_15704,N_15521,N_15380);
nand U15705 (N_15705,N_15329,N_15565);
nand U15706 (N_15706,N_15379,N_15407);
nand U15707 (N_15707,N_15574,N_15277);
nor U15708 (N_15708,N_15552,N_15578);
nor U15709 (N_15709,N_15231,N_15522);
nand U15710 (N_15710,N_15478,N_15515);
xor U15711 (N_15711,N_15433,N_15245);
nand U15712 (N_15712,N_15316,N_15315);
or U15713 (N_15713,N_15365,N_15507);
or U15714 (N_15714,N_15244,N_15305);
nand U15715 (N_15715,N_15528,N_15203);
nor U15716 (N_15716,N_15550,N_15201);
xor U15717 (N_15717,N_15596,N_15557);
xnor U15718 (N_15718,N_15243,N_15259);
xor U15719 (N_15719,N_15328,N_15427);
xor U15720 (N_15720,N_15256,N_15385);
and U15721 (N_15721,N_15290,N_15473);
xor U15722 (N_15722,N_15516,N_15468);
nor U15723 (N_15723,N_15324,N_15276);
nor U15724 (N_15724,N_15496,N_15330);
nor U15725 (N_15725,N_15280,N_15333);
nor U15726 (N_15726,N_15558,N_15361);
and U15727 (N_15727,N_15411,N_15517);
and U15728 (N_15728,N_15559,N_15587);
xor U15729 (N_15729,N_15451,N_15255);
xnor U15730 (N_15730,N_15398,N_15439);
nand U15731 (N_15731,N_15289,N_15462);
and U15732 (N_15732,N_15248,N_15404);
or U15733 (N_15733,N_15389,N_15363);
nor U15734 (N_15734,N_15285,N_15317);
and U15735 (N_15735,N_15595,N_15469);
nor U15736 (N_15736,N_15353,N_15538);
or U15737 (N_15737,N_15217,N_15542);
xor U15738 (N_15738,N_15247,N_15391);
or U15739 (N_15739,N_15270,N_15200);
nor U15740 (N_15740,N_15266,N_15580);
xnor U15741 (N_15741,N_15294,N_15511);
xnor U15742 (N_15742,N_15297,N_15322);
or U15743 (N_15743,N_15224,N_15597);
nor U15744 (N_15744,N_15384,N_15331);
or U15745 (N_15745,N_15284,N_15442);
xor U15746 (N_15746,N_15209,N_15564);
or U15747 (N_15747,N_15495,N_15267);
nor U15748 (N_15748,N_15432,N_15490);
xor U15749 (N_15749,N_15484,N_15527);
nor U15750 (N_15750,N_15275,N_15343);
xor U15751 (N_15751,N_15591,N_15295);
or U15752 (N_15752,N_15304,N_15491);
nand U15753 (N_15753,N_15327,N_15238);
nand U15754 (N_15754,N_15223,N_15594);
or U15755 (N_15755,N_15567,N_15588);
or U15756 (N_15756,N_15208,N_15421);
xor U15757 (N_15757,N_15570,N_15582);
nand U15758 (N_15758,N_15301,N_15458);
nand U15759 (N_15759,N_15262,N_15429);
xor U15760 (N_15760,N_15393,N_15529);
and U15761 (N_15761,N_15366,N_15576);
nor U15762 (N_15762,N_15344,N_15474);
xnor U15763 (N_15763,N_15268,N_15352);
and U15764 (N_15764,N_15299,N_15419);
nor U15765 (N_15765,N_15435,N_15487);
xnor U15766 (N_15766,N_15443,N_15313);
nor U15767 (N_15767,N_15464,N_15560);
or U15768 (N_15768,N_15566,N_15422);
nor U15769 (N_15769,N_15320,N_15498);
nand U15770 (N_15770,N_15351,N_15264);
xor U15771 (N_15771,N_15455,N_15543);
nand U15772 (N_15772,N_15525,N_15220);
xor U15773 (N_15773,N_15358,N_15367);
xnor U15774 (N_15774,N_15218,N_15512);
and U15775 (N_15775,N_15434,N_15354);
nand U15776 (N_15776,N_15205,N_15454);
xnor U15777 (N_15777,N_15355,N_15375);
or U15778 (N_15778,N_15292,N_15214);
nor U15779 (N_15779,N_15402,N_15575);
xor U15780 (N_15780,N_15293,N_15335);
and U15781 (N_15781,N_15334,N_15561);
nand U15782 (N_15782,N_15426,N_15371);
and U15783 (N_15783,N_15235,N_15418);
nor U15784 (N_15784,N_15234,N_15489);
or U15785 (N_15785,N_15417,N_15242);
nand U15786 (N_15786,N_15415,N_15228);
xnor U15787 (N_15787,N_15492,N_15364);
and U15788 (N_15788,N_15437,N_15568);
nand U15789 (N_15789,N_15287,N_15502);
nor U15790 (N_15790,N_15252,N_15547);
nand U15791 (N_15791,N_15210,N_15475);
xnor U15792 (N_15792,N_15221,N_15368);
nor U15793 (N_15793,N_15518,N_15479);
or U15794 (N_15794,N_15296,N_15396);
and U15795 (N_15795,N_15534,N_15307);
nand U15796 (N_15796,N_15577,N_15545);
nand U15797 (N_15797,N_15444,N_15253);
nand U15798 (N_15798,N_15399,N_15282);
nor U15799 (N_15799,N_15274,N_15372);
and U15800 (N_15800,N_15311,N_15538);
and U15801 (N_15801,N_15564,N_15508);
or U15802 (N_15802,N_15374,N_15559);
nor U15803 (N_15803,N_15501,N_15243);
xor U15804 (N_15804,N_15531,N_15353);
nor U15805 (N_15805,N_15379,N_15417);
or U15806 (N_15806,N_15347,N_15330);
nor U15807 (N_15807,N_15488,N_15245);
or U15808 (N_15808,N_15519,N_15547);
xor U15809 (N_15809,N_15399,N_15459);
and U15810 (N_15810,N_15264,N_15217);
xor U15811 (N_15811,N_15221,N_15472);
and U15812 (N_15812,N_15561,N_15230);
xnor U15813 (N_15813,N_15338,N_15459);
xnor U15814 (N_15814,N_15490,N_15503);
nand U15815 (N_15815,N_15499,N_15235);
and U15816 (N_15816,N_15541,N_15547);
and U15817 (N_15817,N_15460,N_15452);
xnor U15818 (N_15818,N_15292,N_15541);
nor U15819 (N_15819,N_15523,N_15421);
xnor U15820 (N_15820,N_15454,N_15465);
nand U15821 (N_15821,N_15392,N_15242);
nor U15822 (N_15822,N_15416,N_15475);
nor U15823 (N_15823,N_15403,N_15236);
nand U15824 (N_15824,N_15573,N_15254);
nor U15825 (N_15825,N_15394,N_15258);
nor U15826 (N_15826,N_15577,N_15451);
xnor U15827 (N_15827,N_15390,N_15354);
nand U15828 (N_15828,N_15451,N_15341);
nor U15829 (N_15829,N_15402,N_15552);
nor U15830 (N_15830,N_15323,N_15533);
nor U15831 (N_15831,N_15379,N_15364);
or U15832 (N_15832,N_15433,N_15599);
xor U15833 (N_15833,N_15552,N_15533);
nor U15834 (N_15834,N_15245,N_15456);
nand U15835 (N_15835,N_15447,N_15503);
or U15836 (N_15836,N_15445,N_15530);
nand U15837 (N_15837,N_15254,N_15596);
nand U15838 (N_15838,N_15426,N_15213);
or U15839 (N_15839,N_15261,N_15541);
nor U15840 (N_15840,N_15562,N_15542);
and U15841 (N_15841,N_15385,N_15320);
nand U15842 (N_15842,N_15421,N_15448);
nand U15843 (N_15843,N_15589,N_15548);
and U15844 (N_15844,N_15389,N_15484);
nand U15845 (N_15845,N_15592,N_15580);
or U15846 (N_15846,N_15414,N_15589);
and U15847 (N_15847,N_15385,N_15294);
and U15848 (N_15848,N_15291,N_15260);
or U15849 (N_15849,N_15406,N_15526);
and U15850 (N_15850,N_15423,N_15294);
nand U15851 (N_15851,N_15564,N_15520);
or U15852 (N_15852,N_15294,N_15311);
nor U15853 (N_15853,N_15533,N_15467);
and U15854 (N_15854,N_15279,N_15459);
nor U15855 (N_15855,N_15464,N_15471);
xor U15856 (N_15856,N_15317,N_15286);
xnor U15857 (N_15857,N_15497,N_15355);
xor U15858 (N_15858,N_15211,N_15236);
xor U15859 (N_15859,N_15366,N_15317);
xor U15860 (N_15860,N_15521,N_15285);
and U15861 (N_15861,N_15508,N_15446);
xor U15862 (N_15862,N_15459,N_15552);
or U15863 (N_15863,N_15300,N_15201);
or U15864 (N_15864,N_15384,N_15349);
nor U15865 (N_15865,N_15241,N_15368);
and U15866 (N_15866,N_15583,N_15300);
or U15867 (N_15867,N_15542,N_15564);
xor U15868 (N_15868,N_15347,N_15586);
xor U15869 (N_15869,N_15539,N_15418);
nand U15870 (N_15870,N_15330,N_15523);
xor U15871 (N_15871,N_15449,N_15590);
nor U15872 (N_15872,N_15241,N_15214);
nor U15873 (N_15873,N_15532,N_15390);
or U15874 (N_15874,N_15476,N_15321);
nand U15875 (N_15875,N_15435,N_15304);
xor U15876 (N_15876,N_15444,N_15270);
xor U15877 (N_15877,N_15495,N_15579);
and U15878 (N_15878,N_15337,N_15346);
xor U15879 (N_15879,N_15235,N_15263);
and U15880 (N_15880,N_15218,N_15234);
and U15881 (N_15881,N_15417,N_15326);
nand U15882 (N_15882,N_15520,N_15424);
xnor U15883 (N_15883,N_15428,N_15400);
nor U15884 (N_15884,N_15285,N_15237);
xnor U15885 (N_15885,N_15494,N_15392);
xnor U15886 (N_15886,N_15387,N_15431);
nand U15887 (N_15887,N_15464,N_15260);
nor U15888 (N_15888,N_15411,N_15567);
and U15889 (N_15889,N_15588,N_15235);
xor U15890 (N_15890,N_15597,N_15331);
and U15891 (N_15891,N_15426,N_15347);
nand U15892 (N_15892,N_15566,N_15417);
or U15893 (N_15893,N_15332,N_15555);
xor U15894 (N_15894,N_15547,N_15309);
nor U15895 (N_15895,N_15426,N_15589);
and U15896 (N_15896,N_15451,N_15278);
xnor U15897 (N_15897,N_15280,N_15371);
xnor U15898 (N_15898,N_15566,N_15236);
xor U15899 (N_15899,N_15255,N_15532);
xnor U15900 (N_15900,N_15287,N_15416);
nand U15901 (N_15901,N_15592,N_15219);
nand U15902 (N_15902,N_15560,N_15243);
xor U15903 (N_15903,N_15311,N_15516);
and U15904 (N_15904,N_15405,N_15342);
or U15905 (N_15905,N_15343,N_15522);
nand U15906 (N_15906,N_15352,N_15375);
nor U15907 (N_15907,N_15502,N_15489);
and U15908 (N_15908,N_15464,N_15392);
nor U15909 (N_15909,N_15595,N_15540);
nand U15910 (N_15910,N_15538,N_15453);
nor U15911 (N_15911,N_15398,N_15456);
nor U15912 (N_15912,N_15355,N_15350);
xnor U15913 (N_15913,N_15283,N_15564);
and U15914 (N_15914,N_15248,N_15399);
nor U15915 (N_15915,N_15590,N_15510);
xnor U15916 (N_15916,N_15377,N_15524);
xnor U15917 (N_15917,N_15408,N_15355);
xnor U15918 (N_15918,N_15305,N_15343);
xor U15919 (N_15919,N_15488,N_15526);
or U15920 (N_15920,N_15245,N_15214);
and U15921 (N_15921,N_15530,N_15250);
and U15922 (N_15922,N_15308,N_15564);
nor U15923 (N_15923,N_15491,N_15314);
or U15924 (N_15924,N_15357,N_15514);
nand U15925 (N_15925,N_15569,N_15572);
or U15926 (N_15926,N_15481,N_15595);
xnor U15927 (N_15927,N_15288,N_15597);
or U15928 (N_15928,N_15513,N_15541);
nor U15929 (N_15929,N_15271,N_15310);
xnor U15930 (N_15930,N_15585,N_15383);
nand U15931 (N_15931,N_15452,N_15347);
nor U15932 (N_15932,N_15423,N_15218);
nor U15933 (N_15933,N_15454,N_15498);
nor U15934 (N_15934,N_15328,N_15437);
nand U15935 (N_15935,N_15396,N_15254);
nor U15936 (N_15936,N_15486,N_15426);
nand U15937 (N_15937,N_15484,N_15203);
nor U15938 (N_15938,N_15547,N_15583);
and U15939 (N_15939,N_15283,N_15472);
xor U15940 (N_15940,N_15231,N_15220);
and U15941 (N_15941,N_15570,N_15549);
and U15942 (N_15942,N_15332,N_15401);
nand U15943 (N_15943,N_15353,N_15414);
and U15944 (N_15944,N_15410,N_15528);
and U15945 (N_15945,N_15595,N_15319);
and U15946 (N_15946,N_15299,N_15225);
and U15947 (N_15947,N_15564,N_15419);
or U15948 (N_15948,N_15279,N_15320);
xor U15949 (N_15949,N_15331,N_15395);
nor U15950 (N_15950,N_15427,N_15461);
xnor U15951 (N_15951,N_15422,N_15215);
and U15952 (N_15952,N_15590,N_15381);
nand U15953 (N_15953,N_15460,N_15359);
xnor U15954 (N_15954,N_15586,N_15224);
and U15955 (N_15955,N_15470,N_15499);
or U15956 (N_15956,N_15554,N_15549);
xor U15957 (N_15957,N_15303,N_15408);
or U15958 (N_15958,N_15289,N_15436);
or U15959 (N_15959,N_15291,N_15442);
nor U15960 (N_15960,N_15531,N_15396);
nor U15961 (N_15961,N_15577,N_15404);
and U15962 (N_15962,N_15298,N_15423);
and U15963 (N_15963,N_15472,N_15318);
nand U15964 (N_15964,N_15214,N_15534);
xnor U15965 (N_15965,N_15529,N_15532);
nand U15966 (N_15966,N_15562,N_15531);
nand U15967 (N_15967,N_15516,N_15505);
nand U15968 (N_15968,N_15268,N_15492);
and U15969 (N_15969,N_15495,N_15502);
xnor U15970 (N_15970,N_15270,N_15336);
and U15971 (N_15971,N_15471,N_15304);
or U15972 (N_15972,N_15510,N_15358);
and U15973 (N_15973,N_15248,N_15480);
or U15974 (N_15974,N_15534,N_15498);
or U15975 (N_15975,N_15437,N_15432);
nand U15976 (N_15976,N_15371,N_15524);
nand U15977 (N_15977,N_15538,N_15228);
nor U15978 (N_15978,N_15413,N_15214);
nand U15979 (N_15979,N_15560,N_15230);
xor U15980 (N_15980,N_15511,N_15442);
xnor U15981 (N_15981,N_15552,N_15564);
nor U15982 (N_15982,N_15472,N_15235);
nor U15983 (N_15983,N_15596,N_15577);
nor U15984 (N_15984,N_15242,N_15539);
nor U15985 (N_15985,N_15478,N_15207);
or U15986 (N_15986,N_15545,N_15527);
nor U15987 (N_15987,N_15467,N_15295);
and U15988 (N_15988,N_15311,N_15271);
or U15989 (N_15989,N_15573,N_15468);
nand U15990 (N_15990,N_15320,N_15359);
nor U15991 (N_15991,N_15305,N_15585);
xor U15992 (N_15992,N_15579,N_15543);
nor U15993 (N_15993,N_15485,N_15547);
and U15994 (N_15994,N_15317,N_15515);
and U15995 (N_15995,N_15567,N_15552);
xnor U15996 (N_15996,N_15252,N_15322);
and U15997 (N_15997,N_15429,N_15535);
nand U15998 (N_15998,N_15317,N_15496);
xor U15999 (N_15999,N_15581,N_15513);
xnor U16000 (N_16000,N_15954,N_15967);
and U16001 (N_16001,N_15883,N_15912);
nand U16002 (N_16002,N_15855,N_15809);
or U16003 (N_16003,N_15679,N_15794);
or U16004 (N_16004,N_15744,N_15639);
nor U16005 (N_16005,N_15745,N_15934);
nand U16006 (N_16006,N_15663,N_15825);
and U16007 (N_16007,N_15801,N_15808);
nand U16008 (N_16008,N_15987,N_15617);
nand U16009 (N_16009,N_15964,N_15765);
nand U16010 (N_16010,N_15637,N_15715);
nand U16011 (N_16011,N_15652,N_15624);
nor U16012 (N_16012,N_15780,N_15916);
nor U16013 (N_16013,N_15755,N_15648);
xnor U16014 (N_16014,N_15775,N_15701);
nand U16015 (N_16015,N_15841,N_15851);
or U16016 (N_16016,N_15820,N_15914);
nor U16017 (N_16017,N_15871,N_15710);
nand U16018 (N_16018,N_15960,N_15785);
nand U16019 (N_16019,N_15731,N_15703);
nand U16020 (N_16020,N_15892,N_15678);
and U16021 (N_16021,N_15897,N_15681);
nor U16022 (N_16022,N_15804,N_15782);
or U16023 (N_16023,N_15640,N_15784);
or U16024 (N_16024,N_15757,N_15880);
xor U16025 (N_16025,N_15781,N_15674);
xor U16026 (N_16026,N_15740,N_15935);
or U16027 (N_16027,N_15969,N_15844);
nor U16028 (N_16028,N_15848,N_15816);
and U16029 (N_16029,N_15933,N_15913);
and U16030 (N_16030,N_15682,N_15923);
xor U16031 (N_16031,N_15872,N_15698);
nand U16032 (N_16032,N_15894,N_15658);
xor U16033 (N_16033,N_15712,N_15833);
nor U16034 (N_16034,N_15846,N_15815);
nand U16035 (N_16035,N_15667,N_15948);
xor U16036 (N_16036,N_15911,N_15902);
xor U16037 (N_16037,N_15649,N_15942);
and U16038 (N_16038,N_15963,N_15749);
or U16039 (N_16039,N_15705,N_15734);
nor U16040 (N_16040,N_15994,N_15862);
nand U16041 (N_16041,N_15845,N_15773);
or U16042 (N_16042,N_15907,N_15647);
or U16043 (N_16043,N_15929,N_15978);
nand U16044 (N_16044,N_15725,N_15992);
nand U16045 (N_16045,N_15881,N_15983);
xnor U16046 (N_16046,N_15918,N_15768);
or U16047 (N_16047,N_15993,N_15664);
nand U16048 (N_16048,N_15909,N_15970);
nand U16049 (N_16049,N_15753,N_15791);
nand U16050 (N_16050,N_15974,N_15771);
xor U16051 (N_16051,N_15830,N_15870);
nor U16052 (N_16052,N_15747,N_15975);
xnor U16053 (N_16053,N_15814,N_15998);
and U16054 (N_16054,N_15899,N_15612);
nand U16055 (N_16055,N_15818,N_15921);
or U16056 (N_16056,N_15888,N_15986);
nor U16057 (N_16057,N_15843,N_15860);
nor U16058 (N_16058,N_15858,N_15671);
or U16059 (N_16059,N_15635,N_15873);
xnor U16060 (N_16060,N_15650,N_15939);
xnor U16061 (N_16061,N_15953,N_15702);
or U16062 (N_16062,N_15875,N_15854);
nor U16063 (N_16063,N_15828,N_15750);
nand U16064 (N_16064,N_15769,N_15767);
nand U16065 (N_16065,N_15877,N_15944);
nor U16066 (N_16066,N_15842,N_15932);
nor U16067 (N_16067,N_15659,N_15824);
and U16068 (N_16068,N_15866,N_15766);
and U16069 (N_16069,N_15996,N_15813);
nor U16070 (N_16070,N_15847,N_15901);
xor U16071 (N_16071,N_15850,N_15645);
nor U16072 (N_16072,N_15925,N_15979);
and U16073 (N_16073,N_15985,N_15661);
or U16074 (N_16074,N_15826,N_15945);
nor U16075 (N_16075,N_15807,N_15924);
or U16076 (N_16076,N_15643,N_15905);
or U16077 (N_16077,N_15764,N_15889);
nand U16078 (N_16078,N_15926,N_15930);
or U16079 (N_16079,N_15642,N_15603);
and U16080 (N_16080,N_15885,N_15922);
or U16081 (N_16081,N_15800,N_15938);
nand U16082 (N_16082,N_15607,N_15687);
and U16083 (N_16083,N_15633,N_15811);
and U16084 (N_16084,N_15779,N_15952);
or U16085 (N_16085,N_15604,N_15746);
or U16086 (N_16086,N_15611,N_15774);
and U16087 (N_16087,N_15721,N_15761);
and U16088 (N_16088,N_15675,N_15708);
nand U16089 (N_16089,N_15946,N_15890);
and U16090 (N_16090,N_15641,N_15623);
nor U16091 (N_16091,N_15874,N_15982);
nor U16092 (N_16092,N_15799,N_15720);
nand U16093 (N_16093,N_15699,N_15829);
and U16094 (N_16094,N_15927,N_15651);
and U16095 (N_16095,N_15758,N_15646);
and U16096 (N_16096,N_15835,N_15893);
and U16097 (N_16097,N_15751,N_15886);
or U16098 (N_16098,N_15827,N_15980);
or U16099 (N_16099,N_15989,N_15821);
nand U16100 (N_16100,N_15903,N_15704);
nand U16101 (N_16101,N_15754,N_15707);
nor U16102 (N_16102,N_15789,N_15865);
nand U16103 (N_16103,N_15692,N_15849);
and U16104 (N_16104,N_15714,N_15798);
xnor U16105 (N_16105,N_15614,N_15666);
xor U16106 (N_16106,N_15931,N_15683);
nand U16107 (N_16107,N_15962,N_15950);
and U16108 (N_16108,N_15615,N_15991);
nand U16109 (N_16109,N_15995,N_15853);
nand U16110 (N_16110,N_15680,N_15803);
or U16111 (N_16111,N_15852,N_15981);
nor U16112 (N_16112,N_15917,N_15718);
nand U16113 (N_16113,N_15997,N_15955);
nand U16114 (N_16114,N_15760,N_15752);
and U16115 (N_16115,N_15616,N_15887);
and U16116 (N_16116,N_15727,N_15920);
xnor U16117 (N_16117,N_15696,N_15786);
nand U16118 (N_16118,N_15906,N_15688);
nor U16119 (N_16119,N_15738,N_15823);
nand U16120 (N_16120,N_15869,N_15857);
nor U16121 (N_16121,N_15795,N_15961);
xor U16122 (N_16122,N_15742,N_15601);
xor U16123 (N_16123,N_15787,N_15728);
and U16124 (N_16124,N_15722,N_15672);
xor U16125 (N_16125,N_15817,N_15741);
or U16126 (N_16126,N_15943,N_15959);
or U16127 (N_16127,N_15763,N_15644);
nand U16128 (N_16128,N_15951,N_15695);
nor U16129 (N_16129,N_15977,N_15910);
nand U16130 (N_16130,N_15631,N_15729);
or U16131 (N_16131,N_15936,N_15940);
or U16132 (N_16132,N_15988,N_15622);
nand U16133 (N_16133,N_15697,N_15733);
nand U16134 (N_16134,N_15802,N_15949);
nor U16135 (N_16135,N_15837,N_15898);
or U16136 (N_16136,N_15730,N_15896);
nor U16137 (N_16137,N_15900,N_15669);
nand U16138 (N_16138,N_15717,N_15836);
xnor U16139 (N_16139,N_15610,N_15999);
and U16140 (N_16140,N_15735,N_15676);
nand U16141 (N_16141,N_15956,N_15810);
and U16142 (N_16142,N_15867,N_15976);
nor U16143 (N_16143,N_15868,N_15971);
nor U16144 (N_16144,N_15736,N_15965);
and U16145 (N_16145,N_15619,N_15632);
xnor U16146 (N_16146,N_15973,N_15891);
nor U16147 (N_16147,N_15834,N_15684);
nand U16148 (N_16148,N_15723,N_15796);
or U16149 (N_16149,N_15822,N_15777);
nand U16150 (N_16150,N_15690,N_15739);
and U16151 (N_16151,N_15693,N_15990);
or U16152 (N_16152,N_15608,N_15879);
or U16153 (N_16153,N_15831,N_15840);
nor U16154 (N_16154,N_15919,N_15762);
or U16155 (N_16155,N_15689,N_15716);
and U16156 (N_16156,N_15972,N_15941);
nor U16157 (N_16157,N_15878,N_15668);
and U16158 (N_16158,N_15605,N_15806);
nor U16159 (N_16159,N_15984,N_15904);
nor U16160 (N_16160,N_15819,N_15737);
and U16161 (N_16161,N_15685,N_15856);
xor U16162 (N_16162,N_15947,N_15620);
or U16163 (N_16163,N_15694,N_15861);
and U16164 (N_16164,N_15621,N_15602);
or U16165 (N_16165,N_15653,N_15662);
or U16166 (N_16166,N_15613,N_15792);
and U16167 (N_16167,N_15609,N_15958);
nand U16168 (N_16168,N_15636,N_15859);
or U16169 (N_16169,N_15719,N_15797);
and U16170 (N_16170,N_15957,N_15638);
xor U16171 (N_16171,N_15625,N_15724);
and U16172 (N_16172,N_15776,N_15627);
or U16173 (N_16173,N_15706,N_15673);
nor U16174 (N_16174,N_15743,N_15634);
or U16175 (N_16175,N_15790,N_15618);
nand U16176 (N_16176,N_15691,N_15838);
and U16177 (N_16177,N_15606,N_15783);
or U16178 (N_16178,N_15772,N_15630);
nor U16179 (N_16179,N_15839,N_15805);
xnor U16180 (N_16180,N_15686,N_15660);
or U16181 (N_16181,N_15793,N_15732);
xnor U16182 (N_16182,N_15968,N_15876);
nor U16183 (N_16183,N_15759,N_15863);
or U16184 (N_16184,N_15928,N_15657);
nor U16185 (N_16185,N_15915,N_15700);
and U16186 (N_16186,N_15756,N_15628);
nor U16187 (N_16187,N_15884,N_15600);
or U16188 (N_16188,N_15670,N_15726);
xor U16189 (N_16189,N_15908,N_15895);
or U16190 (N_16190,N_15812,N_15966);
xor U16191 (N_16191,N_15788,N_15832);
nor U16192 (N_16192,N_15626,N_15770);
xor U16193 (N_16193,N_15677,N_15864);
or U16194 (N_16194,N_15778,N_15748);
nand U16195 (N_16195,N_15711,N_15665);
or U16196 (N_16196,N_15882,N_15656);
nor U16197 (N_16197,N_15713,N_15654);
and U16198 (N_16198,N_15655,N_15629);
xnor U16199 (N_16199,N_15937,N_15709);
xnor U16200 (N_16200,N_15756,N_15856);
xor U16201 (N_16201,N_15748,N_15702);
nand U16202 (N_16202,N_15674,N_15929);
and U16203 (N_16203,N_15934,N_15997);
xor U16204 (N_16204,N_15693,N_15764);
xor U16205 (N_16205,N_15899,N_15735);
nor U16206 (N_16206,N_15794,N_15969);
nand U16207 (N_16207,N_15857,N_15742);
xor U16208 (N_16208,N_15691,N_15745);
xnor U16209 (N_16209,N_15653,N_15903);
nor U16210 (N_16210,N_15839,N_15876);
or U16211 (N_16211,N_15897,N_15785);
and U16212 (N_16212,N_15626,N_15722);
nor U16213 (N_16213,N_15665,N_15765);
and U16214 (N_16214,N_15669,N_15906);
nor U16215 (N_16215,N_15886,N_15749);
or U16216 (N_16216,N_15807,N_15904);
and U16217 (N_16217,N_15967,N_15635);
nand U16218 (N_16218,N_15645,N_15631);
or U16219 (N_16219,N_15623,N_15835);
xor U16220 (N_16220,N_15900,N_15616);
nand U16221 (N_16221,N_15758,N_15608);
nor U16222 (N_16222,N_15803,N_15741);
nand U16223 (N_16223,N_15922,N_15914);
nand U16224 (N_16224,N_15617,N_15867);
nand U16225 (N_16225,N_15622,N_15964);
nor U16226 (N_16226,N_15948,N_15973);
or U16227 (N_16227,N_15608,N_15907);
or U16228 (N_16228,N_15767,N_15825);
or U16229 (N_16229,N_15624,N_15986);
and U16230 (N_16230,N_15955,N_15954);
nand U16231 (N_16231,N_15743,N_15732);
or U16232 (N_16232,N_15614,N_15879);
xnor U16233 (N_16233,N_15712,N_15776);
or U16234 (N_16234,N_15952,N_15733);
or U16235 (N_16235,N_15855,N_15627);
and U16236 (N_16236,N_15759,N_15753);
and U16237 (N_16237,N_15657,N_15897);
xor U16238 (N_16238,N_15930,N_15959);
or U16239 (N_16239,N_15880,N_15756);
or U16240 (N_16240,N_15797,N_15971);
xnor U16241 (N_16241,N_15936,N_15613);
nor U16242 (N_16242,N_15638,N_15662);
xor U16243 (N_16243,N_15934,N_15907);
xor U16244 (N_16244,N_15964,N_15950);
or U16245 (N_16245,N_15899,N_15685);
or U16246 (N_16246,N_15643,N_15960);
xor U16247 (N_16247,N_15755,N_15621);
or U16248 (N_16248,N_15807,N_15894);
nand U16249 (N_16249,N_15611,N_15708);
xnor U16250 (N_16250,N_15841,N_15708);
nor U16251 (N_16251,N_15703,N_15919);
nand U16252 (N_16252,N_15993,N_15758);
nor U16253 (N_16253,N_15890,N_15936);
xor U16254 (N_16254,N_15630,N_15849);
and U16255 (N_16255,N_15733,N_15975);
nor U16256 (N_16256,N_15683,N_15662);
nand U16257 (N_16257,N_15604,N_15945);
nor U16258 (N_16258,N_15933,N_15819);
and U16259 (N_16259,N_15769,N_15793);
nand U16260 (N_16260,N_15642,N_15651);
xor U16261 (N_16261,N_15758,N_15870);
nor U16262 (N_16262,N_15675,N_15827);
nand U16263 (N_16263,N_15741,N_15840);
nand U16264 (N_16264,N_15717,N_15788);
nand U16265 (N_16265,N_15709,N_15958);
xnor U16266 (N_16266,N_15860,N_15676);
and U16267 (N_16267,N_15902,N_15966);
nor U16268 (N_16268,N_15803,N_15907);
or U16269 (N_16269,N_15885,N_15932);
nor U16270 (N_16270,N_15689,N_15690);
or U16271 (N_16271,N_15683,N_15737);
nand U16272 (N_16272,N_15958,N_15887);
and U16273 (N_16273,N_15831,N_15712);
or U16274 (N_16274,N_15808,N_15981);
and U16275 (N_16275,N_15807,N_15952);
and U16276 (N_16276,N_15634,N_15956);
and U16277 (N_16277,N_15786,N_15827);
and U16278 (N_16278,N_15996,N_15935);
or U16279 (N_16279,N_15851,N_15995);
or U16280 (N_16280,N_15923,N_15606);
xnor U16281 (N_16281,N_15626,N_15930);
xnor U16282 (N_16282,N_15979,N_15920);
nand U16283 (N_16283,N_15690,N_15943);
and U16284 (N_16284,N_15628,N_15870);
xor U16285 (N_16285,N_15891,N_15864);
xnor U16286 (N_16286,N_15795,N_15744);
or U16287 (N_16287,N_15891,N_15931);
nor U16288 (N_16288,N_15746,N_15703);
nor U16289 (N_16289,N_15886,N_15721);
xnor U16290 (N_16290,N_15857,N_15660);
nor U16291 (N_16291,N_15968,N_15770);
or U16292 (N_16292,N_15914,N_15713);
or U16293 (N_16293,N_15635,N_15869);
or U16294 (N_16294,N_15861,N_15936);
or U16295 (N_16295,N_15988,N_15803);
or U16296 (N_16296,N_15621,N_15802);
xor U16297 (N_16297,N_15975,N_15636);
nand U16298 (N_16298,N_15938,N_15631);
xnor U16299 (N_16299,N_15753,N_15957);
nor U16300 (N_16300,N_15629,N_15941);
nor U16301 (N_16301,N_15737,N_15930);
xor U16302 (N_16302,N_15995,N_15761);
or U16303 (N_16303,N_15801,N_15932);
and U16304 (N_16304,N_15952,N_15944);
or U16305 (N_16305,N_15781,N_15922);
or U16306 (N_16306,N_15618,N_15878);
nand U16307 (N_16307,N_15747,N_15656);
and U16308 (N_16308,N_15841,N_15799);
or U16309 (N_16309,N_15869,N_15932);
and U16310 (N_16310,N_15820,N_15972);
xor U16311 (N_16311,N_15606,N_15793);
xor U16312 (N_16312,N_15915,N_15724);
and U16313 (N_16313,N_15813,N_15934);
nor U16314 (N_16314,N_15936,N_15826);
nor U16315 (N_16315,N_15838,N_15930);
nor U16316 (N_16316,N_15628,N_15885);
xnor U16317 (N_16317,N_15625,N_15734);
and U16318 (N_16318,N_15961,N_15779);
xor U16319 (N_16319,N_15831,N_15694);
nor U16320 (N_16320,N_15716,N_15910);
and U16321 (N_16321,N_15623,N_15805);
and U16322 (N_16322,N_15658,N_15791);
or U16323 (N_16323,N_15957,N_15844);
xnor U16324 (N_16324,N_15747,N_15701);
xnor U16325 (N_16325,N_15895,N_15727);
nand U16326 (N_16326,N_15701,N_15825);
nand U16327 (N_16327,N_15910,N_15991);
nand U16328 (N_16328,N_15654,N_15956);
and U16329 (N_16329,N_15921,N_15760);
or U16330 (N_16330,N_15776,N_15876);
nor U16331 (N_16331,N_15958,N_15771);
xnor U16332 (N_16332,N_15813,N_15792);
or U16333 (N_16333,N_15877,N_15778);
nand U16334 (N_16334,N_15990,N_15605);
xor U16335 (N_16335,N_15791,N_15879);
nand U16336 (N_16336,N_15861,N_15783);
nor U16337 (N_16337,N_15737,N_15865);
xnor U16338 (N_16338,N_15611,N_15661);
nor U16339 (N_16339,N_15878,N_15917);
nor U16340 (N_16340,N_15692,N_15909);
nand U16341 (N_16341,N_15735,N_15631);
or U16342 (N_16342,N_15822,N_15799);
nand U16343 (N_16343,N_15735,N_15834);
nand U16344 (N_16344,N_15713,N_15784);
nand U16345 (N_16345,N_15696,N_15985);
nand U16346 (N_16346,N_15626,N_15773);
nand U16347 (N_16347,N_15975,N_15658);
or U16348 (N_16348,N_15834,N_15836);
or U16349 (N_16349,N_15634,N_15823);
nand U16350 (N_16350,N_15792,N_15612);
nor U16351 (N_16351,N_15991,N_15697);
and U16352 (N_16352,N_15987,N_15910);
nand U16353 (N_16353,N_15704,N_15707);
nor U16354 (N_16354,N_15884,N_15638);
nand U16355 (N_16355,N_15629,N_15862);
nor U16356 (N_16356,N_15990,N_15831);
nand U16357 (N_16357,N_15714,N_15661);
xnor U16358 (N_16358,N_15776,N_15771);
xor U16359 (N_16359,N_15935,N_15941);
nor U16360 (N_16360,N_15952,N_15712);
or U16361 (N_16361,N_15622,N_15870);
and U16362 (N_16362,N_15940,N_15868);
or U16363 (N_16363,N_15833,N_15834);
nor U16364 (N_16364,N_15644,N_15815);
and U16365 (N_16365,N_15723,N_15645);
or U16366 (N_16366,N_15632,N_15794);
nor U16367 (N_16367,N_15861,N_15623);
nor U16368 (N_16368,N_15860,N_15985);
nor U16369 (N_16369,N_15851,N_15731);
xor U16370 (N_16370,N_15861,N_15699);
nand U16371 (N_16371,N_15630,N_15688);
and U16372 (N_16372,N_15695,N_15730);
xor U16373 (N_16373,N_15666,N_15913);
nor U16374 (N_16374,N_15710,N_15813);
xnor U16375 (N_16375,N_15788,N_15964);
xnor U16376 (N_16376,N_15925,N_15924);
nand U16377 (N_16377,N_15623,N_15893);
nand U16378 (N_16378,N_15838,N_15955);
xor U16379 (N_16379,N_15656,N_15716);
nor U16380 (N_16380,N_15616,N_15994);
nor U16381 (N_16381,N_15766,N_15954);
nand U16382 (N_16382,N_15812,N_15618);
nand U16383 (N_16383,N_15623,N_15833);
nand U16384 (N_16384,N_15786,N_15816);
or U16385 (N_16385,N_15689,N_15958);
nand U16386 (N_16386,N_15627,N_15991);
nand U16387 (N_16387,N_15699,N_15849);
and U16388 (N_16388,N_15885,N_15826);
xnor U16389 (N_16389,N_15951,N_15703);
nor U16390 (N_16390,N_15835,N_15749);
nand U16391 (N_16391,N_15668,N_15792);
xor U16392 (N_16392,N_15917,N_15724);
or U16393 (N_16393,N_15902,N_15760);
xnor U16394 (N_16394,N_15758,N_15975);
and U16395 (N_16395,N_15761,N_15737);
or U16396 (N_16396,N_15807,N_15715);
xor U16397 (N_16397,N_15729,N_15835);
or U16398 (N_16398,N_15744,N_15904);
and U16399 (N_16399,N_15866,N_15797);
and U16400 (N_16400,N_16228,N_16388);
nand U16401 (N_16401,N_16362,N_16106);
and U16402 (N_16402,N_16205,N_16146);
nand U16403 (N_16403,N_16119,N_16132);
nor U16404 (N_16404,N_16216,N_16347);
nand U16405 (N_16405,N_16313,N_16239);
nor U16406 (N_16406,N_16312,N_16316);
nand U16407 (N_16407,N_16217,N_16315);
and U16408 (N_16408,N_16286,N_16369);
xnor U16409 (N_16409,N_16270,N_16298);
xor U16410 (N_16410,N_16066,N_16279);
and U16411 (N_16411,N_16337,N_16248);
and U16412 (N_16412,N_16116,N_16361);
nand U16413 (N_16413,N_16135,N_16189);
xnor U16414 (N_16414,N_16044,N_16301);
or U16415 (N_16415,N_16272,N_16215);
or U16416 (N_16416,N_16084,N_16012);
nand U16417 (N_16417,N_16187,N_16077);
nand U16418 (N_16418,N_16173,N_16280);
xor U16419 (N_16419,N_16114,N_16193);
nor U16420 (N_16420,N_16399,N_16240);
nand U16421 (N_16421,N_16037,N_16092);
nor U16422 (N_16422,N_16054,N_16294);
nor U16423 (N_16423,N_16328,N_16167);
and U16424 (N_16424,N_16107,N_16224);
nand U16425 (N_16425,N_16250,N_16276);
nand U16426 (N_16426,N_16214,N_16262);
xor U16427 (N_16427,N_16039,N_16147);
nand U16428 (N_16428,N_16290,N_16111);
nor U16429 (N_16429,N_16389,N_16023);
nand U16430 (N_16430,N_16178,N_16082);
nor U16431 (N_16431,N_16201,N_16257);
or U16432 (N_16432,N_16245,N_16220);
and U16433 (N_16433,N_16303,N_16018);
nor U16434 (N_16434,N_16297,N_16287);
and U16435 (N_16435,N_16052,N_16199);
or U16436 (N_16436,N_16050,N_16309);
nor U16437 (N_16437,N_16295,N_16035);
and U16438 (N_16438,N_16078,N_16324);
nor U16439 (N_16439,N_16380,N_16058);
xnor U16440 (N_16440,N_16252,N_16184);
nand U16441 (N_16441,N_16273,N_16293);
and U16442 (N_16442,N_16096,N_16393);
and U16443 (N_16443,N_16013,N_16055);
nand U16444 (N_16444,N_16153,N_16382);
and U16445 (N_16445,N_16125,N_16271);
xor U16446 (N_16446,N_16289,N_16182);
and U16447 (N_16447,N_16152,N_16000);
nor U16448 (N_16448,N_16005,N_16233);
xor U16449 (N_16449,N_16376,N_16100);
and U16450 (N_16450,N_16083,N_16129);
or U16451 (N_16451,N_16230,N_16306);
nor U16452 (N_16452,N_16001,N_16069);
xor U16453 (N_16453,N_16063,N_16318);
xor U16454 (N_16454,N_16260,N_16232);
or U16455 (N_16455,N_16340,N_16336);
or U16456 (N_16456,N_16350,N_16198);
xor U16457 (N_16457,N_16317,N_16162);
nand U16458 (N_16458,N_16020,N_16138);
and U16459 (N_16459,N_16086,N_16091);
nand U16460 (N_16460,N_16166,N_16397);
or U16461 (N_16461,N_16164,N_16075);
xnor U16462 (N_16462,N_16131,N_16163);
or U16463 (N_16463,N_16265,N_16379);
or U16464 (N_16464,N_16145,N_16115);
and U16465 (N_16465,N_16211,N_16149);
nor U16466 (N_16466,N_16275,N_16219);
and U16467 (N_16467,N_16103,N_16356);
or U16468 (N_16468,N_16113,N_16081);
and U16469 (N_16469,N_16108,N_16170);
or U16470 (N_16470,N_16383,N_16177);
and U16471 (N_16471,N_16259,N_16367);
nand U16472 (N_16472,N_16057,N_16156);
nor U16473 (N_16473,N_16181,N_16112);
xor U16474 (N_16474,N_16142,N_16266);
nor U16475 (N_16475,N_16141,N_16323);
xor U16476 (N_16476,N_16033,N_16034);
nor U16477 (N_16477,N_16355,N_16067);
or U16478 (N_16478,N_16028,N_16030);
and U16479 (N_16479,N_16253,N_16038);
nor U16480 (N_16480,N_16196,N_16237);
nand U16481 (N_16481,N_16004,N_16386);
xnor U16482 (N_16482,N_16049,N_16352);
and U16483 (N_16483,N_16200,N_16174);
and U16484 (N_16484,N_16026,N_16263);
nor U16485 (N_16485,N_16104,N_16056);
or U16486 (N_16486,N_16311,N_16330);
and U16487 (N_16487,N_16094,N_16226);
nand U16488 (N_16488,N_16148,N_16090);
nor U16489 (N_16489,N_16172,N_16251);
or U16490 (N_16490,N_16321,N_16308);
nand U16491 (N_16491,N_16365,N_16015);
and U16492 (N_16492,N_16314,N_16267);
nand U16493 (N_16493,N_16209,N_16042);
nor U16494 (N_16494,N_16009,N_16274);
nor U16495 (N_16495,N_16025,N_16344);
or U16496 (N_16496,N_16207,N_16333);
nand U16497 (N_16497,N_16045,N_16194);
nand U16498 (N_16498,N_16264,N_16281);
or U16499 (N_16499,N_16068,N_16006);
nor U16500 (N_16500,N_16307,N_16246);
or U16501 (N_16501,N_16368,N_16171);
and U16502 (N_16502,N_16041,N_16351);
and U16503 (N_16503,N_16175,N_16121);
xnor U16504 (N_16504,N_16398,N_16123);
xnor U16505 (N_16505,N_16243,N_16073);
or U16506 (N_16506,N_16032,N_16024);
and U16507 (N_16507,N_16176,N_16169);
nand U16508 (N_16508,N_16190,N_16338);
xnor U16509 (N_16509,N_16059,N_16305);
and U16510 (N_16510,N_16358,N_16047);
or U16511 (N_16511,N_16375,N_16366);
or U16512 (N_16512,N_16016,N_16332);
nor U16513 (N_16513,N_16341,N_16140);
and U16514 (N_16514,N_16359,N_16291);
xor U16515 (N_16515,N_16095,N_16019);
nand U16516 (N_16516,N_16124,N_16097);
or U16517 (N_16517,N_16255,N_16225);
xnor U16518 (N_16518,N_16109,N_16165);
nand U16519 (N_16519,N_16102,N_16343);
nor U16520 (N_16520,N_16364,N_16269);
or U16521 (N_16521,N_16010,N_16371);
or U16522 (N_16522,N_16160,N_16377);
or U16523 (N_16523,N_16210,N_16051);
nand U16524 (N_16524,N_16168,N_16229);
or U16525 (N_16525,N_16322,N_16342);
xor U16526 (N_16526,N_16085,N_16234);
xnor U16527 (N_16527,N_16186,N_16254);
nor U16528 (N_16528,N_16180,N_16285);
nor U16529 (N_16529,N_16335,N_16122);
and U16530 (N_16530,N_16249,N_16278);
nand U16531 (N_16531,N_16161,N_16372);
or U16532 (N_16532,N_16238,N_16325);
or U16533 (N_16533,N_16204,N_16282);
nor U16534 (N_16534,N_16357,N_16076);
nand U16535 (N_16535,N_16284,N_16222);
xnor U16536 (N_16536,N_16060,N_16195);
nor U16537 (N_16537,N_16208,N_16394);
nor U16538 (N_16538,N_16299,N_16391);
xor U16539 (N_16539,N_16021,N_16319);
and U16540 (N_16540,N_16374,N_16370);
nand U16541 (N_16541,N_16070,N_16089);
xor U16542 (N_16542,N_16133,N_16071);
xnor U16543 (N_16543,N_16137,N_16256);
or U16544 (N_16544,N_16191,N_16065);
nand U16545 (N_16545,N_16158,N_16244);
and U16546 (N_16546,N_16247,N_16017);
nor U16547 (N_16547,N_16292,N_16043);
and U16548 (N_16548,N_16353,N_16144);
nor U16549 (N_16549,N_16345,N_16079);
nor U16550 (N_16550,N_16062,N_16188);
nor U16551 (N_16551,N_16088,N_16373);
nor U16552 (N_16552,N_16395,N_16157);
nand U16553 (N_16553,N_16346,N_16130);
or U16554 (N_16554,N_16022,N_16101);
nand U16555 (N_16555,N_16046,N_16212);
nor U16556 (N_16556,N_16304,N_16128);
nor U16557 (N_16557,N_16331,N_16185);
or U16558 (N_16558,N_16011,N_16098);
xor U16559 (N_16559,N_16348,N_16136);
nand U16560 (N_16560,N_16036,N_16258);
nor U16561 (N_16561,N_16143,N_16002);
nand U16562 (N_16562,N_16218,N_16151);
nand U16563 (N_16563,N_16048,N_16320);
nor U16564 (N_16564,N_16003,N_16105);
nor U16565 (N_16565,N_16110,N_16339);
or U16566 (N_16566,N_16392,N_16329);
and U16567 (N_16567,N_16093,N_16014);
nand U16568 (N_16568,N_16213,N_16029);
nand U16569 (N_16569,N_16227,N_16360);
and U16570 (N_16570,N_16235,N_16378);
nor U16571 (N_16571,N_16390,N_16087);
or U16572 (N_16572,N_16288,N_16302);
or U16573 (N_16573,N_16126,N_16007);
or U16574 (N_16574,N_16118,N_16349);
and U16575 (N_16575,N_16064,N_16179);
or U16576 (N_16576,N_16221,N_16242);
nand U16577 (N_16577,N_16202,N_16053);
nor U16578 (N_16578,N_16223,N_16354);
and U16579 (N_16579,N_16327,N_16139);
and U16580 (N_16580,N_16159,N_16261);
xnor U16581 (N_16581,N_16074,N_16150);
nor U16582 (N_16582,N_16206,N_16099);
nand U16583 (N_16583,N_16385,N_16384);
or U16584 (N_16584,N_16236,N_16300);
nor U16585 (N_16585,N_16203,N_16396);
nor U16586 (N_16586,N_16040,N_16197);
or U16587 (N_16587,N_16326,N_16154);
nand U16588 (N_16588,N_16381,N_16155);
nor U16589 (N_16589,N_16387,N_16183);
nor U16590 (N_16590,N_16061,N_16027);
nor U16591 (N_16591,N_16363,N_16231);
and U16592 (N_16592,N_16296,N_16031);
or U16593 (N_16593,N_16127,N_16008);
and U16594 (N_16594,N_16268,N_16080);
xor U16595 (N_16595,N_16283,N_16117);
xor U16596 (N_16596,N_16334,N_16120);
nand U16597 (N_16597,N_16192,N_16072);
and U16598 (N_16598,N_16310,N_16277);
or U16599 (N_16599,N_16241,N_16134);
xor U16600 (N_16600,N_16367,N_16298);
nor U16601 (N_16601,N_16397,N_16034);
nand U16602 (N_16602,N_16351,N_16313);
nand U16603 (N_16603,N_16371,N_16255);
and U16604 (N_16604,N_16115,N_16363);
nor U16605 (N_16605,N_16286,N_16392);
xor U16606 (N_16606,N_16100,N_16005);
and U16607 (N_16607,N_16389,N_16026);
nor U16608 (N_16608,N_16341,N_16295);
and U16609 (N_16609,N_16146,N_16273);
and U16610 (N_16610,N_16226,N_16015);
and U16611 (N_16611,N_16097,N_16296);
nor U16612 (N_16612,N_16281,N_16378);
nor U16613 (N_16613,N_16224,N_16395);
xor U16614 (N_16614,N_16103,N_16168);
or U16615 (N_16615,N_16320,N_16085);
and U16616 (N_16616,N_16179,N_16309);
and U16617 (N_16617,N_16081,N_16287);
xnor U16618 (N_16618,N_16183,N_16312);
or U16619 (N_16619,N_16279,N_16036);
or U16620 (N_16620,N_16029,N_16066);
and U16621 (N_16621,N_16362,N_16147);
or U16622 (N_16622,N_16220,N_16382);
or U16623 (N_16623,N_16014,N_16303);
and U16624 (N_16624,N_16232,N_16209);
xnor U16625 (N_16625,N_16189,N_16026);
and U16626 (N_16626,N_16197,N_16316);
nor U16627 (N_16627,N_16324,N_16390);
or U16628 (N_16628,N_16060,N_16031);
nand U16629 (N_16629,N_16034,N_16024);
and U16630 (N_16630,N_16359,N_16305);
xnor U16631 (N_16631,N_16227,N_16048);
and U16632 (N_16632,N_16083,N_16143);
nand U16633 (N_16633,N_16264,N_16243);
xnor U16634 (N_16634,N_16094,N_16350);
and U16635 (N_16635,N_16152,N_16043);
nand U16636 (N_16636,N_16148,N_16304);
or U16637 (N_16637,N_16373,N_16184);
xor U16638 (N_16638,N_16035,N_16164);
nand U16639 (N_16639,N_16136,N_16176);
xor U16640 (N_16640,N_16390,N_16145);
nor U16641 (N_16641,N_16049,N_16310);
nor U16642 (N_16642,N_16007,N_16257);
nor U16643 (N_16643,N_16291,N_16148);
or U16644 (N_16644,N_16111,N_16351);
xnor U16645 (N_16645,N_16205,N_16196);
nor U16646 (N_16646,N_16084,N_16211);
or U16647 (N_16647,N_16397,N_16172);
nor U16648 (N_16648,N_16172,N_16162);
nand U16649 (N_16649,N_16145,N_16070);
xnor U16650 (N_16650,N_16136,N_16153);
xor U16651 (N_16651,N_16036,N_16029);
nor U16652 (N_16652,N_16300,N_16112);
nor U16653 (N_16653,N_16141,N_16368);
and U16654 (N_16654,N_16242,N_16011);
or U16655 (N_16655,N_16148,N_16294);
nor U16656 (N_16656,N_16394,N_16357);
xor U16657 (N_16657,N_16398,N_16147);
xor U16658 (N_16658,N_16086,N_16093);
nor U16659 (N_16659,N_16336,N_16248);
nand U16660 (N_16660,N_16060,N_16247);
nand U16661 (N_16661,N_16176,N_16364);
and U16662 (N_16662,N_16213,N_16382);
or U16663 (N_16663,N_16164,N_16196);
xor U16664 (N_16664,N_16180,N_16233);
or U16665 (N_16665,N_16235,N_16215);
and U16666 (N_16666,N_16035,N_16155);
or U16667 (N_16667,N_16212,N_16076);
xnor U16668 (N_16668,N_16230,N_16214);
or U16669 (N_16669,N_16035,N_16233);
or U16670 (N_16670,N_16287,N_16289);
or U16671 (N_16671,N_16209,N_16106);
and U16672 (N_16672,N_16283,N_16191);
xnor U16673 (N_16673,N_16080,N_16018);
nor U16674 (N_16674,N_16330,N_16050);
and U16675 (N_16675,N_16002,N_16204);
and U16676 (N_16676,N_16318,N_16202);
nand U16677 (N_16677,N_16136,N_16160);
nand U16678 (N_16678,N_16138,N_16081);
nor U16679 (N_16679,N_16237,N_16101);
nor U16680 (N_16680,N_16369,N_16382);
xor U16681 (N_16681,N_16292,N_16030);
nand U16682 (N_16682,N_16130,N_16273);
nand U16683 (N_16683,N_16352,N_16280);
or U16684 (N_16684,N_16280,N_16186);
or U16685 (N_16685,N_16113,N_16021);
and U16686 (N_16686,N_16247,N_16368);
nand U16687 (N_16687,N_16094,N_16198);
xor U16688 (N_16688,N_16024,N_16019);
xnor U16689 (N_16689,N_16069,N_16396);
and U16690 (N_16690,N_16139,N_16068);
nor U16691 (N_16691,N_16038,N_16087);
or U16692 (N_16692,N_16190,N_16195);
xnor U16693 (N_16693,N_16185,N_16223);
nor U16694 (N_16694,N_16045,N_16238);
or U16695 (N_16695,N_16292,N_16006);
xor U16696 (N_16696,N_16070,N_16020);
or U16697 (N_16697,N_16003,N_16301);
and U16698 (N_16698,N_16170,N_16122);
xnor U16699 (N_16699,N_16049,N_16271);
nor U16700 (N_16700,N_16209,N_16145);
xor U16701 (N_16701,N_16044,N_16345);
nor U16702 (N_16702,N_16194,N_16321);
or U16703 (N_16703,N_16156,N_16113);
or U16704 (N_16704,N_16244,N_16188);
nand U16705 (N_16705,N_16110,N_16234);
or U16706 (N_16706,N_16014,N_16244);
nand U16707 (N_16707,N_16096,N_16368);
nand U16708 (N_16708,N_16046,N_16035);
or U16709 (N_16709,N_16354,N_16102);
or U16710 (N_16710,N_16272,N_16117);
xnor U16711 (N_16711,N_16035,N_16080);
nand U16712 (N_16712,N_16001,N_16058);
nor U16713 (N_16713,N_16169,N_16398);
nand U16714 (N_16714,N_16105,N_16194);
or U16715 (N_16715,N_16335,N_16153);
nand U16716 (N_16716,N_16200,N_16328);
xor U16717 (N_16717,N_16200,N_16111);
xor U16718 (N_16718,N_16022,N_16160);
xor U16719 (N_16719,N_16104,N_16268);
or U16720 (N_16720,N_16080,N_16065);
and U16721 (N_16721,N_16377,N_16262);
nor U16722 (N_16722,N_16171,N_16193);
xnor U16723 (N_16723,N_16104,N_16321);
xnor U16724 (N_16724,N_16347,N_16327);
or U16725 (N_16725,N_16316,N_16307);
or U16726 (N_16726,N_16167,N_16169);
or U16727 (N_16727,N_16358,N_16349);
nand U16728 (N_16728,N_16367,N_16315);
or U16729 (N_16729,N_16328,N_16162);
xnor U16730 (N_16730,N_16344,N_16129);
xnor U16731 (N_16731,N_16239,N_16086);
and U16732 (N_16732,N_16141,N_16146);
xnor U16733 (N_16733,N_16075,N_16190);
nand U16734 (N_16734,N_16193,N_16014);
or U16735 (N_16735,N_16222,N_16231);
and U16736 (N_16736,N_16104,N_16091);
or U16737 (N_16737,N_16316,N_16053);
nand U16738 (N_16738,N_16169,N_16070);
and U16739 (N_16739,N_16069,N_16188);
or U16740 (N_16740,N_16332,N_16305);
nor U16741 (N_16741,N_16286,N_16383);
or U16742 (N_16742,N_16065,N_16368);
nor U16743 (N_16743,N_16138,N_16234);
nand U16744 (N_16744,N_16152,N_16322);
nand U16745 (N_16745,N_16009,N_16257);
or U16746 (N_16746,N_16263,N_16007);
nor U16747 (N_16747,N_16255,N_16132);
and U16748 (N_16748,N_16313,N_16219);
nor U16749 (N_16749,N_16295,N_16005);
and U16750 (N_16750,N_16176,N_16156);
and U16751 (N_16751,N_16200,N_16093);
or U16752 (N_16752,N_16342,N_16183);
nor U16753 (N_16753,N_16010,N_16222);
xnor U16754 (N_16754,N_16099,N_16202);
nand U16755 (N_16755,N_16051,N_16239);
nand U16756 (N_16756,N_16086,N_16032);
or U16757 (N_16757,N_16261,N_16395);
or U16758 (N_16758,N_16182,N_16321);
or U16759 (N_16759,N_16173,N_16377);
or U16760 (N_16760,N_16243,N_16070);
or U16761 (N_16761,N_16314,N_16373);
nor U16762 (N_16762,N_16133,N_16124);
and U16763 (N_16763,N_16252,N_16110);
or U16764 (N_16764,N_16363,N_16118);
nor U16765 (N_16765,N_16175,N_16283);
xor U16766 (N_16766,N_16212,N_16178);
nand U16767 (N_16767,N_16217,N_16231);
or U16768 (N_16768,N_16223,N_16391);
xor U16769 (N_16769,N_16215,N_16024);
or U16770 (N_16770,N_16169,N_16310);
and U16771 (N_16771,N_16317,N_16256);
nand U16772 (N_16772,N_16357,N_16007);
nand U16773 (N_16773,N_16019,N_16109);
xnor U16774 (N_16774,N_16219,N_16260);
nand U16775 (N_16775,N_16027,N_16118);
or U16776 (N_16776,N_16249,N_16361);
nand U16777 (N_16777,N_16020,N_16349);
and U16778 (N_16778,N_16179,N_16368);
nor U16779 (N_16779,N_16045,N_16253);
xnor U16780 (N_16780,N_16210,N_16300);
and U16781 (N_16781,N_16134,N_16159);
nand U16782 (N_16782,N_16117,N_16252);
nor U16783 (N_16783,N_16359,N_16083);
and U16784 (N_16784,N_16354,N_16326);
nand U16785 (N_16785,N_16132,N_16229);
nor U16786 (N_16786,N_16334,N_16056);
nor U16787 (N_16787,N_16137,N_16161);
xor U16788 (N_16788,N_16136,N_16291);
xnor U16789 (N_16789,N_16053,N_16190);
nor U16790 (N_16790,N_16091,N_16024);
and U16791 (N_16791,N_16358,N_16299);
or U16792 (N_16792,N_16197,N_16213);
nor U16793 (N_16793,N_16066,N_16179);
nor U16794 (N_16794,N_16369,N_16053);
nand U16795 (N_16795,N_16287,N_16150);
nand U16796 (N_16796,N_16175,N_16007);
or U16797 (N_16797,N_16165,N_16322);
nor U16798 (N_16798,N_16019,N_16128);
nor U16799 (N_16799,N_16150,N_16024);
nand U16800 (N_16800,N_16749,N_16486);
and U16801 (N_16801,N_16735,N_16445);
nand U16802 (N_16802,N_16415,N_16673);
nand U16803 (N_16803,N_16664,N_16513);
nor U16804 (N_16804,N_16419,N_16411);
nand U16805 (N_16805,N_16765,N_16593);
xnor U16806 (N_16806,N_16492,N_16758);
or U16807 (N_16807,N_16794,N_16518);
or U16808 (N_16808,N_16647,N_16413);
and U16809 (N_16809,N_16434,N_16549);
or U16810 (N_16810,N_16515,N_16533);
and U16811 (N_16811,N_16669,N_16550);
or U16812 (N_16812,N_16630,N_16613);
nand U16813 (N_16813,N_16626,N_16601);
nor U16814 (N_16814,N_16639,N_16611);
nor U16815 (N_16815,N_16562,N_16444);
nor U16816 (N_16816,N_16598,N_16542);
or U16817 (N_16817,N_16602,N_16430);
and U16818 (N_16818,N_16769,N_16487);
xor U16819 (N_16819,N_16529,N_16660);
and U16820 (N_16820,N_16726,N_16584);
nand U16821 (N_16821,N_16485,N_16575);
xor U16822 (N_16822,N_16561,N_16754);
and U16823 (N_16823,N_16753,N_16614);
nand U16824 (N_16824,N_16606,N_16517);
xor U16825 (N_16825,N_16576,N_16510);
or U16826 (N_16826,N_16740,N_16458);
and U16827 (N_16827,N_16460,N_16636);
nand U16828 (N_16828,N_16684,N_16648);
xor U16829 (N_16829,N_16483,N_16424);
or U16830 (N_16830,N_16632,N_16768);
and U16831 (N_16831,N_16704,N_16693);
nor U16832 (N_16832,N_16590,N_16620);
and U16833 (N_16833,N_16428,N_16470);
nor U16834 (N_16834,N_16496,N_16674);
or U16835 (N_16835,N_16642,N_16708);
xnor U16836 (N_16836,N_16464,N_16530);
or U16837 (N_16837,N_16707,N_16761);
nor U16838 (N_16838,N_16503,N_16716);
or U16839 (N_16839,N_16650,N_16617);
nor U16840 (N_16840,N_16763,N_16570);
and U16841 (N_16841,N_16766,N_16622);
or U16842 (N_16842,N_16508,N_16710);
nor U16843 (N_16843,N_16661,N_16556);
or U16844 (N_16844,N_16523,N_16423);
nor U16845 (N_16845,N_16438,N_16668);
nand U16846 (N_16846,N_16791,N_16658);
nor U16847 (N_16847,N_16680,N_16432);
or U16848 (N_16848,N_16696,N_16457);
and U16849 (N_16849,N_16686,N_16488);
and U16850 (N_16850,N_16790,N_16654);
nor U16851 (N_16851,N_16469,N_16634);
nor U16852 (N_16852,N_16578,N_16446);
and U16853 (N_16853,N_16545,N_16795);
nand U16854 (N_16854,N_16745,N_16547);
xor U16855 (N_16855,N_16682,N_16420);
nand U16856 (N_16856,N_16453,N_16551);
xnor U16857 (N_16857,N_16752,N_16425);
nand U16858 (N_16858,N_16638,N_16589);
nor U16859 (N_16859,N_16785,N_16798);
nor U16860 (N_16860,N_16709,N_16456);
or U16861 (N_16861,N_16481,N_16504);
or U16862 (N_16862,N_16454,N_16565);
or U16863 (N_16863,N_16422,N_16512);
xnor U16864 (N_16864,N_16467,N_16466);
xnor U16865 (N_16865,N_16750,N_16649);
and U16866 (N_16866,N_16499,N_16653);
nand U16867 (N_16867,N_16462,N_16706);
or U16868 (N_16868,N_16657,N_16553);
xor U16869 (N_16869,N_16776,N_16566);
xnor U16870 (N_16870,N_16463,N_16737);
xnor U16871 (N_16871,N_16646,N_16494);
or U16872 (N_16872,N_16651,N_16662);
xnor U16873 (N_16873,N_16468,N_16580);
nor U16874 (N_16874,N_16670,N_16521);
and U16875 (N_16875,N_16730,N_16641);
xnor U16876 (N_16876,N_16482,N_16500);
nor U16877 (N_16877,N_16683,N_16679);
nand U16878 (N_16878,N_16782,N_16715);
xnor U16879 (N_16879,N_16563,N_16722);
xnor U16880 (N_16880,N_16607,N_16426);
and U16881 (N_16881,N_16414,N_16448);
and U16882 (N_16882,N_16738,N_16595);
and U16883 (N_16883,N_16672,N_16472);
xor U16884 (N_16884,N_16699,N_16775);
nor U16885 (N_16885,N_16728,N_16451);
or U16886 (N_16886,N_16544,N_16605);
xnor U16887 (N_16887,N_16698,N_16506);
xor U16888 (N_16888,N_16771,N_16690);
nor U16889 (N_16889,N_16573,N_16505);
or U16890 (N_16890,N_16645,N_16748);
and U16891 (N_16891,N_16681,N_16489);
nand U16892 (N_16892,N_16408,N_16747);
nand U16893 (N_16893,N_16741,N_16703);
xor U16894 (N_16894,N_16427,N_16474);
nand U16895 (N_16895,N_16739,N_16729);
xnor U16896 (N_16896,N_16799,N_16537);
xor U16897 (N_16897,N_16461,N_16619);
or U16898 (N_16898,N_16786,N_16628);
nand U16899 (N_16899,N_16541,N_16671);
xnor U16900 (N_16900,N_16447,N_16455);
nand U16901 (N_16901,N_16498,N_16597);
or U16902 (N_16902,N_16571,N_16609);
xnor U16903 (N_16903,N_16538,N_16406);
or U16904 (N_16904,N_16600,N_16407);
xor U16905 (N_16905,N_16635,N_16585);
and U16906 (N_16906,N_16441,N_16443);
nand U16907 (N_16907,N_16519,N_16701);
nand U16908 (N_16908,N_16449,N_16582);
nor U16909 (N_16909,N_16592,N_16437);
and U16910 (N_16910,N_16579,N_16625);
xor U16911 (N_16911,N_16659,N_16450);
nor U16912 (N_16912,N_16760,N_16405);
or U16913 (N_16913,N_16526,N_16631);
and U16914 (N_16914,N_16557,N_16569);
nand U16915 (N_16915,N_16539,N_16724);
xor U16916 (N_16916,N_16478,N_16687);
and U16917 (N_16917,N_16577,N_16792);
nor U16918 (N_16918,N_16501,N_16718);
or U16919 (N_16919,N_16583,N_16689);
nand U16920 (N_16920,N_16685,N_16401);
nor U16921 (N_16921,N_16568,N_16436);
or U16922 (N_16922,N_16656,N_16796);
nor U16923 (N_16923,N_16678,N_16714);
or U16924 (N_16924,N_16743,N_16574);
or U16925 (N_16925,N_16644,N_16480);
or U16926 (N_16926,N_16717,N_16531);
nor U16927 (N_16927,N_16564,N_16552);
nand U16928 (N_16928,N_16410,N_16711);
and U16929 (N_16929,N_16667,N_16621);
xor U16930 (N_16930,N_16502,N_16764);
nor U16931 (N_16931,N_16692,N_16509);
nor U16932 (N_16932,N_16442,N_16591);
and U16933 (N_16933,N_16719,N_16522);
or U16934 (N_16934,N_16514,N_16471);
and U16935 (N_16935,N_16746,N_16532);
xor U16936 (N_16936,N_16546,N_16599);
and U16937 (N_16937,N_16555,N_16623);
nand U16938 (N_16938,N_16507,N_16476);
nand U16939 (N_16939,N_16705,N_16417);
or U16940 (N_16940,N_16787,N_16655);
nand U16941 (N_16941,N_16778,N_16731);
nor U16942 (N_16942,N_16528,N_16633);
and U16943 (N_16943,N_16781,N_16400);
xnor U16944 (N_16944,N_16756,N_16495);
nand U16945 (N_16945,N_16677,N_16643);
nand U16946 (N_16946,N_16525,N_16475);
xor U16947 (N_16947,N_16733,N_16543);
xnor U16948 (N_16948,N_16581,N_16700);
nand U16949 (N_16949,N_16793,N_16663);
nor U16950 (N_16950,N_16789,N_16572);
and U16951 (N_16951,N_16627,N_16762);
and U16952 (N_16952,N_16759,N_16788);
and U16953 (N_16953,N_16548,N_16535);
or U16954 (N_16954,N_16567,N_16757);
or U16955 (N_16955,N_16403,N_16594);
xnor U16956 (N_16956,N_16520,N_16723);
nand U16957 (N_16957,N_16477,N_16612);
and U16958 (N_16958,N_16587,N_16435);
and U16959 (N_16959,N_16459,N_16697);
nor U16960 (N_16960,N_16652,N_16713);
xnor U16961 (N_16961,N_16429,N_16691);
or U16962 (N_16962,N_16732,N_16774);
or U16963 (N_16963,N_16586,N_16721);
nor U16964 (N_16964,N_16431,N_16493);
nor U16965 (N_16965,N_16666,N_16416);
nor U16966 (N_16966,N_16511,N_16421);
or U16967 (N_16967,N_16558,N_16610);
nor U16968 (N_16968,N_16465,N_16665);
nor U16969 (N_16969,N_16603,N_16784);
xnor U16970 (N_16970,N_16479,N_16497);
or U16971 (N_16971,N_16409,N_16688);
nand U16972 (N_16972,N_16734,N_16412);
nand U16973 (N_16973,N_16712,N_16694);
and U16974 (N_16974,N_16524,N_16755);
xor U16975 (N_16975,N_16440,N_16637);
nor U16976 (N_16976,N_16596,N_16516);
nor U16977 (N_16977,N_16588,N_16629);
or U16978 (N_16978,N_16615,N_16725);
and U16979 (N_16979,N_16783,N_16560);
or U16980 (N_16980,N_16402,N_16702);
or U16981 (N_16981,N_16676,N_16618);
or U16982 (N_16982,N_16433,N_16439);
and U16983 (N_16983,N_16540,N_16404);
or U16984 (N_16984,N_16536,N_16418);
nand U16985 (N_16985,N_16640,N_16473);
xor U16986 (N_16986,N_16777,N_16780);
xor U16987 (N_16987,N_16720,N_16554);
and U16988 (N_16988,N_16452,N_16797);
and U16989 (N_16989,N_16773,N_16772);
xnor U16990 (N_16990,N_16770,N_16484);
nand U16991 (N_16991,N_16767,N_16695);
nand U16992 (N_16992,N_16751,N_16736);
and U16993 (N_16993,N_16559,N_16527);
and U16994 (N_16994,N_16604,N_16616);
nand U16995 (N_16995,N_16675,N_16608);
or U16996 (N_16996,N_16624,N_16779);
xnor U16997 (N_16997,N_16491,N_16744);
nand U16998 (N_16998,N_16727,N_16534);
or U16999 (N_16999,N_16490,N_16742);
and U17000 (N_17000,N_16626,N_16616);
or U17001 (N_17001,N_16716,N_16447);
nand U17002 (N_17002,N_16629,N_16633);
nand U17003 (N_17003,N_16778,N_16552);
nand U17004 (N_17004,N_16421,N_16656);
or U17005 (N_17005,N_16434,N_16555);
nor U17006 (N_17006,N_16640,N_16790);
and U17007 (N_17007,N_16526,N_16779);
or U17008 (N_17008,N_16602,N_16499);
and U17009 (N_17009,N_16643,N_16733);
nor U17010 (N_17010,N_16520,N_16421);
or U17011 (N_17011,N_16563,N_16470);
and U17012 (N_17012,N_16571,N_16786);
nor U17013 (N_17013,N_16615,N_16518);
xor U17014 (N_17014,N_16504,N_16785);
and U17015 (N_17015,N_16466,N_16554);
nor U17016 (N_17016,N_16735,N_16717);
or U17017 (N_17017,N_16514,N_16791);
xor U17018 (N_17018,N_16579,N_16601);
xnor U17019 (N_17019,N_16602,N_16790);
and U17020 (N_17020,N_16531,N_16688);
xor U17021 (N_17021,N_16775,N_16750);
xnor U17022 (N_17022,N_16723,N_16582);
xor U17023 (N_17023,N_16773,N_16747);
nand U17024 (N_17024,N_16573,N_16528);
nor U17025 (N_17025,N_16759,N_16557);
nor U17026 (N_17026,N_16772,N_16666);
nand U17027 (N_17027,N_16452,N_16691);
and U17028 (N_17028,N_16639,N_16666);
nor U17029 (N_17029,N_16799,N_16432);
or U17030 (N_17030,N_16578,N_16686);
nand U17031 (N_17031,N_16454,N_16777);
or U17032 (N_17032,N_16674,N_16717);
and U17033 (N_17033,N_16547,N_16585);
nand U17034 (N_17034,N_16789,N_16792);
nand U17035 (N_17035,N_16782,N_16408);
or U17036 (N_17036,N_16766,N_16773);
and U17037 (N_17037,N_16428,N_16417);
nand U17038 (N_17038,N_16649,N_16798);
nor U17039 (N_17039,N_16475,N_16483);
or U17040 (N_17040,N_16426,N_16792);
or U17041 (N_17041,N_16767,N_16639);
nor U17042 (N_17042,N_16543,N_16516);
nor U17043 (N_17043,N_16444,N_16716);
nand U17044 (N_17044,N_16436,N_16647);
and U17045 (N_17045,N_16468,N_16661);
nand U17046 (N_17046,N_16744,N_16457);
and U17047 (N_17047,N_16496,N_16500);
and U17048 (N_17048,N_16745,N_16501);
or U17049 (N_17049,N_16598,N_16621);
and U17050 (N_17050,N_16732,N_16713);
nand U17051 (N_17051,N_16445,N_16433);
or U17052 (N_17052,N_16798,N_16625);
and U17053 (N_17053,N_16629,N_16726);
and U17054 (N_17054,N_16784,N_16401);
nor U17055 (N_17055,N_16607,N_16420);
or U17056 (N_17056,N_16734,N_16744);
or U17057 (N_17057,N_16591,N_16452);
and U17058 (N_17058,N_16690,N_16595);
and U17059 (N_17059,N_16572,N_16593);
nor U17060 (N_17060,N_16499,N_16532);
nand U17061 (N_17061,N_16692,N_16624);
and U17062 (N_17062,N_16723,N_16611);
or U17063 (N_17063,N_16651,N_16598);
xor U17064 (N_17064,N_16637,N_16684);
and U17065 (N_17065,N_16762,N_16577);
xnor U17066 (N_17066,N_16761,N_16592);
xnor U17067 (N_17067,N_16511,N_16720);
or U17068 (N_17068,N_16510,N_16681);
nand U17069 (N_17069,N_16607,N_16721);
or U17070 (N_17070,N_16408,N_16582);
nor U17071 (N_17071,N_16515,N_16564);
xor U17072 (N_17072,N_16596,N_16439);
nor U17073 (N_17073,N_16476,N_16620);
xor U17074 (N_17074,N_16539,N_16625);
nand U17075 (N_17075,N_16521,N_16580);
or U17076 (N_17076,N_16528,N_16602);
or U17077 (N_17077,N_16436,N_16727);
nand U17078 (N_17078,N_16584,N_16548);
nand U17079 (N_17079,N_16565,N_16487);
nor U17080 (N_17080,N_16497,N_16448);
nand U17081 (N_17081,N_16721,N_16417);
xor U17082 (N_17082,N_16762,N_16726);
nor U17083 (N_17083,N_16474,N_16769);
nor U17084 (N_17084,N_16643,N_16623);
and U17085 (N_17085,N_16717,N_16412);
xnor U17086 (N_17086,N_16541,N_16759);
nand U17087 (N_17087,N_16517,N_16601);
nand U17088 (N_17088,N_16493,N_16677);
xor U17089 (N_17089,N_16775,N_16592);
nand U17090 (N_17090,N_16553,N_16799);
xor U17091 (N_17091,N_16505,N_16576);
xor U17092 (N_17092,N_16493,N_16475);
and U17093 (N_17093,N_16497,N_16556);
nand U17094 (N_17094,N_16682,N_16574);
and U17095 (N_17095,N_16604,N_16765);
or U17096 (N_17096,N_16763,N_16569);
nor U17097 (N_17097,N_16511,N_16564);
and U17098 (N_17098,N_16730,N_16751);
or U17099 (N_17099,N_16721,N_16479);
nand U17100 (N_17100,N_16580,N_16586);
and U17101 (N_17101,N_16532,N_16760);
nor U17102 (N_17102,N_16743,N_16762);
or U17103 (N_17103,N_16672,N_16758);
nor U17104 (N_17104,N_16734,N_16711);
nand U17105 (N_17105,N_16432,N_16468);
xor U17106 (N_17106,N_16697,N_16642);
nor U17107 (N_17107,N_16536,N_16689);
and U17108 (N_17108,N_16601,N_16770);
and U17109 (N_17109,N_16721,N_16551);
or U17110 (N_17110,N_16450,N_16616);
nor U17111 (N_17111,N_16602,N_16740);
or U17112 (N_17112,N_16403,N_16624);
nand U17113 (N_17113,N_16484,N_16578);
or U17114 (N_17114,N_16574,N_16649);
nand U17115 (N_17115,N_16664,N_16733);
xor U17116 (N_17116,N_16735,N_16670);
and U17117 (N_17117,N_16676,N_16653);
xor U17118 (N_17118,N_16544,N_16549);
and U17119 (N_17119,N_16441,N_16523);
and U17120 (N_17120,N_16744,N_16466);
and U17121 (N_17121,N_16727,N_16672);
xor U17122 (N_17122,N_16486,N_16716);
or U17123 (N_17123,N_16675,N_16767);
or U17124 (N_17124,N_16590,N_16408);
or U17125 (N_17125,N_16540,N_16532);
nand U17126 (N_17126,N_16406,N_16777);
nor U17127 (N_17127,N_16638,N_16481);
xnor U17128 (N_17128,N_16539,N_16580);
nor U17129 (N_17129,N_16786,N_16452);
xor U17130 (N_17130,N_16498,N_16701);
nor U17131 (N_17131,N_16686,N_16455);
nor U17132 (N_17132,N_16651,N_16415);
or U17133 (N_17133,N_16410,N_16567);
nand U17134 (N_17134,N_16618,N_16756);
xnor U17135 (N_17135,N_16799,N_16452);
nor U17136 (N_17136,N_16553,N_16592);
or U17137 (N_17137,N_16440,N_16790);
or U17138 (N_17138,N_16737,N_16530);
nor U17139 (N_17139,N_16443,N_16553);
xnor U17140 (N_17140,N_16477,N_16711);
xnor U17141 (N_17141,N_16720,N_16402);
or U17142 (N_17142,N_16758,N_16654);
xor U17143 (N_17143,N_16615,N_16498);
or U17144 (N_17144,N_16756,N_16414);
or U17145 (N_17145,N_16719,N_16548);
and U17146 (N_17146,N_16659,N_16658);
or U17147 (N_17147,N_16704,N_16792);
and U17148 (N_17148,N_16659,N_16581);
xnor U17149 (N_17149,N_16429,N_16713);
or U17150 (N_17150,N_16672,N_16748);
nor U17151 (N_17151,N_16403,N_16514);
nand U17152 (N_17152,N_16583,N_16408);
or U17153 (N_17153,N_16406,N_16594);
or U17154 (N_17154,N_16506,N_16620);
and U17155 (N_17155,N_16518,N_16729);
and U17156 (N_17156,N_16711,N_16620);
or U17157 (N_17157,N_16558,N_16448);
and U17158 (N_17158,N_16775,N_16473);
nor U17159 (N_17159,N_16759,N_16605);
nor U17160 (N_17160,N_16797,N_16429);
xor U17161 (N_17161,N_16501,N_16509);
or U17162 (N_17162,N_16457,N_16472);
or U17163 (N_17163,N_16584,N_16649);
and U17164 (N_17164,N_16652,N_16710);
and U17165 (N_17165,N_16620,N_16517);
xnor U17166 (N_17166,N_16792,N_16668);
xnor U17167 (N_17167,N_16565,N_16469);
and U17168 (N_17168,N_16791,N_16589);
or U17169 (N_17169,N_16658,N_16587);
and U17170 (N_17170,N_16652,N_16442);
nor U17171 (N_17171,N_16443,N_16771);
or U17172 (N_17172,N_16661,N_16710);
and U17173 (N_17173,N_16636,N_16589);
xnor U17174 (N_17174,N_16653,N_16679);
and U17175 (N_17175,N_16615,N_16588);
nor U17176 (N_17176,N_16790,N_16506);
nand U17177 (N_17177,N_16689,N_16425);
and U17178 (N_17178,N_16708,N_16563);
and U17179 (N_17179,N_16642,N_16451);
or U17180 (N_17180,N_16481,N_16413);
xor U17181 (N_17181,N_16775,N_16495);
nor U17182 (N_17182,N_16607,N_16634);
or U17183 (N_17183,N_16710,N_16594);
xor U17184 (N_17184,N_16657,N_16501);
and U17185 (N_17185,N_16550,N_16591);
xor U17186 (N_17186,N_16502,N_16592);
nand U17187 (N_17187,N_16507,N_16705);
nor U17188 (N_17188,N_16758,N_16757);
and U17189 (N_17189,N_16403,N_16779);
and U17190 (N_17190,N_16402,N_16560);
nor U17191 (N_17191,N_16753,N_16519);
nand U17192 (N_17192,N_16795,N_16677);
nor U17193 (N_17193,N_16460,N_16563);
nor U17194 (N_17194,N_16557,N_16697);
nor U17195 (N_17195,N_16421,N_16694);
xnor U17196 (N_17196,N_16598,N_16669);
and U17197 (N_17197,N_16577,N_16760);
nor U17198 (N_17198,N_16402,N_16794);
xnor U17199 (N_17199,N_16759,N_16432);
nor U17200 (N_17200,N_17172,N_17100);
xor U17201 (N_17201,N_17083,N_17106);
nand U17202 (N_17202,N_17065,N_17051);
or U17203 (N_17203,N_17017,N_17014);
and U17204 (N_17204,N_16960,N_16941);
nand U17205 (N_17205,N_16936,N_16982);
xnor U17206 (N_17206,N_16828,N_16923);
and U17207 (N_17207,N_17026,N_16933);
nor U17208 (N_17208,N_16878,N_17029);
and U17209 (N_17209,N_17179,N_16928);
nor U17210 (N_17210,N_16940,N_16932);
and U17211 (N_17211,N_17150,N_16974);
nand U17212 (N_17212,N_17174,N_16883);
xor U17213 (N_17213,N_16935,N_16890);
xor U17214 (N_17214,N_17192,N_17187);
nand U17215 (N_17215,N_17069,N_16863);
and U17216 (N_17216,N_16814,N_17163);
and U17217 (N_17217,N_16919,N_17068);
and U17218 (N_17218,N_16918,N_17115);
nand U17219 (N_17219,N_17198,N_16897);
and U17220 (N_17220,N_17104,N_17166);
nor U17221 (N_17221,N_16976,N_17058);
nor U17222 (N_17222,N_17008,N_17040);
nand U17223 (N_17223,N_16999,N_16859);
nor U17224 (N_17224,N_16856,N_16849);
and U17225 (N_17225,N_16830,N_17047);
nor U17226 (N_17226,N_16874,N_17018);
and U17227 (N_17227,N_16857,N_17062);
and U17228 (N_17228,N_17139,N_17171);
and U17229 (N_17229,N_16892,N_17054);
xor U17230 (N_17230,N_16804,N_16971);
nor U17231 (N_17231,N_17036,N_17035);
or U17232 (N_17232,N_17034,N_17123);
and U17233 (N_17233,N_17095,N_16959);
and U17234 (N_17234,N_16805,N_17120);
nor U17235 (N_17235,N_17070,N_16884);
xnor U17236 (N_17236,N_17101,N_16870);
xnor U17237 (N_17237,N_17019,N_17170);
nor U17238 (N_17238,N_16901,N_16984);
and U17239 (N_17239,N_17025,N_16835);
xor U17240 (N_17240,N_16893,N_17168);
xor U17241 (N_17241,N_17154,N_17005);
xnor U17242 (N_17242,N_16930,N_17199);
or U17243 (N_17243,N_16986,N_17081);
xnor U17244 (N_17244,N_16860,N_17001);
nand U17245 (N_17245,N_17114,N_16946);
nor U17246 (N_17246,N_16827,N_17184);
nand U17247 (N_17247,N_17108,N_17066);
or U17248 (N_17248,N_16871,N_16836);
nor U17249 (N_17249,N_16925,N_17117);
or U17250 (N_17250,N_16990,N_17151);
and U17251 (N_17251,N_17041,N_17128);
xnor U17252 (N_17252,N_16907,N_16978);
or U17253 (N_17253,N_16981,N_17090);
and U17254 (N_17254,N_16848,N_17191);
nor U17255 (N_17255,N_16894,N_16800);
xnor U17256 (N_17256,N_17122,N_16916);
xor U17257 (N_17257,N_17024,N_16954);
or U17258 (N_17258,N_17189,N_16912);
nor U17259 (N_17259,N_16845,N_16812);
and U17260 (N_17260,N_16921,N_17010);
and U17261 (N_17261,N_16866,N_17099);
or U17262 (N_17262,N_16972,N_16858);
xor U17263 (N_17263,N_17022,N_16815);
nand U17264 (N_17264,N_17177,N_16802);
nand U17265 (N_17265,N_16917,N_17109);
or U17266 (N_17266,N_17105,N_16962);
or U17267 (N_17267,N_16904,N_17000);
or U17268 (N_17268,N_16869,N_16979);
nand U17269 (N_17269,N_17007,N_17031);
or U17270 (N_17270,N_16996,N_17178);
nor U17271 (N_17271,N_17021,N_17063);
nand U17272 (N_17272,N_17015,N_17078);
and U17273 (N_17273,N_16843,N_16810);
nand U17274 (N_17274,N_17003,N_17030);
and U17275 (N_17275,N_16942,N_16876);
and U17276 (N_17276,N_17190,N_17145);
nand U17277 (N_17277,N_16943,N_16807);
and U17278 (N_17278,N_16998,N_17148);
and U17279 (N_17279,N_16834,N_16953);
xor U17280 (N_17280,N_16862,N_16886);
and U17281 (N_17281,N_17084,N_17142);
nand U17282 (N_17282,N_17131,N_17134);
nor U17283 (N_17283,N_16947,N_16840);
nor U17284 (N_17284,N_16839,N_16889);
nand U17285 (N_17285,N_17049,N_16842);
and U17286 (N_17286,N_16929,N_17195);
and U17287 (N_17287,N_16826,N_17155);
and U17288 (N_17288,N_16949,N_17044);
and U17289 (N_17289,N_17085,N_16872);
or U17290 (N_17290,N_17033,N_16838);
xnor U17291 (N_17291,N_16868,N_16822);
and U17292 (N_17292,N_16934,N_16969);
nand U17293 (N_17293,N_16994,N_16948);
xnor U17294 (N_17294,N_16823,N_17112);
and U17295 (N_17295,N_16813,N_17077);
xnor U17296 (N_17296,N_17159,N_17130);
or U17297 (N_17297,N_17175,N_16809);
and U17298 (N_17298,N_17169,N_17056);
nand U17299 (N_17299,N_16875,N_17053);
xor U17300 (N_17300,N_17004,N_16989);
and U17301 (N_17301,N_17097,N_17197);
and U17302 (N_17302,N_16854,N_17127);
xor U17303 (N_17303,N_16899,N_17135);
nor U17304 (N_17304,N_17129,N_17074);
xnor U17305 (N_17305,N_16885,N_17091);
or U17306 (N_17306,N_17032,N_17048);
and U17307 (N_17307,N_16903,N_17028);
and U17308 (N_17308,N_16977,N_16995);
or U17309 (N_17309,N_17143,N_17089);
nor U17310 (N_17310,N_17167,N_17088);
xnor U17311 (N_17311,N_17102,N_17020);
and U17312 (N_17312,N_16816,N_16980);
or U17313 (N_17313,N_16865,N_17045);
nor U17314 (N_17314,N_17093,N_16945);
nand U17315 (N_17315,N_17042,N_17194);
nor U17316 (N_17316,N_16993,N_16846);
or U17317 (N_17317,N_17061,N_16864);
or U17318 (N_17318,N_16831,N_16881);
and U17319 (N_17319,N_17055,N_16801);
and U17320 (N_17320,N_16950,N_16965);
and U17321 (N_17321,N_16915,N_17125);
or U17322 (N_17322,N_16902,N_16852);
xnor U17323 (N_17323,N_17147,N_16825);
nor U17324 (N_17324,N_16829,N_17118);
or U17325 (N_17325,N_17176,N_17016);
nor U17326 (N_17326,N_17116,N_17080);
and U17327 (N_17327,N_16821,N_17113);
xor U17328 (N_17328,N_17165,N_17076);
and U17329 (N_17329,N_17013,N_16888);
and U17330 (N_17330,N_16853,N_17027);
xor U17331 (N_17331,N_16898,N_16819);
and U17332 (N_17332,N_16939,N_17071);
xor U17333 (N_17333,N_17059,N_17132);
and U17334 (N_17334,N_17133,N_16975);
and U17335 (N_17335,N_17094,N_17011);
nand U17336 (N_17336,N_17064,N_16970);
nor U17337 (N_17337,N_17023,N_16924);
and U17338 (N_17338,N_17107,N_16910);
xnor U17339 (N_17339,N_16958,N_16882);
xnor U17340 (N_17340,N_16817,N_17124);
xnor U17341 (N_17341,N_17039,N_16992);
xor U17342 (N_17342,N_17138,N_16879);
nand U17343 (N_17343,N_16914,N_16938);
nand U17344 (N_17344,N_17149,N_16867);
nand U17345 (N_17345,N_16944,N_17043);
nor U17346 (N_17346,N_17086,N_16967);
or U17347 (N_17347,N_17183,N_17067);
nand U17348 (N_17348,N_17046,N_16832);
nand U17349 (N_17349,N_17153,N_16905);
nand U17350 (N_17350,N_17156,N_16926);
xnor U17351 (N_17351,N_16880,N_17119);
or U17352 (N_17352,N_16955,N_17103);
and U17353 (N_17353,N_16991,N_17141);
or U17354 (N_17354,N_17087,N_16811);
and U17355 (N_17355,N_16891,N_17126);
xor U17356 (N_17356,N_17073,N_17188);
nor U17357 (N_17357,N_16952,N_16803);
or U17358 (N_17358,N_16906,N_17181);
xnor U17359 (N_17359,N_16837,N_17152);
nor U17360 (N_17360,N_17137,N_16961);
nand U17361 (N_17361,N_17164,N_16861);
and U17362 (N_17362,N_17161,N_16847);
nor U17363 (N_17363,N_16851,N_17038);
xnor U17364 (N_17364,N_16951,N_17037);
nor U17365 (N_17365,N_17111,N_16896);
nor U17366 (N_17366,N_16895,N_17157);
or U17367 (N_17367,N_16983,N_16833);
and U17368 (N_17368,N_16808,N_17185);
or U17369 (N_17369,N_17182,N_16824);
and U17370 (N_17370,N_17075,N_17092);
or U17371 (N_17371,N_16927,N_16922);
xnor U17372 (N_17372,N_17012,N_17144);
nor U17373 (N_17373,N_16900,N_16887);
and U17374 (N_17374,N_16937,N_16841);
xor U17375 (N_17375,N_17096,N_17009);
xor U17376 (N_17376,N_16985,N_16931);
and U17377 (N_17377,N_16913,N_16988);
or U17378 (N_17378,N_16911,N_17136);
and U17379 (N_17379,N_17006,N_16966);
nand U17380 (N_17380,N_17173,N_17186);
and U17381 (N_17381,N_17121,N_17079);
or U17382 (N_17382,N_16818,N_17082);
xor U17383 (N_17383,N_16908,N_17193);
nand U17384 (N_17384,N_16850,N_17146);
and U17385 (N_17385,N_16973,N_17050);
and U17386 (N_17386,N_17160,N_16968);
or U17387 (N_17387,N_17002,N_17098);
and U17388 (N_17388,N_17180,N_16963);
and U17389 (N_17389,N_16909,N_16844);
nor U17390 (N_17390,N_16956,N_17052);
nand U17391 (N_17391,N_17196,N_17057);
nor U17392 (N_17392,N_16855,N_16877);
nand U17393 (N_17393,N_16806,N_17140);
or U17394 (N_17394,N_17060,N_16957);
nor U17395 (N_17395,N_17158,N_16873);
xor U17396 (N_17396,N_16820,N_16920);
or U17397 (N_17397,N_17110,N_17072);
or U17398 (N_17398,N_17162,N_16997);
nand U17399 (N_17399,N_16964,N_16987);
and U17400 (N_17400,N_17154,N_17101);
xnor U17401 (N_17401,N_16972,N_17103);
or U17402 (N_17402,N_16968,N_16921);
nor U17403 (N_17403,N_16968,N_16935);
and U17404 (N_17404,N_17033,N_16960);
xnor U17405 (N_17405,N_16889,N_16924);
and U17406 (N_17406,N_17174,N_17081);
nand U17407 (N_17407,N_17057,N_16897);
nor U17408 (N_17408,N_17198,N_16986);
nand U17409 (N_17409,N_16914,N_16811);
or U17410 (N_17410,N_17058,N_16820);
and U17411 (N_17411,N_16973,N_16998);
and U17412 (N_17412,N_17140,N_17181);
nor U17413 (N_17413,N_16946,N_17067);
nand U17414 (N_17414,N_16935,N_17049);
xor U17415 (N_17415,N_16993,N_17155);
xnor U17416 (N_17416,N_17060,N_17015);
and U17417 (N_17417,N_16874,N_17182);
or U17418 (N_17418,N_16958,N_16947);
xor U17419 (N_17419,N_16964,N_17002);
nor U17420 (N_17420,N_17094,N_16842);
nor U17421 (N_17421,N_17091,N_17183);
nand U17422 (N_17422,N_17006,N_16869);
nor U17423 (N_17423,N_17162,N_16897);
nand U17424 (N_17424,N_17113,N_16808);
xor U17425 (N_17425,N_16982,N_16958);
or U17426 (N_17426,N_16892,N_17107);
nor U17427 (N_17427,N_16986,N_16911);
xnor U17428 (N_17428,N_16967,N_17031);
xor U17429 (N_17429,N_17064,N_17159);
and U17430 (N_17430,N_17069,N_16837);
xor U17431 (N_17431,N_16942,N_16964);
and U17432 (N_17432,N_16873,N_16972);
xnor U17433 (N_17433,N_16873,N_17010);
and U17434 (N_17434,N_16814,N_17183);
nand U17435 (N_17435,N_17185,N_17144);
nand U17436 (N_17436,N_16929,N_16827);
nor U17437 (N_17437,N_16960,N_17184);
xor U17438 (N_17438,N_16847,N_16998);
nor U17439 (N_17439,N_17131,N_16853);
nor U17440 (N_17440,N_16950,N_16809);
or U17441 (N_17441,N_17112,N_17199);
and U17442 (N_17442,N_16890,N_16929);
nand U17443 (N_17443,N_17064,N_17146);
xnor U17444 (N_17444,N_16881,N_16933);
xnor U17445 (N_17445,N_17065,N_17148);
nand U17446 (N_17446,N_16805,N_16989);
or U17447 (N_17447,N_17008,N_16840);
xnor U17448 (N_17448,N_16828,N_17189);
xor U17449 (N_17449,N_16848,N_16880);
nor U17450 (N_17450,N_16806,N_16992);
and U17451 (N_17451,N_16973,N_16946);
nor U17452 (N_17452,N_16833,N_17072);
or U17453 (N_17453,N_16980,N_16860);
nor U17454 (N_17454,N_17165,N_17178);
nand U17455 (N_17455,N_17142,N_16830);
and U17456 (N_17456,N_17112,N_16836);
or U17457 (N_17457,N_17002,N_16995);
nor U17458 (N_17458,N_16959,N_17158);
xnor U17459 (N_17459,N_16849,N_16845);
and U17460 (N_17460,N_17100,N_16863);
nand U17461 (N_17461,N_17173,N_16975);
and U17462 (N_17462,N_16845,N_17193);
nand U17463 (N_17463,N_16818,N_17108);
xor U17464 (N_17464,N_16834,N_17058);
nor U17465 (N_17465,N_17153,N_16956);
or U17466 (N_17466,N_16808,N_17081);
nor U17467 (N_17467,N_16977,N_17117);
xnor U17468 (N_17468,N_17154,N_17036);
nor U17469 (N_17469,N_17128,N_17000);
nor U17470 (N_17470,N_17155,N_17050);
or U17471 (N_17471,N_17118,N_16986);
nand U17472 (N_17472,N_17149,N_16941);
or U17473 (N_17473,N_16983,N_16976);
nand U17474 (N_17474,N_16825,N_16873);
nand U17475 (N_17475,N_16830,N_16831);
nand U17476 (N_17476,N_17138,N_17133);
or U17477 (N_17477,N_17014,N_17042);
nand U17478 (N_17478,N_17180,N_17184);
nor U17479 (N_17479,N_16901,N_16914);
and U17480 (N_17480,N_17163,N_16903);
or U17481 (N_17481,N_16808,N_16935);
and U17482 (N_17482,N_17028,N_16929);
xor U17483 (N_17483,N_16870,N_17070);
nor U17484 (N_17484,N_17073,N_17147);
nand U17485 (N_17485,N_17080,N_16992);
xnor U17486 (N_17486,N_17029,N_17054);
xnor U17487 (N_17487,N_17032,N_16965);
nor U17488 (N_17488,N_16982,N_16946);
nor U17489 (N_17489,N_17021,N_17139);
and U17490 (N_17490,N_16836,N_16969);
nor U17491 (N_17491,N_17197,N_17067);
and U17492 (N_17492,N_17017,N_17188);
or U17493 (N_17493,N_16935,N_16916);
or U17494 (N_17494,N_17153,N_16883);
and U17495 (N_17495,N_17183,N_17106);
xor U17496 (N_17496,N_17166,N_16942);
or U17497 (N_17497,N_16996,N_17104);
nand U17498 (N_17498,N_17174,N_17069);
and U17499 (N_17499,N_17175,N_17195);
xor U17500 (N_17500,N_16946,N_17047);
and U17501 (N_17501,N_16979,N_16943);
xor U17502 (N_17502,N_17199,N_17127);
xor U17503 (N_17503,N_17036,N_16871);
nor U17504 (N_17504,N_17050,N_16958);
nand U17505 (N_17505,N_17086,N_16831);
and U17506 (N_17506,N_16947,N_16965);
or U17507 (N_17507,N_17070,N_17106);
xor U17508 (N_17508,N_16837,N_16939);
xor U17509 (N_17509,N_16969,N_17068);
nand U17510 (N_17510,N_16870,N_16898);
nor U17511 (N_17511,N_16904,N_17189);
or U17512 (N_17512,N_16889,N_16874);
nor U17513 (N_17513,N_16970,N_16937);
nor U17514 (N_17514,N_17047,N_16988);
nand U17515 (N_17515,N_16942,N_17138);
and U17516 (N_17516,N_16913,N_16892);
xnor U17517 (N_17517,N_16894,N_16906);
or U17518 (N_17518,N_17040,N_17063);
xnor U17519 (N_17519,N_16870,N_16955);
nor U17520 (N_17520,N_17124,N_17086);
xnor U17521 (N_17521,N_16881,N_16909);
xor U17522 (N_17522,N_17193,N_17149);
nor U17523 (N_17523,N_17198,N_17161);
and U17524 (N_17524,N_17113,N_16835);
xor U17525 (N_17525,N_17050,N_16933);
xnor U17526 (N_17526,N_16801,N_16833);
or U17527 (N_17527,N_17104,N_17025);
nor U17528 (N_17528,N_17086,N_17020);
xnor U17529 (N_17529,N_16920,N_17111);
xnor U17530 (N_17530,N_17107,N_17002);
or U17531 (N_17531,N_16991,N_16844);
or U17532 (N_17532,N_16892,N_16919);
or U17533 (N_17533,N_16975,N_16808);
nand U17534 (N_17534,N_16844,N_16885);
nand U17535 (N_17535,N_16891,N_16855);
xor U17536 (N_17536,N_17145,N_17002);
nand U17537 (N_17537,N_17101,N_17150);
and U17538 (N_17538,N_16859,N_16927);
or U17539 (N_17539,N_16897,N_17074);
nor U17540 (N_17540,N_17109,N_17128);
nand U17541 (N_17541,N_17193,N_16999);
nor U17542 (N_17542,N_17140,N_17166);
nor U17543 (N_17543,N_16848,N_17118);
xnor U17544 (N_17544,N_17056,N_16918);
xor U17545 (N_17545,N_17128,N_17186);
nor U17546 (N_17546,N_16886,N_16855);
xor U17547 (N_17547,N_17120,N_17179);
and U17548 (N_17548,N_17181,N_16862);
xor U17549 (N_17549,N_16861,N_16814);
xnor U17550 (N_17550,N_16983,N_17155);
nor U17551 (N_17551,N_16934,N_16939);
nand U17552 (N_17552,N_16987,N_17003);
or U17553 (N_17553,N_17033,N_16934);
xnor U17554 (N_17554,N_17097,N_16908);
xor U17555 (N_17555,N_16884,N_17033);
and U17556 (N_17556,N_17049,N_17005);
nor U17557 (N_17557,N_17187,N_17179);
nor U17558 (N_17558,N_17044,N_17190);
xor U17559 (N_17559,N_17064,N_16847);
xnor U17560 (N_17560,N_17009,N_17133);
nor U17561 (N_17561,N_16862,N_16914);
or U17562 (N_17562,N_16800,N_16992);
xnor U17563 (N_17563,N_17060,N_16881);
xor U17564 (N_17564,N_17178,N_17153);
xor U17565 (N_17565,N_17116,N_17177);
xor U17566 (N_17566,N_17023,N_16906);
or U17567 (N_17567,N_16976,N_17141);
nor U17568 (N_17568,N_16930,N_16989);
nor U17569 (N_17569,N_17062,N_16811);
xor U17570 (N_17570,N_17182,N_17056);
xor U17571 (N_17571,N_16887,N_16822);
nor U17572 (N_17572,N_16971,N_17040);
or U17573 (N_17573,N_16843,N_17194);
or U17574 (N_17574,N_17093,N_16862);
and U17575 (N_17575,N_16979,N_16930);
xor U17576 (N_17576,N_17001,N_16931);
xnor U17577 (N_17577,N_17104,N_17004);
and U17578 (N_17578,N_16858,N_17051);
or U17579 (N_17579,N_17076,N_16802);
or U17580 (N_17580,N_16997,N_17024);
nor U17581 (N_17581,N_17090,N_17193);
and U17582 (N_17582,N_16893,N_16837);
nand U17583 (N_17583,N_17025,N_16902);
and U17584 (N_17584,N_16920,N_17113);
or U17585 (N_17585,N_16812,N_16974);
nand U17586 (N_17586,N_17134,N_16943);
xnor U17587 (N_17587,N_16862,N_16929);
xor U17588 (N_17588,N_17145,N_17054);
nor U17589 (N_17589,N_16829,N_17149);
nand U17590 (N_17590,N_16860,N_17127);
and U17591 (N_17591,N_16802,N_17164);
or U17592 (N_17592,N_16816,N_17114);
xor U17593 (N_17593,N_17039,N_16926);
xnor U17594 (N_17594,N_16921,N_17134);
nand U17595 (N_17595,N_16841,N_17181);
and U17596 (N_17596,N_16855,N_16984);
and U17597 (N_17597,N_17155,N_17076);
nand U17598 (N_17598,N_16979,N_17046);
or U17599 (N_17599,N_17028,N_17196);
nand U17600 (N_17600,N_17311,N_17280);
or U17601 (N_17601,N_17443,N_17463);
nor U17602 (N_17602,N_17351,N_17365);
nand U17603 (N_17603,N_17230,N_17349);
or U17604 (N_17604,N_17386,N_17557);
or U17605 (N_17605,N_17314,N_17266);
xnor U17606 (N_17606,N_17539,N_17300);
nor U17607 (N_17607,N_17387,N_17451);
or U17608 (N_17608,N_17220,N_17570);
nor U17609 (N_17609,N_17565,N_17242);
nor U17610 (N_17610,N_17375,N_17363);
nand U17611 (N_17611,N_17518,N_17355);
nand U17612 (N_17612,N_17503,N_17405);
nand U17613 (N_17613,N_17307,N_17323);
and U17614 (N_17614,N_17338,N_17221);
and U17615 (N_17615,N_17337,N_17301);
nand U17616 (N_17616,N_17473,N_17373);
or U17617 (N_17617,N_17331,N_17596);
nor U17618 (N_17618,N_17594,N_17422);
nand U17619 (N_17619,N_17385,N_17219);
xnor U17620 (N_17620,N_17392,N_17203);
nand U17621 (N_17621,N_17345,N_17315);
or U17622 (N_17622,N_17213,N_17420);
and U17623 (N_17623,N_17553,N_17474);
xnor U17624 (N_17624,N_17329,N_17429);
or U17625 (N_17625,N_17306,N_17528);
and U17626 (N_17626,N_17568,N_17454);
or U17627 (N_17627,N_17292,N_17340);
nand U17628 (N_17628,N_17441,N_17299);
and U17629 (N_17629,N_17237,N_17509);
xor U17630 (N_17630,N_17212,N_17467);
and U17631 (N_17631,N_17464,N_17452);
nand U17632 (N_17632,N_17332,N_17293);
and U17633 (N_17633,N_17354,N_17379);
and U17634 (N_17634,N_17364,N_17590);
nand U17635 (N_17635,N_17303,N_17589);
and U17636 (N_17636,N_17318,N_17324);
or U17637 (N_17637,N_17457,N_17361);
and U17638 (N_17638,N_17481,N_17426);
nor U17639 (N_17639,N_17341,N_17333);
xnor U17640 (N_17640,N_17583,N_17538);
xnor U17641 (N_17641,N_17547,N_17261);
nor U17642 (N_17642,N_17475,N_17384);
nand U17643 (N_17643,N_17563,N_17211);
or U17644 (N_17644,N_17419,N_17357);
or U17645 (N_17645,N_17433,N_17552);
xor U17646 (N_17646,N_17448,N_17418);
and U17647 (N_17647,N_17291,N_17245);
nor U17648 (N_17648,N_17572,N_17410);
nand U17649 (N_17649,N_17421,N_17284);
and U17650 (N_17650,N_17223,N_17297);
xor U17651 (N_17651,N_17328,N_17541);
nand U17652 (N_17652,N_17330,N_17296);
or U17653 (N_17653,N_17466,N_17522);
and U17654 (N_17654,N_17368,N_17478);
or U17655 (N_17655,N_17346,N_17581);
nor U17656 (N_17656,N_17586,N_17304);
or U17657 (N_17657,N_17305,N_17445);
and U17658 (N_17658,N_17582,N_17550);
nor U17659 (N_17659,N_17523,N_17277);
nand U17660 (N_17660,N_17512,N_17453);
nand U17661 (N_17661,N_17575,N_17286);
nand U17662 (N_17662,N_17372,N_17390);
nand U17663 (N_17663,N_17336,N_17484);
or U17664 (N_17664,N_17444,N_17207);
nor U17665 (N_17665,N_17486,N_17377);
and U17666 (N_17666,N_17252,N_17487);
and U17667 (N_17667,N_17413,N_17432);
nor U17668 (N_17668,N_17241,N_17571);
nand U17669 (N_17669,N_17489,N_17485);
nand U17670 (N_17670,N_17551,N_17248);
nand U17671 (N_17671,N_17506,N_17455);
nor U17672 (N_17672,N_17504,N_17289);
nor U17673 (N_17673,N_17356,N_17555);
nor U17674 (N_17674,N_17529,N_17263);
xor U17675 (N_17675,N_17210,N_17224);
xnor U17676 (N_17676,N_17281,N_17469);
and U17677 (N_17677,N_17206,N_17273);
nand U17678 (N_17678,N_17200,N_17470);
nor U17679 (N_17679,N_17597,N_17450);
and U17680 (N_17680,N_17348,N_17309);
and U17681 (N_17681,N_17326,N_17217);
nand U17682 (N_17682,N_17515,N_17576);
xnor U17683 (N_17683,N_17317,N_17558);
nor U17684 (N_17684,N_17517,N_17440);
and U17685 (N_17685,N_17371,N_17415);
or U17686 (N_17686,N_17577,N_17430);
and U17687 (N_17687,N_17446,N_17257);
xnor U17688 (N_17688,N_17508,N_17388);
and U17689 (N_17689,N_17228,N_17358);
nand U17690 (N_17690,N_17393,N_17262);
xnor U17691 (N_17691,N_17229,N_17254);
and U17692 (N_17692,N_17549,N_17412);
nor U17693 (N_17693,N_17434,N_17431);
nor U17694 (N_17694,N_17414,N_17408);
nor U17695 (N_17695,N_17535,N_17216);
nand U17696 (N_17696,N_17239,N_17598);
nand U17697 (N_17697,N_17599,N_17510);
nor U17698 (N_17698,N_17437,N_17505);
nor U17699 (N_17699,N_17573,N_17246);
nand U17700 (N_17700,N_17240,N_17471);
and U17701 (N_17701,N_17580,N_17268);
or U17702 (N_17702,N_17425,N_17302);
nand U17703 (N_17703,N_17271,N_17497);
xor U17704 (N_17704,N_17278,N_17516);
and U17705 (N_17705,N_17399,N_17397);
nor U17706 (N_17706,N_17209,N_17592);
xor U17707 (N_17707,N_17423,N_17335);
and U17708 (N_17708,N_17359,N_17526);
or U17709 (N_17709,N_17436,N_17205);
nand U17710 (N_17710,N_17283,N_17537);
or U17711 (N_17711,N_17476,N_17267);
xnor U17712 (N_17712,N_17574,N_17591);
or U17713 (N_17713,N_17428,N_17204);
nor U17714 (N_17714,N_17310,N_17491);
xnor U17715 (N_17715,N_17493,N_17394);
nand U17716 (N_17716,N_17514,N_17380);
or U17717 (N_17717,N_17334,N_17322);
and U17718 (N_17718,N_17227,N_17498);
and U17719 (N_17719,N_17294,N_17513);
and U17720 (N_17720,N_17339,N_17370);
nand U17721 (N_17721,N_17403,N_17232);
or U17722 (N_17722,N_17265,N_17215);
or U17723 (N_17723,N_17459,N_17439);
and U17724 (N_17724,N_17319,N_17507);
and U17725 (N_17725,N_17567,N_17308);
nor U17726 (N_17726,N_17561,N_17381);
xor U17727 (N_17727,N_17218,N_17544);
and U17728 (N_17728,N_17417,N_17238);
and U17729 (N_17729,N_17427,N_17519);
nand U17730 (N_17730,N_17347,N_17531);
or U17731 (N_17731,N_17276,N_17396);
nor U17732 (N_17732,N_17411,N_17226);
nand U17733 (N_17733,N_17530,N_17543);
nand U17734 (N_17734,N_17559,N_17480);
or U17735 (N_17735,N_17548,N_17374);
nand U17736 (N_17736,N_17442,N_17472);
and U17737 (N_17737,N_17536,N_17401);
xor U17738 (N_17738,N_17595,N_17542);
xnor U17739 (N_17739,N_17479,N_17342);
nor U17740 (N_17740,N_17495,N_17593);
nor U17741 (N_17741,N_17462,N_17406);
nand U17742 (N_17742,N_17316,N_17260);
xnor U17743 (N_17743,N_17579,N_17527);
and U17744 (N_17744,N_17369,N_17201);
nand U17745 (N_17745,N_17521,N_17400);
nor U17746 (N_17746,N_17447,N_17222);
xor U17747 (N_17747,N_17424,N_17458);
or U17748 (N_17748,N_17494,N_17244);
nand U17749 (N_17749,N_17264,N_17416);
nor U17750 (N_17750,N_17554,N_17350);
nor U17751 (N_17751,N_17465,N_17540);
and U17752 (N_17752,N_17325,N_17320);
nand U17753 (N_17753,N_17279,N_17435);
nor U17754 (N_17754,N_17389,N_17569);
and U17755 (N_17755,N_17295,N_17362);
or U17756 (N_17756,N_17492,N_17270);
and U17757 (N_17757,N_17499,N_17312);
nand U17758 (N_17758,N_17327,N_17460);
xor U17759 (N_17759,N_17376,N_17438);
xnor U17760 (N_17760,N_17225,N_17556);
or U17761 (N_17761,N_17449,N_17236);
nor U17762 (N_17762,N_17407,N_17382);
nand U17763 (N_17763,N_17398,N_17461);
or U17764 (N_17764,N_17546,N_17456);
or U17765 (N_17765,N_17287,N_17500);
nand U17766 (N_17766,N_17247,N_17490);
and U17767 (N_17767,N_17468,N_17532);
or U17768 (N_17768,N_17395,N_17496);
or U17769 (N_17769,N_17243,N_17313);
xor U17770 (N_17770,N_17391,N_17255);
or U17771 (N_17771,N_17564,N_17383);
and U17772 (N_17772,N_17202,N_17343);
or U17773 (N_17773,N_17366,N_17249);
xnor U17774 (N_17774,N_17562,N_17208);
nor U17775 (N_17775,N_17214,N_17234);
xor U17776 (N_17776,N_17483,N_17524);
nor U17777 (N_17777,N_17501,N_17298);
xor U17778 (N_17778,N_17290,N_17344);
and U17779 (N_17779,N_17352,N_17288);
xor U17780 (N_17780,N_17259,N_17235);
and U17781 (N_17781,N_17285,N_17282);
nor U17782 (N_17782,N_17231,N_17404);
nand U17783 (N_17783,N_17378,N_17533);
nand U17784 (N_17784,N_17321,N_17367);
or U17785 (N_17785,N_17587,N_17253);
nand U17786 (N_17786,N_17584,N_17353);
xnor U17787 (N_17787,N_17566,N_17251);
or U17788 (N_17788,N_17258,N_17409);
xnor U17789 (N_17789,N_17560,N_17585);
and U17790 (N_17790,N_17250,N_17511);
nand U17791 (N_17791,N_17272,N_17578);
nor U17792 (N_17792,N_17545,N_17360);
nand U17793 (N_17793,N_17488,N_17275);
and U17794 (N_17794,N_17477,N_17502);
or U17795 (N_17795,N_17269,N_17534);
xor U17796 (N_17796,N_17588,N_17402);
and U17797 (N_17797,N_17525,N_17520);
xnor U17798 (N_17798,N_17233,N_17256);
nor U17799 (N_17799,N_17274,N_17482);
nor U17800 (N_17800,N_17352,N_17354);
or U17801 (N_17801,N_17533,N_17231);
nor U17802 (N_17802,N_17237,N_17406);
xnor U17803 (N_17803,N_17369,N_17456);
xnor U17804 (N_17804,N_17469,N_17275);
and U17805 (N_17805,N_17436,N_17306);
xnor U17806 (N_17806,N_17581,N_17332);
and U17807 (N_17807,N_17281,N_17313);
xnor U17808 (N_17808,N_17312,N_17303);
or U17809 (N_17809,N_17377,N_17570);
nor U17810 (N_17810,N_17207,N_17263);
and U17811 (N_17811,N_17248,N_17400);
nand U17812 (N_17812,N_17271,N_17442);
xor U17813 (N_17813,N_17482,N_17593);
xnor U17814 (N_17814,N_17576,N_17331);
xnor U17815 (N_17815,N_17570,N_17437);
and U17816 (N_17816,N_17464,N_17470);
nor U17817 (N_17817,N_17222,N_17506);
nand U17818 (N_17818,N_17498,N_17511);
nand U17819 (N_17819,N_17599,N_17351);
xnor U17820 (N_17820,N_17396,N_17475);
or U17821 (N_17821,N_17226,N_17266);
xor U17822 (N_17822,N_17200,N_17320);
nand U17823 (N_17823,N_17263,N_17562);
nand U17824 (N_17824,N_17357,N_17412);
xnor U17825 (N_17825,N_17288,N_17201);
nor U17826 (N_17826,N_17219,N_17360);
xnor U17827 (N_17827,N_17517,N_17243);
xnor U17828 (N_17828,N_17398,N_17509);
nor U17829 (N_17829,N_17321,N_17484);
or U17830 (N_17830,N_17257,N_17523);
nor U17831 (N_17831,N_17411,N_17360);
nor U17832 (N_17832,N_17222,N_17352);
nor U17833 (N_17833,N_17417,N_17325);
and U17834 (N_17834,N_17478,N_17395);
and U17835 (N_17835,N_17298,N_17535);
or U17836 (N_17836,N_17585,N_17394);
nand U17837 (N_17837,N_17548,N_17238);
or U17838 (N_17838,N_17409,N_17530);
nor U17839 (N_17839,N_17403,N_17435);
and U17840 (N_17840,N_17496,N_17400);
nand U17841 (N_17841,N_17437,N_17549);
and U17842 (N_17842,N_17427,N_17557);
nand U17843 (N_17843,N_17521,N_17351);
or U17844 (N_17844,N_17488,N_17254);
or U17845 (N_17845,N_17555,N_17574);
or U17846 (N_17846,N_17591,N_17599);
xnor U17847 (N_17847,N_17403,N_17553);
nor U17848 (N_17848,N_17573,N_17302);
and U17849 (N_17849,N_17468,N_17218);
and U17850 (N_17850,N_17387,N_17269);
nand U17851 (N_17851,N_17560,N_17429);
nor U17852 (N_17852,N_17460,N_17267);
xor U17853 (N_17853,N_17523,N_17351);
nand U17854 (N_17854,N_17446,N_17523);
and U17855 (N_17855,N_17423,N_17571);
nand U17856 (N_17856,N_17587,N_17389);
nor U17857 (N_17857,N_17243,N_17402);
or U17858 (N_17858,N_17502,N_17538);
nand U17859 (N_17859,N_17583,N_17432);
nor U17860 (N_17860,N_17346,N_17397);
and U17861 (N_17861,N_17450,N_17289);
and U17862 (N_17862,N_17234,N_17565);
xor U17863 (N_17863,N_17380,N_17304);
or U17864 (N_17864,N_17515,N_17364);
nand U17865 (N_17865,N_17427,N_17356);
xor U17866 (N_17866,N_17582,N_17568);
and U17867 (N_17867,N_17485,N_17211);
and U17868 (N_17868,N_17357,N_17537);
nor U17869 (N_17869,N_17553,N_17573);
nor U17870 (N_17870,N_17200,N_17288);
and U17871 (N_17871,N_17430,N_17367);
nand U17872 (N_17872,N_17419,N_17536);
nor U17873 (N_17873,N_17586,N_17292);
or U17874 (N_17874,N_17362,N_17533);
xnor U17875 (N_17875,N_17561,N_17342);
nor U17876 (N_17876,N_17452,N_17441);
nand U17877 (N_17877,N_17359,N_17200);
nand U17878 (N_17878,N_17399,N_17377);
nor U17879 (N_17879,N_17370,N_17333);
nor U17880 (N_17880,N_17388,N_17334);
nor U17881 (N_17881,N_17504,N_17448);
xnor U17882 (N_17882,N_17552,N_17536);
nand U17883 (N_17883,N_17422,N_17353);
or U17884 (N_17884,N_17361,N_17242);
xnor U17885 (N_17885,N_17256,N_17495);
nor U17886 (N_17886,N_17405,N_17578);
nand U17887 (N_17887,N_17540,N_17265);
nor U17888 (N_17888,N_17572,N_17466);
nor U17889 (N_17889,N_17498,N_17506);
nand U17890 (N_17890,N_17304,N_17290);
xnor U17891 (N_17891,N_17261,N_17528);
xnor U17892 (N_17892,N_17590,N_17218);
nand U17893 (N_17893,N_17393,N_17236);
nand U17894 (N_17894,N_17531,N_17266);
or U17895 (N_17895,N_17538,N_17491);
and U17896 (N_17896,N_17581,N_17448);
and U17897 (N_17897,N_17257,N_17216);
xnor U17898 (N_17898,N_17296,N_17348);
nand U17899 (N_17899,N_17243,N_17315);
and U17900 (N_17900,N_17292,N_17475);
nand U17901 (N_17901,N_17325,N_17462);
nor U17902 (N_17902,N_17347,N_17450);
nand U17903 (N_17903,N_17450,N_17454);
xor U17904 (N_17904,N_17219,N_17585);
nand U17905 (N_17905,N_17334,N_17579);
or U17906 (N_17906,N_17452,N_17375);
nand U17907 (N_17907,N_17331,N_17285);
nor U17908 (N_17908,N_17392,N_17596);
xnor U17909 (N_17909,N_17397,N_17486);
nor U17910 (N_17910,N_17289,N_17556);
or U17911 (N_17911,N_17452,N_17501);
nand U17912 (N_17912,N_17499,N_17349);
and U17913 (N_17913,N_17353,N_17285);
nor U17914 (N_17914,N_17559,N_17579);
nor U17915 (N_17915,N_17379,N_17439);
and U17916 (N_17916,N_17323,N_17447);
xor U17917 (N_17917,N_17516,N_17369);
nand U17918 (N_17918,N_17566,N_17201);
nand U17919 (N_17919,N_17416,N_17205);
nand U17920 (N_17920,N_17332,N_17289);
nor U17921 (N_17921,N_17593,N_17496);
and U17922 (N_17922,N_17418,N_17305);
nand U17923 (N_17923,N_17577,N_17201);
or U17924 (N_17924,N_17322,N_17391);
and U17925 (N_17925,N_17388,N_17599);
nand U17926 (N_17926,N_17515,N_17217);
nand U17927 (N_17927,N_17459,N_17264);
nand U17928 (N_17928,N_17447,N_17366);
and U17929 (N_17929,N_17432,N_17317);
xor U17930 (N_17930,N_17578,N_17543);
nand U17931 (N_17931,N_17388,N_17337);
and U17932 (N_17932,N_17520,N_17363);
nor U17933 (N_17933,N_17365,N_17405);
or U17934 (N_17934,N_17365,N_17294);
xor U17935 (N_17935,N_17589,N_17456);
nand U17936 (N_17936,N_17540,N_17497);
xor U17937 (N_17937,N_17249,N_17392);
nor U17938 (N_17938,N_17334,N_17440);
and U17939 (N_17939,N_17489,N_17526);
and U17940 (N_17940,N_17267,N_17280);
xor U17941 (N_17941,N_17318,N_17281);
nand U17942 (N_17942,N_17287,N_17209);
xnor U17943 (N_17943,N_17393,N_17496);
and U17944 (N_17944,N_17571,N_17452);
nor U17945 (N_17945,N_17229,N_17221);
nand U17946 (N_17946,N_17430,N_17482);
nand U17947 (N_17947,N_17208,N_17264);
nor U17948 (N_17948,N_17443,N_17385);
or U17949 (N_17949,N_17256,N_17544);
or U17950 (N_17950,N_17262,N_17296);
nor U17951 (N_17951,N_17393,N_17408);
nand U17952 (N_17952,N_17303,N_17419);
and U17953 (N_17953,N_17476,N_17265);
nand U17954 (N_17954,N_17270,N_17517);
and U17955 (N_17955,N_17415,N_17345);
and U17956 (N_17956,N_17541,N_17327);
or U17957 (N_17957,N_17260,N_17378);
nor U17958 (N_17958,N_17279,N_17596);
and U17959 (N_17959,N_17275,N_17417);
nand U17960 (N_17960,N_17566,N_17490);
xnor U17961 (N_17961,N_17381,N_17525);
xnor U17962 (N_17962,N_17301,N_17221);
xnor U17963 (N_17963,N_17534,N_17263);
xnor U17964 (N_17964,N_17477,N_17414);
and U17965 (N_17965,N_17579,N_17319);
nor U17966 (N_17966,N_17428,N_17532);
or U17967 (N_17967,N_17227,N_17229);
nand U17968 (N_17968,N_17580,N_17513);
xnor U17969 (N_17969,N_17508,N_17380);
xnor U17970 (N_17970,N_17463,N_17250);
or U17971 (N_17971,N_17239,N_17211);
nor U17972 (N_17972,N_17207,N_17585);
nand U17973 (N_17973,N_17256,N_17360);
nand U17974 (N_17974,N_17359,N_17292);
nor U17975 (N_17975,N_17514,N_17262);
or U17976 (N_17976,N_17396,N_17342);
nand U17977 (N_17977,N_17323,N_17456);
or U17978 (N_17978,N_17598,N_17396);
nand U17979 (N_17979,N_17379,N_17339);
nor U17980 (N_17980,N_17518,N_17393);
nand U17981 (N_17981,N_17401,N_17240);
and U17982 (N_17982,N_17464,N_17226);
and U17983 (N_17983,N_17407,N_17393);
nand U17984 (N_17984,N_17467,N_17527);
or U17985 (N_17985,N_17380,N_17443);
or U17986 (N_17986,N_17309,N_17240);
or U17987 (N_17987,N_17260,N_17285);
xnor U17988 (N_17988,N_17260,N_17547);
and U17989 (N_17989,N_17218,N_17479);
nand U17990 (N_17990,N_17215,N_17478);
nand U17991 (N_17991,N_17550,N_17217);
nand U17992 (N_17992,N_17270,N_17343);
nor U17993 (N_17993,N_17297,N_17549);
xor U17994 (N_17994,N_17434,N_17547);
and U17995 (N_17995,N_17412,N_17342);
and U17996 (N_17996,N_17297,N_17391);
and U17997 (N_17997,N_17267,N_17495);
nor U17998 (N_17998,N_17296,N_17430);
xnor U17999 (N_17999,N_17211,N_17372);
nand U18000 (N_18000,N_17844,N_17742);
nand U18001 (N_18001,N_17995,N_17609);
nor U18002 (N_18002,N_17600,N_17746);
or U18003 (N_18003,N_17998,N_17829);
xor U18004 (N_18004,N_17902,N_17707);
and U18005 (N_18005,N_17868,N_17643);
nor U18006 (N_18006,N_17860,N_17627);
or U18007 (N_18007,N_17881,N_17685);
nor U18008 (N_18008,N_17726,N_17740);
or U18009 (N_18009,N_17852,N_17831);
nand U18010 (N_18010,N_17745,N_17792);
nand U18011 (N_18011,N_17678,N_17786);
xor U18012 (N_18012,N_17640,N_17946);
nor U18013 (N_18013,N_17862,N_17762);
nor U18014 (N_18014,N_17624,N_17700);
or U18015 (N_18015,N_17670,N_17933);
xnor U18016 (N_18016,N_17602,N_17721);
and U18017 (N_18017,N_17833,N_17729);
nand U18018 (N_18018,N_17992,N_17774);
nand U18019 (N_18019,N_17922,N_17848);
xnor U18020 (N_18020,N_17728,N_17855);
or U18021 (N_18021,N_17814,N_17790);
xor U18022 (N_18022,N_17949,N_17921);
nor U18023 (N_18023,N_17972,N_17611);
and U18024 (N_18024,N_17645,N_17706);
xor U18025 (N_18025,N_17626,N_17966);
nor U18026 (N_18026,N_17675,N_17895);
xnor U18027 (N_18027,N_17928,N_17925);
xor U18028 (N_18028,N_17956,N_17771);
and U18029 (N_18029,N_17867,N_17646);
xnor U18030 (N_18030,N_17899,N_17840);
or U18031 (N_18031,N_17976,N_17770);
nand U18032 (N_18032,N_17942,N_17669);
xnor U18033 (N_18033,N_17847,N_17871);
nand U18034 (N_18034,N_17679,N_17621);
nor U18035 (N_18035,N_17781,N_17690);
nand U18036 (N_18036,N_17959,N_17967);
nor U18037 (N_18037,N_17761,N_17910);
xor U18038 (N_18038,N_17904,N_17725);
nor U18039 (N_18039,N_17633,N_17658);
nand U18040 (N_18040,N_17912,N_17744);
nor U18041 (N_18041,N_17913,N_17751);
or U18042 (N_18042,N_17954,N_17653);
nor U18043 (N_18043,N_17684,N_17939);
and U18044 (N_18044,N_17615,N_17769);
and U18045 (N_18045,N_17806,N_17782);
xor U18046 (N_18046,N_17756,N_17656);
nand U18047 (N_18047,N_17681,N_17632);
and U18048 (N_18048,N_17758,N_17647);
and U18049 (N_18049,N_17808,N_17642);
or U18050 (N_18050,N_17957,N_17962);
nor U18051 (N_18051,N_17672,N_17694);
nand U18052 (N_18052,N_17735,N_17733);
or U18053 (N_18053,N_17858,N_17603);
nand U18054 (N_18054,N_17613,N_17631);
xnor U18055 (N_18055,N_17724,N_17630);
nand U18056 (N_18056,N_17604,N_17826);
nor U18057 (N_18057,N_17837,N_17650);
xor U18058 (N_18058,N_17897,N_17971);
and U18059 (N_18059,N_17827,N_17709);
and U18060 (N_18060,N_17951,N_17661);
nor U18061 (N_18061,N_17984,N_17736);
xnor U18062 (N_18062,N_17809,N_17875);
xor U18063 (N_18063,N_17961,N_17828);
nand U18064 (N_18064,N_17916,N_17749);
xnor U18065 (N_18065,N_17815,N_17686);
nor U18066 (N_18066,N_17738,N_17702);
or U18067 (N_18067,N_17993,N_17796);
nand U18068 (N_18068,N_17698,N_17877);
nand U18069 (N_18069,N_17915,N_17789);
nor U18070 (N_18070,N_17955,N_17964);
xor U18071 (N_18071,N_17682,N_17811);
nand U18072 (N_18072,N_17989,N_17885);
xor U18073 (N_18073,N_17919,N_17773);
and U18074 (N_18074,N_17823,N_17715);
nand U18075 (N_18075,N_17768,N_17930);
xor U18076 (N_18076,N_17937,N_17605);
nor U18077 (N_18077,N_17798,N_17634);
or U18078 (N_18078,N_17987,N_17772);
nand U18079 (N_18079,N_17610,N_17824);
xor U18080 (N_18080,N_17652,N_17854);
or U18081 (N_18081,N_17960,N_17657);
nand U18082 (N_18082,N_17635,N_17775);
and U18083 (N_18083,N_17607,N_17932);
xor U18084 (N_18084,N_17812,N_17842);
xnor U18085 (N_18085,N_17759,N_17901);
or U18086 (N_18086,N_17861,N_17628);
and U18087 (N_18087,N_17799,N_17648);
nor U18088 (N_18088,N_17903,N_17780);
and U18089 (N_18089,N_17760,N_17801);
and U18090 (N_18090,N_17950,N_17712);
and U18091 (N_18091,N_17920,N_17965);
nand U18092 (N_18092,N_17870,N_17890);
or U18093 (N_18093,N_17716,N_17680);
and U18094 (N_18094,N_17893,N_17739);
nor U18095 (N_18095,N_17664,N_17662);
nor U18096 (N_18096,N_17636,N_17825);
or U18097 (N_18097,N_17934,N_17718);
xnor U18098 (N_18098,N_17654,N_17838);
nor U18099 (N_18099,N_17800,N_17975);
and U18100 (N_18100,N_17918,N_17791);
xnor U18101 (N_18101,N_17804,N_17817);
and U18102 (N_18102,N_17834,N_17793);
nor U18103 (N_18103,N_17730,N_17889);
nor U18104 (N_18104,N_17944,N_17639);
and U18105 (N_18105,N_17969,N_17671);
nand U18106 (N_18106,N_17990,N_17754);
nor U18107 (N_18107,N_17908,N_17982);
or U18108 (N_18108,N_17708,N_17601);
and U18109 (N_18109,N_17963,N_17689);
or U18110 (N_18110,N_17991,N_17649);
nor U18111 (N_18111,N_17637,N_17620);
xnor U18112 (N_18112,N_17926,N_17734);
and U18113 (N_18113,N_17765,N_17947);
xnor U18114 (N_18114,N_17936,N_17673);
or U18115 (N_18115,N_17625,N_17722);
xnor U18116 (N_18116,N_17898,N_17999);
nand U18117 (N_18117,N_17803,N_17612);
and U18118 (N_18118,N_17900,N_17695);
xor U18119 (N_18119,N_17731,N_17785);
nor U18120 (N_18120,N_17835,N_17667);
and U18121 (N_18121,N_17927,N_17655);
or U18122 (N_18122,N_17948,N_17952);
or U18123 (N_18123,N_17874,N_17914);
or U18124 (N_18124,N_17713,N_17660);
and U18125 (N_18125,N_17909,N_17979);
nor U18126 (N_18126,N_17651,N_17906);
nor U18127 (N_18127,N_17880,N_17720);
xnor U18128 (N_18128,N_17986,N_17691);
xnor U18129 (N_18129,N_17978,N_17666);
nor U18130 (N_18130,N_17816,N_17813);
or U18131 (N_18131,N_17894,N_17851);
xor U18132 (N_18132,N_17787,N_17614);
xor U18133 (N_18133,N_17766,N_17940);
nand U18134 (N_18134,N_17763,N_17703);
nand U18135 (N_18135,N_17767,N_17832);
nand U18136 (N_18136,N_17737,N_17981);
nand U18137 (N_18137,N_17887,N_17616);
nand U18138 (N_18138,N_17714,N_17841);
nand U18139 (N_18139,N_17983,N_17710);
nand U18140 (N_18140,N_17997,N_17864);
nor U18141 (N_18141,N_17866,N_17846);
nand U18142 (N_18142,N_17917,N_17687);
nand U18143 (N_18143,N_17886,N_17968);
nor U18144 (N_18144,N_17757,N_17945);
nor U18145 (N_18145,N_17820,N_17723);
and U18146 (N_18146,N_17872,N_17873);
nor U18147 (N_18147,N_17638,N_17704);
and U18148 (N_18148,N_17911,N_17974);
nand U18149 (N_18149,N_17629,N_17929);
and U18150 (N_18150,N_17705,N_17802);
nand U18151 (N_18151,N_17943,N_17663);
and U18152 (N_18152,N_17849,N_17797);
and U18153 (N_18153,N_17891,N_17821);
or U18154 (N_18154,N_17699,N_17924);
or U18155 (N_18155,N_17883,N_17853);
xnor U18156 (N_18156,N_17985,N_17884);
nand U18157 (N_18157,N_17779,N_17750);
and U18158 (N_18158,N_17810,N_17644);
or U18159 (N_18159,N_17784,N_17953);
or U18160 (N_18160,N_17980,N_17727);
nor U18161 (N_18161,N_17988,N_17896);
and U18162 (N_18162,N_17958,N_17683);
xnor U18163 (N_18163,N_17677,N_17776);
or U18164 (N_18164,N_17973,N_17888);
or U18165 (N_18165,N_17859,N_17818);
xnor U18166 (N_18166,N_17619,N_17819);
nand U18167 (N_18167,N_17606,N_17665);
or U18168 (N_18168,N_17905,N_17747);
xnor U18169 (N_18169,N_17892,N_17688);
or U18170 (N_18170,N_17623,N_17830);
xnor U18171 (N_18171,N_17996,N_17676);
xor U18172 (N_18172,N_17836,N_17882);
or U18173 (N_18173,N_17674,N_17805);
nand U18174 (N_18174,N_17641,N_17907);
xor U18175 (N_18175,N_17923,N_17783);
or U18176 (N_18176,N_17743,N_17931);
or U18177 (N_18177,N_17618,N_17701);
and U18178 (N_18178,N_17879,N_17970);
and U18179 (N_18179,N_17935,N_17845);
or U18180 (N_18180,N_17697,N_17807);
nor U18181 (N_18181,N_17764,N_17693);
xnor U18182 (N_18182,N_17696,N_17732);
or U18183 (N_18183,N_17857,N_17994);
xor U18184 (N_18184,N_17752,N_17748);
and U18185 (N_18185,N_17822,N_17692);
nor U18186 (N_18186,N_17876,N_17795);
nand U18187 (N_18187,N_17977,N_17711);
nor U18188 (N_18188,N_17878,N_17869);
and U18189 (N_18189,N_17753,N_17608);
xnor U18190 (N_18190,N_17863,N_17622);
xnor U18191 (N_18191,N_17719,N_17777);
or U18192 (N_18192,N_17850,N_17938);
or U18193 (N_18193,N_17788,N_17755);
nand U18194 (N_18194,N_17717,N_17659);
nor U18195 (N_18195,N_17856,N_17843);
xor U18196 (N_18196,N_17778,N_17668);
xor U18197 (N_18197,N_17839,N_17741);
or U18198 (N_18198,N_17794,N_17941);
nor U18199 (N_18199,N_17865,N_17617);
nor U18200 (N_18200,N_17719,N_17960);
nand U18201 (N_18201,N_17809,N_17601);
xnor U18202 (N_18202,N_17938,N_17728);
and U18203 (N_18203,N_17806,N_17855);
nor U18204 (N_18204,N_17861,N_17743);
and U18205 (N_18205,N_17921,N_17641);
nand U18206 (N_18206,N_17956,N_17938);
nor U18207 (N_18207,N_17926,N_17777);
and U18208 (N_18208,N_17702,N_17654);
or U18209 (N_18209,N_17806,N_17822);
and U18210 (N_18210,N_17819,N_17631);
xor U18211 (N_18211,N_17999,N_17830);
nor U18212 (N_18212,N_17831,N_17795);
or U18213 (N_18213,N_17669,N_17876);
or U18214 (N_18214,N_17977,N_17820);
nand U18215 (N_18215,N_17621,N_17743);
nor U18216 (N_18216,N_17723,N_17900);
or U18217 (N_18217,N_17683,N_17909);
xor U18218 (N_18218,N_17907,N_17730);
nand U18219 (N_18219,N_17815,N_17813);
nor U18220 (N_18220,N_17829,N_17706);
and U18221 (N_18221,N_17769,N_17788);
nor U18222 (N_18222,N_17770,N_17920);
xnor U18223 (N_18223,N_17998,N_17852);
xor U18224 (N_18224,N_17715,N_17884);
nor U18225 (N_18225,N_17836,N_17997);
xnor U18226 (N_18226,N_17872,N_17790);
xor U18227 (N_18227,N_17691,N_17796);
and U18228 (N_18228,N_17862,N_17730);
and U18229 (N_18229,N_17772,N_17907);
nand U18230 (N_18230,N_17931,N_17939);
nor U18231 (N_18231,N_17902,N_17746);
xor U18232 (N_18232,N_17606,N_17745);
xnor U18233 (N_18233,N_17755,N_17957);
xor U18234 (N_18234,N_17722,N_17612);
nand U18235 (N_18235,N_17818,N_17788);
or U18236 (N_18236,N_17709,N_17626);
and U18237 (N_18237,N_17683,N_17647);
or U18238 (N_18238,N_17603,N_17794);
nor U18239 (N_18239,N_17845,N_17700);
xnor U18240 (N_18240,N_17727,N_17659);
nor U18241 (N_18241,N_17658,N_17750);
or U18242 (N_18242,N_17606,N_17816);
and U18243 (N_18243,N_17905,N_17801);
and U18244 (N_18244,N_17604,N_17789);
nor U18245 (N_18245,N_17855,N_17835);
and U18246 (N_18246,N_17656,N_17939);
or U18247 (N_18247,N_17778,N_17864);
nor U18248 (N_18248,N_17984,N_17783);
nor U18249 (N_18249,N_17893,N_17871);
and U18250 (N_18250,N_17794,N_17776);
and U18251 (N_18251,N_17966,N_17625);
or U18252 (N_18252,N_17668,N_17745);
nand U18253 (N_18253,N_17954,N_17830);
or U18254 (N_18254,N_17771,N_17916);
and U18255 (N_18255,N_17736,N_17877);
or U18256 (N_18256,N_17630,N_17662);
and U18257 (N_18257,N_17752,N_17670);
nand U18258 (N_18258,N_17610,N_17643);
or U18259 (N_18259,N_17969,N_17680);
nor U18260 (N_18260,N_17764,N_17839);
nand U18261 (N_18261,N_17905,N_17806);
xor U18262 (N_18262,N_17799,N_17793);
and U18263 (N_18263,N_17908,N_17985);
nor U18264 (N_18264,N_17668,N_17713);
nor U18265 (N_18265,N_17991,N_17777);
xor U18266 (N_18266,N_17812,N_17719);
nor U18267 (N_18267,N_17758,N_17896);
xor U18268 (N_18268,N_17657,N_17951);
nor U18269 (N_18269,N_17951,N_17730);
xor U18270 (N_18270,N_17950,N_17776);
nor U18271 (N_18271,N_17604,N_17610);
nand U18272 (N_18272,N_17639,N_17770);
or U18273 (N_18273,N_17747,N_17659);
and U18274 (N_18274,N_17965,N_17781);
or U18275 (N_18275,N_17628,N_17970);
nand U18276 (N_18276,N_17754,N_17789);
nor U18277 (N_18277,N_17636,N_17811);
and U18278 (N_18278,N_17838,N_17986);
nand U18279 (N_18279,N_17669,N_17625);
or U18280 (N_18280,N_17729,N_17697);
xor U18281 (N_18281,N_17994,N_17610);
nand U18282 (N_18282,N_17853,N_17805);
xnor U18283 (N_18283,N_17659,N_17627);
nand U18284 (N_18284,N_17693,N_17909);
and U18285 (N_18285,N_17746,N_17702);
xnor U18286 (N_18286,N_17824,N_17646);
or U18287 (N_18287,N_17617,N_17812);
nor U18288 (N_18288,N_17779,N_17860);
nor U18289 (N_18289,N_17940,N_17661);
xor U18290 (N_18290,N_17649,N_17787);
xor U18291 (N_18291,N_17772,N_17798);
nand U18292 (N_18292,N_17979,N_17612);
nand U18293 (N_18293,N_17937,N_17918);
or U18294 (N_18294,N_17767,N_17725);
xor U18295 (N_18295,N_17626,N_17954);
nor U18296 (N_18296,N_17927,N_17751);
nor U18297 (N_18297,N_17677,N_17796);
xor U18298 (N_18298,N_17892,N_17653);
xor U18299 (N_18299,N_17723,N_17630);
and U18300 (N_18300,N_17612,N_17689);
or U18301 (N_18301,N_17877,N_17963);
nand U18302 (N_18302,N_17795,N_17725);
and U18303 (N_18303,N_17913,N_17958);
nor U18304 (N_18304,N_17697,N_17847);
and U18305 (N_18305,N_17833,N_17675);
nor U18306 (N_18306,N_17834,N_17669);
or U18307 (N_18307,N_17779,N_17678);
nor U18308 (N_18308,N_17672,N_17707);
or U18309 (N_18309,N_17777,N_17723);
xnor U18310 (N_18310,N_17910,N_17992);
nand U18311 (N_18311,N_17827,N_17933);
xor U18312 (N_18312,N_17669,N_17771);
or U18313 (N_18313,N_17939,N_17651);
nand U18314 (N_18314,N_17985,N_17890);
xor U18315 (N_18315,N_17616,N_17877);
and U18316 (N_18316,N_17843,N_17834);
and U18317 (N_18317,N_17918,N_17969);
nand U18318 (N_18318,N_17706,N_17880);
or U18319 (N_18319,N_17814,N_17609);
or U18320 (N_18320,N_17744,N_17860);
and U18321 (N_18321,N_17826,N_17692);
or U18322 (N_18322,N_17732,N_17679);
xnor U18323 (N_18323,N_17917,N_17885);
nor U18324 (N_18324,N_17606,N_17608);
xnor U18325 (N_18325,N_17727,N_17895);
or U18326 (N_18326,N_17846,N_17770);
or U18327 (N_18327,N_17736,N_17743);
or U18328 (N_18328,N_17692,N_17735);
nand U18329 (N_18329,N_17947,N_17935);
nor U18330 (N_18330,N_17795,N_17890);
and U18331 (N_18331,N_17715,N_17814);
or U18332 (N_18332,N_17650,N_17918);
and U18333 (N_18333,N_17748,N_17638);
and U18334 (N_18334,N_17703,N_17880);
or U18335 (N_18335,N_17646,N_17854);
nor U18336 (N_18336,N_17985,N_17943);
or U18337 (N_18337,N_17686,N_17729);
and U18338 (N_18338,N_17898,N_17701);
and U18339 (N_18339,N_17799,N_17697);
xor U18340 (N_18340,N_17989,N_17873);
or U18341 (N_18341,N_17828,N_17752);
nand U18342 (N_18342,N_17618,N_17844);
or U18343 (N_18343,N_17626,N_17881);
and U18344 (N_18344,N_17723,N_17946);
or U18345 (N_18345,N_17929,N_17993);
and U18346 (N_18346,N_17627,N_17960);
nand U18347 (N_18347,N_17716,N_17857);
or U18348 (N_18348,N_17681,N_17877);
nor U18349 (N_18349,N_17669,N_17630);
and U18350 (N_18350,N_17772,N_17638);
nand U18351 (N_18351,N_17966,N_17933);
xor U18352 (N_18352,N_17849,N_17606);
nand U18353 (N_18353,N_17952,N_17826);
nand U18354 (N_18354,N_17772,N_17942);
nor U18355 (N_18355,N_17839,N_17612);
and U18356 (N_18356,N_17775,N_17874);
and U18357 (N_18357,N_17941,N_17782);
xor U18358 (N_18358,N_17676,N_17871);
xor U18359 (N_18359,N_17744,N_17958);
or U18360 (N_18360,N_17962,N_17987);
xor U18361 (N_18361,N_17819,N_17830);
nand U18362 (N_18362,N_17654,N_17624);
and U18363 (N_18363,N_17654,N_17628);
xor U18364 (N_18364,N_17836,N_17887);
and U18365 (N_18365,N_17993,N_17818);
or U18366 (N_18366,N_17683,N_17752);
or U18367 (N_18367,N_17647,N_17760);
and U18368 (N_18368,N_17718,N_17838);
nand U18369 (N_18369,N_17607,N_17990);
xor U18370 (N_18370,N_17617,N_17627);
nand U18371 (N_18371,N_17712,N_17780);
and U18372 (N_18372,N_17833,N_17996);
xor U18373 (N_18373,N_17612,N_17772);
nor U18374 (N_18374,N_17702,N_17634);
and U18375 (N_18375,N_17775,N_17814);
nand U18376 (N_18376,N_17858,N_17985);
xor U18377 (N_18377,N_17643,N_17658);
xnor U18378 (N_18378,N_17622,N_17811);
xor U18379 (N_18379,N_17694,N_17893);
nand U18380 (N_18380,N_17945,N_17762);
nor U18381 (N_18381,N_17731,N_17621);
xnor U18382 (N_18382,N_17946,N_17692);
and U18383 (N_18383,N_17823,N_17721);
nor U18384 (N_18384,N_17709,N_17776);
xor U18385 (N_18385,N_17811,N_17915);
and U18386 (N_18386,N_17757,N_17813);
nor U18387 (N_18387,N_17826,N_17957);
nand U18388 (N_18388,N_17833,N_17888);
or U18389 (N_18389,N_17679,N_17717);
and U18390 (N_18390,N_17775,N_17994);
nor U18391 (N_18391,N_17971,N_17759);
xnor U18392 (N_18392,N_17789,N_17649);
nor U18393 (N_18393,N_17722,N_17946);
and U18394 (N_18394,N_17753,N_17874);
or U18395 (N_18395,N_17930,N_17912);
or U18396 (N_18396,N_17981,N_17921);
xnor U18397 (N_18397,N_17803,N_17990);
or U18398 (N_18398,N_17762,N_17715);
and U18399 (N_18399,N_17906,N_17927);
and U18400 (N_18400,N_18118,N_18363);
or U18401 (N_18401,N_18180,N_18396);
nor U18402 (N_18402,N_18083,N_18288);
or U18403 (N_18403,N_18240,N_18225);
or U18404 (N_18404,N_18060,N_18094);
and U18405 (N_18405,N_18297,N_18177);
xor U18406 (N_18406,N_18127,N_18069);
or U18407 (N_18407,N_18107,N_18277);
nand U18408 (N_18408,N_18052,N_18167);
nor U18409 (N_18409,N_18186,N_18384);
and U18410 (N_18410,N_18054,N_18019);
nand U18411 (N_18411,N_18174,N_18124);
or U18412 (N_18412,N_18189,N_18279);
xnor U18413 (N_18413,N_18151,N_18373);
or U18414 (N_18414,N_18275,N_18294);
xnor U18415 (N_18415,N_18222,N_18377);
nor U18416 (N_18416,N_18047,N_18133);
or U18417 (N_18417,N_18257,N_18205);
or U18418 (N_18418,N_18187,N_18261);
xnor U18419 (N_18419,N_18276,N_18059);
or U18420 (N_18420,N_18335,N_18082);
nand U18421 (N_18421,N_18101,N_18226);
xor U18422 (N_18422,N_18175,N_18330);
or U18423 (N_18423,N_18302,N_18134);
or U18424 (N_18424,N_18185,N_18049);
nand U18425 (N_18425,N_18084,N_18166);
xnor U18426 (N_18426,N_18280,N_18221);
or U18427 (N_18427,N_18292,N_18295);
and U18428 (N_18428,N_18285,N_18190);
or U18429 (N_18429,N_18372,N_18150);
xor U18430 (N_18430,N_18341,N_18308);
or U18431 (N_18431,N_18304,N_18154);
or U18432 (N_18432,N_18013,N_18207);
nor U18433 (N_18433,N_18228,N_18326);
or U18434 (N_18434,N_18340,N_18345);
and U18435 (N_18435,N_18193,N_18259);
nor U18436 (N_18436,N_18130,N_18145);
xor U18437 (N_18437,N_18367,N_18290);
xnor U18438 (N_18438,N_18212,N_18022);
nor U18439 (N_18439,N_18119,N_18202);
nand U18440 (N_18440,N_18139,N_18243);
or U18441 (N_18441,N_18195,N_18293);
and U18442 (N_18442,N_18040,N_18080);
xor U18443 (N_18443,N_18048,N_18036);
and U18444 (N_18444,N_18244,N_18178);
or U18445 (N_18445,N_18387,N_18067);
nand U18446 (N_18446,N_18092,N_18135);
nand U18447 (N_18447,N_18374,N_18351);
xnor U18448 (N_18448,N_18254,N_18021);
xnor U18449 (N_18449,N_18283,N_18129);
nor U18450 (N_18450,N_18072,N_18126);
xnor U18451 (N_18451,N_18332,N_18336);
and U18452 (N_18452,N_18016,N_18309);
and U18453 (N_18453,N_18220,N_18123);
and U18454 (N_18454,N_18322,N_18039);
and U18455 (N_18455,N_18306,N_18331);
nor U18456 (N_18456,N_18091,N_18256);
and U18457 (N_18457,N_18110,N_18089);
xnor U18458 (N_18458,N_18201,N_18017);
nand U18459 (N_18459,N_18375,N_18313);
nor U18460 (N_18460,N_18081,N_18246);
nor U18461 (N_18461,N_18128,N_18064);
and U18462 (N_18462,N_18090,N_18149);
or U18463 (N_18463,N_18323,N_18156);
and U18464 (N_18464,N_18355,N_18338);
xnor U18465 (N_18465,N_18038,N_18024);
nand U18466 (N_18466,N_18380,N_18362);
nor U18467 (N_18467,N_18142,N_18321);
nor U18468 (N_18468,N_18121,N_18171);
xor U18469 (N_18469,N_18028,N_18043);
and U18470 (N_18470,N_18381,N_18312);
nor U18471 (N_18471,N_18366,N_18242);
xor U18472 (N_18472,N_18271,N_18010);
nor U18473 (N_18473,N_18162,N_18211);
nor U18474 (N_18474,N_18389,N_18347);
or U18475 (N_18475,N_18179,N_18291);
nor U18476 (N_18476,N_18216,N_18266);
nand U18477 (N_18477,N_18392,N_18305);
xnor U18478 (N_18478,N_18289,N_18164);
nand U18479 (N_18479,N_18074,N_18388);
nand U18480 (N_18480,N_18298,N_18001);
xor U18481 (N_18481,N_18035,N_18192);
and U18482 (N_18482,N_18329,N_18217);
or U18483 (N_18483,N_18112,N_18364);
or U18484 (N_18484,N_18109,N_18100);
nor U18485 (N_18485,N_18070,N_18218);
or U18486 (N_18486,N_18147,N_18353);
xnor U18487 (N_18487,N_18268,N_18030);
nor U18488 (N_18488,N_18004,N_18324);
or U18489 (N_18489,N_18394,N_18042);
nor U18490 (N_18490,N_18311,N_18235);
nand U18491 (N_18491,N_18209,N_18037);
or U18492 (N_18492,N_18076,N_18066);
nor U18493 (N_18493,N_18265,N_18344);
and U18494 (N_18494,N_18114,N_18391);
and U18495 (N_18495,N_18029,N_18386);
and U18496 (N_18496,N_18231,N_18223);
nand U18497 (N_18497,N_18073,N_18262);
nand U18498 (N_18498,N_18153,N_18095);
xnor U18499 (N_18499,N_18328,N_18274);
or U18500 (N_18500,N_18077,N_18249);
xor U18501 (N_18501,N_18005,N_18334);
nor U18502 (N_18502,N_18346,N_18104);
nand U18503 (N_18503,N_18361,N_18057);
nand U18504 (N_18504,N_18120,N_18342);
nor U18505 (N_18505,N_18065,N_18356);
or U18506 (N_18506,N_18273,N_18315);
or U18507 (N_18507,N_18034,N_18371);
or U18508 (N_18508,N_18258,N_18234);
nand U18509 (N_18509,N_18337,N_18333);
xnor U18510 (N_18510,N_18055,N_18011);
or U18511 (N_18511,N_18284,N_18317);
and U18512 (N_18512,N_18318,N_18208);
and U18513 (N_18513,N_18003,N_18354);
or U18514 (N_18514,N_18339,N_18390);
nor U18515 (N_18515,N_18232,N_18163);
nand U18516 (N_18516,N_18105,N_18172);
nand U18517 (N_18517,N_18161,N_18320);
and U18518 (N_18518,N_18141,N_18278);
or U18519 (N_18519,N_18009,N_18097);
and U18520 (N_18520,N_18044,N_18236);
nor U18521 (N_18521,N_18144,N_18146);
nand U18522 (N_18522,N_18008,N_18007);
xor U18523 (N_18523,N_18058,N_18379);
and U18524 (N_18524,N_18111,N_18224);
or U18525 (N_18525,N_18018,N_18108);
and U18526 (N_18526,N_18238,N_18117);
nor U18527 (N_18527,N_18296,N_18061);
nand U18528 (N_18528,N_18071,N_18300);
nor U18529 (N_18529,N_18382,N_18113);
nand U18530 (N_18530,N_18213,N_18376);
nand U18531 (N_18531,N_18173,N_18203);
or U18532 (N_18532,N_18063,N_18184);
nor U18533 (N_18533,N_18196,N_18319);
or U18534 (N_18534,N_18033,N_18310);
or U18535 (N_18535,N_18160,N_18079);
xor U18536 (N_18536,N_18357,N_18012);
and U18537 (N_18537,N_18015,N_18031);
xor U18538 (N_18538,N_18096,N_18350);
nor U18539 (N_18539,N_18358,N_18181);
and U18540 (N_18540,N_18002,N_18360);
xnor U18541 (N_18541,N_18398,N_18014);
or U18542 (N_18542,N_18045,N_18253);
nand U18543 (N_18543,N_18085,N_18098);
nor U18544 (N_18544,N_18314,N_18348);
xor U18545 (N_18545,N_18365,N_18020);
and U18546 (N_18546,N_18027,N_18197);
nand U18547 (N_18547,N_18199,N_18282);
nor U18548 (N_18548,N_18032,N_18131);
nand U18549 (N_18549,N_18272,N_18251);
or U18550 (N_18550,N_18183,N_18239);
nand U18551 (N_18551,N_18327,N_18260);
or U18552 (N_18552,N_18237,N_18041);
xor U18553 (N_18553,N_18385,N_18368);
xor U18554 (N_18554,N_18343,N_18158);
or U18555 (N_18555,N_18287,N_18169);
nor U18556 (N_18556,N_18399,N_18397);
nand U18557 (N_18557,N_18281,N_18369);
or U18558 (N_18558,N_18138,N_18026);
nor U18559 (N_18559,N_18349,N_18263);
and U18560 (N_18560,N_18301,N_18157);
xor U18561 (N_18561,N_18269,N_18286);
nand U18562 (N_18562,N_18307,N_18215);
or U18563 (N_18563,N_18198,N_18088);
xnor U18564 (N_18564,N_18191,N_18006);
xnor U18565 (N_18565,N_18250,N_18383);
xor U18566 (N_18566,N_18182,N_18168);
or U18567 (N_18567,N_18206,N_18053);
xor U18568 (N_18568,N_18267,N_18270);
nand U18569 (N_18569,N_18132,N_18099);
or U18570 (N_18570,N_18370,N_18087);
xor U18571 (N_18571,N_18148,N_18075);
xor U18572 (N_18572,N_18159,N_18204);
or U18573 (N_18573,N_18176,N_18106);
xor U18574 (N_18574,N_18255,N_18247);
or U18575 (N_18575,N_18102,N_18188);
or U18576 (N_18576,N_18068,N_18393);
and U18577 (N_18577,N_18025,N_18325);
xor U18578 (N_18578,N_18116,N_18056);
nand U18579 (N_18579,N_18264,N_18230);
nor U18580 (N_18580,N_18137,N_18210);
and U18581 (N_18581,N_18219,N_18143);
or U18582 (N_18582,N_18050,N_18395);
nand U18583 (N_18583,N_18103,N_18299);
or U18584 (N_18584,N_18152,N_18170);
nor U18585 (N_18585,N_18245,N_18378);
and U18586 (N_18586,N_18214,N_18200);
xnor U18587 (N_18587,N_18252,N_18023);
xor U18588 (N_18588,N_18062,N_18046);
nor U18589 (N_18589,N_18136,N_18352);
nor U18590 (N_18590,N_18086,N_18303);
and U18591 (N_18591,N_18359,N_18155);
or U18592 (N_18592,N_18078,N_18122);
xor U18593 (N_18593,N_18125,N_18229);
or U18594 (N_18594,N_18140,N_18000);
nand U18595 (N_18595,N_18194,N_18051);
xnor U18596 (N_18596,N_18227,N_18248);
xnor U18597 (N_18597,N_18233,N_18115);
and U18598 (N_18598,N_18093,N_18165);
nand U18599 (N_18599,N_18241,N_18316);
xnor U18600 (N_18600,N_18199,N_18095);
or U18601 (N_18601,N_18290,N_18164);
nand U18602 (N_18602,N_18303,N_18206);
and U18603 (N_18603,N_18160,N_18131);
xor U18604 (N_18604,N_18265,N_18020);
or U18605 (N_18605,N_18232,N_18131);
nand U18606 (N_18606,N_18373,N_18168);
nand U18607 (N_18607,N_18336,N_18199);
xnor U18608 (N_18608,N_18316,N_18360);
xor U18609 (N_18609,N_18098,N_18385);
xnor U18610 (N_18610,N_18219,N_18191);
nand U18611 (N_18611,N_18119,N_18201);
nand U18612 (N_18612,N_18351,N_18119);
nand U18613 (N_18613,N_18389,N_18281);
nor U18614 (N_18614,N_18199,N_18195);
or U18615 (N_18615,N_18116,N_18203);
or U18616 (N_18616,N_18029,N_18164);
and U18617 (N_18617,N_18222,N_18284);
and U18618 (N_18618,N_18044,N_18066);
xnor U18619 (N_18619,N_18323,N_18009);
or U18620 (N_18620,N_18110,N_18016);
nor U18621 (N_18621,N_18075,N_18102);
nor U18622 (N_18622,N_18232,N_18329);
nand U18623 (N_18623,N_18121,N_18149);
nor U18624 (N_18624,N_18225,N_18166);
nor U18625 (N_18625,N_18078,N_18380);
nand U18626 (N_18626,N_18380,N_18277);
nor U18627 (N_18627,N_18297,N_18016);
nor U18628 (N_18628,N_18207,N_18349);
and U18629 (N_18629,N_18052,N_18304);
xnor U18630 (N_18630,N_18127,N_18028);
or U18631 (N_18631,N_18198,N_18280);
nor U18632 (N_18632,N_18010,N_18330);
or U18633 (N_18633,N_18161,N_18006);
nand U18634 (N_18634,N_18359,N_18334);
nor U18635 (N_18635,N_18335,N_18027);
nor U18636 (N_18636,N_18187,N_18355);
nand U18637 (N_18637,N_18295,N_18237);
or U18638 (N_18638,N_18229,N_18264);
and U18639 (N_18639,N_18025,N_18340);
nor U18640 (N_18640,N_18173,N_18329);
nor U18641 (N_18641,N_18207,N_18274);
nand U18642 (N_18642,N_18330,N_18162);
or U18643 (N_18643,N_18021,N_18090);
nand U18644 (N_18644,N_18041,N_18178);
nor U18645 (N_18645,N_18200,N_18259);
nand U18646 (N_18646,N_18043,N_18233);
nor U18647 (N_18647,N_18288,N_18034);
nor U18648 (N_18648,N_18383,N_18263);
nand U18649 (N_18649,N_18338,N_18353);
or U18650 (N_18650,N_18222,N_18038);
nand U18651 (N_18651,N_18218,N_18127);
and U18652 (N_18652,N_18091,N_18175);
or U18653 (N_18653,N_18206,N_18064);
xnor U18654 (N_18654,N_18304,N_18379);
nand U18655 (N_18655,N_18246,N_18329);
and U18656 (N_18656,N_18308,N_18375);
or U18657 (N_18657,N_18392,N_18243);
nand U18658 (N_18658,N_18066,N_18074);
nand U18659 (N_18659,N_18046,N_18322);
or U18660 (N_18660,N_18116,N_18254);
or U18661 (N_18661,N_18295,N_18327);
or U18662 (N_18662,N_18111,N_18028);
and U18663 (N_18663,N_18279,N_18001);
nor U18664 (N_18664,N_18066,N_18230);
or U18665 (N_18665,N_18348,N_18050);
and U18666 (N_18666,N_18270,N_18038);
nor U18667 (N_18667,N_18005,N_18165);
nor U18668 (N_18668,N_18049,N_18394);
and U18669 (N_18669,N_18145,N_18076);
nor U18670 (N_18670,N_18316,N_18221);
or U18671 (N_18671,N_18338,N_18218);
nor U18672 (N_18672,N_18304,N_18137);
xor U18673 (N_18673,N_18382,N_18047);
nor U18674 (N_18674,N_18397,N_18033);
or U18675 (N_18675,N_18352,N_18128);
and U18676 (N_18676,N_18040,N_18372);
nand U18677 (N_18677,N_18263,N_18079);
nor U18678 (N_18678,N_18253,N_18008);
or U18679 (N_18679,N_18170,N_18181);
nand U18680 (N_18680,N_18060,N_18384);
xnor U18681 (N_18681,N_18242,N_18191);
nand U18682 (N_18682,N_18338,N_18132);
xor U18683 (N_18683,N_18383,N_18249);
nand U18684 (N_18684,N_18336,N_18283);
nand U18685 (N_18685,N_18114,N_18316);
nor U18686 (N_18686,N_18170,N_18325);
nand U18687 (N_18687,N_18107,N_18096);
nor U18688 (N_18688,N_18387,N_18259);
xnor U18689 (N_18689,N_18258,N_18114);
xnor U18690 (N_18690,N_18143,N_18173);
and U18691 (N_18691,N_18393,N_18097);
nor U18692 (N_18692,N_18321,N_18286);
and U18693 (N_18693,N_18348,N_18343);
nor U18694 (N_18694,N_18160,N_18238);
and U18695 (N_18695,N_18230,N_18012);
nand U18696 (N_18696,N_18162,N_18088);
xnor U18697 (N_18697,N_18233,N_18373);
or U18698 (N_18698,N_18202,N_18075);
or U18699 (N_18699,N_18203,N_18038);
or U18700 (N_18700,N_18025,N_18010);
or U18701 (N_18701,N_18152,N_18203);
nand U18702 (N_18702,N_18319,N_18326);
nor U18703 (N_18703,N_18309,N_18296);
or U18704 (N_18704,N_18132,N_18275);
nor U18705 (N_18705,N_18209,N_18019);
nor U18706 (N_18706,N_18212,N_18124);
nand U18707 (N_18707,N_18122,N_18376);
nor U18708 (N_18708,N_18147,N_18250);
or U18709 (N_18709,N_18067,N_18028);
nand U18710 (N_18710,N_18160,N_18219);
xnor U18711 (N_18711,N_18281,N_18342);
nand U18712 (N_18712,N_18383,N_18092);
nand U18713 (N_18713,N_18293,N_18022);
or U18714 (N_18714,N_18195,N_18097);
or U18715 (N_18715,N_18162,N_18046);
nor U18716 (N_18716,N_18371,N_18192);
or U18717 (N_18717,N_18014,N_18315);
nand U18718 (N_18718,N_18170,N_18368);
xor U18719 (N_18719,N_18130,N_18376);
nand U18720 (N_18720,N_18164,N_18265);
nand U18721 (N_18721,N_18145,N_18017);
and U18722 (N_18722,N_18013,N_18255);
and U18723 (N_18723,N_18107,N_18284);
and U18724 (N_18724,N_18199,N_18342);
xor U18725 (N_18725,N_18215,N_18333);
and U18726 (N_18726,N_18284,N_18088);
nand U18727 (N_18727,N_18319,N_18163);
and U18728 (N_18728,N_18092,N_18318);
or U18729 (N_18729,N_18123,N_18253);
nand U18730 (N_18730,N_18304,N_18247);
or U18731 (N_18731,N_18270,N_18368);
and U18732 (N_18732,N_18275,N_18326);
nor U18733 (N_18733,N_18096,N_18170);
and U18734 (N_18734,N_18139,N_18267);
nor U18735 (N_18735,N_18351,N_18079);
nor U18736 (N_18736,N_18224,N_18379);
nand U18737 (N_18737,N_18270,N_18282);
nor U18738 (N_18738,N_18204,N_18016);
nand U18739 (N_18739,N_18146,N_18045);
nor U18740 (N_18740,N_18029,N_18030);
nor U18741 (N_18741,N_18113,N_18143);
nor U18742 (N_18742,N_18339,N_18260);
nand U18743 (N_18743,N_18190,N_18318);
xnor U18744 (N_18744,N_18275,N_18271);
nand U18745 (N_18745,N_18042,N_18274);
nand U18746 (N_18746,N_18310,N_18003);
nand U18747 (N_18747,N_18276,N_18090);
nor U18748 (N_18748,N_18097,N_18061);
or U18749 (N_18749,N_18351,N_18176);
and U18750 (N_18750,N_18085,N_18009);
nand U18751 (N_18751,N_18115,N_18337);
nand U18752 (N_18752,N_18082,N_18179);
nor U18753 (N_18753,N_18299,N_18238);
xor U18754 (N_18754,N_18130,N_18199);
xnor U18755 (N_18755,N_18260,N_18301);
and U18756 (N_18756,N_18393,N_18049);
xor U18757 (N_18757,N_18308,N_18390);
nand U18758 (N_18758,N_18144,N_18170);
nand U18759 (N_18759,N_18320,N_18273);
nand U18760 (N_18760,N_18184,N_18253);
and U18761 (N_18761,N_18154,N_18327);
and U18762 (N_18762,N_18364,N_18021);
xor U18763 (N_18763,N_18055,N_18207);
nand U18764 (N_18764,N_18379,N_18199);
xnor U18765 (N_18765,N_18386,N_18275);
and U18766 (N_18766,N_18326,N_18044);
nand U18767 (N_18767,N_18278,N_18335);
or U18768 (N_18768,N_18143,N_18333);
and U18769 (N_18769,N_18164,N_18210);
or U18770 (N_18770,N_18054,N_18262);
or U18771 (N_18771,N_18039,N_18008);
xor U18772 (N_18772,N_18194,N_18142);
nand U18773 (N_18773,N_18058,N_18367);
nor U18774 (N_18774,N_18033,N_18368);
xor U18775 (N_18775,N_18244,N_18275);
or U18776 (N_18776,N_18283,N_18271);
or U18777 (N_18777,N_18013,N_18308);
and U18778 (N_18778,N_18192,N_18284);
nand U18779 (N_18779,N_18126,N_18108);
xor U18780 (N_18780,N_18295,N_18040);
xnor U18781 (N_18781,N_18336,N_18208);
nor U18782 (N_18782,N_18318,N_18000);
and U18783 (N_18783,N_18177,N_18347);
xnor U18784 (N_18784,N_18087,N_18081);
and U18785 (N_18785,N_18166,N_18272);
or U18786 (N_18786,N_18049,N_18052);
nand U18787 (N_18787,N_18019,N_18260);
or U18788 (N_18788,N_18275,N_18323);
nor U18789 (N_18789,N_18001,N_18064);
and U18790 (N_18790,N_18379,N_18129);
nor U18791 (N_18791,N_18383,N_18054);
nor U18792 (N_18792,N_18105,N_18244);
and U18793 (N_18793,N_18291,N_18113);
or U18794 (N_18794,N_18290,N_18099);
nor U18795 (N_18795,N_18251,N_18207);
nand U18796 (N_18796,N_18277,N_18140);
nor U18797 (N_18797,N_18113,N_18135);
xnor U18798 (N_18798,N_18283,N_18326);
nand U18799 (N_18799,N_18077,N_18255);
nor U18800 (N_18800,N_18782,N_18640);
xnor U18801 (N_18801,N_18409,N_18772);
and U18802 (N_18802,N_18797,N_18606);
xor U18803 (N_18803,N_18495,N_18438);
nor U18804 (N_18804,N_18710,N_18751);
nand U18805 (N_18805,N_18449,N_18633);
or U18806 (N_18806,N_18530,N_18542);
or U18807 (N_18807,N_18484,N_18647);
and U18808 (N_18808,N_18416,N_18568);
xor U18809 (N_18809,N_18659,N_18716);
nor U18810 (N_18810,N_18417,N_18497);
or U18811 (N_18811,N_18569,N_18550);
nor U18812 (N_18812,N_18776,N_18470);
xor U18813 (N_18813,N_18713,N_18591);
or U18814 (N_18814,N_18551,N_18791);
and U18815 (N_18815,N_18717,N_18467);
and U18816 (N_18816,N_18586,N_18627);
and U18817 (N_18817,N_18456,N_18486);
or U18818 (N_18818,N_18441,N_18476);
or U18819 (N_18819,N_18735,N_18726);
nor U18820 (N_18820,N_18614,N_18738);
and U18821 (N_18821,N_18460,N_18549);
or U18822 (N_18822,N_18660,N_18469);
nor U18823 (N_18823,N_18752,N_18464);
nand U18824 (N_18824,N_18674,N_18458);
nor U18825 (N_18825,N_18434,N_18618);
and U18826 (N_18826,N_18418,N_18679);
nand U18827 (N_18827,N_18421,N_18553);
or U18828 (N_18828,N_18462,N_18795);
nand U18829 (N_18829,N_18755,N_18663);
nand U18830 (N_18830,N_18767,N_18559);
and U18831 (N_18831,N_18668,N_18637);
and U18832 (N_18832,N_18787,N_18743);
nand U18833 (N_18833,N_18638,N_18571);
nor U18834 (N_18834,N_18683,N_18731);
nand U18835 (N_18835,N_18623,N_18646);
xnor U18836 (N_18836,N_18565,N_18561);
or U18837 (N_18837,N_18471,N_18667);
nand U18838 (N_18838,N_18781,N_18715);
nor U18839 (N_18839,N_18711,N_18415);
nand U18840 (N_18840,N_18773,N_18461);
nor U18841 (N_18841,N_18406,N_18630);
nand U18842 (N_18842,N_18475,N_18436);
xor U18843 (N_18843,N_18770,N_18563);
nor U18844 (N_18844,N_18651,N_18560);
nor U18845 (N_18845,N_18574,N_18611);
nand U18846 (N_18846,N_18478,N_18511);
or U18847 (N_18847,N_18708,N_18496);
nand U18848 (N_18848,N_18639,N_18404);
and U18849 (N_18849,N_18665,N_18485);
and U18850 (N_18850,N_18468,N_18420);
nand U18851 (N_18851,N_18675,N_18526);
nand U18852 (N_18852,N_18603,N_18727);
nand U18853 (N_18853,N_18671,N_18691);
or U18854 (N_18854,N_18629,N_18473);
nor U18855 (N_18855,N_18670,N_18457);
and U18856 (N_18856,N_18589,N_18535);
and U18857 (N_18857,N_18539,N_18402);
xnor U18858 (N_18858,N_18707,N_18554);
nand U18859 (N_18859,N_18548,N_18523);
nand U18860 (N_18860,N_18613,N_18537);
xor U18861 (N_18861,N_18666,N_18519);
or U18862 (N_18862,N_18578,N_18493);
xor U18863 (N_18863,N_18642,N_18512);
nor U18864 (N_18864,N_18628,N_18562);
nor U18865 (N_18865,N_18545,N_18435);
and U18866 (N_18866,N_18426,N_18446);
and U18867 (N_18867,N_18728,N_18693);
and U18868 (N_18868,N_18520,N_18699);
nand U18869 (N_18869,N_18598,N_18531);
nor U18870 (N_18870,N_18766,N_18483);
xnor U18871 (N_18871,N_18798,N_18769);
nor U18872 (N_18872,N_18465,N_18445);
nor U18873 (N_18873,N_18590,N_18427);
nand U18874 (N_18874,N_18479,N_18734);
nand U18875 (N_18875,N_18701,N_18600);
and U18876 (N_18876,N_18570,N_18662);
and U18877 (N_18877,N_18780,N_18422);
and U18878 (N_18878,N_18431,N_18487);
xor U18879 (N_18879,N_18747,N_18596);
nand U18880 (N_18880,N_18527,N_18423);
nand U18881 (N_18881,N_18739,N_18786);
or U18882 (N_18882,N_18583,N_18430);
or U18883 (N_18883,N_18736,N_18758);
nand U18884 (N_18884,N_18609,N_18690);
nor U18885 (N_18885,N_18759,N_18622);
nand U18886 (N_18886,N_18792,N_18405);
and U18887 (N_18887,N_18518,N_18489);
and U18888 (N_18888,N_18654,N_18411);
nand U18889 (N_18889,N_18625,N_18543);
and U18890 (N_18890,N_18607,N_18472);
nor U18891 (N_18891,N_18677,N_18525);
nand U18892 (N_18892,N_18580,N_18601);
or U18893 (N_18893,N_18706,N_18702);
and U18894 (N_18894,N_18746,N_18587);
nand U18895 (N_18895,N_18432,N_18740);
and U18896 (N_18896,N_18621,N_18724);
or U18897 (N_18897,N_18558,N_18745);
or U18898 (N_18898,N_18788,N_18692);
or U18899 (N_18899,N_18612,N_18721);
nand U18900 (N_18900,N_18761,N_18703);
or U18901 (N_18901,N_18730,N_18547);
xor U18902 (N_18902,N_18641,N_18424);
or U18903 (N_18903,N_18556,N_18529);
nor U18904 (N_18904,N_18648,N_18695);
and U18905 (N_18905,N_18491,N_18437);
or U18906 (N_18906,N_18459,N_18451);
and U18907 (N_18907,N_18794,N_18452);
nand U18908 (N_18908,N_18722,N_18765);
nor U18909 (N_18909,N_18644,N_18729);
nor U18910 (N_18910,N_18610,N_18506);
nor U18911 (N_18911,N_18669,N_18604);
nor U18912 (N_18912,N_18777,N_18725);
nor U18913 (N_18913,N_18676,N_18748);
or U18914 (N_18914,N_18709,N_18419);
and U18915 (N_18915,N_18785,N_18634);
nand U18916 (N_18916,N_18649,N_18588);
or U18917 (N_18917,N_18661,N_18594);
or U18918 (N_18918,N_18686,N_18510);
or U18919 (N_18919,N_18582,N_18741);
nand U18920 (N_18920,N_18577,N_18635);
nand U18921 (N_18921,N_18689,N_18680);
and U18922 (N_18922,N_18768,N_18515);
or U18923 (N_18923,N_18775,N_18517);
xor U18924 (N_18924,N_18499,N_18608);
nor U18925 (N_18925,N_18442,N_18756);
nor U18926 (N_18926,N_18737,N_18657);
xnor U18927 (N_18927,N_18753,N_18439);
and U18928 (N_18928,N_18750,N_18521);
nor U18929 (N_18929,N_18448,N_18454);
nor U18930 (N_18930,N_18744,N_18494);
and U18931 (N_18931,N_18507,N_18605);
and U18932 (N_18932,N_18593,N_18575);
nand U18933 (N_18933,N_18488,N_18455);
or U18934 (N_18934,N_18643,N_18616);
or U18935 (N_18935,N_18567,N_18617);
nor U18936 (N_18936,N_18732,N_18664);
xor U18937 (N_18937,N_18723,N_18754);
or U18938 (N_18938,N_18500,N_18650);
nand U18939 (N_18939,N_18763,N_18536);
nor U18940 (N_18940,N_18619,N_18490);
nand U18941 (N_18941,N_18790,N_18760);
nand U18942 (N_18942,N_18685,N_18698);
or U18943 (N_18943,N_18672,N_18764);
or U18944 (N_18944,N_18762,N_18514);
nor U18945 (N_18945,N_18408,N_18688);
and U18946 (N_18946,N_18656,N_18771);
xor U18947 (N_18947,N_18429,N_18503);
xnor U18948 (N_18948,N_18516,N_18433);
nand U18949 (N_18949,N_18564,N_18626);
or U18950 (N_18950,N_18742,N_18620);
or U18951 (N_18951,N_18783,N_18774);
and U18952 (N_18952,N_18733,N_18504);
nor U18953 (N_18953,N_18632,N_18793);
and U18954 (N_18954,N_18538,N_18541);
nor U18955 (N_18955,N_18573,N_18480);
or U18956 (N_18956,N_18533,N_18796);
xnor U18957 (N_18957,N_18576,N_18555);
and U18958 (N_18958,N_18700,N_18789);
xnor U18959 (N_18959,N_18509,N_18624);
nor U18960 (N_18960,N_18524,N_18528);
nand U18961 (N_18961,N_18697,N_18522);
nand U18962 (N_18962,N_18599,N_18655);
and U18963 (N_18963,N_18428,N_18652);
and U18964 (N_18964,N_18502,N_18532);
xor U18965 (N_18965,N_18681,N_18714);
and U18966 (N_18966,N_18410,N_18401);
nand U18967 (N_18967,N_18645,N_18585);
xnor U18968 (N_18968,N_18602,N_18505);
and U18969 (N_18969,N_18407,N_18720);
xnor U18970 (N_18970,N_18719,N_18498);
nor U18971 (N_18971,N_18678,N_18540);
nor U18972 (N_18972,N_18400,N_18466);
or U18973 (N_18973,N_18544,N_18682);
nor U18974 (N_18974,N_18463,N_18492);
nand U18975 (N_18975,N_18566,N_18481);
nor U18976 (N_18976,N_18778,N_18414);
or U18977 (N_18977,N_18597,N_18653);
nand U18978 (N_18978,N_18615,N_18513);
nor U18979 (N_18979,N_18687,N_18508);
nor U18980 (N_18980,N_18453,N_18658);
or U18981 (N_18981,N_18474,N_18696);
nor U18982 (N_18982,N_18705,N_18477);
nor U18983 (N_18983,N_18403,N_18447);
nand U18984 (N_18984,N_18712,N_18694);
or U18985 (N_18985,N_18581,N_18572);
xor U18986 (N_18986,N_18718,N_18546);
nor U18987 (N_18987,N_18749,N_18631);
and U18988 (N_18988,N_18450,N_18482);
xor U18989 (N_18989,N_18584,N_18444);
or U18990 (N_18990,N_18443,N_18579);
and U18991 (N_18991,N_18757,N_18704);
and U18992 (N_18992,N_18412,N_18779);
nor U18993 (N_18993,N_18636,N_18595);
nor U18994 (N_18994,N_18799,N_18592);
nor U18995 (N_18995,N_18552,N_18534);
nor U18996 (N_18996,N_18425,N_18673);
or U18997 (N_18997,N_18413,N_18501);
and U18998 (N_18998,N_18557,N_18784);
or U18999 (N_18999,N_18440,N_18684);
xor U19000 (N_19000,N_18764,N_18574);
nor U19001 (N_19001,N_18772,N_18663);
xnor U19002 (N_19002,N_18535,N_18616);
and U19003 (N_19003,N_18778,N_18483);
or U19004 (N_19004,N_18586,N_18667);
and U19005 (N_19005,N_18531,N_18418);
nor U19006 (N_19006,N_18448,N_18547);
nor U19007 (N_19007,N_18416,N_18516);
nor U19008 (N_19008,N_18517,N_18562);
nand U19009 (N_19009,N_18450,N_18578);
nand U19010 (N_19010,N_18697,N_18409);
xnor U19011 (N_19011,N_18601,N_18796);
and U19012 (N_19012,N_18633,N_18713);
nor U19013 (N_19013,N_18705,N_18431);
and U19014 (N_19014,N_18697,N_18776);
xnor U19015 (N_19015,N_18735,N_18699);
or U19016 (N_19016,N_18640,N_18621);
xnor U19017 (N_19017,N_18636,N_18488);
and U19018 (N_19018,N_18464,N_18519);
or U19019 (N_19019,N_18524,N_18507);
nand U19020 (N_19020,N_18460,N_18615);
and U19021 (N_19021,N_18506,N_18714);
or U19022 (N_19022,N_18537,N_18764);
xor U19023 (N_19023,N_18410,N_18521);
and U19024 (N_19024,N_18735,N_18640);
or U19025 (N_19025,N_18524,N_18541);
xor U19026 (N_19026,N_18562,N_18643);
and U19027 (N_19027,N_18712,N_18613);
nand U19028 (N_19028,N_18663,N_18594);
or U19029 (N_19029,N_18575,N_18604);
and U19030 (N_19030,N_18405,N_18799);
or U19031 (N_19031,N_18630,N_18544);
nor U19032 (N_19032,N_18401,N_18670);
nand U19033 (N_19033,N_18697,N_18690);
xor U19034 (N_19034,N_18425,N_18648);
nand U19035 (N_19035,N_18691,N_18796);
or U19036 (N_19036,N_18544,N_18416);
and U19037 (N_19037,N_18479,N_18760);
nor U19038 (N_19038,N_18664,N_18484);
xnor U19039 (N_19039,N_18488,N_18669);
nand U19040 (N_19040,N_18758,N_18742);
nor U19041 (N_19041,N_18760,N_18746);
or U19042 (N_19042,N_18795,N_18775);
nor U19043 (N_19043,N_18578,N_18429);
or U19044 (N_19044,N_18432,N_18486);
or U19045 (N_19045,N_18765,N_18644);
xor U19046 (N_19046,N_18484,N_18402);
nor U19047 (N_19047,N_18601,N_18628);
nor U19048 (N_19048,N_18570,N_18459);
xnor U19049 (N_19049,N_18670,N_18435);
and U19050 (N_19050,N_18560,N_18448);
or U19051 (N_19051,N_18448,N_18646);
or U19052 (N_19052,N_18439,N_18482);
nand U19053 (N_19053,N_18715,N_18466);
nor U19054 (N_19054,N_18489,N_18521);
nand U19055 (N_19055,N_18708,N_18719);
or U19056 (N_19056,N_18645,N_18728);
xnor U19057 (N_19057,N_18722,N_18754);
xnor U19058 (N_19058,N_18742,N_18725);
xor U19059 (N_19059,N_18625,N_18434);
and U19060 (N_19060,N_18465,N_18486);
xnor U19061 (N_19061,N_18561,N_18637);
and U19062 (N_19062,N_18520,N_18603);
nor U19063 (N_19063,N_18573,N_18592);
nand U19064 (N_19064,N_18442,N_18609);
and U19065 (N_19065,N_18503,N_18414);
and U19066 (N_19066,N_18644,N_18476);
nand U19067 (N_19067,N_18791,N_18665);
and U19068 (N_19068,N_18531,N_18495);
and U19069 (N_19069,N_18771,N_18674);
nor U19070 (N_19070,N_18663,N_18415);
nand U19071 (N_19071,N_18649,N_18415);
or U19072 (N_19072,N_18682,N_18626);
or U19073 (N_19073,N_18489,N_18581);
nor U19074 (N_19074,N_18501,N_18647);
and U19075 (N_19075,N_18424,N_18523);
and U19076 (N_19076,N_18741,N_18725);
xor U19077 (N_19077,N_18500,N_18421);
nor U19078 (N_19078,N_18574,N_18588);
nor U19079 (N_19079,N_18579,N_18504);
or U19080 (N_19080,N_18496,N_18539);
or U19081 (N_19081,N_18466,N_18497);
and U19082 (N_19082,N_18561,N_18479);
nor U19083 (N_19083,N_18543,N_18424);
or U19084 (N_19084,N_18697,N_18749);
nor U19085 (N_19085,N_18708,N_18795);
xnor U19086 (N_19086,N_18724,N_18442);
or U19087 (N_19087,N_18536,N_18681);
nor U19088 (N_19088,N_18783,N_18426);
nand U19089 (N_19089,N_18428,N_18633);
or U19090 (N_19090,N_18787,N_18785);
or U19091 (N_19091,N_18642,N_18754);
xor U19092 (N_19092,N_18592,N_18624);
nand U19093 (N_19093,N_18506,N_18661);
or U19094 (N_19094,N_18469,N_18563);
or U19095 (N_19095,N_18755,N_18506);
nand U19096 (N_19096,N_18577,N_18451);
and U19097 (N_19097,N_18456,N_18492);
and U19098 (N_19098,N_18759,N_18793);
xnor U19099 (N_19099,N_18507,N_18513);
xor U19100 (N_19100,N_18626,N_18402);
nand U19101 (N_19101,N_18765,N_18534);
xor U19102 (N_19102,N_18574,N_18511);
xnor U19103 (N_19103,N_18578,N_18669);
nor U19104 (N_19104,N_18609,N_18573);
xnor U19105 (N_19105,N_18425,N_18619);
nand U19106 (N_19106,N_18487,N_18586);
or U19107 (N_19107,N_18673,N_18582);
xnor U19108 (N_19108,N_18456,N_18751);
xnor U19109 (N_19109,N_18429,N_18550);
xor U19110 (N_19110,N_18450,N_18609);
xnor U19111 (N_19111,N_18434,N_18777);
nand U19112 (N_19112,N_18721,N_18744);
or U19113 (N_19113,N_18419,N_18781);
and U19114 (N_19114,N_18725,N_18454);
xor U19115 (N_19115,N_18584,N_18586);
and U19116 (N_19116,N_18439,N_18563);
and U19117 (N_19117,N_18674,N_18779);
and U19118 (N_19118,N_18754,N_18591);
xor U19119 (N_19119,N_18788,N_18511);
and U19120 (N_19120,N_18718,N_18659);
nor U19121 (N_19121,N_18772,N_18732);
and U19122 (N_19122,N_18602,N_18501);
xor U19123 (N_19123,N_18667,N_18598);
nor U19124 (N_19124,N_18463,N_18588);
or U19125 (N_19125,N_18688,N_18571);
xor U19126 (N_19126,N_18522,N_18477);
nand U19127 (N_19127,N_18591,N_18441);
xnor U19128 (N_19128,N_18471,N_18586);
and U19129 (N_19129,N_18702,N_18695);
xor U19130 (N_19130,N_18422,N_18554);
nor U19131 (N_19131,N_18458,N_18429);
or U19132 (N_19132,N_18631,N_18684);
and U19133 (N_19133,N_18777,N_18511);
xnor U19134 (N_19134,N_18582,N_18546);
xnor U19135 (N_19135,N_18728,N_18643);
nor U19136 (N_19136,N_18577,N_18665);
nor U19137 (N_19137,N_18436,N_18776);
nand U19138 (N_19138,N_18718,N_18446);
and U19139 (N_19139,N_18456,N_18440);
or U19140 (N_19140,N_18554,N_18428);
xor U19141 (N_19141,N_18557,N_18472);
nand U19142 (N_19142,N_18626,N_18405);
nand U19143 (N_19143,N_18738,N_18776);
nor U19144 (N_19144,N_18643,N_18766);
nor U19145 (N_19145,N_18414,N_18413);
nor U19146 (N_19146,N_18659,N_18433);
xor U19147 (N_19147,N_18515,N_18576);
or U19148 (N_19148,N_18487,N_18442);
nand U19149 (N_19149,N_18633,N_18580);
xor U19150 (N_19150,N_18533,N_18542);
or U19151 (N_19151,N_18789,N_18525);
xnor U19152 (N_19152,N_18617,N_18716);
nand U19153 (N_19153,N_18514,N_18434);
or U19154 (N_19154,N_18797,N_18508);
and U19155 (N_19155,N_18744,N_18552);
and U19156 (N_19156,N_18774,N_18765);
nor U19157 (N_19157,N_18785,N_18541);
nor U19158 (N_19158,N_18485,N_18656);
and U19159 (N_19159,N_18603,N_18661);
and U19160 (N_19160,N_18571,N_18593);
and U19161 (N_19161,N_18758,N_18434);
nor U19162 (N_19162,N_18504,N_18609);
or U19163 (N_19163,N_18666,N_18537);
and U19164 (N_19164,N_18475,N_18671);
nand U19165 (N_19165,N_18543,N_18470);
nand U19166 (N_19166,N_18726,N_18641);
nor U19167 (N_19167,N_18586,N_18553);
or U19168 (N_19168,N_18404,N_18553);
and U19169 (N_19169,N_18560,N_18550);
nand U19170 (N_19170,N_18782,N_18409);
nor U19171 (N_19171,N_18463,N_18659);
nor U19172 (N_19172,N_18679,N_18441);
or U19173 (N_19173,N_18556,N_18763);
or U19174 (N_19174,N_18691,N_18424);
and U19175 (N_19175,N_18678,N_18599);
nand U19176 (N_19176,N_18429,N_18541);
xor U19177 (N_19177,N_18558,N_18499);
or U19178 (N_19178,N_18570,N_18522);
and U19179 (N_19179,N_18731,N_18621);
nor U19180 (N_19180,N_18576,N_18605);
xor U19181 (N_19181,N_18527,N_18577);
and U19182 (N_19182,N_18787,N_18469);
or U19183 (N_19183,N_18457,N_18728);
nand U19184 (N_19184,N_18424,N_18709);
and U19185 (N_19185,N_18484,N_18643);
or U19186 (N_19186,N_18401,N_18488);
nand U19187 (N_19187,N_18606,N_18522);
or U19188 (N_19188,N_18690,N_18468);
nand U19189 (N_19189,N_18602,N_18570);
nor U19190 (N_19190,N_18450,N_18672);
and U19191 (N_19191,N_18795,N_18420);
nand U19192 (N_19192,N_18519,N_18592);
nand U19193 (N_19193,N_18658,N_18577);
and U19194 (N_19194,N_18646,N_18727);
and U19195 (N_19195,N_18686,N_18731);
xor U19196 (N_19196,N_18428,N_18471);
xor U19197 (N_19197,N_18572,N_18686);
and U19198 (N_19198,N_18677,N_18614);
xnor U19199 (N_19199,N_18764,N_18549);
nor U19200 (N_19200,N_19109,N_18913);
xor U19201 (N_19201,N_18852,N_19049);
xor U19202 (N_19202,N_19141,N_19008);
nand U19203 (N_19203,N_18972,N_19099);
or U19204 (N_19204,N_19195,N_19169);
nand U19205 (N_19205,N_19120,N_18901);
and U19206 (N_19206,N_18824,N_19007);
or U19207 (N_19207,N_19020,N_19065);
and U19208 (N_19208,N_19115,N_19085);
and U19209 (N_19209,N_19146,N_18989);
nor U19210 (N_19210,N_18930,N_18874);
xor U19211 (N_19211,N_19196,N_19100);
nand U19212 (N_19212,N_19063,N_18821);
or U19213 (N_19213,N_18830,N_18802);
or U19214 (N_19214,N_18812,N_19143);
nand U19215 (N_19215,N_19199,N_18856);
or U19216 (N_19216,N_18940,N_19108);
or U19217 (N_19217,N_19009,N_19047);
and U19218 (N_19218,N_18900,N_18911);
and U19219 (N_19219,N_19044,N_19095);
or U19220 (N_19220,N_18937,N_18988);
xnor U19221 (N_19221,N_18890,N_19075);
nand U19222 (N_19222,N_19061,N_18967);
and U19223 (N_19223,N_19062,N_18983);
nor U19224 (N_19224,N_19104,N_18892);
nand U19225 (N_19225,N_19129,N_19121);
and U19226 (N_19226,N_18834,N_19154);
xnor U19227 (N_19227,N_19032,N_18800);
nand U19228 (N_19228,N_19091,N_18957);
and U19229 (N_19229,N_18837,N_18979);
and U19230 (N_19230,N_19170,N_18903);
nor U19231 (N_19231,N_18853,N_19168);
nor U19232 (N_19232,N_18994,N_19135);
xnor U19233 (N_19233,N_18814,N_18843);
nor U19234 (N_19234,N_18970,N_18859);
nand U19235 (N_19235,N_19015,N_19092);
or U19236 (N_19236,N_18858,N_19084);
or U19237 (N_19237,N_18872,N_18904);
or U19238 (N_19238,N_18891,N_19145);
nand U19239 (N_19239,N_18813,N_19161);
nor U19240 (N_19240,N_19174,N_18823);
nand U19241 (N_19241,N_18923,N_18946);
nand U19242 (N_19242,N_18985,N_19024);
and U19243 (N_19243,N_19040,N_18982);
nor U19244 (N_19244,N_18819,N_18966);
and U19245 (N_19245,N_19149,N_19182);
nor U19246 (N_19246,N_19112,N_19031);
nand U19247 (N_19247,N_18999,N_18849);
nand U19248 (N_19248,N_18841,N_19124);
nand U19249 (N_19249,N_18854,N_19012);
nand U19250 (N_19250,N_18918,N_18862);
and U19251 (N_19251,N_19119,N_18878);
or U19252 (N_19252,N_18959,N_18861);
and U19253 (N_19253,N_18873,N_19076);
nand U19254 (N_19254,N_18955,N_18984);
or U19255 (N_19255,N_18997,N_19153);
nor U19256 (N_19256,N_18816,N_18950);
or U19257 (N_19257,N_18990,N_19177);
nor U19258 (N_19258,N_18805,N_19029);
and U19259 (N_19259,N_19017,N_19064);
nor U19260 (N_19260,N_19056,N_18956);
xnor U19261 (N_19261,N_19002,N_18939);
xnor U19262 (N_19262,N_18870,N_18839);
and U19263 (N_19263,N_19074,N_18825);
or U19264 (N_19264,N_18905,N_18807);
and U19265 (N_19265,N_18871,N_18860);
nand U19266 (N_19266,N_19046,N_19133);
nand U19267 (N_19267,N_19068,N_18920);
or U19268 (N_19268,N_18826,N_19082);
xnor U19269 (N_19269,N_19172,N_18818);
nand U19270 (N_19270,N_18943,N_19137);
or U19271 (N_19271,N_18949,N_19050);
nor U19272 (N_19272,N_18995,N_18914);
nand U19273 (N_19273,N_19114,N_19001);
nor U19274 (N_19274,N_18842,N_18962);
nand U19275 (N_19275,N_18875,N_19126);
nor U19276 (N_19276,N_18969,N_18971);
xor U19277 (N_19277,N_18811,N_18836);
or U19278 (N_19278,N_19081,N_19151);
nand U19279 (N_19279,N_19144,N_18936);
nand U19280 (N_19280,N_19045,N_19198);
nand U19281 (N_19281,N_18980,N_18898);
nor U19282 (N_19282,N_18881,N_18879);
or U19283 (N_19283,N_18965,N_18976);
or U19284 (N_19284,N_18864,N_18916);
nor U19285 (N_19285,N_18835,N_19043);
nor U19286 (N_19286,N_19034,N_18922);
and U19287 (N_19287,N_18876,N_18869);
nor U19288 (N_19288,N_19014,N_19163);
nand U19289 (N_19289,N_18838,N_18895);
xnor U19290 (N_19290,N_19021,N_19123);
nand U19291 (N_19291,N_18897,N_18929);
and U19292 (N_19292,N_19103,N_19194);
xnor U19293 (N_19293,N_18927,N_19131);
nand U19294 (N_19294,N_19110,N_18865);
xnor U19295 (N_19295,N_19058,N_18817);
xnor U19296 (N_19296,N_18938,N_19080);
nor U19297 (N_19297,N_18902,N_18993);
nor U19298 (N_19298,N_19057,N_19132);
nor U19299 (N_19299,N_19054,N_18910);
and U19300 (N_19300,N_18880,N_18991);
xor U19301 (N_19301,N_19113,N_18915);
nor U19302 (N_19302,N_19083,N_18931);
xnor U19303 (N_19303,N_18844,N_19093);
or U19304 (N_19304,N_18953,N_18951);
nor U19305 (N_19305,N_19060,N_18935);
xnor U19306 (N_19306,N_19184,N_19088);
nor U19307 (N_19307,N_19019,N_19025);
or U19308 (N_19308,N_18942,N_18963);
and U19309 (N_19309,N_18925,N_19142);
nand U19310 (N_19310,N_19000,N_19152);
nor U19311 (N_19311,N_19087,N_19086);
nor U19312 (N_19312,N_19011,N_19193);
or U19313 (N_19313,N_18899,N_19090);
nor U19314 (N_19314,N_18909,N_19185);
nor U19315 (N_19315,N_19097,N_18921);
or U19316 (N_19316,N_18986,N_19010);
nand U19317 (N_19317,N_19166,N_19181);
nor U19318 (N_19318,N_19134,N_18867);
and U19319 (N_19319,N_19173,N_18992);
nor U19320 (N_19320,N_18884,N_18893);
nor U19321 (N_19321,N_18882,N_18919);
and U19322 (N_19322,N_18809,N_18964);
or U19323 (N_19323,N_18952,N_18987);
nand U19324 (N_19324,N_19036,N_18894);
and U19325 (N_19325,N_18954,N_19077);
nor U19326 (N_19326,N_19018,N_18977);
and U19327 (N_19327,N_18847,N_19162);
nand U19328 (N_19328,N_19171,N_19038);
nor U19329 (N_19329,N_19187,N_19128);
or U19330 (N_19330,N_18887,N_18855);
or U19331 (N_19331,N_19102,N_18815);
nor U19332 (N_19332,N_19186,N_19160);
nand U19333 (N_19333,N_19101,N_19138);
nand U19334 (N_19334,N_18832,N_18801);
and U19335 (N_19335,N_19042,N_19176);
xnor U19336 (N_19336,N_19127,N_19055);
nand U19337 (N_19337,N_19107,N_19122);
nand U19338 (N_19338,N_18803,N_18808);
nor U19339 (N_19339,N_18851,N_19188);
nor U19340 (N_19340,N_18889,N_18885);
nand U19341 (N_19341,N_18883,N_18917);
and U19342 (N_19342,N_18968,N_19130);
and U19343 (N_19343,N_19179,N_18960);
and U19344 (N_19344,N_18924,N_19004);
xnor U19345 (N_19345,N_19136,N_18948);
or U19346 (N_19346,N_19183,N_18840);
and U19347 (N_19347,N_19013,N_19165);
nand U19348 (N_19348,N_19139,N_19106);
nand U19349 (N_19349,N_18822,N_19158);
or U19350 (N_19350,N_19030,N_18866);
or U19351 (N_19351,N_19117,N_18848);
and U19352 (N_19352,N_19052,N_19189);
nor U19353 (N_19353,N_18941,N_18981);
or U19354 (N_19354,N_19059,N_19037);
nand U19355 (N_19355,N_19005,N_18806);
nand U19356 (N_19356,N_18998,N_18896);
xor U19357 (N_19357,N_19167,N_19022);
and U19358 (N_19358,N_19006,N_19028);
nor U19359 (N_19359,N_19067,N_19071);
and U19360 (N_19360,N_19072,N_18833);
or U19361 (N_19361,N_19159,N_19147);
nor U19362 (N_19362,N_19180,N_18804);
nor U19363 (N_19363,N_18926,N_18828);
nor U19364 (N_19364,N_19164,N_18868);
xor U19365 (N_19365,N_19035,N_19041);
and U19366 (N_19366,N_18850,N_19192);
nand U19367 (N_19367,N_19197,N_18908);
nand U19368 (N_19368,N_19078,N_18810);
and U19369 (N_19369,N_19033,N_18996);
nand U19370 (N_19370,N_18888,N_18827);
and U19371 (N_19371,N_19089,N_18932);
xnor U19372 (N_19372,N_18857,N_18978);
or U19373 (N_19373,N_18886,N_18928);
xnor U19374 (N_19374,N_18947,N_19026);
xnor U19375 (N_19375,N_18820,N_19155);
xor U19376 (N_19376,N_18944,N_19094);
nor U19377 (N_19377,N_19157,N_18974);
nand U19378 (N_19378,N_19178,N_19070);
nor U19379 (N_19379,N_18877,N_19053);
nand U19380 (N_19380,N_19023,N_19073);
nor U19381 (N_19381,N_19140,N_19016);
nor U19382 (N_19382,N_19098,N_18907);
and U19383 (N_19383,N_19003,N_18906);
nor U19384 (N_19384,N_18945,N_19190);
nand U19385 (N_19385,N_19156,N_19105);
nand U19386 (N_19386,N_18961,N_18845);
xnor U19387 (N_19387,N_19175,N_18933);
nand U19388 (N_19388,N_19048,N_19069);
xnor U19389 (N_19389,N_19027,N_18831);
nor U19390 (N_19390,N_19066,N_19079);
nor U19391 (N_19391,N_19096,N_18846);
nand U19392 (N_19392,N_18973,N_19150);
xor U19393 (N_19393,N_19148,N_18975);
or U19394 (N_19394,N_19051,N_19125);
or U19395 (N_19395,N_19118,N_18958);
xnor U19396 (N_19396,N_18934,N_19191);
or U19397 (N_19397,N_19116,N_19111);
and U19398 (N_19398,N_19039,N_18912);
nand U19399 (N_19399,N_18863,N_18829);
xor U19400 (N_19400,N_19045,N_18936);
and U19401 (N_19401,N_18916,N_18878);
nand U19402 (N_19402,N_18935,N_19140);
nand U19403 (N_19403,N_19134,N_18897);
nand U19404 (N_19404,N_18911,N_18959);
nor U19405 (N_19405,N_18841,N_19002);
or U19406 (N_19406,N_19055,N_18929);
or U19407 (N_19407,N_18889,N_19134);
nand U19408 (N_19408,N_19128,N_18863);
nand U19409 (N_19409,N_18856,N_18801);
nor U19410 (N_19410,N_18922,N_19142);
nand U19411 (N_19411,N_18844,N_19167);
nor U19412 (N_19412,N_18972,N_18836);
or U19413 (N_19413,N_19137,N_18960);
or U19414 (N_19414,N_18967,N_19157);
nand U19415 (N_19415,N_19006,N_19139);
and U19416 (N_19416,N_19036,N_18967);
and U19417 (N_19417,N_19073,N_18839);
or U19418 (N_19418,N_18905,N_19107);
xor U19419 (N_19419,N_19144,N_19042);
and U19420 (N_19420,N_19075,N_18808);
xnor U19421 (N_19421,N_18854,N_19053);
nand U19422 (N_19422,N_19198,N_18979);
xor U19423 (N_19423,N_18869,N_18893);
xnor U19424 (N_19424,N_19178,N_19043);
xnor U19425 (N_19425,N_19086,N_19026);
xor U19426 (N_19426,N_18814,N_18984);
nor U19427 (N_19427,N_19066,N_19115);
nand U19428 (N_19428,N_19160,N_19051);
and U19429 (N_19429,N_18892,N_19140);
nor U19430 (N_19430,N_19092,N_19183);
xor U19431 (N_19431,N_19010,N_19181);
nand U19432 (N_19432,N_18957,N_19020);
nand U19433 (N_19433,N_19088,N_18955);
nor U19434 (N_19434,N_18971,N_18844);
nand U19435 (N_19435,N_18874,N_18968);
nor U19436 (N_19436,N_18893,N_18851);
xnor U19437 (N_19437,N_19099,N_19056);
nand U19438 (N_19438,N_18845,N_19108);
or U19439 (N_19439,N_19029,N_18964);
or U19440 (N_19440,N_19111,N_18983);
or U19441 (N_19441,N_19045,N_19118);
nor U19442 (N_19442,N_18805,N_19069);
and U19443 (N_19443,N_18892,N_18977);
or U19444 (N_19444,N_18932,N_19169);
and U19445 (N_19445,N_18912,N_18871);
xnor U19446 (N_19446,N_19052,N_18977);
and U19447 (N_19447,N_19165,N_18801);
xor U19448 (N_19448,N_19072,N_19121);
xnor U19449 (N_19449,N_19056,N_19112);
xnor U19450 (N_19450,N_18833,N_19137);
and U19451 (N_19451,N_18895,N_19040);
or U19452 (N_19452,N_18989,N_19032);
nand U19453 (N_19453,N_18836,N_19145);
nor U19454 (N_19454,N_18853,N_18804);
nand U19455 (N_19455,N_19155,N_19152);
nand U19456 (N_19456,N_18910,N_19132);
nand U19457 (N_19457,N_19166,N_18952);
and U19458 (N_19458,N_18979,N_19079);
nor U19459 (N_19459,N_18972,N_18856);
xor U19460 (N_19460,N_19124,N_19180);
nand U19461 (N_19461,N_18929,N_19090);
and U19462 (N_19462,N_19136,N_19011);
and U19463 (N_19463,N_19194,N_19143);
and U19464 (N_19464,N_18891,N_19073);
and U19465 (N_19465,N_19000,N_18825);
xor U19466 (N_19466,N_18875,N_19034);
nand U19467 (N_19467,N_18835,N_18858);
xor U19468 (N_19468,N_18959,N_18817);
xor U19469 (N_19469,N_19149,N_19025);
or U19470 (N_19470,N_19017,N_18954);
nand U19471 (N_19471,N_19042,N_18860);
or U19472 (N_19472,N_19032,N_19070);
nor U19473 (N_19473,N_19060,N_18867);
or U19474 (N_19474,N_19003,N_19049);
xnor U19475 (N_19475,N_18904,N_18963);
and U19476 (N_19476,N_18861,N_19063);
nand U19477 (N_19477,N_18801,N_18800);
nor U19478 (N_19478,N_18942,N_18889);
nand U19479 (N_19479,N_18820,N_19160);
or U19480 (N_19480,N_18814,N_18810);
or U19481 (N_19481,N_19002,N_19118);
nand U19482 (N_19482,N_18990,N_19052);
nor U19483 (N_19483,N_18978,N_19036);
nor U19484 (N_19484,N_19129,N_19192);
nand U19485 (N_19485,N_19002,N_19164);
nor U19486 (N_19486,N_18862,N_19185);
nand U19487 (N_19487,N_19159,N_19010);
and U19488 (N_19488,N_19032,N_19080);
and U19489 (N_19489,N_18995,N_19192);
and U19490 (N_19490,N_18906,N_18834);
nand U19491 (N_19491,N_19121,N_18951);
nand U19492 (N_19492,N_18897,N_18869);
nand U19493 (N_19493,N_18847,N_18843);
or U19494 (N_19494,N_19154,N_18899);
nand U19495 (N_19495,N_19189,N_18946);
xnor U19496 (N_19496,N_18964,N_18939);
nand U19497 (N_19497,N_18893,N_18917);
or U19498 (N_19498,N_19044,N_18800);
xnor U19499 (N_19499,N_18877,N_18834);
nor U19500 (N_19500,N_18871,N_19031);
xor U19501 (N_19501,N_18911,N_19176);
nand U19502 (N_19502,N_18899,N_18890);
and U19503 (N_19503,N_18956,N_19144);
nand U19504 (N_19504,N_19120,N_19024);
xnor U19505 (N_19505,N_19077,N_19017);
or U19506 (N_19506,N_19023,N_19007);
nor U19507 (N_19507,N_19188,N_18999);
nand U19508 (N_19508,N_18819,N_19132);
xor U19509 (N_19509,N_19132,N_19159);
xnor U19510 (N_19510,N_19096,N_18823);
or U19511 (N_19511,N_18806,N_19163);
xor U19512 (N_19512,N_18844,N_18926);
or U19513 (N_19513,N_18924,N_19188);
nand U19514 (N_19514,N_18898,N_19108);
nor U19515 (N_19515,N_18817,N_18949);
nand U19516 (N_19516,N_19044,N_19173);
nand U19517 (N_19517,N_19100,N_18869);
xor U19518 (N_19518,N_19134,N_18854);
and U19519 (N_19519,N_19145,N_18914);
or U19520 (N_19520,N_19185,N_18816);
nand U19521 (N_19521,N_18862,N_18847);
xor U19522 (N_19522,N_18952,N_19129);
or U19523 (N_19523,N_19133,N_18847);
xnor U19524 (N_19524,N_19146,N_19133);
or U19525 (N_19525,N_18935,N_19116);
nand U19526 (N_19526,N_18833,N_19180);
nor U19527 (N_19527,N_19158,N_19152);
or U19528 (N_19528,N_19026,N_18907);
nand U19529 (N_19529,N_19013,N_19050);
xnor U19530 (N_19530,N_18853,N_19142);
and U19531 (N_19531,N_19039,N_19170);
nand U19532 (N_19532,N_18843,N_18986);
nand U19533 (N_19533,N_18980,N_19167);
xnor U19534 (N_19534,N_18960,N_18814);
nand U19535 (N_19535,N_19116,N_19108);
xnor U19536 (N_19536,N_19047,N_19060);
and U19537 (N_19537,N_18960,N_18805);
nand U19538 (N_19538,N_19132,N_19155);
or U19539 (N_19539,N_18857,N_19060);
nand U19540 (N_19540,N_19057,N_18913);
nor U19541 (N_19541,N_18967,N_19181);
nor U19542 (N_19542,N_18843,N_18808);
nor U19543 (N_19543,N_18892,N_19012);
and U19544 (N_19544,N_18912,N_18889);
nand U19545 (N_19545,N_19080,N_18863);
xnor U19546 (N_19546,N_19034,N_19065);
nor U19547 (N_19547,N_18918,N_19022);
or U19548 (N_19548,N_19107,N_18940);
nand U19549 (N_19549,N_19132,N_18867);
and U19550 (N_19550,N_18849,N_18884);
or U19551 (N_19551,N_18960,N_19011);
or U19552 (N_19552,N_19121,N_18960);
or U19553 (N_19553,N_19104,N_19028);
nand U19554 (N_19554,N_18899,N_18866);
or U19555 (N_19555,N_18880,N_18874);
and U19556 (N_19556,N_19043,N_18813);
nand U19557 (N_19557,N_19018,N_18928);
xor U19558 (N_19558,N_18892,N_18996);
nand U19559 (N_19559,N_18848,N_18811);
nand U19560 (N_19560,N_19061,N_18884);
or U19561 (N_19561,N_19102,N_19042);
and U19562 (N_19562,N_19172,N_19123);
xnor U19563 (N_19563,N_19182,N_18872);
or U19564 (N_19564,N_18857,N_18894);
or U19565 (N_19565,N_18858,N_18992);
or U19566 (N_19566,N_18812,N_19062);
and U19567 (N_19567,N_19106,N_19118);
nor U19568 (N_19568,N_18897,N_19060);
xnor U19569 (N_19569,N_19165,N_18854);
or U19570 (N_19570,N_19128,N_18931);
and U19571 (N_19571,N_18962,N_18870);
xor U19572 (N_19572,N_18803,N_19098);
nand U19573 (N_19573,N_18816,N_18867);
nor U19574 (N_19574,N_19065,N_19194);
nor U19575 (N_19575,N_18901,N_18876);
nor U19576 (N_19576,N_18894,N_19130);
nand U19577 (N_19577,N_19070,N_18960);
xor U19578 (N_19578,N_19004,N_18948);
or U19579 (N_19579,N_18970,N_19158);
nor U19580 (N_19580,N_19123,N_18844);
nand U19581 (N_19581,N_18888,N_18945);
or U19582 (N_19582,N_18980,N_18816);
or U19583 (N_19583,N_18854,N_18932);
xor U19584 (N_19584,N_19042,N_19155);
nand U19585 (N_19585,N_18920,N_18894);
or U19586 (N_19586,N_18919,N_18888);
nand U19587 (N_19587,N_18913,N_18915);
xor U19588 (N_19588,N_19170,N_19160);
and U19589 (N_19589,N_19076,N_18952);
and U19590 (N_19590,N_19082,N_19035);
xor U19591 (N_19591,N_19171,N_19079);
xor U19592 (N_19592,N_18825,N_18998);
nand U19593 (N_19593,N_19194,N_18887);
or U19594 (N_19594,N_19191,N_19108);
and U19595 (N_19595,N_18965,N_18884);
nand U19596 (N_19596,N_18994,N_18848);
or U19597 (N_19597,N_19035,N_18902);
xnor U19598 (N_19598,N_19194,N_19107);
and U19599 (N_19599,N_18994,N_18889);
or U19600 (N_19600,N_19391,N_19564);
nand U19601 (N_19601,N_19398,N_19572);
and U19602 (N_19602,N_19592,N_19545);
and U19603 (N_19603,N_19473,N_19229);
nor U19604 (N_19604,N_19361,N_19461);
xor U19605 (N_19605,N_19454,N_19569);
nand U19606 (N_19606,N_19577,N_19415);
nor U19607 (N_19607,N_19281,N_19340);
nand U19608 (N_19608,N_19242,N_19286);
or U19609 (N_19609,N_19432,N_19587);
nand U19610 (N_19610,N_19452,N_19335);
xor U19611 (N_19611,N_19384,N_19480);
or U19612 (N_19612,N_19259,N_19322);
nand U19613 (N_19613,N_19389,N_19532);
nor U19614 (N_19614,N_19568,N_19505);
xor U19615 (N_19615,N_19582,N_19515);
xor U19616 (N_19616,N_19268,N_19299);
or U19617 (N_19617,N_19284,N_19500);
and U19618 (N_19618,N_19430,N_19449);
and U19619 (N_19619,N_19504,N_19513);
and U19620 (N_19620,N_19221,N_19485);
xnor U19621 (N_19621,N_19364,N_19344);
nand U19622 (N_19622,N_19293,N_19230);
xnor U19623 (N_19623,N_19424,N_19362);
or U19624 (N_19624,N_19235,N_19524);
and U19625 (N_19625,N_19556,N_19442);
xnor U19626 (N_19626,N_19542,N_19216);
or U19627 (N_19627,N_19292,N_19204);
and U19628 (N_19628,N_19538,N_19313);
or U19629 (N_19629,N_19414,N_19451);
or U19630 (N_19630,N_19254,N_19366);
nand U19631 (N_19631,N_19525,N_19381);
nor U19632 (N_19632,N_19291,N_19327);
or U19633 (N_19633,N_19319,N_19562);
and U19634 (N_19634,N_19326,N_19595);
nor U19635 (N_19635,N_19285,N_19390);
and U19636 (N_19636,N_19571,N_19288);
xnor U19637 (N_19637,N_19527,N_19289);
nor U19638 (N_19638,N_19447,N_19201);
xnor U19639 (N_19639,N_19223,N_19502);
nor U19640 (N_19640,N_19388,N_19420);
nand U19641 (N_19641,N_19565,N_19533);
or U19642 (N_19642,N_19343,N_19401);
and U19643 (N_19643,N_19383,N_19446);
nor U19644 (N_19644,N_19591,N_19549);
nor U19645 (N_19645,N_19471,N_19200);
nand U19646 (N_19646,N_19375,N_19330);
and U19647 (N_19647,N_19596,N_19489);
nand U19648 (N_19648,N_19438,N_19528);
nor U19649 (N_19649,N_19211,N_19484);
xnor U19650 (N_19650,N_19298,N_19474);
nor U19651 (N_19651,N_19400,N_19363);
and U19652 (N_19652,N_19555,N_19481);
and U19653 (N_19653,N_19546,N_19277);
xor U19654 (N_19654,N_19354,N_19437);
nand U19655 (N_19655,N_19550,N_19411);
nand U19656 (N_19656,N_19267,N_19333);
xor U19657 (N_19657,N_19419,N_19578);
or U19658 (N_19658,N_19305,N_19331);
nand U19659 (N_19659,N_19580,N_19355);
nand U19660 (N_19660,N_19219,N_19205);
nand U19661 (N_19661,N_19439,N_19537);
or U19662 (N_19662,N_19349,N_19249);
and U19663 (N_19663,N_19307,N_19251);
nand U19664 (N_19664,N_19493,N_19306);
and U19665 (N_19665,N_19462,N_19244);
xor U19666 (N_19666,N_19283,N_19226);
nand U19667 (N_19667,N_19234,N_19339);
xnor U19668 (N_19668,N_19412,N_19310);
or U19669 (N_19669,N_19212,N_19560);
nor U19670 (N_19670,N_19463,N_19522);
and U19671 (N_19671,N_19465,N_19269);
nor U19672 (N_19672,N_19370,N_19365);
nor U19673 (N_19673,N_19265,N_19236);
xnor U19674 (N_19674,N_19264,N_19338);
xor U19675 (N_19675,N_19599,N_19585);
nor U19676 (N_19676,N_19252,N_19466);
nor U19677 (N_19677,N_19325,N_19294);
or U19678 (N_19678,N_19297,N_19581);
and U19679 (N_19679,N_19351,N_19304);
and U19680 (N_19680,N_19460,N_19455);
or U19681 (N_19681,N_19261,N_19290);
or U19682 (N_19682,N_19272,N_19309);
nor U19683 (N_19683,N_19404,N_19588);
or U19684 (N_19684,N_19329,N_19494);
xor U19685 (N_19685,N_19250,N_19535);
xnor U19686 (N_19686,N_19512,N_19282);
xor U19687 (N_19687,N_19403,N_19457);
xnor U19688 (N_19688,N_19429,N_19589);
xnor U19689 (N_19689,N_19213,N_19518);
xor U19690 (N_19690,N_19440,N_19217);
xor U19691 (N_19691,N_19300,N_19316);
nor U19692 (N_19692,N_19256,N_19367);
xor U19693 (N_19693,N_19237,N_19315);
nor U19694 (N_19694,N_19516,N_19397);
xnor U19695 (N_19695,N_19434,N_19496);
and U19696 (N_19696,N_19245,N_19579);
and U19697 (N_19697,N_19422,N_19436);
nand U19698 (N_19698,N_19425,N_19257);
nor U19699 (N_19699,N_19202,N_19559);
nor U19700 (N_19700,N_19413,N_19356);
and U19701 (N_19701,N_19406,N_19492);
xnor U19702 (N_19702,N_19233,N_19407);
and U19703 (N_19703,N_19220,N_19276);
xnor U19704 (N_19704,N_19321,N_19240);
or U19705 (N_19705,N_19308,N_19260);
nor U19706 (N_19706,N_19273,N_19262);
nor U19707 (N_19707,N_19295,N_19476);
nor U19708 (N_19708,N_19382,N_19453);
or U19709 (N_19709,N_19544,N_19215);
nor U19710 (N_19710,N_19408,N_19311);
nor U19711 (N_19711,N_19598,N_19353);
and U19712 (N_19712,N_19360,N_19570);
and U19713 (N_19713,N_19371,N_19593);
nand U19714 (N_19714,N_19483,N_19507);
nor U19715 (N_19715,N_19266,N_19506);
and U19716 (N_19716,N_19469,N_19405);
nor U19717 (N_19717,N_19318,N_19498);
nor U19718 (N_19718,N_19431,N_19594);
or U19719 (N_19719,N_19334,N_19279);
and U19720 (N_19720,N_19526,N_19336);
and U19721 (N_19721,N_19551,N_19418);
or U19722 (N_19722,N_19486,N_19248);
xnor U19723 (N_19723,N_19296,N_19558);
nor U19724 (N_19724,N_19369,N_19227);
nor U19725 (N_19725,N_19274,N_19243);
nand U19726 (N_19726,N_19534,N_19359);
xor U19727 (N_19727,N_19380,N_19399);
nand U19728 (N_19728,N_19239,N_19287);
and U19729 (N_19729,N_19402,N_19557);
nand U19730 (N_19730,N_19539,N_19554);
xnor U19731 (N_19731,N_19563,N_19519);
nor U19732 (N_19732,N_19443,N_19323);
or U19733 (N_19733,N_19225,N_19337);
xnor U19734 (N_19734,N_19495,N_19464);
nand U19735 (N_19735,N_19448,N_19232);
xnor U19736 (N_19736,N_19421,N_19328);
nor U19737 (N_19737,N_19458,N_19583);
nand U19738 (N_19738,N_19263,N_19520);
and U19739 (N_19739,N_19255,N_19246);
nand U19740 (N_19740,N_19553,N_19392);
nor U19741 (N_19741,N_19517,N_19374);
xnor U19742 (N_19742,N_19499,N_19586);
and U19743 (N_19743,N_19450,N_19378);
nor U19744 (N_19744,N_19433,N_19358);
nand U19745 (N_19745,N_19324,N_19428);
xnor U19746 (N_19746,N_19503,N_19491);
or U19747 (N_19747,N_19470,N_19342);
and U19748 (N_19748,N_19222,N_19472);
nor U19749 (N_19749,N_19341,N_19258);
xor U19750 (N_19750,N_19488,N_19206);
nor U19751 (N_19751,N_19314,N_19497);
xnor U19752 (N_19752,N_19467,N_19253);
nor U19753 (N_19753,N_19444,N_19247);
nand U19754 (N_19754,N_19478,N_19459);
nor U19755 (N_19755,N_19487,N_19214);
xor U19756 (N_19756,N_19270,N_19373);
nor U19757 (N_19757,N_19590,N_19409);
nor U19758 (N_19758,N_19379,N_19435);
nor U19759 (N_19759,N_19547,N_19529);
nor U19760 (N_19760,N_19368,N_19575);
or U19761 (N_19761,N_19385,N_19275);
or U19762 (N_19762,N_19301,N_19468);
nand U19763 (N_19763,N_19372,N_19548);
or U19764 (N_19764,N_19231,N_19521);
xor U19765 (N_19765,N_19543,N_19395);
nand U19766 (N_19766,N_19224,N_19376);
nor U19767 (N_19767,N_19238,N_19394);
xnor U19768 (N_19768,N_19208,N_19386);
and U19769 (N_19769,N_19576,N_19241);
and U19770 (N_19770,N_19278,N_19574);
and U19771 (N_19771,N_19584,N_19203);
and U19772 (N_19772,N_19352,N_19312);
or U19773 (N_19773,N_19477,N_19423);
or U19774 (N_19774,N_19207,N_19597);
and U19775 (N_19775,N_19302,N_19445);
or U19776 (N_19776,N_19303,N_19456);
xnor U19777 (N_19777,N_19417,N_19490);
nand U19778 (N_19778,N_19540,N_19531);
and U19779 (N_19779,N_19320,N_19511);
xor U19780 (N_19780,N_19210,N_19396);
nand U19781 (N_19781,N_19573,N_19393);
nand U19782 (N_19782,N_19410,N_19479);
and U19783 (N_19783,N_19332,N_19350);
or U19784 (N_19784,N_19348,N_19482);
and U19785 (N_19785,N_19501,N_19218);
and U19786 (N_19786,N_19552,N_19541);
or U19787 (N_19787,N_19510,N_19567);
and U19788 (N_19788,N_19317,N_19530);
and U19789 (N_19789,N_19347,N_19209);
nor U19790 (N_19790,N_19561,N_19377);
or U19791 (N_19791,N_19566,N_19271);
and U19792 (N_19792,N_19346,N_19387);
or U19793 (N_19793,N_19509,N_19280);
xor U19794 (N_19794,N_19514,N_19475);
nor U19795 (N_19795,N_19508,N_19523);
nand U19796 (N_19796,N_19345,N_19357);
xor U19797 (N_19797,N_19427,N_19228);
and U19798 (N_19798,N_19416,N_19426);
nand U19799 (N_19799,N_19441,N_19536);
nor U19800 (N_19800,N_19467,N_19596);
nand U19801 (N_19801,N_19221,N_19554);
nand U19802 (N_19802,N_19279,N_19359);
xnor U19803 (N_19803,N_19358,N_19520);
nor U19804 (N_19804,N_19417,N_19298);
and U19805 (N_19805,N_19309,N_19546);
and U19806 (N_19806,N_19386,N_19215);
nand U19807 (N_19807,N_19506,N_19383);
or U19808 (N_19808,N_19469,N_19223);
nor U19809 (N_19809,N_19222,N_19466);
nor U19810 (N_19810,N_19347,N_19316);
and U19811 (N_19811,N_19504,N_19312);
and U19812 (N_19812,N_19311,N_19264);
and U19813 (N_19813,N_19241,N_19466);
nand U19814 (N_19814,N_19228,N_19510);
nor U19815 (N_19815,N_19542,N_19496);
xor U19816 (N_19816,N_19563,N_19205);
and U19817 (N_19817,N_19337,N_19232);
and U19818 (N_19818,N_19352,N_19295);
xor U19819 (N_19819,N_19571,N_19510);
or U19820 (N_19820,N_19473,N_19321);
xor U19821 (N_19821,N_19427,N_19345);
or U19822 (N_19822,N_19556,N_19445);
and U19823 (N_19823,N_19592,N_19451);
nand U19824 (N_19824,N_19243,N_19595);
and U19825 (N_19825,N_19489,N_19506);
xnor U19826 (N_19826,N_19324,N_19210);
xnor U19827 (N_19827,N_19253,N_19338);
xnor U19828 (N_19828,N_19298,N_19335);
nand U19829 (N_19829,N_19538,N_19412);
nand U19830 (N_19830,N_19511,N_19275);
nor U19831 (N_19831,N_19332,N_19428);
nor U19832 (N_19832,N_19208,N_19366);
nor U19833 (N_19833,N_19339,N_19225);
and U19834 (N_19834,N_19553,N_19294);
nor U19835 (N_19835,N_19576,N_19380);
or U19836 (N_19836,N_19233,N_19498);
nand U19837 (N_19837,N_19557,N_19440);
xor U19838 (N_19838,N_19562,N_19387);
and U19839 (N_19839,N_19574,N_19345);
nor U19840 (N_19840,N_19327,N_19345);
nor U19841 (N_19841,N_19329,N_19522);
nor U19842 (N_19842,N_19384,N_19404);
or U19843 (N_19843,N_19303,N_19489);
and U19844 (N_19844,N_19285,N_19465);
nor U19845 (N_19845,N_19314,N_19406);
and U19846 (N_19846,N_19413,N_19436);
nor U19847 (N_19847,N_19317,N_19532);
and U19848 (N_19848,N_19438,N_19417);
xnor U19849 (N_19849,N_19421,N_19256);
nand U19850 (N_19850,N_19283,N_19252);
and U19851 (N_19851,N_19436,N_19369);
nor U19852 (N_19852,N_19555,N_19405);
xnor U19853 (N_19853,N_19406,N_19367);
nand U19854 (N_19854,N_19479,N_19580);
nor U19855 (N_19855,N_19370,N_19389);
or U19856 (N_19856,N_19306,N_19410);
and U19857 (N_19857,N_19554,N_19545);
nor U19858 (N_19858,N_19598,N_19222);
nor U19859 (N_19859,N_19448,N_19374);
and U19860 (N_19860,N_19594,N_19337);
xor U19861 (N_19861,N_19304,N_19470);
nand U19862 (N_19862,N_19322,N_19489);
and U19863 (N_19863,N_19338,N_19391);
nand U19864 (N_19864,N_19291,N_19559);
nor U19865 (N_19865,N_19435,N_19363);
nand U19866 (N_19866,N_19469,N_19541);
nor U19867 (N_19867,N_19465,N_19545);
and U19868 (N_19868,N_19339,N_19583);
or U19869 (N_19869,N_19211,N_19264);
nor U19870 (N_19870,N_19438,N_19357);
and U19871 (N_19871,N_19376,N_19338);
nand U19872 (N_19872,N_19468,N_19453);
or U19873 (N_19873,N_19576,N_19425);
or U19874 (N_19874,N_19417,N_19364);
nor U19875 (N_19875,N_19450,N_19282);
nor U19876 (N_19876,N_19367,N_19228);
nand U19877 (N_19877,N_19364,N_19286);
nand U19878 (N_19878,N_19279,N_19537);
xor U19879 (N_19879,N_19416,N_19384);
and U19880 (N_19880,N_19402,N_19417);
or U19881 (N_19881,N_19426,N_19567);
nand U19882 (N_19882,N_19393,N_19586);
or U19883 (N_19883,N_19524,N_19284);
xnor U19884 (N_19884,N_19599,N_19451);
or U19885 (N_19885,N_19554,N_19462);
xor U19886 (N_19886,N_19332,N_19483);
or U19887 (N_19887,N_19564,N_19532);
nor U19888 (N_19888,N_19560,N_19291);
xnor U19889 (N_19889,N_19338,N_19462);
nor U19890 (N_19890,N_19530,N_19473);
nand U19891 (N_19891,N_19425,N_19254);
and U19892 (N_19892,N_19543,N_19582);
xor U19893 (N_19893,N_19486,N_19528);
nor U19894 (N_19894,N_19585,N_19223);
nand U19895 (N_19895,N_19266,N_19285);
nor U19896 (N_19896,N_19523,N_19518);
nor U19897 (N_19897,N_19488,N_19537);
nor U19898 (N_19898,N_19415,N_19262);
nor U19899 (N_19899,N_19455,N_19313);
nand U19900 (N_19900,N_19385,N_19367);
or U19901 (N_19901,N_19248,N_19548);
or U19902 (N_19902,N_19535,N_19363);
xor U19903 (N_19903,N_19273,N_19258);
nand U19904 (N_19904,N_19226,N_19244);
nor U19905 (N_19905,N_19562,N_19212);
and U19906 (N_19906,N_19236,N_19411);
nand U19907 (N_19907,N_19433,N_19455);
nand U19908 (N_19908,N_19499,N_19297);
and U19909 (N_19909,N_19539,N_19335);
xnor U19910 (N_19910,N_19563,N_19363);
and U19911 (N_19911,N_19533,N_19324);
and U19912 (N_19912,N_19354,N_19235);
xor U19913 (N_19913,N_19494,N_19385);
or U19914 (N_19914,N_19361,N_19370);
nor U19915 (N_19915,N_19503,N_19596);
xor U19916 (N_19916,N_19571,N_19596);
xnor U19917 (N_19917,N_19528,N_19374);
nand U19918 (N_19918,N_19381,N_19538);
xnor U19919 (N_19919,N_19208,N_19307);
and U19920 (N_19920,N_19309,N_19505);
xor U19921 (N_19921,N_19543,N_19277);
xor U19922 (N_19922,N_19475,N_19244);
and U19923 (N_19923,N_19384,N_19261);
or U19924 (N_19924,N_19313,N_19491);
nor U19925 (N_19925,N_19417,N_19429);
or U19926 (N_19926,N_19489,N_19335);
nand U19927 (N_19927,N_19344,N_19399);
nand U19928 (N_19928,N_19221,N_19567);
nor U19929 (N_19929,N_19280,N_19447);
and U19930 (N_19930,N_19524,N_19394);
xnor U19931 (N_19931,N_19291,N_19296);
and U19932 (N_19932,N_19377,N_19457);
nand U19933 (N_19933,N_19518,N_19426);
xnor U19934 (N_19934,N_19296,N_19509);
and U19935 (N_19935,N_19224,N_19368);
nor U19936 (N_19936,N_19253,N_19371);
nor U19937 (N_19937,N_19565,N_19418);
and U19938 (N_19938,N_19490,N_19315);
nand U19939 (N_19939,N_19235,N_19405);
nand U19940 (N_19940,N_19302,N_19337);
xnor U19941 (N_19941,N_19329,N_19251);
and U19942 (N_19942,N_19490,N_19564);
nand U19943 (N_19943,N_19213,N_19366);
nand U19944 (N_19944,N_19564,N_19255);
and U19945 (N_19945,N_19532,N_19230);
nor U19946 (N_19946,N_19335,N_19483);
nor U19947 (N_19947,N_19412,N_19301);
or U19948 (N_19948,N_19221,N_19210);
nand U19949 (N_19949,N_19401,N_19279);
and U19950 (N_19950,N_19526,N_19317);
nor U19951 (N_19951,N_19443,N_19290);
nor U19952 (N_19952,N_19513,N_19250);
and U19953 (N_19953,N_19537,N_19563);
xnor U19954 (N_19954,N_19331,N_19395);
or U19955 (N_19955,N_19263,N_19363);
and U19956 (N_19956,N_19241,N_19389);
xor U19957 (N_19957,N_19529,N_19456);
xnor U19958 (N_19958,N_19338,N_19466);
xor U19959 (N_19959,N_19405,N_19436);
nand U19960 (N_19960,N_19472,N_19219);
xor U19961 (N_19961,N_19262,N_19495);
and U19962 (N_19962,N_19374,N_19336);
nand U19963 (N_19963,N_19270,N_19393);
xor U19964 (N_19964,N_19507,N_19220);
or U19965 (N_19965,N_19534,N_19235);
nor U19966 (N_19966,N_19368,N_19391);
nor U19967 (N_19967,N_19368,N_19397);
and U19968 (N_19968,N_19259,N_19320);
and U19969 (N_19969,N_19235,N_19325);
and U19970 (N_19970,N_19218,N_19505);
xnor U19971 (N_19971,N_19432,N_19234);
nor U19972 (N_19972,N_19224,N_19474);
nor U19973 (N_19973,N_19523,N_19473);
xnor U19974 (N_19974,N_19302,N_19577);
xnor U19975 (N_19975,N_19273,N_19299);
and U19976 (N_19976,N_19298,N_19236);
xnor U19977 (N_19977,N_19492,N_19205);
or U19978 (N_19978,N_19404,N_19591);
nor U19979 (N_19979,N_19413,N_19305);
nand U19980 (N_19980,N_19220,N_19297);
nand U19981 (N_19981,N_19379,N_19250);
and U19982 (N_19982,N_19279,N_19293);
and U19983 (N_19983,N_19572,N_19502);
and U19984 (N_19984,N_19226,N_19230);
or U19985 (N_19985,N_19303,N_19439);
xnor U19986 (N_19986,N_19358,N_19258);
or U19987 (N_19987,N_19250,N_19478);
nand U19988 (N_19988,N_19429,N_19503);
or U19989 (N_19989,N_19416,N_19285);
and U19990 (N_19990,N_19285,N_19493);
or U19991 (N_19991,N_19222,N_19304);
nor U19992 (N_19992,N_19547,N_19440);
nand U19993 (N_19993,N_19494,N_19470);
or U19994 (N_19994,N_19291,N_19307);
and U19995 (N_19995,N_19312,N_19226);
or U19996 (N_19996,N_19452,N_19466);
or U19997 (N_19997,N_19438,N_19590);
nor U19998 (N_19998,N_19472,N_19224);
xnor U19999 (N_19999,N_19268,N_19321);
or UO_0 (O_0,N_19664,N_19966);
nand UO_1 (O_1,N_19703,N_19820);
nor UO_2 (O_2,N_19997,N_19620);
nand UO_3 (O_3,N_19771,N_19626);
nand UO_4 (O_4,N_19780,N_19706);
nand UO_5 (O_5,N_19674,N_19775);
or UO_6 (O_6,N_19690,N_19833);
xnor UO_7 (O_7,N_19750,N_19684);
nand UO_8 (O_8,N_19954,N_19976);
and UO_9 (O_9,N_19808,N_19752);
or UO_10 (O_10,N_19759,N_19678);
nor UO_11 (O_11,N_19985,N_19854);
or UO_12 (O_12,N_19915,N_19831);
nand UO_13 (O_13,N_19799,N_19961);
nand UO_14 (O_14,N_19712,N_19627);
and UO_15 (O_15,N_19959,N_19872);
and UO_16 (O_16,N_19785,N_19629);
or UO_17 (O_17,N_19903,N_19718);
or UO_18 (O_18,N_19793,N_19933);
nor UO_19 (O_19,N_19797,N_19601);
nand UO_20 (O_20,N_19930,N_19751);
xnor UO_21 (O_21,N_19823,N_19864);
or UO_22 (O_22,N_19732,N_19618);
or UO_23 (O_23,N_19858,N_19708);
nand UO_24 (O_24,N_19981,N_19711);
nor UO_25 (O_25,N_19757,N_19746);
and UO_26 (O_26,N_19975,N_19801);
nand UO_27 (O_27,N_19779,N_19825);
xnor UO_28 (O_28,N_19972,N_19683);
xnor UO_29 (O_29,N_19624,N_19867);
nor UO_30 (O_30,N_19869,N_19804);
and UO_31 (O_31,N_19646,N_19693);
xnor UO_32 (O_32,N_19896,N_19717);
nor UO_33 (O_33,N_19734,N_19743);
or UO_34 (O_34,N_19821,N_19947);
or UO_35 (O_35,N_19698,N_19894);
and UO_36 (O_36,N_19829,N_19689);
nand UO_37 (O_37,N_19950,N_19639);
or UO_38 (O_38,N_19605,N_19745);
or UO_39 (O_39,N_19748,N_19739);
nand UO_40 (O_40,N_19974,N_19670);
nor UO_41 (O_41,N_19921,N_19982);
or UO_42 (O_42,N_19967,N_19811);
xor UO_43 (O_43,N_19849,N_19892);
and UO_44 (O_44,N_19875,N_19819);
or UO_45 (O_45,N_19913,N_19705);
or UO_46 (O_46,N_19891,N_19859);
xnor UO_47 (O_47,N_19616,N_19932);
nor UO_48 (O_48,N_19955,N_19958);
xnor UO_49 (O_49,N_19792,N_19747);
xnor UO_50 (O_50,N_19699,N_19986);
nor UO_51 (O_51,N_19978,N_19631);
and UO_52 (O_52,N_19787,N_19878);
or UO_53 (O_53,N_19687,N_19672);
xnor UO_54 (O_54,N_19650,N_19742);
nand UO_55 (O_55,N_19905,N_19802);
nor UO_56 (O_56,N_19635,N_19874);
or UO_57 (O_57,N_19862,N_19924);
or UO_58 (O_58,N_19965,N_19740);
and UO_59 (O_59,N_19764,N_19991);
and UO_60 (O_60,N_19604,N_19756);
and UO_61 (O_61,N_19658,N_19656);
nor UO_62 (O_62,N_19918,N_19938);
xnor UO_63 (O_63,N_19637,N_19948);
xnor UO_64 (O_64,N_19715,N_19619);
nand UO_65 (O_65,N_19931,N_19939);
nor UO_66 (O_66,N_19716,N_19815);
xnor UO_67 (O_67,N_19813,N_19912);
nand UO_68 (O_68,N_19881,N_19884);
nand UO_69 (O_69,N_19988,N_19774);
xnor UO_70 (O_70,N_19890,N_19606);
nand UO_71 (O_71,N_19856,N_19807);
or UO_72 (O_72,N_19772,N_19790);
xor UO_73 (O_73,N_19843,N_19979);
nor UO_74 (O_74,N_19614,N_19769);
and UO_75 (O_75,N_19659,N_19640);
or UO_76 (O_76,N_19749,N_19704);
or UO_77 (O_77,N_19860,N_19852);
nand UO_78 (O_78,N_19876,N_19902);
nand UO_79 (O_79,N_19638,N_19855);
nand UO_80 (O_80,N_19861,N_19673);
or UO_81 (O_81,N_19736,N_19617);
or UO_82 (O_82,N_19697,N_19768);
nor UO_83 (O_83,N_19720,N_19865);
and UO_84 (O_84,N_19755,N_19761);
xnor UO_85 (O_85,N_19642,N_19953);
nand UO_86 (O_86,N_19655,N_19737);
xor UO_87 (O_87,N_19844,N_19887);
or UO_88 (O_88,N_19733,N_19773);
and UO_89 (O_89,N_19866,N_19900);
or UO_90 (O_90,N_19814,N_19722);
and UO_91 (O_91,N_19798,N_19879);
or UO_92 (O_92,N_19968,N_19994);
nor UO_93 (O_93,N_19837,N_19923);
nand UO_94 (O_94,N_19665,N_19653);
nor UO_95 (O_95,N_19870,N_19803);
xor UO_96 (O_96,N_19694,N_19692);
nor UO_97 (O_97,N_19645,N_19731);
nand UO_98 (O_98,N_19990,N_19877);
or UO_99 (O_99,N_19971,N_19662);
nor UO_100 (O_100,N_19758,N_19842);
nor UO_101 (O_101,N_19857,N_19969);
nor UO_102 (O_102,N_19784,N_19984);
nand UO_103 (O_103,N_19663,N_19686);
nor UO_104 (O_104,N_19666,N_19956);
xnor UO_105 (O_105,N_19911,N_19841);
nor UO_106 (O_106,N_19753,N_19928);
nor UO_107 (O_107,N_19776,N_19936);
nand UO_108 (O_108,N_19868,N_19770);
and UO_109 (O_109,N_19993,N_19871);
nor UO_110 (O_110,N_19783,N_19895);
nor UO_111 (O_111,N_19839,N_19727);
nor UO_112 (O_112,N_19679,N_19945);
nor UO_113 (O_113,N_19644,N_19735);
nor UO_114 (O_114,N_19880,N_19760);
xor UO_115 (O_115,N_19724,N_19778);
and UO_116 (O_116,N_19987,N_19668);
nor UO_117 (O_117,N_19602,N_19794);
xor UO_118 (O_118,N_19763,N_19669);
nor UO_119 (O_119,N_19942,N_19889);
nand UO_120 (O_120,N_19714,N_19719);
xnor UO_121 (O_121,N_19782,N_19973);
or UO_122 (O_122,N_19647,N_19651);
nand UO_123 (O_123,N_19998,N_19701);
nor UO_124 (O_124,N_19847,N_19846);
xor UO_125 (O_125,N_19609,N_19922);
nand UO_126 (O_126,N_19634,N_19927);
nor UO_127 (O_127,N_19612,N_19713);
or UO_128 (O_128,N_19741,N_19685);
xnor UO_129 (O_129,N_19816,N_19677);
xnor UO_130 (O_130,N_19957,N_19652);
xnor UO_131 (O_131,N_19929,N_19691);
nor UO_132 (O_132,N_19788,N_19886);
xor UO_133 (O_133,N_19630,N_19908);
and UO_134 (O_134,N_19850,N_19700);
and UO_135 (O_135,N_19901,N_19834);
xor UO_136 (O_136,N_19611,N_19920);
and UO_137 (O_137,N_19723,N_19996);
nor UO_138 (O_138,N_19962,N_19657);
nor UO_139 (O_139,N_19963,N_19628);
nor UO_140 (O_140,N_19688,N_19800);
nor UO_141 (O_141,N_19934,N_19682);
xor UO_142 (O_142,N_19730,N_19809);
or UO_143 (O_143,N_19964,N_19989);
or UO_144 (O_144,N_19835,N_19840);
and UO_145 (O_145,N_19943,N_19710);
nor UO_146 (O_146,N_19944,N_19925);
and UO_147 (O_147,N_19853,N_19941);
nor UO_148 (O_148,N_19952,N_19812);
nor UO_149 (O_149,N_19643,N_19830);
nand UO_150 (O_150,N_19951,N_19926);
nor UO_151 (O_151,N_19897,N_19882);
nor UO_152 (O_152,N_19600,N_19827);
and UO_153 (O_153,N_19649,N_19828);
xnor UO_154 (O_154,N_19603,N_19786);
or UO_155 (O_155,N_19695,N_19725);
nand UO_156 (O_156,N_19817,N_19818);
nand UO_157 (O_157,N_19940,N_19671);
xnor UO_158 (O_158,N_19781,N_19980);
nand UO_159 (O_159,N_19765,N_19917);
nor UO_160 (O_160,N_19910,N_19851);
nor UO_161 (O_161,N_19661,N_19762);
nand UO_162 (O_162,N_19960,N_19622);
xnor UO_163 (O_163,N_19625,N_19623);
nand UO_164 (O_164,N_19914,N_19728);
xor UO_165 (O_165,N_19767,N_19909);
nand UO_166 (O_166,N_19777,N_19709);
and UO_167 (O_167,N_19806,N_19796);
or UO_168 (O_168,N_19907,N_19893);
and UO_169 (O_169,N_19845,N_19633);
and UO_170 (O_170,N_19826,N_19848);
nand UO_171 (O_171,N_19977,N_19729);
or UO_172 (O_172,N_19999,N_19754);
nand UO_173 (O_173,N_19791,N_19738);
or UO_174 (O_174,N_19681,N_19883);
or UO_175 (O_175,N_19899,N_19824);
xor UO_176 (O_176,N_19946,N_19995);
nand UO_177 (O_177,N_19766,N_19744);
or UO_178 (O_178,N_19696,N_19832);
nand UO_179 (O_179,N_19675,N_19726);
or UO_180 (O_180,N_19885,N_19937);
or UO_181 (O_181,N_19707,N_19836);
nand UO_182 (O_182,N_19919,N_19992);
and UO_183 (O_183,N_19805,N_19654);
nor UO_184 (O_184,N_19607,N_19680);
nor UO_185 (O_185,N_19610,N_19904);
or UO_186 (O_186,N_19608,N_19838);
or UO_187 (O_187,N_19873,N_19916);
nor UO_188 (O_188,N_19702,N_19898);
and UO_189 (O_189,N_19863,N_19983);
xor UO_190 (O_190,N_19810,N_19906);
and UO_191 (O_191,N_19648,N_19935);
xnor UO_192 (O_192,N_19636,N_19970);
nor UO_193 (O_193,N_19615,N_19795);
and UO_194 (O_194,N_19949,N_19621);
nand UO_195 (O_195,N_19721,N_19641);
nor UO_196 (O_196,N_19667,N_19789);
nand UO_197 (O_197,N_19888,N_19660);
nor UO_198 (O_198,N_19822,N_19613);
xnor UO_199 (O_199,N_19632,N_19676);
nand UO_200 (O_200,N_19870,N_19865);
nand UO_201 (O_201,N_19719,N_19834);
or UO_202 (O_202,N_19922,N_19814);
or UO_203 (O_203,N_19694,N_19948);
xnor UO_204 (O_204,N_19864,N_19685);
or UO_205 (O_205,N_19921,N_19672);
or UO_206 (O_206,N_19824,N_19895);
and UO_207 (O_207,N_19930,N_19947);
xor UO_208 (O_208,N_19865,N_19960);
nand UO_209 (O_209,N_19703,N_19928);
and UO_210 (O_210,N_19879,N_19975);
and UO_211 (O_211,N_19941,N_19919);
xnor UO_212 (O_212,N_19855,N_19870);
nand UO_213 (O_213,N_19620,N_19945);
and UO_214 (O_214,N_19932,N_19959);
xnor UO_215 (O_215,N_19769,N_19880);
or UO_216 (O_216,N_19735,N_19698);
and UO_217 (O_217,N_19666,N_19779);
nor UO_218 (O_218,N_19629,N_19602);
nand UO_219 (O_219,N_19881,N_19792);
xnor UO_220 (O_220,N_19779,N_19604);
xor UO_221 (O_221,N_19994,N_19700);
nor UO_222 (O_222,N_19994,N_19987);
nor UO_223 (O_223,N_19666,N_19853);
and UO_224 (O_224,N_19920,N_19834);
and UO_225 (O_225,N_19882,N_19895);
and UO_226 (O_226,N_19913,N_19726);
and UO_227 (O_227,N_19943,N_19828);
nand UO_228 (O_228,N_19867,N_19727);
and UO_229 (O_229,N_19619,N_19610);
and UO_230 (O_230,N_19842,N_19998);
nand UO_231 (O_231,N_19612,N_19741);
nor UO_232 (O_232,N_19811,N_19882);
and UO_233 (O_233,N_19873,N_19761);
and UO_234 (O_234,N_19906,N_19741);
nor UO_235 (O_235,N_19947,N_19774);
nor UO_236 (O_236,N_19915,N_19617);
nor UO_237 (O_237,N_19784,N_19855);
and UO_238 (O_238,N_19860,N_19687);
nor UO_239 (O_239,N_19755,N_19787);
nand UO_240 (O_240,N_19952,N_19749);
nand UO_241 (O_241,N_19945,N_19777);
xnor UO_242 (O_242,N_19724,N_19647);
or UO_243 (O_243,N_19837,N_19807);
xor UO_244 (O_244,N_19711,N_19855);
or UO_245 (O_245,N_19758,N_19974);
nand UO_246 (O_246,N_19951,N_19899);
and UO_247 (O_247,N_19852,N_19767);
xnor UO_248 (O_248,N_19890,N_19801);
xor UO_249 (O_249,N_19664,N_19750);
xnor UO_250 (O_250,N_19843,N_19986);
or UO_251 (O_251,N_19902,N_19841);
or UO_252 (O_252,N_19673,N_19988);
nand UO_253 (O_253,N_19924,N_19728);
or UO_254 (O_254,N_19732,N_19846);
nand UO_255 (O_255,N_19940,N_19761);
nor UO_256 (O_256,N_19635,N_19863);
xnor UO_257 (O_257,N_19697,N_19602);
nand UO_258 (O_258,N_19659,N_19944);
or UO_259 (O_259,N_19611,N_19878);
and UO_260 (O_260,N_19703,N_19640);
xnor UO_261 (O_261,N_19707,N_19727);
nor UO_262 (O_262,N_19913,N_19968);
or UO_263 (O_263,N_19613,N_19782);
xor UO_264 (O_264,N_19894,N_19826);
nand UO_265 (O_265,N_19817,N_19911);
or UO_266 (O_266,N_19699,N_19670);
xnor UO_267 (O_267,N_19806,N_19844);
or UO_268 (O_268,N_19724,N_19666);
xor UO_269 (O_269,N_19850,N_19783);
and UO_270 (O_270,N_19778,N_19638);
or UO_271 (O_271,N_19975,N_19629);
nand UO_272 (O_272,N_19956,N_19662);
nand UO_273 (O_273,N_19645,N_19774);
nor UO_274 (O_274,N_19688,N_19723);
and UO_275 (O_275,N_19781,N_19649);
and UO_276 (O_276,N_19692,N_19748);
and UO_277 (O_277,N_19925,N_19707);
xnor UO_278 (O_278,N_19775,N_19632);
and UO_279 (O_279,N_19994,N_19966);
nor UO_280 (O_280,N_19636,N_19994);
xor UO_281 (O_281,N_19783,N_19845);
or UO_282 (O_282,N_19808,N_19848);
or UO_283 (O_283,N_19621,N_19723);
nor UO_284 (O_284,N_19847,N_19620);
and UO_285 (O_285,N_19748,N_19687);
and UO_286 (O_286,N_19712,N_19783);
nor UO_287 (O_287,N_19835,N_19759);
and UO_288 (O_288,N_19909,N_19746);
and UO_289 (O_289,N_19639,N_19728);
xnor UO_290 (O_290,N_19729,N_19875);
and UO_291 (O_291,N_19932,N_19808);
and UO_292 (O_292,N_19884,N_19727);
and UO_293 (O_293,N_19689,N_19997);
nand UO_294 (O_294,N_19967,N_19657);
and UO_295 (O_295,N_19851,N_19722);
nand UO_296 (O_296,N_19954,N_19625);
or UO_297 (O_297,N_19612,N_19684);
nand UO_298 (O_298,N_19665,N_19682);
or UO_299 (O_299,N_19761,N_19626);
nor UO_300 (O_300,N_19999,N_19807);
nand UO_301 (O_301,N_19660,N_19919);
nor UO_302 (O_302,N_19954,N_19915);
and UO_303 (O_303,N_19779,N_19988);
xnor UO_304 (O_304,N_19745,N_19782);
or UO_305 (O_305,N_19663,N_19895);
or UO_306 (O_306,N_19606,N_19782);
xnor UO_307 (O_307,N_19894,N_19939);
and UO_308 (O_308,N_19817,N_19847);
or UO_309 (O_309,N_19745,N_19731);
or UO_310 (O_310,N_19924,N_19622);
nor UO_311 (O_311,N_19967,N_19659);
nand UO_312 (O_312,N_19607,N_19609);
nand UO_313 (O_313,N_19795,N_19831);
xnor UO_314 (O_314,N_19943,N_19910);
and UO_315 (O_315,N_19921,N_19783);
or UO_316 (O_316,N_19729,N_19827);
nand UO_317 (O_317,N_19811,N_19890);
xor UO_318 (O_318,N_19980,N_19899);
nand UO_319 (O_319,N_19966,N_19952);
nor UO_320 (O_320,N_19789,N_19601);
nor UO_321 (O_321,N_19700,N_19703);
and UO_322 (O_322,N_19748,N_19975);
or UO_323 (O_323,N_19706,N_19776);
nor UO_324 (O_324,N_19792,N_19659);
and UO_325 (O_325,N_19902,N_19798);
and UO_326 (O_326,N_19952,N_19685);
nand UO_327 (O_327,N_19627,N_19867);
nor UO_328 (O_328,N_19919,N_19824);
nor UO_329 (O_329,N_19806,N_19786);
or UO_330 (O_330,N_19749,N_19767);
nand UO_331 (O_331,N_19874,N_19861);
and UO_332 (O_332,N_19614,N_19921);
or UO_333 (O_333,N_19778,N_19926);
and UO_334 (O_334,N_19717,N_19630);
nor UO_335 (O_335,N_19864,N_19679);
xnor UO_336 (O_336,N_19732,N_19839);
xnor UO_337 (O_337,N_19943,N_19956);
nand UO_338 (O_338,N_19712,N_19637);
nand UO_339 (O_339,N_19620,N_19826);
nand UO_340 (O_340,N_19636,N_19991);
nor UO_341 (O_341,N_19833,N_19932);
and UO_342 (O_342,N_19798,N_19833);
or UO_343 (O_343,N_19645,N_19851);
nor UO_344 (O_344,N_19947,N_19885);
nor UO_345 (O_345,N_19826,N_19634);
and UO_346 (O_346,N_19940,N_19654);
and UO_347 (O_347,N_19759,N_19747);
xor UO_348 (O_348,N_19930,N_19999);
or UO_349 (O_349,N_19804,N_19710);
xor UO_350 (O_350,N_19839,N_19602);
or UO_351 (O_351,N_19982,N_19631);
nand UO_352 (O_352,N_19844,N_19759);
nand UO_353 (O_353,N_19889,N_19776);
xnor UO_354 (O_354,N_19955,N_19659);
xnor UO_355 (O_355,N_19750,N_19889);
or UO_356 (O_356,N_19689,N_19993);
xnor UO_357 (O_357,N_19893,N_19938);
and UO_358 (O_358,N_19867,N_19855);
nand UO_359 (O_359,N_19882,N_19876);
nand UO_360 (O_360,N_19607,N_19894);
and UO_361 (O_361,N_19795,N_19694);
nor UO_362 (O_362,N_19606,N_19757);
xor UO_363 (O_363,N_19967,N_19685);
and UO_364 (O_364,N_19704,N_19679);
nand UO_365 (O_365,N_19666,N_19649);
nand UO_366 (O_366,N_19606,N_19876);
nor UO_367 (O_367,N_19856,N_19819);
nand UO_368 (O_368,N_19603,N_19772);
nand UO_369 (O_369,N_19961,N_19866);
or UO_370 (O_370,N_19723,N_19808);
xnor UO_371 (O_371,N_19982,N_19637);
xnor UO_372 (O_372,N_19907,N_19743);
nor UO_373 (O_373,N_19944,N_19928);
nor UO_374 (O_374,N_19761,N_19779);
or UO_375 (O_375,N_19785,N_19839);
nand UO_376 (O_376,N_19752,N_19904);
xnor UO_377 (O_377,N_19828,N_19827);
nand UO_378 (O_378,N_19889,N_19819);
nor UO_379 (O_379,N_19870,N_19971);
nand UO_380 (O_380,N_19704,N_19965);
and UO_381 (O_381,N_19932,N_19873);
or UO_382 (O_382,N_19855,N_19787);
nand UO_383 (O_383,N_19873,N_19970);
and UO_384 (O_384,N_19775,N_19615);
nor UO_385 (O_385,N_19624,N_19669);
nand UO_386 (O_386,N_19961,N_19817);
or UO_387 (O_387,N_19653,N_19820);
nand UO_388 (O_388,N_19609,N_19869);
or UO_389 (O_389,N_19657,N_19770);
nor UO_390 (O_390,N_19824,N_19709);
nor UO_391 (O_391,N_19708,N_19820);
or UO_392 (O_392,N_19973,N_19698);
nand UO_393 (O_393,N_19800,N_19999);
nand UO_394 (O_394,N_19745,N_19730);
and UO_395 (O_395,N_19703,N_19752);
or UO_396 (O_396,N_19927,N_19813);
or UO_397 (O_397,N_19662,N_19722);
or UO_398 (O_398,N_19763,N_19636);
nor UO_399 (O_399,N_19708,N_19633);
nand UO_400 (O_400,N_19873,N_19674);
or UO_401 (O_401,N_19959,N_19647);
nand UO_402 (O_402,N_19917,N_19641);
nand UO_403 (O_403,N_19918,N_19799);
or UO_404 (O_404,N_19746,N_19626);
or UO_405 (O_405,N_19673,N_19724);
nor UO_406 (O_406,N_19834,N_19876);
nand UO_407 (O_407,N_19827,N_19932);
xnor UO_408 (O_408,N_19606,N_19621);
nor UO_409 (O_409,N_19845,N_19744);
or UO_410 (O_410,N_19793,N_19637);
nand UO_411 (O_411,N_19741,N_19609);
nand UO_412 (O_412,N_19919,N_19821);
nor UO_413 (O_413,N_19635,N_19885);
nor UO_414 (O_414,N_19936,N_19737);
nor UO_415 (O_415,N_19671,N_19983);
and UO_416 (O_416,N_19773,N_19641);
nand UO_417 (O_417,N_19889,N_19884);
nor UO_418 (O_418,N_19939,N_19750);
nor UO_419 (O_419,N_19627,N_19694);
xnor UO_420 (O_420,N_19714,N_19967);
xor UO_421 (O_421,N_19847,N_19926);
nand UO_422 (O_422,N_19613,N_19915);
nand UO_423 (O_423,N_19700,N_19781);
nor UO_424 (O_424,N_19679,N_19778);
nor UO_425 (O_425,N_19995,N_19758);
xnor UO_426 (O_426,N_19664,N_19860);
or UO_427 (O_427,N_19851,N_19745);
nand UO_428 (O_428,N_19999,N_19971);
nor UO_429 (O_429,N_19654,N_19890);
or UO_430 (O_430,N_19896,N_19716);
nor UO_431 (O_431,N_19770,N_19998);
or UO_432 (O_432,N_19750,N_19609);
xor UO_433 (O_433,N_19845,N_19846);
and UO_434 (O_434,N_19706,N_19688);
nand UO_435 (O_435,N_19840,N_19637);
or UO_436 (O_436,N_19607,N_19788);
or UO_437 (O_437,N_19927,N_19609);
nor UO_438 (O_438,N_19953,N_19980);
xor UO_439 (O_439,N_19880,N_19817);
and UO_440 (O_440,N_19936,N_19621);
nor UO_441 (O_441,N_19844,N_19825);
xor UO_442 (O_442,N_19976,N_19712);
or UO_443 (O_443,N_19608,N_19996);
and UO_444 (O_444,N_19671,N_19669);
xnor UO_445 (O_445,N_19797,N_19965);
and UO_446 (O_446,N_19890,N_19918);
and UO_447 (O_447,N_19626,N_19894);
and UO_448 (O_448,N_19644,N_19969);
nand UO_449 (O_449,N_19628,N_19790);
and UO_450 (O_450,N_19890,N_19802);
xnor UO_451 (O_451,N_19670,N_19734);
or UO_452 (O_452,N_19971,N_19931);
and UO_453 (O_453,N_19780,N_19796);
nand UO_454 (O_454,N_19631,N_19758);
nand UO_455 (O_455,N_19742,N_19989);
or UO_456 (O_456,N_19742,N_19775);
nand UO_457 (O_457,N_19893,N_19844);
nor UO_458 (O_458,N_19792,N_19647);
xnor UO_459 (O_459,N_19749,N_19680);
nor UO_460 (O_460,N_19649,N_19794);
nand UO_461 (O_461,N_19828,N_19830);
and UO_462 (O_462,N_19790,N_19714);
nand UO_463 (O_463,N_19786,N_19902);
or UO_464 (O_464,N_19831,N_19712);
xnor UO_465 (O_465,N_19743,N_19933);
nand UO_466 (O_466,N_19923,N_19815);
nand UO_467 (O_467,N_19956,N_19716);
nand UO_468 (O_468,N_19897,N_19718);
or UO_469 (O_469,N_19708,N_19729);
and UO_470 (O_470,N_19848,N_19806);
xor UO_471 (O_471,N_19916,N_19930);
nand UO_472 (O_472,N_19825,N_19924);
or UO_473 (O_473,N_19632,N_19604);
and UO_474 (O_474,N_19675,N_19658);
xnor UO_475 (O_475,N_19822,N_19730);
xor UO_476 (O_476,N_19845,N_19714);
and UO_477 (O_477,N_19967,N_19655);
or UO_478 (O_478,N_19930,N_19900);
or UO_479 (O_479,N_19747,N_19995);
nor UO_480 (O_480,N_19999,N_19687);
nand UO_481 (O_481,N_19741,N_19716);
nor UO_482 (O_482,N_19767,N_19943);
nor UO_483 (O_483,N_19826,N_19999);
nor UO_484 (O_484,N_19898,N_19654);
xnor UO_485 (O_485,N_19970,N_19849);
nand UO_486 (O_486,N_19882,N_19612);
nor UO_487 (O_487,N_19931,N_19896);
nor UO_488 (O_488,N_19658,N_19774);
or UO_489 (O_489,N_19987,N_19806);
nand UO_490 (O_490,N_19674,N_19907);
nand UO_491 (O_491,N_19602,N_19937);
nand UO_492 (O_492,N_19616,N_19867);
or UO_493 (O_493,N_19853,N_19738);
xor UO_494 (O_494,N_19926,N_19945);
and UO_495 (O_495,N_19812,N_19806);
nand UO_496 (O_496,N_19624,N_19941);
nor UO_497 (O_497,N_19650,N_19977);
nor UO_498 (O_498,N_19652,N_19986);
or UO_499 (O_499,N_19643,N_19722);
and UO_500 (O_500,N_19778,N_19688);
and UO_501 (O_501,N_19750,N_19739);
nor UO_502 (O_502,N_19626,N_19971);
nor UO_503 (O_503,N_19946,N_19668);
nand UO_504 (O_504,N_19982,N_19776);
xnor UO_505 (O_505,N_19745,N_19896);
nand UO_506 (O_506,N_19952,N_19860);
and UO_507 (O_507,N_19836,N_19633);
nor UO_508 (O_508,N_19891,N_19973);
or UO_509 (O_509,N_19977,N_19616);
nor UO_510 (O_510,N_19895,N_19709);
xnor UO_511 (O_511,N_19819,N_19912);
or UO_512 (O_512,N_19885,N_19912);
nor UO_513 (O_513,N_19814,N_19745);
or UO_514 (O_514,N_19669,N_19860);
or UO_515 (O_515,N_19977,N_19922);
or UO_516 (O_516,N_19624,N_19946);
nand UO_517 (O_517,N_19856,N_19846);
nor UO_518 (O_518,N_19803,N_19887);
or UO_519 (O_519,N_19694,N_19944);
or UO_520 (O_520,N_19899,N_19691);
nand UO_521 (O_521,N_19711,N_19789);
and UO_522 (O_522,N_19652,N_19611);
or UO_523 (O_523,N_19637,N_19925);
xnor UO_524 (O_524,N_19886,N_19696);
xor UO_525 (O_525,N_19888,N_19702);
nor UO_526 (O_526,N_19685,N_19673);
xnor UO_527 (O_527,N_19727,N_19639);
and UO_528 (O_528,N_19996,N_19650);
xor UO_529 (O_529,N_19701,N_19933);
or UO_530 (O_530,N_19878,N_19853);
nor UO_531 (O_531,N_19806,N_19822);
or UO_532 (O_532,N_19674,N_19745);
xnor UO_533 (O_533,N_19734,N_19993);
nand UO_534 (O_534,N_19883,N_19987);
or UO_535 (O_535,N_19945,N_19654);
xnor UO_536 (O_536,N_19662,N_19869);
and UO_537 (O_537,N_19831,N_19987);
nand UO_538 (O_538,N_19815,N_19830);
xnor UO_539 (O_539,N_19776,N_19677);
nor UO_540 (O_540,N_19834,N_19877);
and UO_541 (O_541,N_19682,N_19611);
xor UO_542 (O_542,N_19677,N_19637);
or UO_543 (O_543,N_19898,N_19715);
or UO_544 (O_544,N_19669,N_19767);
xor UO_545 (O_545,N_19719,N_19871);
nor UO_546 (O_546,N_19968,N_19677);
and UO_547 (O_547,N_19605,N_19974);
nor UO_548 (O_548,N_19856,N_19958);
nand UO_549 (O_549,N_19703,N_19761);
or UO_550 (O_550,N_19666,N_19628);
xor UO_551 (O_551,N_19651,N_19710);
nor UO_552 (O_552,N_19814,N_19897);
nor UO_553 (O_553,N_19990,N_19806);
and UO_554 (O_554,N_19860,N_19896);
xnor UO_555 (O_555,N_19739,N_19699);
nor UO_556 (O_556,N_19962,N_19997);
nand UO_557 (O_557,N_19895,N_19681);
and UO_558 (O_558,N_19820,N_19924);
nor UO_559 (O_559,N_19666,N_19658);
or UO_560 (O_560,N_19658,N_19881);
nand UO_561 (O_561,N_19749,N_19632);
or UO_562 (O_562,N_19903,N_19805);
nor UO_563 (O_563,N_19616,N_19730);
or UO_564 (O_564,N_19860,N_19949);
nand UO_565 (O_565,N_19780,N_19966);
nor UO_566 (O_566,N_19989,N_19630);
xor UO_567 (O_567,N_19702,N_19681);
or UO_568 (O_568,N_19894,N_19871);
xor UO_569 (O_569,N_19834,N_19843);
nor UO_570 (O_570,N_19933,N_19866);
nand UO_571 (O_571,N_19682,N_19827);
xnor UO_572 (O_572,N_19923,N_19945);
nand UO_573 (O_573,N_19826,N_19856);
or UO_574 (O_574,N_19956,N_19984);
nor UO_575 (O_575,N_19859,N_19917);
nand UO_576 (O_576,N_19647,N_19754);
or UO_577 (O_577,N_19951,N_19600);
xor UO_578 (O_578,N_19752,N_19693);
or UO_579 (O_579,N_19908,N_19937);
xor UO_580 (O_580,N_19941,N_19908);
nand UO_581 (O_581,N_19601,N_19929);
xor UO_582 (O_582,N_19674,N_19956);
xor UO_583 (O_583,N_19646,N_19833);
nor UO_584 (O_584,N_19953,N_19698);
nor UO_585 (O_585,N_19741,N_19631);
nand UO_586 (O_586,N_19969,N_19673);
or UO_587 (O_587,N_19632,N_19726);
nand UO_588 (O_588,N_19661,N_19977);
or UO_589 (O_589,N_19661,N_19645);
or UO_590 (O_590,N_19623,N_19859);
or UO_591 (O_591,N_19861,N_19667);
nand UO_592 (O_592,N_19911,N_19902);
or UO_593 (O_593,N_19899,N_19986);
or UO_594 (O_594,N_19747,N_19890);
nor UO_595 (O_595,N_19950,N_19940);
xnor UO_596 (O_596,N_19656,N_19879);
or UO_597 (O_597,N_19834,N_19689);
nor UO_598 (O_598,N_19767,N_19652);
xnor UO_599 (O_599,N_19815,N_19795);
and UO_600 (O_600,N_19799,N_19765);
or UO_601 (O_601,N_19713,N_19653);
nand UO_602 (O_602,N_19862,N_19731);
or UO_603 (O_603,N_19912,N_19880);
xor UO_604 (O_604,N_19924,N_19823);
xor UO_605 (O_605,N_19743,N_19987);
xor UO_606 (O_606,N_19821,N_19970);
nor UO_607 (O_607,N_19706,N_19787);
nor UO_608 (O_608,N_19685,N_19727);
and UO_609 (O_609,N_19761,N_19692);
xor UO_610 (O_610,N_19812,N_19689);
nor UO_611 (O_611,N_19601,N_19689);
nor UO_612 (O_612,N_19676,N_19997);
nand UO_613 (O_613,N_19636,N_19899);
or UO_614 (O_614,N_19936,N_19695);
nand UO_615 (O_615,N_19947,N_19753);
nor UO_616 (O_616,N_19784,N_19913);
nand UO_617 (O_617,N_19868,N_19857);
and UO_618 (O_618,N_19705,N_19852);
nand UO_619 (O_619,N_19751,N_19759);
and UO_620 (O_620,N_19794,N_19680);
nor UO_621 (O_621,N_19726,N_19750);
nor UO_622 (O_622,N_19978,N_19850);
nand UO_623 (O_623,N_19633,N_19841);
or UO_624 (O_624,N_19995,N_19656);
nand UO_625 (O_625,N_19872,N_19612);
xnor UO_626 (O_626,N_19677,N_19745);
xnor UO_627 (O_627,N_19909,N_19639);
xor UO_628 (O_628,N_19811,N_19788);
or UO_629 (O_629,N_19637,N_19857);
and UO_630 (O_630,N_19913,N_19651);
or UO_631 (O_631,N_19605,N_19896);
nor UO_632 (O_632,N_19831,N_19912);
or UO_633 (O_633,N_19762,N_19897);
xnor UO_634 (O_634,N_19997,N_19630);
and UO_635 (O_635,N_19786,N_19626);
xnor UO_636 (O_636,N_19974,N_19845);
xor UO_637 (O_637,N_19977,N_19871);
nand UO_638 (O_638,N_19853,N_19611);
and UO_639 (O_639,N_19634,N_19755);
or UO_640 (O_640,N_19616,N_19967);
nand UO_641 (O_641,N_19725,N_19967);
nor UO_642 (O_642,N_19733,N_19965);
xor UO_643 (O_643,N_19892,N_19878);
xnor UO_644 (O_644,N_19665,N_19655);
xnor UO_645 (O_645,N_19659,N_19648);
and UO_646 (O_646,N_19746,N_19604);
and UO_647 (O_647,N_19885,N_19816);
nor UO_648 (O_648,N_19932,N_19980);
xor UO_649 (O_649,N_19608,N_19607);
and UO_650 (O_650,N_19708,N_19780);
or UO_651 (O_651,N_19773,N_19997);
xnor UO_652 (O_652,N_19713,N_19718);
xnor UO_653 (O_653,N_19960,N_19844);
nand UO_654 (O_654,N_19606,N_19835);
nand UO_655 (O_655,N_19907,N_19899);
or UO_656 (O_656,N_19833,N_19686);
or UO_657 (O_657,N_19750,N_19984);
and UO_658 (O_658,N_19808,N_19695);
xor UO_659 (O_659,N_19748,N_19953);
or UO_660 (O_660,N_19959,N_19982);
nor UO_661 (O_661,N_19790,N_19689);
nor UO_662 (O_662,N_19730,N_19894);
and UO_663 (O_663,N_19759,N_19937);
and UO_664 (O_664,N_19761,N_19649);
or UO_665 (O_665,N_19988,N_19949);
nor UO_666 (O_666,N_19737,N_19685);
or UO_667 (O_667,N_19702,N_19959);
and UO_668 (O_668,N_19609,N_19804);
nand UO_669 (O_669,N_19817,N_19621);
and UO_670 (O_670,N_19743,N_19993);
and UO_671 (O_671,N_19755,N_19826);
nand UO_672 (O_672,N_19645,N_19868);
or UO_673 (O_673,N_19617,N_19811);
or UO_674 (O_674,N_19800,N_19860);
nand UO_675 (O_675,N_19849,N_19705);
xnor UO_676 (O_676,N_19906,N_19728);
or UO_677 (O_677,N_19600,N_19930);
nor UO_678 (O_678,N_19770,N_19747);
or UO_679 (O_679,N_19798,N_19996);
nand UO_680 (O_680,N_19738,N_19983);
nor UO_681 (O_681,N_19668,N_19739);
and UO_682 (O_682,N_19791,N_19774);
nor UO_683 (O_683,N_19946,N_19666);
or UO_684 (O_684,N_19859,N_19601);
or UO_685 (O_685,N_19835,N_19757);
or UO_686 (O_686,N_19948,N_19885);
or UO_687 (O_687,N_19752,N_19623);
nor UO_688 (O_688,N_19751,N_19820);
nor UO_689 (O_689,N_19630,N_19839);
nor UO_690 (O_690,N_19977,N_19960);
and UO_691 (O_691,N_19809,N_19794);
nor UO_692 (O_692,N_19925,N_19814);
and UO_693 (O_693,N_19995,N_19895);
nand UO_694 (O_694,N_19841,N_19605);
and UO_695 (O_695,N_19860,N_19666);
xnor UO_696 (O_696,N_19610,N_19917);
or UO_697 (O_697,N_19603,N_19673);
or UO_698 (O_698,N_19994,N_19702);
nand UO_699 (O_699,N_19840,N_19739);
xor UO_700 (O_700,N_19706,N_19980);
nand UO_701 (O_701,N_19717,N_19857);
or UO_702 (O_702,N_19652,N_19860);
nor UO_703 (O_703,N_19939,N_19715);
and UO_704 (O_704,N_19844,N_19848);
or UO_705 (O_705,N_19985,N_19645);
nand UO_706 (O_706,N_19777,N_19933);
or UO_707 (O_707,N_19672,N_19760);
xor UO_708 (O_708,N_19912,N_19629);
nand UO_709 (O_709,N_19963,N_19894);
nand UO_710 (O_710,N_19948,N_19695);
xor UO_711 (O_711,N_19994,N_19603);
nand UO_712 (O_712,N_19744,N_19736);
and UO_713 (O_713,N_19809,N_19897);
nor UO_714 (O_714,N_19782,N_19938);
xor UO_715 (O_715,N_19826,N_19883);
or UO_716 (O_716,N_19666,N_19973);
and UO_717 (O_717,N_19767,N_19955);
nor UO_718 (O_718,N_19725,N_19845);
nand UO_719 (O_719,N_19983,N_19873);
nand UO_720 (O_720,N_19816,N_19951);
xor UO_721 (O_721,N_19781,N_19787);
and UO_722 (O_722,N_19959,N_19777);
nand UO_723 (O_723,N_19672,N_19970);
nor UO_724 (O_724,N_19911,N_19863);
and UO_725 (O_725,N_19731,N_19686);
nor UO_726 (O_726,N_19713,N_19627);
and UO_727 (O_727,N_19908,N_19753);
nand UO_728 (O_728,N_19903,N_19669);
nand UO_729 (O_729,N_19810,N_19749);
nor UO_730 (O_730,N_19886,N_19650);
and UO_731 (O_731,N_19800,N_19856);
nor UO_732 (O_732,N_19849,N_19695);
or UO_733 (O_733,N_19773,N_19606);
and UO_734 (O_734,N_19930,N_19606);
nand UO_735 (O_735,N_19741,N_19858);
xnor UO_736 (O_736,N_19764,N_19624);
nor UO_737 (O_737,N_19631,N_19867);
xnor UO_738 (O_738,N_19989,N_19730);
or UO_739 (O_739,N_19720,N_19986);
nand UO_740 (O_740,N_19635,N_19971);
xor UO_741 (O_741,N_19777,N_19839);
xor UO_742 (O_742,N_19737,N_19881);
and UO_743 (O_743,N_19751,N_19980);
or UO_744 (O_744,N_19667,N_19853);
nor UO_745 (O_745,N_19723,N_19788);
nand UO_746 (O_746,N_19908,N_19730);
nor UO_747 (O_747,N_19864,N_19937);
nand UO_748 (O_748,N_19929,N_19663);
or UO_749 (O_749,N_19863,N_19877);
nand UO_750 (O_750,N_19648,N_19951);
xor UO_751 (O_751,N_19790,N_19797);
xnor UO_752 (O_752,N_19935,N_19852);
nand UO_753 (O_753,N_19647,N_19683);
xnor UO_754 (O_754,N_19687,N_19664);
and UO_755 (O_755,N_19642,N_19998);
nor UO_756 (O_756,N_19911,N_19912);
nor UO_757 (O_757,N_19990,N_19669);
xnor UO_758 (O_758,N_19840,N_19924);
and UO_759 (O_759,N_19780,N_19784);
xnor UO_760 (O_760,N_19857,N_19753);
xnor UO_761 (O_761,N_19781,N_19871);
nand UO_762 (O_762,N_19634,N_19877);
xor UO_763 (O_763,N_19612,N_19873);
nor UO_764 (O_764,N_19600,N_19808);
or UO_765 (O_765,N_19620,N_19704);
nand UO_766 (O_766,N_19931,N_19928);
or UO_767 (O_767,N_19692,N_19976);
xnor UO_768 (O_768,N_19826,N_19854);
or UO_769 (O_769,N_19968,N_19779);
or UO_770 (O_770,N_19771,N_19796);
or UO_771 (O_771,N_19866,N_19817);
nor UO_772 (O_772,N_19644,N_19813);
nor UO_773 (O_773,N_19616,N_19964);
and UO_774 (O_774,N_19832,N_19989);
or UO_775 (O_775,N_19977,N_19685);
nand UO_776 (O_776,N_19812,N_19809);
xor UO_777 (O_777,N_19883,N_19905);
xnor UO_778 (O_778,N_19757,N_19795);
nor UO_779 (O_779,N_19733,N_19844);
nor UO_780 (O_780,N_19734,N_19673);
nand UO_781 (O_781,N_19961,N_19906);
nand UO_782 (O_782,N_19639,N_19759);
nor UO_783 (O_783,N_19962,N_19694);
or UO_784 (O_784,N_19873,N_19609);
and UO_785 (O_785,N_19765,N_19740);
or UO_786 (O_786,N_19748,N_19639);
and UO_787 (O_787,N_19992,N_19632);
xor UO_788 (O_788,N_19994,N_19710);
xor UO_789 (O_789,N_19885,N_19750);
nand UO_790 (O_790,N_19866,N_19878);
nor UO_791 (O_791,N_19857,N_19745);
or UO_792 (O_792,N_19753,N_19892);
nand UO_793 (O_793,N_19677,N_19932);
nand UO_794 (O_794,N_19929,N_19604);
nor UO_795 (O_795,N_19808,N_19844);
nand UO_796 (O_796,N_19681,N_19795);
nor UO_797 (O_797,N_19743,N_19915);
nor UO_798 (O_798,N_19759,N_19672);
nand UO_799 (O_799,N_19770,N_19713);
nor UO_800 (O_800,N_19741,N_19952);
xnor UO_801 (O_801,N_19669,N_19920);
nand UO_802 (O_802,N_19987,N_19788);
or UO_803 (O_803,N_19813,N_19695);
nor UO_804 (O_804,N_19931,N_19992);
and UO_805 (O_805,N_19612,N_19614);
nand UO_806 (O_806,N_19837,N_19607);
nor UO_807 (O_807,N_19955,N_19877);
xor UO_808 (O_808,N_19874,N_19693);
or UO_809 (O_809,N_19792,N_19815);
or UO_810 (O_810,N_19920,N_19972);
or UO_811 (O_811,N_19945,N_19830);
xor UO_812 (O_812,N_19713,N_19753);
xnor UO_813 (O_813,N_19939,N_19978);
nor UO_814 (O_814,N_19932,N_19624);
and UO_815 (O_815,N_19801,N_19746);
and UO_816 (O_816,N_19638,N_19908);
and UO_817 (O_817,N_19964,N_19787);
and UO_818 (O_818,N_19623,N_19643);
xnor UO_819 (O_819,N_19612,N_19743);
nand UO_820 (O_820,N_19947,N_19667);
and UO_821 (O_821,N_19981,N_19752);
and UO_822 (O_822,N_19673,N_19694);
nor UO_823 (O_823,N_19626,N_19898);
nand UO_824 (O_824,N_19683,N_19869);
xnor UO_825 (O_825,N_19683,N_19994);
nor UO_826 (O_826,N_19974,N_19999);
nand UO_827 (O_827,N_19605,N_19739);
nand UO_828 (O_828,N_19920,N_19874);
xnor UO_829 (O_829,N_19796,N_19660);
xnor UO_830 (O_830,N_19895,N_19751);
xnor UO_831 (O_831,N_19828,N_19647);
and UO_832 (O_832,N_19648,N_19756);
nand UO_833 (O_833,N_19807,N_19779);
xnor UO_834 (O_834,N_19883,N_19739);
xor UO_835 (O_835,N_19779,N_19766);
and UO_836 (O_836,N_19810,N_19795);
and UO_837 (O_837,N_19647,N_19760);
xnor UO_838 (O_838,N_19973,N_19653);
and UO_839 (O_839,N_19817,N_19944);
and UO_840 (O_840,N_19940,N_19653);
nand UO_841 (O_841,N_19846,N_19743);
and UO_842 (O_842,N_19960,N_19893);
and UO_843 (O_843,N_19624,N_19780);
nand UO_844 (O_844,N_19720,N_19823);
nand UO_845 (O_845,N_19858,N_19946);
and UO_846 (O_846,N_19626,N_19885);
xor UO_847 (O_847,N_19847,N_19806);
nor UO_848 (O_848,N_19722,N_19654);
xor UO_849 (O_849,N_19729,N_19604);
xnor UO_850 (O_850,N_19736,N_19894);
xor UO_851 (O_851,N_19695,N_19737);
xnor UO_852 (O_852,N_19857,N_19843);
nor UO_853 (O_853,N_19726,N_19890);
xor UO_854 (O_854,N_19995,N_19892);
xor UO_855 (O_855,N_19976,N_19758);
and UO_856 (O_856,N_19714,N_19994);
and UO_857 (O_857,N_19802,N_19738);
nand UO_858 (O_858,N_19790,N_19932);
nand UO_859 (O_859,N_19900,N_19998);
nand UO_860 (O_860,N_19708,N_19781);
or UO_861 (O_861,N_19863,N_19837);
xnor UO_862 (O_862,N_19826,N_19940);
xor UO_863 (O_863,N_19676,N_19796);
nand UO_864 (O_864,N_19625,N_19852);
nor UO_865 (O_865,N_19769,N_19858);
nor UO_866 (O_866,N_19976,N_19784);
or UO_867 (O_867,N_19937,N_19943);
nand UO_868 (O_868,N_19733,N_19688);
nor UO_869 (O_869,N_19693,N_19801);
xnor UO_870 (O_870,N_19945,N_19910);
nand UO_871 (O_871,N_19975,N_19685);
or UO_872 (O_872,N_19795,N_19802);
nand UO_873 (O_873,N_19975,N_19658);
nand UO_874 (O_874,N_19986,N_19797);
and UO_875 (O_875,N_19846,N_19636);
or UO_876 (O_876,N_19920,N_19815);
nand UO_877 (O_877,N_19755,N_19886);
and UO_878 (O_878,N_19980,N_19938);
nor UO_879 (O_879,N_19944,N_19993);
nor UO_880 (O_880,N_19788,N_19972);
xnor UO_881 (O_881,N_19630,N_19982);
nand UO_882 (O_882,N_19906,N_19749);
or UO_883 (O_883,N_19861,N_19756);
xor UO_884 (O_884,N_19843,N_19944);
nor UO_885 (O_885,N_19686,N_19740);
xnor UO_886 (O_886,N_19848,N_19940);
nand UO_887 (O_887,N_19656,N_19669);
and UO_888 (O_888,N_19730,N_19719);
or UO_889 (O_889,N_19776,N_19759);
and UO_890 (O_890,N_19854,N_19636);
nand UO_891 (O_891,N_19996,N_19616);
and UO_892 (O_892,N_19755,N_19767);
xor UO_893 (O_893,N_19647,N_19952);
xnor UO_894 (O_894,N_19935,N_19818);
xor UO_895 (O_895,N_19720,N_19916);
or UO_896 (O_896,N_19948,N_19792);
and UO_897 (O_897,N_19866,N_19627);
nand UO_898 (O_898,N_19609,N_19714);
nand UO_899 (O_899,N_19966,N_19934);
nor UO_900 (O_900,N_19783,N_19954);
nor UO_901 (O_901,N_19752,N_19740);
nand UO_902 (O_902,N_19611,N_19721);
or UO_903 (O_903,N_19962,N_19944);
or UO_904 (O_904,N_19746,N_19943);
nor UO_905 (O_905,N_19932,N_19815);
and UO_906 (O_906,N_19641,N_19634);
nor UO_907 (O_907,N_19944,N_19750);
nand UO_908 (O_908,N_19770,N_19775);
or UO_909 (O_909,N_19656,N_19673);
xnor UO_910 (O_910,N_19630,N_19715);
nand UO_911 (O_911,N_19717,N_19983);
nor UO_912 (O_912,N_19629,N_19647);
or UO_913 (O_913,N_19996,N_19970);
and UO_914 (O_914,N_19851,N_19973);
or UO_915 (O_915,N_19857,N_19628);
xnor UO_916 (O_916,N_19808,N_19716);
xor UO_917 (O_917,N_19692,N_19963);
nor UO_918 (O_918,N_19809,N_19995);
and UO_919 (O_919,N_19791,N_19968);
xor UO_920 (O_920,N_19635,N_19692);
nor UO_921 (O_921,N_19708,N_19785);
and UO_922 (O_922,N_19831,N_19676);
or UO_923 (O_923,N_19723,N_19812);
or UO_924 (O_924,N_19809,N_19603);
nand UO_925 (O_925,N_19894,N_19962);
xor UO_926 (O_926,N_19640,N_19903);
xor UO_927 (O_927,N_19895,N_19937);
xor UO_928 (O_928,N_19748,N_19933);
nand UO_929 (O_929,N_19681,N_19778);
or UO_930 (O_930,N_19731,N_19924);
or UO_931 (O_931,N_19795,N_19989);
nor UO_932 (O_932,N_19703,N_19937);
nor UO_933 (O_933,N_19938,N_19868);
xor UO_934 (O_934,N_19811,N_19688);
or UO_935 (O_935,N_19759,N_19818);
and UO_936 (O_936,N_19839,N_19800);
and UO_937 (O_937,N_19652,N_19742);
or UO_938 (O_938,N_19931,N_19875);
nor UO_939 (O_939,N_19750,N_19745);
or UO_940 (O_940,N_19607,N_19953);
nand UO_941 (O_941,N_19773,N_19850);
nor UO_942 (O_942,N_19975,N_19855);
or UO_943 (O_943,N_19678,N_19947);
xnor UO_944 (O_944,N_19760,N_19615);
or UO_945 (O_945,N_19772,N_19854);
xnor UO_946 (O_946,N_19787,N_19854);
and UO_947 (O_947,N_19953,N_19829);
nand UO_948 (O_948,N_19852,N_19813);
and UO_949 (O_949,N_19879,N_19688);
and UO_950 (O_950,N_19638,N_19680);
xor UO_951 (O_951,N_19854,N_19632);
xor UO_952 (O_952,N_19933,N_19758);
and UO_953 (O_953,N_19872,N_19819);
nor UO_954 (O_954,N_19659,N_19863);
nand UO_955 (O_955,N_19836,N_19603);
or UO_956 (O_956,N_19699,N_19888);
nor UO_957 (O_957,N_19921,N_19885);
xor UO_958 (O_958,N_19733,N_19914);
xnor UO_959 (O_959,N_19614,N_19790);
xnor UO_960 (O_960,N_19744,N_19729);
or UO_961 (O_961,N_19717,N_19611);
and UO_962 (O_962,N_19709,N_19918);
nand UO_963 (O_963,N_19763,N_19617);
or UO_964 (O_964,N_19872,N_19682);
nor UO_965 (O_965,N_19632,N_19973);
nor UO_966 (O_966,N_19815,N_19878);
and UO_967 (O_967,N_19873,N_19947);
and UO_968 (O_968,N_19859,N_19753);
nor UO_969 (O_969,N_19621,N_19867);
nor UO_970 (O_970,N_19629,N_19997);
and UO_971 (O_971,N_19608,N_19945);
xnor UO_972 (O_972,N_19880,N_19653);
and UO_973 (O_973,N_19902,N_19755);
xnor UO_974 (O_974,N_19733,N_19780);
xnor UO_975 (O_975,N_19821,N_19932);
xnor UO_976 (O_976,N_19691,N_19644);
nor UO_977 (O_977,N_19639,N_19764);
nor UO_978 (O_978,N_19918,N_19623);
xor UO_979 (O_979,N_19767,N_19997);
or UO_980 (O_980,N_19792,N_19657);
or UO_981 (O_981,N_19988,N_19617);
nand UO_982 (O_982,N_19693,N_19848);
and UO_983 (O_983,N_19994,N_19633);
nand UO_984 (O_984,N_19611,N_19775);
nand UO_985 (O_985,N_19627,N_19767);
xor UO_986 (O_986,N_19656,N_19836);
and UO_987 (O_987,N_19788,N_19897);
or UO_988 (O_988,N_19755,N_19951);
nor UO_989 (O_989,N_19873,N_19729);
xnor UO_990 (O_990,N_19746,N_19753);
nor UO_991 (O_991,N_19658,N_19718);
nand UO_992 (O_992,N_19718,N_19926);
xor UO_993 (O_993,N_19694,N_19773);
nand UO_994 (O_994,N_19872,N_19681);
xnor UO_995 (O_995,N_19870,N_19950);
and UO_996 (O_996,N_19836,N_19773);
or UO_997 (O_997,N_19792,N_19718);
xor UO_998 (O_998,N_19631,N_19819);
xnor UO_999 (O_999,N_19923,N_19807);
nor UO_1000 (O_1000,N_19673,N_19742);
nand UO_1001 (O_1001,N_19849,N_19640);
nor UO_1002 (O_1002,N_19748,N_19864);
or UO_1003 (O_1003,N_19697,N_19728);
or UO_1004 (O_1004,N_19618,N_19726);
nand UO_1005 (O_1005,N_19886,N_19940);
nand UO_1006 (O_1006,N_19951,N_19823);
xnor UO_1007 (O_1007,N_19761,N_19758);
nand UO_1008 (O_1008,N_19754,N_19665);
or UO_1009 (O_1009,N_19996,N_19818);
nand UO_1010 (O_1010,N_19671,N_19993);
and UO_1011 (O_1011,N_19742,N_19643);
nor UO_1012 (O_1012,N_19798,N_19685);
xor UO_1013 (O_1013,N_19908,N_19907);
nand UO_1014 (O_1014,N_19990,N_19735);
nand UO_1015 (O_1015,N_19629,N_19746);
nor UO_1016 (O_1016,N_19772,N_19838);
xor UO_1017 (O_1017,N_19850,N_19976);
nand UO_1018 (O_1018,N_19655,N_19822);
and UO_1019 (O_1019,N_19991,N_19632);
and UO_1020 (O_1020,N_19809,N_19817);
nor UO_1021 (O_1021,N_19960,N_19668);
nand UO_1022 (O_1022,N_19938,N_19617);
nand UO_1023 (O_1023,N_19897,N_19918);
xnor UO_1024 (O_1024,N_19810,N_19732);
xor UO_1025 (O_1025,N_19849,N_19871);
nand UO_1026 (O_1026,N_19601,N_19622);
nand UO_1027 (O_1027,N_19691,N_19938);
nand UO_1028 (O_1028,N_19758,N_19741);
nor UO_1029 (O_1029,N_19836,N_19988);
nor UO_1030 (O_1030,N_19980,N_19746);
nand UO_1031 (O_1031,N_19994,N_19826);
or UO_1032 (O_1032,N_19934,N_19992);
xor UO_1033 (O_1033,N_19689,N_19690);
nand UO_1034 (O_1034,N_19808,N_19769);
nand UO_1035 (O_1035,N_19867,N_19685);
nor UO_1036 (O_1036,N_19995,N_19648);
and UO_1037 (O_1037,N_19828,N_19987);
xnor UO_1038 (O_1038,N_19690,N_19746);
xnor UO_1039 (O_1039,N_19753,N_19686);
nand UO_1040 (O_1040,N_19878,N_19903);
and UO_1041 (O_1041,N_19741,N_19738);
xnor UO_1042 (O_1042,N_19932,N_19755);
or UO_1043 (O_1043,N_19717,N_19757);
xor UO_1044 (O_1044,N_19723,N_19971);
nand UO_1045 (O_1045,N_19829,N_19905);
and UO_1046 (O_1046,N_19707,N_19662);
xor UO_1047 (O_1047,N_19631,N_19659);
nor UO_1048 (O_1048,N_19700,N_19949);
xor UO_1049 (O_1049,N_19766,N_19761);
or UO_1050 (O_1050,N_19756,N_19761);
or UO_1051 (O_1051,N_19632,N_19936);
nor UO_1052 (O_1052,N_19609,N_19735);
and UO_1053 (O_1053,N_19838,N_19980);
and UO_1054 (O_1054,N_19899,N_19841);
nor UO_1055 (O_1055,N_19958,N_19620);
or UO_1056 (O_1056,N_19761,N_19850);
or UO_1057 (O_1057,N_19735,N_19673);
nor UO_1058 (O_1058,N_19694,N_19762);
and UO_1059 (O_1059,N_19652,N_19806);
nand UO_1060 (O_1060,N_19772,N_19924);
xor UO_1061 (O_1061,N_19684,N_19933);
or UO_1062 (O_1062,N_19826,N_19730);
or UO_1063 (O_1063,N_19694,N_19609);
and UO_1064 (O_1064,N_19657,N_19691);
nor UO_1065 (O_1065,N_19622,N_19785);
and UO_1066 (O_1066,N_19823,N_19631);
nand UO_1067 (O_1067,N_19759,N_19939);
and UO_1068 (O_1068,N_19776,N_19941);
nand UO_1069 (O_1069,N_19847,N_19749);
xor UO_1070 (O_1070,N_19885,N_19623);
xor UO_1071 (O_1071,N_19957,N_19775);
xnor UO_1072 (O_1072,N_19961,N_19932);
nor UO_1073 (O_1073,N_19662,N_19872);
xnor UO_1074 (O_1074,N_19824,N_19851);
nand UO_1075 (O_1075,N_19874,N_19937);
xnor UO_1076 (O_1076,N_19626,N_19707);
and UO_1077 (O_1077,N_19894,N_19896);
or UO_1078 (O_1078,N_19716,N_19753);
xnor UO_1079 (O_1079,N_19947,N_19844);
nor UO_1080 (O_1080,N_19706,N_19672);
nand UO_1081 (O_1081,N_19701,N_19861);
nand UO_1082 (O_1082,N_19801,N_19807);
and UO_1083 (O_1083,N_19994,N_19805);
and UO_1084 (O_1084,N_19715,N_19997);
nor UO_1085 (O_1085,N_19776,N_19665);
xor UO_1086 (O_1086,N_19669,N_19664);
nand UO_1087 (O_1087,N_19689,N_19797);
nand UO_1088 (O_1088,N_19993,N_19921);
and UO_1089 (O_1089,N_19907,N_19927);
and UO_1090 (O_1090,N_19955,N_19934);
or UO_1091 (O_1091,N_19747,N_19834);
nand UO_1092 (O_1092,N_19834,N_19768);
and UO_1093 (O_1093,N_19886,N_19667);
or UO_1094 (O_1094,N_19861,N_19738);
nor UO_1095 (O_1095,N_19654,N_19925);
and UO_1096 (O_1096,N_19999,N_19758);
nor UO_1097 (O_1097,N_19660,N_19626);
nor UO_1098 (O_1098,N_19921,N_19835);
nand UO_1099 (O_1099,N_19852,N_19919);
nand UO_1100 (O_1100,N_19987,N_19692);
nor UO_1101 (O_1101,N_19698,N_19736);
xor UO_1102 (O_1102,N_19962,N_19927);
nand UO_1103 (O_1103,N_19992,N_19936);
and UO_1104 (O_1104,N_19817,N_19713);
nor UO_1105 (O_1105,N_19933,N_19685);
and UO_1106 (O_1106,N_19928,N_19689);
nor UO_1107 (O_1107,N_19703,N_19897);
or UO_1108 (O_1108,N_19660,N_19920);
xnor UO_1109 (O_1109,N_19636,N_19855);
and UO_1110 (O_1110,N_19955,N_19843);
xnor UO_1111 (O_1111,N_19758,N_19885);
or UO_1112 (O_1112,N_19938,N_19924);
nor UO_1113 (O_1113,N_19818,N_19863);
nand UO_1114 (O_1114,N_19616,N_19896);
or UO_1115 (O_1115,N_19892,N_19974);
nor UO_1116 (O_1116,N_19633,N_19612);
nor UO_1117 (O_1117,N_19980,N_19697);
nor UO_1118 (O_1118,N_19953,N_19808);
and UO_1119 (O_1119,N_19840,N_19941);
and UO_1120 (O_1120,N_19698,N_19982);
or UO_1121 (O_1121,N_19908,N_19916);
or UO_1122 (O_1122,N_19794,N_19711);
xor UO_1123 (O_1123,N_19657,N_19957);
nand UO_1124 (O_1124,N_19998,N_19992);
and UO_1125 (O_1125,N_19975,N_19698);
nor UO_1126 (O_1126,N_19799,N_19976);
nand UO_1127 (O_1127,N_19714,N_19610);
nor UO_1128 (O_1128,N_19641,N_19646);
or UO_1129 (O_1129,N_19847,N_19971);
and UO_1130 (O_1130,N_19679,N_19863);
and UO_1131 (O_1131,N_19824,N_19807);
nor UO_1132 (O_1132,N_19697,N_19950);
and UO_1133 (O_1133,N_19688,N_19793);
or UO_1134 (O_1134,N_19809,N_19841);
and UO_1135 (O_1135,N_19949,N_19849);
and UO_1136 (O_1136,N_19756,N_19726);
xor UO_1137 (O_1137,N_19947,N_19600);
nor UO_1138 (O_1138,N_19921,N_19861);
xor UO_1139 (O_1139,N_19767,N_19913);
nor UO_1140 (O_1140,N_19801,N_19803);
or UO_1141 (O_1141,N_19711,N_19983);
and UO_1142 (O_1142,N_19726,N_19733);
and UO_1143 (O_1143,N_19784,N_19642);
or UO_1144 (O_1144,N_19742,N_19777);
nor UO_1145 (O_1145,N_19682,N_19989);
nand UO_1146 (O_1146,N_19601,N_19628);
nor UO_1147 (O_1147,N_19865,N_19854);
xnor UO_1148 (O_1148,N_19962,N_19732);
nor UO_1149 (O_1149,N_19722,N_19904);
or UO_1150 (O_1150,N_19934,N_19675);
nor UO_1151 (O_1151,N_19791,N_19891);
and UO_1152 (O_1152,N_19887,N_19770);
or UO_1153 (O_1153,N_19850,N_19816);
xor UO_1154 (O_1154,N_19902,N_19821);
and UO_1155 (O_1155,N_19724,N_19783);
nand UO_1156 (O_1156,N_19676,N_19722);
xor UO_1157 (O_1157,N_19792,N_19852);
or UO_1158 (O_1158,N_19688,N_19947);
xor UO_1159 (O_1159,N_19731,N_19616);
nand UO_1160 (O_1160,N_19893,N_19766);
xnor UO_1161 (O_1161,N_19875,N_19910);
and UO_1162 (O_1162,N_19763,N_19606);
or UO_1163 (O_1163,N_19840,N_19725);
xor UO_1164 (O_1164,N_19877,N_19971);
nor UO_1165 (O_1165,N_19768,N_19654);
nor UO_1166 (O_1166,N_19639,N_19691);
and UO_1167 (O_1167,N_19957,N_19995);
nor UO_1168 (O_1168,N_19667,N_19677);
nand UO_1169 (O_1169,N_19770,N_19992);
nor UO_1170 (O_1170,N_19958,N_19606);
or UO_1171 (O_1171,N_19992,N_19670);
xnor UO_1172 (O_1172,N_19830,N_19776);
xnor UO_1173 (O_1173,N_19717,N_19620);
xor UO_1174 (O_1174,N_19666,N_19807);
xnor UO_1175 (O_1175,N_19701,N_19696);
nor UO_1176 (O_1176,N_19671,N_19705);
and UO_1177 (O_1177,N_19739,N_19687);
xnor UO_1178 (O_1178,N_19864,N_19711);
nand UO_1179 (O_1179,N_19705,N_19945);
xnor UO_1180 (O_1180,N_19843,N_19923);
xnor UO_1181 (O_1181,N_19703,N_19624);
and UO_1182 (O_1182,N_19932,N_19736);
nor UO_1183 (O_1183,N_19702,N_19826);
nor UO_1184 (O_1184,N_19857,N_19619);
and UO_1185 (O_1185,N_19732,N_19682);
nor UO_1186 (O_1186,N_19883,N_19980);
xor UO_1187 (O_1187,N_19883,N_19715);
or UO_1188 (O_1188,N_19738,N_19947);
nor UO_1189 (O_1189,N_19918,N_19811);
or UO_1190 (O_1190,N_19776,N_19757);
nand UO_1191 (O_1191,N_19731,N_19997);
nand UO_1192 (O_1192,N_19926,N_19636);
nand UO_1193 (O_1193,N_19655,N_19871);
nand UO_1194 (O_1194,N_19917,N_19984);
nor UO_1195 (O_1195,N_19705,N_19976);
and UO_1196 (O_1196,N_19604,N_19888);
and UO_1197 (O_1197,N_19691,N_19752);
nand UO_1198 (O_1198,N_19695,N_19898);
nand UO_1199 (O_1199,N_19955,N_19845);
and UO_1200 (O_1200,N_19722,N_19601);
xnor UO_1201 (O_1201,N_19600,N_19901);
nand UO_1202 (O_1202,N_19937,N_19729);
or UO_1203 (O_1203,N_19832,N_19947);
xor UO_1204 (O_1204,N_19625,N_19816);
nor UO_1205 (O_1205,N_19701,N_19813);
xnor UO_1206 (O_1206,N_19738,N_19692);
and UO_1207 (O_1207,N_19752,N_19625);
or UO_1208 (O_1208,N_19976,N_19871);
nand UO_1209 (O_1209,N_19923,N_19893);
xor UO_1210 (O_1210,N_19623,N_19651);
nor UO_1211 (O_1211,N_19615,N_19627);
and UO_1212 (O_1212,N_19994,N_19920);
nand UO_1213 (O_1213,N_19755,N_19638);
and UO_1214 (O_1214,N_19925,N_19949);
nand UO_1215 (O_1215,N_19886,N_19926);
or UO_1216 (O_1216,N_19704,N_19622);
or UO_1217 (O_1217,N_19610,N_19786);
xor UO_1218 (O_1218,N_19796,N_19971);
and UO_1219 (O_1219,N_19693,N_19989);
and UO_1220 (O_1220,N_19844,N_19784);
nand UO_1221 (O_1221,N_19713,N_19939);
and UO_1222 (O_1222,N_19967,N_19723);
or UO_1223 (O_1223,N_19707,N_19806);
nand UO_1224 (O_1224,N_19778,N_19648);
xor UO_1225 (O_1225,N_19673,N_19805);
nand UO_1226 (O_1226,N_19696,N_19800);
nand UO_1227 (O_1227,N_19615,N_19883);
or UO_1228 (O_1228,N_19843,N_19659);
nand UO_1229 (O_1229,N_19824,N_19829);
and UO_1230 (O_1230,N_19814,N_19899);
or UO_1231 (O_1231,N_19903,N_19981);
xnor UO_1232 (O_1232,N_19768,N_19790);
nor UO_1233 (O_1233,N_19799,N_19767);
nor UO_1234 (O_1234,N_19811,N_19880);
nor UO_1235 (O_1235,N_19913,N_19735);
nor UO_1236 (O_1236,N_19612,N_19761);
or UO_1237 (O_1237,N_19802,N_19618);
and UO_1238 (O_1238,N_19828,N_19923);
xnor UO_1239 (O_1239,N_19844,N_19609);
nor UO_1240 (O_1240,N_19875,N_19798);
nor UO_1241 (O_1241,N_19649,N_19784);
and UO_1242 (O_1242,N_19787,N_19698);
nor UO_1243 (O_1243,N_19884,N_19932);
xnor UO_1244 (O_1244,N_19779,N_19990);
nand UO_1245 (O_1245,N_19710,N_19658);
and UO_1246 (O_1246,N_19866,N_19823);
nor UO_1247 (O_1247,N_19861,N_19725);
nand UO_1248 (O_1248,N_19862,N_19769);
nor UO_1249 (O_1249,N_19680,N_19793);
or UO_1250 (O_1250,N_19723,N_19934);
nand UO_1251 (O_1251,N_19615,N_19840);
nand UO_1252 (O_1252,N_19867,N_19697);
xor UO_1253 (O_1253,N_19909,N_19716);
or UO_1254 (O_1254,N_19929,N_19829);
nor UO_1255 (O_1255,N_19615,N_19853);
xnor UO_1256 (O_1256,N_19970,N_19886);
xnor UO_1257 (O_1257,N_19864,N_19634);
xor UO_1258 (O_1258,N_19924,N_19950);
xnor UO_1259 (O_1259,N_19851,N_19733);
or UO_1260 (O_1260,N_19846,N_19784);
and UO_1261 (O_1261,N_19797,N_19738);
or UO_1262 (O_1262,N_19713,N_19844);
nand UO_1263 (O_1263,N_19605,N_19824);
nor UO_1264 (O_1264,N_19690,N_19762);
or UO_1265 (O_1265,N_19650,N_19870);
xnor UO_1266 (O_1266,N_19701,N_19779);
nand UO_1267 (O_1267,N_19612,N_19733);
nor UO_1268 (O_1268,N_19901,N_19980);
nor UO_1269 (O_1269,N_19952,N_19644);
nand UO_1270 (O_1270,N_19818,N_19957);
xor UO_1271 (O_1271,N_19787,N_19852);
and UO_1272 (O_1272,N_19912,N_19900);
nand UO_1273 (O_1273,N_19679,N_19963);
nor UO_1274 (O_1274,N_19619,N_19732);
xnor UO_1275 (O_1275,N_19631,N_19935);
nand UO_1276 (O_1276,N_19983,N_19866);
xnor UO_1277 (O_1277,N_19892,N_19647);
nor UO_1278 (O_1278,N_19766,N_19700);
and UO_1279 (O_1279,N_19849,N_19979);
xor UO_1280 (O_1280,N_19667,N_19822);
xor UO_1281 (O_1281,N_19669,N_19722);
nand UO_1282 (O_1282,N_19782,N_19763);
or UO_1283 (O_1283,N_19630,N_19757);
nand UO_1284 (O_1284,N_19673,N_19650);
nand UO_1285 (O_1285,N_19706,N_19828);
xnor UO_1286 (O_1286,N_19680,N_19773);
xnor UO_1287 (O_1287,N_19971,N_19756);
nand UO_1288 (O_1288,N_19610,N_19656);
xnor UO_1289 (O_1289,N_19923,N_19663);
or UO_1290 (O_1290,N_19633,N_19702);
and UO_1291 (O_1291,N_19748,N_19836);
and UO_1292 (O_1292,N_19971,N_19899);
or UO_1293 (O_1293,N_19779,N_19667);
and UO_1294 (O_1294,N_19614,N_19943);
and UO_1295 (O_1295,N_19929,N_19694);
nand UO_1296 (O_1296,N_19634,N_19819);
or UO_1297 (O_1297,N_19806,N_19618);
and UO_1298 (O_1298,N_19818,N_19886);
and UO_1299 (O_1299,N_19965,N_19692);
nor UO_1300 (O_1300,N_19774,N_19664);
xor UO_1301 (O_1301,N_19785,N_19642);
xnor UO_1302 (O_1302,N_19787,N_19797);
nand UO_1303 (O_1303,N_19917,N_19940);
xnor UO_1304 (O_1304,N_19751,N_19616);
xnor UO_1305 (O_1305,N_19833,N_19855);
nor UO_1306 (O_1306,N_19634,N_19823);
and UO_1307 (O_1307,N_19992,N_19874);
nor UO_1308 (O_1308,N_19668,N_19601);
xor UO_1309 (O_1309,N_19936,N_19731);
nor UO_1310 (O_1310,N_19759,N_19736);
xnor UO_1311 (O_1311,N_19673,N_19999);
nor UO_1312 (O_1312,N_19655,N_19820);
and UO_1313 (O_1313,N_19691,N_19959);
xnor UO_1314 (O_1314,N_19865,N_19770);
nor UO_1315 (O_1315,N_19805,N_19738);
nor UO_1316 (O_1316,N_19884,N_19765);
nand UO_1317 (O_1317,N_19656,N_19917);
or UO_1318 (O_1318,N_19767,N_19807);
and UO_1319 (O_1319,N_19695,N_19703);
nor UO_1320 (O_1320,N_19891,N_19977);
nor UO_1321 (O_1321,N_19874,N_19803);
nand UO_1322 (O_1322,N_19757,N_19914);
nand UO_1323 (O_1323,N_19673,N_19863);
and UO_1324 (O_1324,N_19857,N_19817);
and UO_1325 (O_1325,N_19672,N_19644);
xnor UO_1326 (O_1326,N_19684,N_19811);
and UO_1327 (O_1327,N_19967,N_19866);
nand UO_1328 (O_1328,N_19635,N_19680);
nand UO_1329 (O_1329,N_19689,N_19700);
xnor UO_1330 (O_1330,N_19938,N_19653);
xnor UO_1331 (O_1331,N_19998,N_19897);
and UO_1332 (O_1332,N_19825,N_19910);
nor UO_1333 (O_1333,N_19746,N_19756);
xnor UO_1334 (O_1334,N_19734,N_19777);
and UO_1335 (O_1335,N_19840,N_19650);
nand UO_1336 (O_1336,N_19845,N_19743);
nand UO_1337 (O_1337,N_19984,N_19882);
nor UO_1338 (O_1338,N_19892,N_19841);
or UO_1339 (O_1339,N_19755,N_19884);
or UO_1340 (O_1340,N_19986,N_19987);
xnor UO_1341 (O_1341,N_19747,N_19836);
nand UO_1342 (O_1342,N_19906,N_19696);
or UO_1343 (O_1343,N_19685,N_19865);
or UO_1344 (O_1344,N_19709,N_19719);
xor UO_1345 (O_1345,N_19835,N_19603);
and UO_1346 (O_1346,N_19824,N_19903);
nor UO_1347 (O_1347,N_19629,N_19887);
xnor UO_1348 (O_1348,N_19650,N_19618);
xor UO_1349 (O_1349,N_19767,N_19818);
or UO_1350 (O_1350,N_19967,N_19684);
and UO_1351 (O_1351,N_19982,N_19756);
nor UO_1352 (O_1352,N_19847,N_19663);
nand UO_1353 (O_1353,N_19704,N_19993);
or UO_1354 (O_1354,N_19989,N_19744);
xor UO_1355 (O_1355,N_19762,N_19616);
and UO_1356 (O_1356,N_19815,N_19952);
and UO_1357 (O_1357,N_19929,N_19931);
xor UO_1358 (O_1358,N_19726,N_19813);
or UO_1359 (O_1359,N_19779,N_19739);
nor UO_1360 (O_1360,N_19896,N_19790);
nor UO_1361 (O_1361,N_19779,N_19822);
xnor UO_1362 (O_1362,N_19609,N_19782);
and UO_1363 (O_1363,N_19872,N_19952);
xor UO_1364 (O_1364,N_19645,N_19993);
nand UO_1365 (O_1365,N_19931,N_19944);
xnor UO_1366 (O_1366,N_19876,N_19689);
or UO_1367 (O_1367,N_19823,N_19940);
and UO_1368 (O_1368,N_19956,N_19772);
and UO_1369 (O_1369,N_19622,N_19830);
nand UO_1370 (O_1370,N_19853,N_19913);
nand UO_1371 (O_1371,N_19923,N_19980);
or UO_1372 (O_1372,N_19868,N_19724);
nand UO_1373 (O_1373,N_19868,N_19870);
nand UO_1374 (O_1374,N_19932,N_19996);
and UO_1375 (O_1375,N_19957,N_19787);
and UO_1376 (O_1376,N_19724,N_19967);
nand UO_1377 (O_1377,N_19785,N_19700);
or UO_1378 (O_1378,N_19608,N_19660);
and UO_1379 (O_1379,N_19927,N_19731);
nand UO_1380 (O_1380,N_19633,N_19705);
or UO_1381 (O_1381,N_19807,N_19863);
and UO_1382 (O_1382,N_19884,N_19960);
or UO_1383 (O_1383,N_19706,N_19784);
or UO_1384 (O_1384,N_19771,N_19878);
xor UO_1385 (O_1385,N_19912,N_19618);
nand UO_1386 (O_1386,N_19865,N_19739);
or UO_1387 (O_1387,N_19609,N_19824);
or UO_1388 (O_1388,N_19849,N_19658);
and UO_1389 (O_1389,N_19815,N_19680);
and UO_1390 (O_1390,N_19749,N_19819);
nand UO_1391 (O_1391,N_19939,N_19937);
or UO_1392 (O_1392,N_19733,N_19701);
nor UO_1393 (O_1393,N_19933,N_19882);
nor UO_1394 (O_1394,N_19927,N_19980);
nand UO_1395 (O_1395,N_19604,N_19945);
and UO_1396 (O_1396,N_19959,N_19787);
xnor UO_1397 (O_1397,N_19860,N_19809);
and UO_1398 (O_1398,N_19671,N_19894);
nand UO_1399 (O_1399,N_19804,N_19864);
nand UO_1400 (O_1400,N_19904,N_19631);
or UO_1401 (O_1401,N_19934,N_19919);
and UO_1402 (O_1402,N_19814,N_19791);
and UO_1403 (O_1403,N_19697,N_19685);
nand UO_1404 (O_1404,N_19723,N_19957);
and UO_1405 (O_1405,N_19702,N_19852);
xnor UO_1406 (O_1406,N_19640,N_19798);
xor UO_1407 (O_1407,N_19784,N_19861);
nor UO_1408 (O_1408,N_19757,N_19909);
xor UO_1409 (O_1409,N_19781,N_19612);
and UO_1410 (O_1410,N_19717,N_19905);
nand UO_1411 (O_1411,N_19750,N_19736);
and UO_1412 (O_1412,N_19795,N_19952);
or UO_1413 (O_1413,N_19963,N_19840);
or UO_1414 (O_1414,N_19834,N_19957);
xnor UO_1415 (O_1415,N_19677,N_19846);
or UO_1416 (O_1416,N_19896,N_19776);
nor UO_1417 (O_1417,N_19915,N_19895);
xnor UO_1418 (O_1418,N_19611,N_19796);
nand UO_1419 (O_1419,N_19753,N_19735);
nand UO_1420 (O_1420,N_19746,N_19988);
xor UO_1421 (O_1421,N_19749,N_19800);
or UO_1422 (O_1422,N_19882,N_19687);
nor UO_1423 (O_1423,N_19619,N_19963);
xnor UO_1424 (O_1424,N_19617,N_19615);
nand UO_1425 (O_1425,N_19993,N_19869);
or UO_1426 (O_1426,N_19920,N_19804);
or UO_1427 (O_1427,N_19825,N_19925);
and UO_1428 (O_1428,N_19718,N_19959);
and UO_1429 (O_1429,N_19764,N_19888);
xor UO_1430 (O_1430,N_19809,N_19755);
and UO_1431 (O_1431,N_19835,N_19985);
and UO_1432 (O_1432,N_19689,N_19905);
nand UO_1433 (O_1433,N_19692,N_19788);
or UO_1434 (O_1434,N_19760,N_19945);
and UO_1435 (O_1435,N_19913,N_19907);
xor UO_1436 (O_1436,N_19942,N_19906);
nor UO_1437 (O_1437,N_19823,N_19729);
or UO_1438 (O_1438,N_19946,N_19920);
nand UO_1439 (O_1439,N_19689,N_19847);
and UO_1440 (O_1440,N_19768,N_19609);
or UO_1441 (O_1441,N_19972,N_19866);
nand UO_1442 (O_1442,N_19644,N_19773);
nor UO_1443 (O_1443,N_19949,N_19659);
and UO_1444 (O_1444,N_19622,N_19683);
nand UO_1445 (O_1445,N_19639,N_19655);
nor UO_1446 (O_1446,N_19886,N_19620);
and UO_1447 (O_1447,N_19673,N_19918);
nor UO_1448 (O_1448,N_19685,N_19609);
nand UO_1449 (O_1449,N_19975,N_19934);
or UO_1450 (O_1450,N_19717,N_19872);
nand UO_1451 (O_1451,N_19793,N_19850);
xor UO_1452 (O_1452,N_19803,N_19774);
xnor UO_1453 (O_1453,N_19830,N_19971);
or UO_1454 (O_1454,N_19811,N_19946);
nand UO_1455 (O_1455,N_19701,N_19802);
nand UO_1456 (O_1456,N_19705,N_19751);
nor UO_1457 (O_1457,N_19980,N_19607);
and UO_1458 (O_1458,N_19967,N_19903);
nand UO_1459 (O_1459,N_19670,N_19979);
xnor UO_1460 (O_1460,N_19800,N_19913);
xnor UO_1461 (O_1461,N_19968,N_19979);
and UO_1462 (O_1462,N_19604,N_19896);
nor UO_1463 (O_1463,N_19993,N_19768);
xnor UO_1464 (O_1464,N_19712,N_19600);
nand UO_1465 (O_1465,N_19797,N_19614);
and UO_1466 (O_1466,N_19924,N_19624);
nor UO_1467 (O_1467,N_19814,N_19651);
xnor UO_1468 (O_1468,N_19990,N_19773);
and UO_1469 (O_1469,N_19919,N_19872);
nor UO_1470 (O_1470,N_19901,N_19946);
and UO_1471 (O_1471,N_19831,N_19965);
and UO_1472 (O_1472,N_19674,N_19871);
nand UO_1473 (O_1473,N_19643,N_19991);
or UO_1474 (O_1474,N_19887,N_19794);
xor UO_1475 (O_1475,N_19658,N_19968);
xor UO_1476 (O_1476,N_19847,N_19839);
and UO_1477 (O_1477,N_19731,N_19839);
nand UO_1478 (O_1478,N_19643,N_19797);
xnor UO_1479 (O_1479,N_19867,N_19760);
or UO_1480 (O_1480,N_19673,N_19789);
nor UO_1481 (O_1481,N_19839,N_19634);
and UO_1482 (O_1482,N_19814,N_19923);
xnor UO_1483 (O_1483,N_19846,N_19728);
or UO_1484 (O_1484,N_19923,N_19836);
or UO_1485 (O_1485,N_19839,N_19843);
nand UO_1486 (O_1486,N_19888,N_19781);
or UO_1487 (O_1487,N_19931,N_19629);
xnor UO_1488 (O_1488,N_19864,N_19764);
and UO_1489 (O_1489,N_19630,N_19655);
xor UO_1490 (O_1490,N_19674,N_19874);
nor UO_1491 (O_1491,N_19954,N_19679);
nor UO_1492 (O_1492,N_19675,N_19660);
or UO_1493 (O_1493,N_19668,N_19901);
nor UO_1494 (O_1494,N_19782,N_19601);
and UO_1495 (O_1495,N_19615,N_19783);
nand UO_1496 (O_1496,N_19933,N_19697);
and UO_1497 (O_1497,N_19745,N_19917);
xor UO_1498 (O_1498,N_19808,N_19842);
nand UO_1499 (O_1499,N_19687,N_19766);
xor UO_1500 (O_1500,N_19971,N_19666);
or UO_1501 (O_1501,N_19883,N_19952);
nand UO_1502 (O_1502,N_19643,N_19669);
xor UO_1503 (O_1503,N_19689,N_19758);
nand UO_1504 (O_1504,N_19838,N_19760);
or UO_1505 (O_1505,N_19723,N_19983);
or UO_1506 (O_1506,N_19604,N_19770);
nand UO_1507 (O_1507,N_19991,N_19670);
nand UO_1508 (O_1508,N_19993,N_19725);
xor UO_1509 (O_1509,N_19761,N_19825);
or UO_1510 (O_1510,N_19980,N_19993);
or UO_1511 (O_1511,N_19978,N_19758);
or UO_1512 (O_1512,N_19912,N_19660);
nor UO_1513 (O_1513,N_19757,N_19912);
nand UO_1514 (O_1514,N_19790,N_19875);
xnor UO_1515 (O_1515,N_19782,N_19861);
xnor UO_1516 (O_1516,N_19713,N_19947);
nor UO_1517 (O_1517,N_19944,N_19696);
xnor UO_1518 (O_1518,N_19673,N_19852);
nor UO_1519 (O_1519,N_19635,N_19657);
nor UO_1520 (O_1520,N_19615,N_19648);
and UO_1521 (O_1521,N_19872,N_19645);
and UO_1522 (O_1522,N_19950,N_19956);
and UO_1523 (O_1523,N_19967,N_19648);
nor UO_1524 (O_1524,N_19642,N_19738);
xnor UO_1525 (O_1525,N_19877,N_19894);
nand UO_1526 (O_1526,N_19964,N_19740);
xor UO_1527 (O_1527,N_19609,N_19970);
or UO_1528 (O_1528,N_19969,N_19735);
or UO_1529 (O_1529,N_19929,N_19828);
and UO_1530 (O_1530,N_19881,N_19837);
or UO_1531 (O_1531,N_19982,N_19992);
and UO_1532 (O_1532,N_19809,N_19691);
nand UO_1533 (O_1533,N_19773,N_19655);
and UO_1534 (O_1534,N_19698,N_19705);
or UO_1535 (O_1535,N_19832,N_19938);
nand UO_1536 (O_1536,N_19665,N_19628);
nor UO_1537 (O_1537,N_19701,N_19709);
nand UO_1538 (O_1538,N_19750,N_19604);
or UO_1539 (O_1539,N_19894,N_19882);
and UO_1540 (O_1540,N_19850,N_19843);
xnor UO_1541 (O_1541,N_19626,N_19909);
or UO_1542 (O_1542,N_19880,N_19606);
xnor UO_1543 (O_1543,N_19973,N_19739);
nand UO_1544 (O_1544,N_19610,N_19989);
or UO_1545 (O_1545,N_19898,N_19788);
or UO_1546 (O_1546,N_19720,N_19864);
nor UO_1547 (O_1547,N_19927,N_19994);
or UO_1548 (O_1548,N_19614,N_19742);
xnor UO_1549 (O_1549,N_19916,N_19867);
nand UO_1550 (O_1550,N_19720,N_19953);
nand UO_1551 (O_1551,N_19788,N_19727);
nand UO_1552 (O_1552,N_19659,N_19627);
nor UO_1553 (O_1553,N_19968,N_19649);
nand UO_1554 (O_1554,N_19915,N_19871);
and UO_1555 (O_1555,N_19844,N_19778);
or UO_1556 (O_1556,N_19705,N_19898);
xnor UO_1557 (O_1557,N_19760,N_19830);
xor UO_1558 (O_1558,N_19847,N_19907);
and UO_1559 (O_1559,N_19610,N_19639);
and UO_1560 (O_1560,N_19651,N_19934);
nor UO_1561 (O_1561,N_19999,N_19747);
nor UO_1562 (O_1562,N_19636,N_19605);
nor UO_1563 (O_1563,N_19649,N_19906);
or UO_1564 (O_1564,N_19931,N_19792);
and UO_1565 (O_1565,N_19663,N_19798);
and UO_1566 (O_1566,N_19932,N_19948);
or UO_1567 (O_1567,N_19676,N_19701);
xor UO_1568 (O_1568,N_19641,N_19865);
xnor UO_1569 (O_1569,N_19758,N_19746);
and UO_1570 (O_1570,N_19858,N_19940);
nor UO_1571 (O_1571,N_19752,N_19651);
or UO_1572 (O_1572,N_19722,N_19947);
or UO_1573 (O_1573,N_19649,N_19805);
and UO_1574 (O_1574,N_19607,N_19666);
nand UO_1575 (O_1575,N_19995,N_19777);
nand UO_1576 (O_1576,N_19699,N_19650);
nor UO_1577 (O_1577,N_19827,N_19999);
or UO_1578 (O_1578,N_19701,N_19980);
nand UO_1579 (O_1579,N_19984,N_19787);
xnor UO_1580 (O_1580,N_19643,N_19899);
or UO_1581 (O_1581,N_19825,N_19955);
nand UO_1582 (O_1582,N_19992,N_19652);
xnor UO_1583 (O_1583,N_19678,N_19939);
nor UO_1584 (O_1584,N_19853,N_19670);
and UO_1585 (O_1585,N_19989,N_19993);
xnor UO_1586 (O_1586,N_19831,N_19903);
nand UO_1587 (O_1587,N_19639,N_19757);
nor UO_1588 (O_1588,N_19854,N_19976);
nor UO_1589 (O_1589,N_19710,N_19820);
xnor UO_1590 (O_1590,N_19601,N_19733);
or UO_1591 (O_1591,N_19840,N_19622);
and UO_1592 (O_1592,N_19969,N_19806);
nor UO_1593 (O_1593,N_19678,N_19975);
nand UO_1594 (O_1594,N_19962,N_19901);
or UO_1595 (O_1595,N_19652,N_19612);
nor UO_1596 (O_1596,N_19614,N_19944);
or UO_1597 (O_1597,N_19678,N_19874);
or UO_1598 (O_1598,N_19629,N_19807);
nand UO_1599 (O_1599,N_19807,N_19937);
xnor UO_1600 (O_1600,N_19743,N_19699);
or UO_1601 (O_1601,N_19622,N_19875);
or UO_1602 (O_1602,N_19727,N_19750);
nor UO_1603 (O_1603,N_19657,N_19887);
xnor UO_1604 (O_1604,N_19803,N_19601);
nand UO_1605 (O_1605,N_19874,N_19721);
or UO_1606 (O_1606,N_19915,N_19833);
nand UO_1607 (O_1607,N_19706,N_19824);
nand UO_1608 (O_1608,N_19967,N_19620);
nor UO_1609 (O_1609,N_19931,N_19934);
nor UO_1610 (O_1610,N_19623,N_19753);
or UO_1611 (O_1611,N_19821,N_19694);
nand UO_1612 (O_1612,N_19625,N_19894);
nor UO_1613 (O_1613,N_19809,N_19961);
nand UO_1614 (O_1614,N_19613,N_19850);
and UO_1615 (O_1615,N_19755,N_19905);
or UO_1616 (O_1616,N_19692,N_19609);
xor UO_1617 (O_1617,N_19760,N_19723);
xnor UO_1618 (O_1618,N_19966,N_19668);
xor UO_1619 (O_1619,N_19793,N_19830);
nor UO_1620 (O_1620,N_19724,N_19608);
nor UO_1621 (O_1621,N_19865,N_19696);
or UO_1622 (O_1622,N_19647,N_19725);
nand UO_1623 (O_1623,N_19748,N_19810);
nand UO_1624 (O_1624,N_19865,N_19918);
and UO_1625 (O_1625,N_19741,N_19647);
and UO_1626 (O_1626,N_19945,N_19646);
nand UO_1627 (O_1627,N_19871,N_19962);
nor UO_1628 (O_1628,N_19661,N_19833);
nor UO_1629 (O_1629,N_19750,N_19661);
or UO_1630 (O_1630,N_19603,N_19672);
xor UO_1631 (O_1631,N_19834,N_19873);
nand UO_1632 (O_1632,N_19609,N_19749);
and UO_1633 (O_1633,N_19600,N_19717);
or UO_1634 (O_1634,N_19937,N_19611);
or UO_1635 (O_1635,N_19832,N_19794);
xor UO_1636 (O_1636,N_19737,N_19768);
or UO_1637 (O_1637,N_19727,N_19815);
nand UO_1638 (O_1638,N_19645,N_19936);
or UO_1639 (O_1639,N_19748,N_19979);
and UO_1640 (O_1640,N_19744,N_19922);
nor UO_1641 (O_1641,N_19674,N_19909);
nand UO_1642 (O_1642,N_19801,N_19959);
nor UO_1643 (O_1643,N_19732,N_19738);
xnor UO_1644 (O_1644,N_19716,N_19679);
and UO_1645 (O_1645,N_19638,N_19996);
nor UO_1646 (O_1646,N_19665,N_19879);
xnor UO_1647 (O_1647,N_19682,N_19740);
or UO_1648 (O_1648,N_19786,N_19920);
or UO_1649 (O_1649,N_19852,N_19684);
or UO_1650 (O_1650,N_19651,N_19845);
or UO_1651 (O_1651,N_19660,N_19713);
and UO_1652 (O_1652,N_19911,N_19838);
nor UO_1653 (O_1653,N_19873,N_19979);
nand UO_1654 (O_1654,N_19830,N_19850);
and UO_1655 (O_1655,N_19954,N_19809);
xnor UO_1656 (O_1656,N_19842,N_19645);
xnor UO_1657 (O_1657,N_19710,N_19634);
nand UO_1658 (O_1658,N_19939,N_19742);
or UO_1659 (O_1659,N_19732,N_19952);
and UO_1660 (O_1660,N_19908,N_19921);
and UO_1661 (O_1661,N_19791,N_19853);
nand UO_1662 (O_1662,N_19844,N_19739);
and UO_1663 (O_1663,N_19883,N_19744);
or UO_1664 (O_1664,N_19650,N_19807);
nand UO_1665 (O_1665,N_19937,N_19846);
nand UO_1666 (O_1666,N_19686,N_19742);
and UO_1667 (O_1667,N_19816,N_19788);
and UO_1668 (O_1668,N_19687,N_19952);
xor UO_1669 (O_1669,N_19680,N_19663);
xnor UO_1670 (O_1670,N_19745,N_19981);
or UO_1671 (O_1671,N_19967,N_19667);
nand UO_1672 (O_1672,N_19740,N_19697);
nand UO_1673 (O_1673,N_19661,N_19697);
nand UO_1674 (O_1674,N_19835,N_19912);
xor UO_1675 (O_1675,N_19689,N_19970);
nor UO_1676 (O_1676,N_19749,N_19979);
or UO_1677 (O_1677,N_19860,N_19749);
and UO_1678 (O_1678,N_19989,N_19736);
and UO_1679 (O_1679,N_19718,N_19779);
or UO_1680 (O_1680,N_19973,N_19748);
and UO_1681 (O_1681,N_19808,N_19957);
nand UO_1682 (O_1682,N_19786,N_19968);
xor UO_1683 (O_1683,N_19804,N_19849);
and UO_1684 (O_1684,N_19854,N_19765);
xnor UO_1685 (O_1685,N_19998,N_19719);
xor UO_1686 (O_1686,N_19984,N_19976);
and UO_1687 (O_1687,N_19653,N_19612);
nor UO_1688 (O_1688,N_19781,N_19827);
nor UO_1689 (O_1689,N_19914,N_19686);
or UO_1690 (O_1690,N_19969,N_19789);
and UO_1691 (O_1691,N_19800,N_19867);
and UO_1692 (O_1692,N_19617,N_19864);
nand UO_1693 (O_1693,N_19854,N_19805);
or UO_1694 (O_1694,N_19666,N_19753);
nor UO_1695 (O_1695,N_19979,N_19833);
or UO_1696 (O_1696,N_19744,N_19669);
nor UO_1697 (O_1697,N_19800,N_19828);
nor UO_1698 (O_1698,N_19759,N_19631);
nor UO_1699 (O_1699,N_19706,N_19647);
xnor UO_1700 (O_1700,N_19808,N_19755);
and UO_1701 (O_1701,N_19996,N_19888);
xor UO_1702 (O_1702,N_19711,N_19813);
xor UO_1703 (O_1703,N_19827,N_19880);
nor UO_1704 (O_1704,N_19750,N_19723);
nor UO_1705 (O_1705,N_19611,N_19791);
nor UO_1706 (O_1706,N_19638,N_19702);
or UO_1707 (O_1707,N_19786,N_19888);
and UO_1708 (O_1708,N_19710,N_19957);
and UO_1709 (O_1709,N_19621,N_19622);
and UO_1710 (O_1710,N_19975,N_19861);
nor UO_1711 (O_1711,N_19911,N_19782);
or UO_1712 (O_1712,N_19620,N_19996);
or UO_1713 (O_1713,N_19833,N_19628);
or UO_1714 (O_1714,N_19923,N_19686);
nor UO_1715 (O_1715,N_19899,N_19645);
and UO_1716 (O_1716,N_19732,N_19954);
or UO_1717 (O_1717,N_19888,N_19710);
nand UO_1718 (O_1718,N_19918,N_19699);
xnor UO_1719 (O_1719,N_19605,N_19718);
nand UO_1720 (O_1720,N_19976,N_19624);
nand UO_1721 (O_1721,N_19885,N_19609);
xor UO_1722 (O_1722,N_19765,N_19824);
xor UO_1723 (O_1723,N_19898,N_19919);
and UO_1724 (O_1724,N_19630,N_19693);
xor UO_1725 (O_1725,N_19643,N_19656);
xnor UO_1726 (O_1726,N_19726,N_19985);
or UO_1727 (O_1727,N_19600,N_19894);
and UO_1728 (O_1728,N_19679,N_19857);
nor UO_1729 (O_1729,N_19904,N_19879);
xnor UO_1730 (O_1730,N_19630,N_19809);
or UO_1731 (O_1731,N_19642,N_19669);
or UO_1732 (O_1732,N_19854,N_19868);
nor UO_1733 (O_1733,N_19655,N_19732);
nor UO_1734 (O_1734,N_19994,N_19678);
or UO_1735 (O_1735,N_19956,N_19605);
or UO_1736 (O_1736,N_19849,N_19959);
xnor UO_1737 (O_1737,N_19893,N_19685);
or UO_1738 (O_1738,N_19608,N_19745);
nand UO_1739 (O_1739,N_19934,N_19602);
xor UO_1740 (O_1740,N_19870,N_19962);
nor UO_1741 (O_1741,N_19710,N_19882);
nand UO_1742 (O_1742,N_19640,N_19958);
xnor UO_1743 (O_1743,N_19998,N_19928);
nand UO_1744 (O_1744,N_19884,N_19891);
xor UO_1745 (O_1745,N_19673,N_19912);
xnor UO_1746 (O_1746,N_19905,N_19644);
nand UO_1747 (O_1747,N_19727,N_19746);
or UO_1748 (O_1748,N_19790,N_19670);
nand UO_1749 (O_1749,N_19717,N_19695);
xor UO_1750 (O_1750,N_19823,N_19771);
xnor UO_1751 (O_1751,N_19820,N_19775);
and UO_1752 (O_1752,N_19734,N_19700);
and UO_1753 (O_1753,N_19675,N_19657);
xor UO_1754 (O_1754,N_19989,N_19728);
xor UO_1755 (O_1755,N_19869,N_19724);
nor UO_1756 (O_1756,N_19613,N_19841);
or UO_1757 (O_1757,N_19797,N_19953);
nor UO_1758 (O_1758,N_19917,N_19685);
nor UO_1759 (O_1759,N_19895,N_19614);
xnor UO_1760 (O_1760,N_19615,N_19738);
xor UO_1761 (O_1761,N_19970,N_19977);
nand UO_1762 (O_1762,N_19775,N_19714);
xor UO_1763 (O_1763,N_19919,N_19782);
nor UO_1764 (O_1764,N_19609,N_19959);
or UO_1765 (O_1765,N_19623,N_19749);
or UO_1766 (O_1766,N_19680,N_19973);
nand UO_1767 (O_1767,N_19721,N_19889);
and UO_1768 (O_1768,N_19809,N_19681);
nand UO_1769 (O_1769,N_19670,N_19920);
nor UO_1770 (O_1770,N_19966,N_19980);
nand UO_1771 (O_1771,N_19971,N_19733);
and UO_1772 (O_1772,N_19993,N_19783);
or UO_1773 (O_1773,N_19654,N_19606);
nand UO_1774 (O_1774,N_19620,N_19883);
or UO_1775 (O_1775,N_19777,N_19613);
nor UO_1776 (O_1776,N_19758,N_19948);
nor UO_1777 (O_1777,N_19917,N_19739);
or UO_1778 (O_1778,N_19714,N_19666);
nand UO_1779 (O_1779,N_19608,N_19722);
or UO_1780 (O_1780,N_19604,N_19628);
xnor UO_1781 (O_1781,N_19959,N_19640);
and UO_1782 (O_1782,N_19676,N_19772);
or UO_1783 (O_1783,N_19831,N_19655);
xnor UO_1784 (O_1784,N_19864,N_19822);
and UO_1785 (O_1785,N_19928,N_19993);
and UO_1786 (O_1786,N_19774,N_19629);
nor UO_1787 (O_1787,N_19619,N_19896);
nor UO_1788 (O_1788,N_19809,N_19964);
nor UO_1789 (O_1789,N_19898,N_19751);
xor UO_1790 (O_1790,N_19651,N_19610);
and UO_1791 (O_1791,N_19723,N_19972);
nor UO_1792 (O_1792,N_19729,N_19787);
or UO_1793 (O_1793,N_19970,N_19990);
nand UO_1794 (O_1794,N_19640,N_19633);
and UO_1795 (O_1795,N_19834,N_19631);
nor UO_1796 (O_1796,N_19965,N_19643);
nor UO_1797 (O_1797,N_19888,N_19676);
and UO_1798 (O_1798,N_19855,N_19694);
nor UO_1799 (O_1799,N_19843,N_19778);
xor UO_1800 (O_1800,N_19854,N_19723);
nand UO_1801 (O_1801,N_19650,N_19604);
or UO_1802 (O_1802,N_19888,N_19939);
xnor UO_1803 (O_1803,N_19747,N_19863);
xnor UO_1804 (O_1804,N_19989,N_19663);
or UO_1805 (O_1805,N_19986,N_19976);
xor UO_1806 (O_1806,N_19870,N_19753);
xor UO_1807 (O_1807,N_19840,N_19695);
nor UO_1808 (O_1808,N_19819,N_19802);
nand UO_1809 (O_1809,N_19619,N_19671);
nand UO_1810 (O_1810,N_19803,N_19883);
and UO_1811 (O_1811,N_19819,N_19645);
nor UO_1812 (O_1812,N_19844,N_19820);
nand UO_1813 (O_1813,N_19652,N_19757);
xor UO_1814 (O_1814,N_19947,N_19895);
and UO_1815 (O_1815,N_19790,N_19700);
or UO_1816 (O_1816,N_19902,N_19958);
or UO_1817 (O_1817,N_19629,N_19707);
or UO_1818 (O_1818,N_19969,N_19643);
nor UO_1819 (O_1819,N_19999,N_19911);
xor UO_1820 (O_1820,N_19748,N_19674);
xor UO_1821 (O_1821,N_19797,N_19998);
or UO_1822 (O_1822,N_19951,N_19785);
and UO_1823 (O_1823,N_19673,N_19784);
nor UO_1824 (O_1824,N_19788,N_19849);
nor UO_1825 (O_1825,N_19723,N_19955);
and UO_1826 (O_1826,N_19930,N_19860);
and UO_1827 (O_1827,N_19660,N_19624);
nand UO_1828 (O_1828,N_19902,N_19646);
nor UO_1829 (O_1829,N_19936,N_19845);
nand UO_1830 (O_1830,N_19707,N_19984);
nor UO_1831 (O_1831,N_19829,N_19765);
or UO_1832 (O_1832,N_19708,N_19957);
and UO_1833 (O_1833,N_19669,N_19867);
nor UO_1834 (O_1834,N_19921,N_19988);
nand UO_1835 (O_1835,N_19729,N_19703);
nor UO_1836 (O_1836,N_19714,N_19965);
xnor UO_1837 (O_1837,N_19802,N_19800);
or UO_1838 (O_1838,N_19972,N_19642);
nor UO_1839 (O_1839,N_19635,N_19826);
nor UO_1840 (O_1840,N_19961,N_19700);
nand UO_1841 (O_1841,N_19929,N_19908);
and UO_1842 (O_1842,N_19819,N_19897);
xor UO_1843 (O_1843,N_19976,N_19888);
nand UO_1844 (O_1844,N_19639,N_19865);
or UO_1845 (O_1845,N_19616,N_19721);
nor UO_1846 (O_1846,N_19795,N_19921);
nor UO_1847 (O_1847,N_19963,N_19678);
or UO_1848 (O_1848,N_19737,N_19879);
or UO_1849 (O_1849,N_19723,N_19729);
or UO_1850 (O_1850,N_19716,N_19995);
or UO_1851 (O_1851,N_19631,N_19886);
nor UO_1852 (O_1852,N_19645,N_19973);
and UO_1853 (O_1853,N_19711,N_19654);
nor UO_1854 (O_1854,N_19696,N_19692);
nand UO_1855 (O_1855,N_19772,N_19961);
or UO_1856 (O_1856,N_19968,N_19719);
nand UO_1857 (O_1857,N_19823,N_19891);
and UO_1858 (O_1858,N_19677,N_19903);
xnor UO_1859 (O_1859,N_19723,N_19647);
and UO_1860 (O_1860,N_19985,N_19997);
and UO_1861 (O_1861,N_19661,N_19832);
nand UO_1862 (O_1862,N_19681,N_19805);
xnor UO_1863 (O_1863,N_19805,N_19808);
xnor UO_1864 (O_1864,N_19844,N_19716);
nand UO_1865 (O_1865,N_19923,N_19832);
and UO_1866 (O_1866,N_19697,N_19777);
xnor UO_1867 (O_1867,N_19751,N_19880);
or UO_1868 (O_1868,N_19640,N_19888);
nor UO_1869 (O_1869,N_19726,N_19797);
xnor UO_1870 (O_1870,N_19642,N_19956);
xnor UO_1871 (O_1871,N_19973,N_19981);
nor UO_1872 (O_1872,N_19787,N_19770);
nor UO_1873 (O_1873,N_19610,N_19718);
or UO_1874 (O_1874,N_19837,N_19878);
and UO_1875 (O_1875,N_19977,N_19696);
or UO_1876 (O_1876,N_19671,N_19864);
nor UO_1877 (O_1877,N_19707,N_19632);
xnor UO_1878 (O_1878,N_19829,N_19726);
xor UO_1879 (O_1879,N_19752,N_19618);
or UO_1880 (O_1880,N_19710,N_19892);
or UO_1881 (O_1881,N_19658,N_19654);
and UO_1882 (O_1882,N_19652,N_19905);
and UO_1883 (O_1883,N_19943,N_19917);
nand UO_1884 (O_1884,N_19763,N_19881);
and UO_1885 (O_1885,N_19845,N_19895);
and UO_1886 (O_1886,N_19693,N_19719);
or UO_1887 (O_1887,N_19735,N_19652);
xor UO_1888 (O_1888,N_19951,N_19774);
nand UO_1889 (O_1889,N_19799,N_19910);
and UO_1890 (O_1890,N_19847,N_19860);
xor UO_1891 (O_1891,N_19688,N_19926);
and UO_1892 (O_1892,N_19943,N_19626);
nor UO_1893 (O_1893,N_19794,N_19889);
nand UO_1894 (O_1894,N_19669,N_19940);
xor UO_1895 (O_1895,N_19914,N_19645);
nor UO_1896 (O_1896,N_19788,N_19653);
xor UO_1897 (O_1897,N_19930,N_19904);
xor UO_1898 (O_1898,N_19693,N_19717);
nand UO_1899 (O_1899,N_19625,N_19928);
and UO_1900 (O_1900,N_19901,N_19741);
nand UO_1901 (O_1901,N_19616,N_19931);
nand UO_1902 (O_1902,N_19636,N_19639);
nor UO_1903 (O_1903,N_19985,N_19890);
or UO_1904 (O_1904,N_19682,N_19856);
or UO_1905 (O_1905,N_19600,N_19635);
or UO_1906 (O_1906,N_19607,N_19713);
nand UO_1907 (O_1907,N_19851,N_19795);
nand UO_1908 (O_1908,N_19820,N_19909);
or UO_1909 (O_1909,N_19781,N_19950);
or UO_1910 (O_1910,N_19854,N_19712);
nor UO_1911 (O_1911,N_19723,N_19703);
or UO_1912 (O_1912,N_19933,N_19611);
nand UO_1913 (O_1913,N_19932,N_19879);
nand UO_1914 (O_1914,N_19628,N_19651);
nor UO_1915 (O_1915,N_19775,N_19942);
and UO_1916 (O_1916,N_19717,N_19784);
nand UO_1917 (O_1917,N_19929,N_19643);
and UO_1918 (O_1918,N_19825,N_19765);
or UO_1919 (O_1919,N_19807,N_19689);
or UO_1920 (O_1920,N_19649,N_19969);
or UO_1921 (O_1921,N_19605,N_19997);
or UO_1922 (O_1922,N_19601,N_19819);
or UO_1923 (O_1923,N_19976,N_19621);
xor UO_1924 (O_1924,N_19963,N_19655);
nand UO_1925 (O_1925,N_19860,N_19616);
xor UO_1926 (O_1926,N_19892,N_19888);
xor UO_1927 (O_1927,N_19694,N_19648);
nor UO_1928 (O_1928,N_19897,N_19743);
xor UO_1929 (O_1929,N_19695,N_19623);
nor UO_1930 (O_1930,N_19896,N_19876);
nand UO_1931 (O_1931,N_19956,N_19676);
and UO_1932 (O_1932,N_19687,N_19818);
nor UO_1933 (O_1933,N_19821,N_19855);
and UO_1934 (O_1934,N_19629,N_19756);
xor UO_1935 (O_1935,N_19904,N_19731);
nor UO_1936 (O_1936,N_19783,N_19964);
nor UO_1937 (O_1937,N_19835,N_19687);
and UO_1938 (O_1938,N_19937,N_19982);
nor UO_1939 (O_1939,N_19865,N_19715);
nand UO_1940 (O_1940,N_19698,N_19799);
xnor UO_1941 (O_1941,N_19671,N_19719);
xnor UO_1942 (O_1942,N_19868,N_19874);
nand UO_1943 (O_1943,N_19757,N_19849);
xor UO_1944 (O_1944,N_19919,N_19737);
nor UO_1945 (O_1945,N_19600,N_19673);
nand UO_1946 (O_1946,N_19803,N_19839);
nor UO_1947 (O_1947,N_19967,N_19869);
and UO_1948 (O_1948,N_19726,N_19612);
or UO_1949 (O_1949,N_19641,N_19966);
or UO_1950 (O_1950,N_19691,N_19695);
xor UO_1951 (O_1951,N_19911,N_19869);
xnor UO_1952 (O_1952,N_19865,N_19882);
and UO_1953 (O_1953,N_19923,N_19740);
or UO_1954 (O_1954,N_19629,N_19706);
or UO_1955 (O_1955,N_19805,N_19672);
nand UO_1956 (O_1956,N_19965,N_19961);
nand UO_1957 (O_1957,N_19958,N_19690);
nand UO_1958 (O_1958,N_19932,N_19655);
xnor UO_1959 (O_1959,N_19750,N_19753);
nand UO_1960 (O_1960,N_19899,N_19903);
xor UO_1961 (O_1961,N_19606,N_19893);
nand UO_1962 (O_1962,N_19689,N_19729);
and UO_1963 (O_1963,N_19932,N_19923);
and UO_1964 (O_1964,N_19907,N_19799);
xor UO_1965 (O_1965,N_19934,N_19917);
or UO_1966 (O_1966,N_19825,N_19889);
nand UO_1967 (O_1967,N_19628,N_19832);
or UO_1968 (O_1968,N_19777,N_19665);
nand UO_1969 (O_1969,N_19733,N_19969);
nor UO_1970 (O_1970,N_19886,N_19914);
xnor UO_1971 (O_1971,N_19602,N_19679);
nor UO_1972 (O_1972,N_19933,N_19842);
nand UO_1973 (O_1973,N_19848,N_19733);
and UO_1974 (O_1974,N_19995,N_19652);
or UO_1975 (O_1975,N_19784,N_19633);
and UO_1976 (O_1976,N_19983,N_19837);
xnor UO_1977 (O_1977,N_19688,N_19739);
or UO_1978 (O_1978,N_19989,N_19602);
or UO_1979 (O_1979,N_19668,N_19900);
xnor UO_1980 (O_1980,N_19805,N_19618);
nand UO_1981 (O_1981,N_19855,N_19844);
nor UO_1982 (O_1982,N_19622,N_19691);
nand UO_1983 (O_1983,N_19877,N_19729);
nor UO_1984 (O_1984,N_19821,N_19939);
nand UO_1985 (O_1985,N_19813,N_19702);
or UO_1986 (O_1986,N_19863,N_19947);
nor UO_1987 (O_1987,N_19887,N_19682);
nor UO_1988 (O_1988,N_19743,N_19866);
and UO_1989 (O_1989,N_19943,N_19669);
nand UO_1990 (O_1990,N_19919,N_19618);
xnor UO_1991 (O_1991,N_19691,N_19694);
and UO_1992 (O_1992,N_19797,N_19642);
and UO_1993 (O_1993,N_19902,N_19700);
and UO_1994 (O_1994,N_19855,N_19738);
nand UO_1995 (O_1995,N_19831,N_19600);
or UO_1996 (O_1996,N_19721,N_19912);
nor UO_1997 (O_1997,N_19601,N_19604);
or UO_1998 (O_1998,N_19784,N_19774);
xnor UO_1999 (O_1999,N_19768,N_19917);
xnor UO_2000 (O_2000,N_19703,N_19620);
and UO_2001 (O_2001,N_19984,N_19832);
and UO_2002 (O_2002,N_19721,N_19807);
nor UO_2003 (O_2003,N_19947,N_19613);
nor UO_2004 (O_2004,N_19705,N_19835);
xor UO_2005 (O_2005,N_19670,N_19922);
nor UO_2006 (O_2006,N_19946,N_19843);
and UO_2007 (O_2007,N_19856,N_19945);
and UO_2008 (O_2008,N_19767,N_19611);
nor UO_2009 (O_2009,N_19951,N_19700);
or UO_2010 (O_2010,N_19950,N_19894);
xnor UO_2011 (O_2011,N_19809,N_19733);
nor UO_2012 (O_2012,N_19705,N_19647);
xnor UO_2013 (O_2013,N_19600,N_19605);
xnor UO_2014 (O_2014,N_19912,N_19638);
xnor UO_2015 (O_2015,N_19882,N_19945);
and UO_2016 (O_2016,N_19687,N_19807);
and UO_2017 (O_2017,N_19989,N_19635);
nor UO_2018 (O_2018,N_19812,N_19617);
nand UO_2019 (O_2019,N_19952,N_19768);
nand UO_2020 (O_2020,N_19604,N_19922);
or UO_2021 (O_2021,N_19816,N_19606);
and UO_2022 (O_2022,N_19633,N_19917);
nor UO_2023 (O_2023,N_19961,N_19864);
and UO_2024 (O_2024,N_19768,N_19699);
xor UO_2025 (O_2025,N_19833,N_19668);
nor UO_2026 (O_2026,N_19817,N_19609);
and UO_2027 (O_2027,N_19988,N_19792);
nor UO_2028 (O_2028,N_19893,N_19958);
nand UO_2029 (O_2029,N_19852,N_19726);
nand UO_2030 (O_2030,N_19862,N_19999);
and UO_2031 (O_2031,N_19954,N_19695);
xor UO_2032 (O_2032,N_19790,N_19876);
xnor UO_2033 (O_2033,N_19959,N_19693);
xor UO_2034 (O_2034,N_19765,N_19678);
or UO_2035 (O_2035,N_19760,N_19856);
or UO_2036 (O_2036,N_19896,N_19840);
nand UO_2037 (O_2037,N_19826,N_19615);
nand UO_2038 (O_2038,N_19824,N_19874);
xnor UO_2039 (O_2039,N_19658,N_19735);
or UO_2040 (O_2040,N_19604,N_19618);
nand UO_2041 (O_2041,N_19782,N_19952);
nor UO_2042 (O_2042,N_19874,N_19644);
and UO_2043 (O_2043,N_19674,N_19707);
or UO_2044 (O_2044,N_19919,N_19888);
or UO_2045 (O_2045,N_19620,N_19607);
nand UO_2046 (O_2046,N_19982,N_19868);
or UO_2047 (O_2047,N_19630,N_19975);
or UO_2048 (O_2048,N_19806,N_19827);
nor UO_2049 (O_2049,N_19794,N_19766);
xnor UO_2050 (O_2050,N_19935,N_19758);
nand UO_2051 (O_2051,N_19892,N_19827);
nor UO_2052 (O_2052,N_19762,N_19942);
nand UO_2053 (O_2053,N_19791,N_19608);
and UO_2054 (O_2054,N_19986,N_19879);
or UO_2055 (O_2055,N_19833,N_19821);
nor UO_2056 (O_2056,N_19826,N_19773);
nand UO_2057 (O_2057,N_19710,N_19841);
or UO_2058 (O_2058,N_19860,N_19999);
nor UO_2059 (O_2059,N_19968,N_19757);
nand UO_2060 (O_2060,N_19989,N_19978);
nor UO_2061 (O_2061,N_19930,N_19971);
nor UO_2062 (O_2062,N_19908,N_19707);
and UO_2063 (O_2063,N_19636,N_19840);
or UO_2064 (O_2064,N_19952,N_19676);
xnor UO_2065 (O_2065,N_19815,N_19904);
and UO_2066 (O_2066,N_19757,N_19809);
xnor UO_2067 (O_2067,N_19825,N_19759);
and UO_2068 (O_2068,N_19668,N_19697);
nand UO_2069 (O_2069,N_19648,N_19706);
nand UO_2070 (O_2070,N_19964,N_19886);
xor UO_2071 (O_2071,N_19794,N_19685);
nor UO_2072 (O_2072,N_19798,N_19793);
nand UO_2073 (O_2073,N_19841,N_19667);
nor UO_2074 (O_2074,N_19973,N_19810);
or UO_2075 (O_2075,N_19708,N_19910);
nand UO_2076 (O_2076,N_19834,N_19796);
nand UO_2077 (O_2077,N_19714,N_19679);
or UO_2078 (O_2078,N_19700,N_19668);
or UO_2079 (O_2079,N_19784,N_19600);
xor UO_2080 (O_2080,N_19715,N_19833);
and UO_2081 (O_2081,N_19675,N_19683);
or UO_2082 (O_2082,N_19764,N_19923);
xnor UO_2083 (O_2083,N_19683,N_19815);
xor UO_2084 (O_2084,N_19908,N_19622);
nand UO_2085 (O_2085,N_19924,N_19681);
and UO_2086 (O_2086,N_19972,N_19821);
nand UO_2087 (O_2087,N_19757,N_19640);
xor UO_2088 (O_2088,N_19918,N_19966);
nor UO_2089 (O_2089,N_19943,N_19818);
xor UO_2090 (O_2090,N_19996,N_19823);
and UO_2091 (O_2091,N_19968,N_19618);
and UO_2092 (O_2092,N_19714,N_19607);
xnor UO_2093 (O_2093,N_19979,N_19800);
nand UO_2094 (O_2094,N_19671,N_19964);
nor UO_2095 (O_2095,N_19913,N_19864);
or UO_2096 (O_2096,N_19713,N_19954);
and UO_2097 (O_2097,N_19736,N_19793);
nand UO_2098 (O_2098,N_19748,N_19662);
nor UO_2099 (O_2099,N_19981,N_19758);
nor UO_2100 (O_2100,N_19967,N_19623);
nand UO_2101 (O_2101,N_19700,N_19666);
or UO_2102 (O_2102,N_19614,N_19844);
nand UO_2103 (O_2103,N_19721,N_19921);
nand UO_2104 (O_2104,N_19676,N_19926);
xnor UO_2105 (O_2105,N_19659,N_19700);
and UO_2106 (O_2106,N_19924,N_19923);
or UO_2107 (O_2107,N_19886,N_19937);
xnor UO_2108 (O_2108,N_19813,N_19725);
nand UO_2109 (O_2109,N_19844,N_19630);
nor UO_2110 (O_2110,N_19716,N_19907);
and UO_2111 (O_2111,N_19931,N_19994);
and UO_2112 (O_2112,N_19750,N_19942);
and UO_2113 (O_2113,N_19967,N_19885);
and UO_2114 (O_2114,N_19663,N_19840);
nand UO_2115 (O_2115,N_19968,N_19761);
and UO_2116 (O_2116,N_19737,N_19686);
nand UO_2117 (O_2117,N_19891,N_19624);
or UO_2118 (O_2118,N_19963,N_19676);
nor UO_2119 (O_2119,N_19642,N_19692);
xnor UO_2120 (O_2120,N_19891,N_19747);
or UO_2121 (O_2121,N_19733,N_19727);
or UO_2122 (O_2122,N_19975,N_19765);
nand UO_2123 (O_2123,N_19803,N_19798);
nand UO_2124 (O_2124,N_19727,N_19604);
nand UO_2125 (O_2125,N_19713,N_19905);
nand UO_2126 (O_2126,N_19788,N_19899);
nor UO_2127 (O_2127,N_19716,N_19806);
nand UO_2128 (O_2128,N_19722,N_19927);
nand UO_2129 (O_2129,N_19872,N_19846);
xnor UO_2130 (O_2130,N_19660,N_19795);
nand UO_2131 (O_2131,N_19907,N_19926);
nor UO_2132 (O_2132,N_19815,N_19908);
nor UO_2133 (O_2133,N_19801,N_19740);
nand UO_2134 (O_2134,N_19683,N_19767);
xor UO_2135 (O_2135,N_19911,N_19754);
nor UO_2136 (O_2136,N_19960,N_19773);
xnor UO_2137 (O_2137,N_19832,N_19622);
xnor UO_2138 (O_2138,N_19991,N_19685);
xor UO_2139 (O_2139,N_19775,N_19858);
nor UO_2140 (O_2140,N_19811,N_19610);
nand UO_2141 (O_2141,N_19969,N_19715);
xnor UO_2142 (O_2142,N_19845,N_19775);
or UO_2143 (O_2143,N_19675,N_19606);
nand UO_2144 (O_2144,N_19962,N_19885);
and UO_2145 (O_2145,N_19705,N_19737);
xor UO_2146 (O_2146,N_19938,N_19643);
and UO_2147 (O_2147,N_19702,N_19822);
nand UO_2148 (O_2148,N_19858,N_19777);
nor UO_2149 (O_2149,N_19690,N_19934);
xor UO_2150 (O_2150,N_19930,N_19764);
nand UO_2151 (O_2151,N_19865,N_19856);
nand UO_2152 (O_2152,N_19775,N_19889);
xnor UO_2153 (O_2153,N_19877,N_19708);
and UO_2154 (O_2154,N_19772,N_19655);
xnor UO_2155 (O_2155,N_19794,N_19746);
and UO_2156 (O_2156,N_19658,N_19805);
nand UO_2157 (O_2157,N_19927,N_19762);
xor UO_2158 (O_2158,N_19710,N_19731);
nand UO_2159 (O_2159,N_19821,N_19906);
and UO_2160 (O_2160,N_19623,N_19848);
nor UO_2161 (O_2161,N_19917,N_19972);
xor UO_2162 (O_2162,N_19969,N_19702);
xor UO_2163 (O_2163,N_19675,N_19702);
nand UO_2164 (O_2164,N_19795,N_19941);
xnor UO_2165 (O_2165,N_19820,N_19853);
nor UO_2166 (O_2166,N_19967,N_19856);
and UO_2167 (O_2167,N_19689,N_19774);
nor UO_2168 (O_2168,N_19685,N_19812);
or UO_2169 (O_2169,N_19690,N_19831);
nand UO_2170 (O_2170,N_19765,N_19754);
nand UO_2171 (O_2171,N_19983,N_19919);
or UO_2172 (O_2172,N_19756,N_19651);
or UO_2173 (O_2173,N_19805,N_19741);
nand UO_2174 (O_2174,N_19985,N_19712);
xnor UO_2175 (O_2175,N_19715,N_19813);
or UO_2176 (O_2176,N_19714,N_19635);
and UO_2177 (O_2177,N_19695,N_19804);
or UO_2178 (O_2178,N_19964,N_19970);
and UO_2179 (O_2179,N_19670,N_19680);
or UO_2180 (O_2180,N_19792,N_19870);
and UO_2181 (O_2181,N_19645,N_19779);
and UO_2182 (O_2182,N_19954,N_19911);
xor UO_2183 (O_2183,N_19896,N_19679);
xor UO_2184 (O_2184,N_19659,N_19849);
xnor UO_2185 (O_2185,N_19991,N_19868);
xor UO_2186 (O_2186,N_19893,N_19963);
or UO_2187 (O_2187,N_19992,N_19820);
and UO_2188 (O_2188,N_19823,N_19791);
nor UO_2189 (O_2189,N_19952,N_19661);
and UO_2190 (O_2190,N_19624,N_19790);
or UO_2191 (O_2191,N_19981,N_19776);
xnor UO_2192 (O_2192,N_19910,N_19993);
or UO_2193 (O_2193,N_19691,N_19814);
xor UO_2194 (O_2194,N_19653,N_19772);
and UO_2195 (O_2195,N_19985,N_19984);
and UO_2196 (O_2196,N_19808,N_19667);
nor UO_2197 (O_2197,N_19925,N_19846);
xor UO_2198 (O_2198,N_19694,N_19943);
nor UO_2199 (O_2199,N_19705,N_19684);
nor UO_2200 (O_2200,N_19909,N_19677);
xor UO_2201 (O_2201,N_19615,N_19757);
nor UO_2202 (O_2202,N_19680,N_19899);
or UO_2203 (O_2203,N_19923,N_19651);
and UO_2204 (O_2204,N_19909,N_19724);
nand UO_2205 (O_2205,N_19748,N_19747);
or UO_2206 (O_2206,N_19886,N_19601);
nand UO_2207 (O_2207,N_19642,N_19763);
nand UO_2208 (O_2208,N_19693,N_19759);
or UO_2209 (O_2209,N_19954,N_19888);
nand UO_2210 (O_2210,N_19763,N_19911);
xor UO_2211 (O_2211,N_19862,N_19773);
nand UO_2212 (O_2212,N_19699,N_19638);
xor UO_2213 (O_2213,N_19683,N_19746);
or UO_2214 (O_2214,N_19742,N_19709);
or UO_2215 (O_2215,N_19827,N_19613);
xnor UO_2216 (O_2216,N_19921,N_19860);
and UO_2217 (O_2217,N_19828,N_19845);
and UO_2218 (O_2218,N_19838,N_19926);
nor UO_2219 (O_2219,N_19900,N_19936);
xor UO_2220 (O_2220,N_19973,N_19895);
xnor UO_2221 (O_2221,N_19720,N_19821);
and UO_2222 (O_2222,N_19746,N_19660);
nor UO_2223 (O_2223,N_19731,N_19847);
xor UO_2224 (O_2224,N_19761,N_19770);
nor UO_2225 (O_2225,N_19964,N_19642);
xnor UO_2226 (O_2226,N_19716,N_19706);
nor UO_2227 (O_2227,N_19795,N_19653);
nand UO_2228 (O_2228,N_19721,N_19956);
nand UO_2229 (O_2229,N_19997,N_19680);
and UO_2230 (O_2230,N_19750,N_19692);
nor UO_2231 (O_2231,N_19858,N_19722);
and UO_2232 (O_2232,N_19782,N_19603);
or UO_2233 (O_2233,N_19647,N_19920);
xnor UO_2234 (O_2234,N_19906,N_19639);
and UO_2235 (O_2235,N_19607,N_19738);
nor UO_2236 (O_2236,N_19825,N_19944);
or UO_2237 (O_2237,N_19997,N_19947);
xor UO_2238 (O_2238,N_19885,N_19959);
and UO_2239 (O_2239,N_19973,N_19930);
and UO_2240 (O_2240,N_19640,N_19613);
or UO_2241 (O_2241,N_19858,N_19754);
or UO_2242 (O_2242,N_19919,N_19692);
and UO_2243 (O_2243,N_19661,N_19740);
xor UO_2244 (O_2244,N_19918,N_19735);
and UO_2245 (O_2245,N_19942,N_19727);
or UO_2246 (O_2246,N_19662,N_19997);
xnor UO_2247 (O_2247,N_19740,N_19831);
nor UO_2248 (O_2248,N_19866,N_19834);
nor UO_2249 (O_2249,N_19915,N_19991);
nand UO_2250 (O_2250,N_19922,N_19884);
xor UO_2251 (O_2251,N_19723,N_19970);
nor UO_2252 (O_2252,N_19829,N_19672);
and UO_2253 (O_2253,N_19901,N_19757);
nor UO_2254 (O_2254,N_19976,N_19659);
or UO_2255 (O_2255,N_19947,N_19626);
and UO_2256 (O_2256,N_19901,N_19608);
nand UO_2257 (O_2257,N_19768,N_19733);
nand UO_2258 (O_2258,N_19974,N_19973);
nand UO_2259 (O_2259,N_19981,N_19742);
or UO_2260 (O_2260,N_19816,N_19738);
xnor UO_2261 (O_2261,N_19621,N_19825);
nor UO_2262 (O_2262,N_19736,N_19875);
or UO_2263 (O_2263,N_19771,N_19903);
xnor UO_2264 (O_2264,N_19734,N_19923);
and UO_2265 (O_2265,N_19642,N_19818);
or UO_2266 (O_2266,N_19701,N_19755);
xnor UO_2267 (O_2267,N_19640,N_19643);
nor UO_2268 (O_2268,N_19786,N_19799);
nand UO_2269 (O_2269,N_19702,N_19685);
nor UO_2270 (O_2270,N_19799,N_19825);
nand UO_2271 (O_2271,N_19890,N_19976);
xnor UO_2272 (O_2272,N_19921,N_19819);
or UO_2273 (O_2273,N_19955,N_19667);
nor UO_2274 (O_2274,N_19683,N_19910);
xor UO_2275 (O_2275,N_19878,N_19999);
xor UO_2276 (O_2276,N_19687,N_19880);
or UO_2277 (O_2277,N_19828,N_19758);
xnor UO_2278 (O_2278,N_19897,N_19854);
xnor UO_2279 (O_2279,N_19624,N_19850);
nand UO_2280 (O_2280,N_19879,N_19842);
xnor UO_2281 (O_2281,N_19891,N_19696);
nor UO_2282 (O_2282,N_19618,N_19931);
xnor UO_2283 (O_2283,N_19812,N_19667);
nor UO_2284 (O_2284,N_19772,N_19602);
nor UO_2285 (O_2285,N_19864,N_19920);
xor UO_2286 (O_2286,N_19910,N_19712);
or UO_2287 (O_2287,N_19624,N_19841);
and UO_2288 (O_2288,N_19995,N_19760);
or UO_2289 (O_2289,N_19839,N_19970);
xnor UO_2290 (O_2290,N_19933,N_19652);
xor UO_2291 (O_2291,N_19808,N_19647);
and UO_2292 (O_2292,N_19637,N_19753);
and UO_2293 (O_2293,N_19995,N_19733);
xor UO_2294 (O_2294,N_19969,N_19690);
nor UO_2295 (O_2295,N_19818,N_19968);
and UO_2296 (O_2296,N_19754,N_19706);
or UO_2297 (O_2297,N_19613,N_19700);
nand UO_2298 (O_2298,N_19694,N_19851);
xnor UO_2299 (O_2299,N_19905,N_19963);
nor UO_2300 (O_2300,N_19917,N_19939);
nor UO_2301 (O_2301,N_19851,N_19628);
or UO_2302 (O_2302,N_19878,N_19734);
nand UO_2303 (O_2303,N_19690,N_19782);
and UO_2304 (O_2304,N_19932,N_19960);
nor UO_2305 (O_2305,N_19840,N_19747);
nand UO_2306 (O_2306,N_19692,N_19630);
nand UO_2307 (O_2307,N_19883,N_19747);
xnor UO_2308 (O_2308,N_19678,N_19776);
nor UO_2309 (O_2309,N_19779,N_19764);
nor UO_2310 (O_2310,N_19863,N_19857);
nand UO_2311 (O_2311,N_19858,N_19687);
or UO_2312 (O_2312,N_19643,N_19762);
and UO_2313 (O_2313,N_19782,N_19872);
and UO_2314 (O_2314,N_19625,N_19925);
nor UO_2315 (O_2315,N_19673,N_19699);
and UO_2316 (O_2316,N_19605,N_19675);
or UO_2317 (O_2317,N_19859,N_19769);
nor UO_2318 (O_2318,N_19933,N_19945);
xor UO_2319 (O_2319,N_19624,N_19682);
xnor UO_2320 (O_2320,N_19865,N_19754);
nor UO_2321 (O_2321,N_19920,N_19751);
nor UO_2322 (O_2322,N_19655,N_19694);
xnor UO_2323 (O_2323,N_19840,N_19986);
and UO_2324 (O_2324,N_19708,N_19627);
or UO_2325 (O_2325,N_19634,N_19618);
xnor UO_2326 (O_2326,N_19868,N_19821);
xnor UO_2327 (O_2327,N_19693,N_19886);
or UO_2328 (O_2328,N_19633,N_19701);
or UO_2329 (O_2329,N_19792,N_19909);
or UO_2330 (O_2330,N_19695,N_19713);
and UO_2331 (O_2331,N_19770,N_19635);
nor UO_2332 (O_2332,N_19767,N_19914);
xor UO_2333 (O_2333,N_19885,N_19805);
or UO_2334 (O_2334,N_19811,N_19926);
xnor UO_2335 (O_2335,N_19857,N_19919);
xnor UO_2336 (O_2336,N_19778,N_19678);
or UO_2337 (O_2337,N_19635,N_19765);
nand UO_2338 (O_2338,N_19922,N_19758);
nand UO_2339 (O_2339,N_19713,N_19809);
xor UO_2340 (O_2340,N_19860,N_19950);
or UO_2341 (O_2341,N_19741,N_19686);
xnor UO_2342 (O_2342,N_19724,N_19746);
or UO_2343 (O_2343,N_19976,N_19733);
or UO_2344 (O_2344,N_19781,N_19792);
and UO_2345 (O_2345,N_19651,N_19782);
nor UO_2346 (O_2346,N_19991,N_19681);
nor UO_2347 (O_2347,N_19626,N_19718);
or UO_2348 (O_2348,N_19813,N_19844);
or UO_2349 (O_2349,N_19742,N_19786);
and UO_2350 (O_2350,N_19727,N_19654);
xnor UO_2351 (O_2351,N_19903,N_19612);
nand UO_2352 (O_2352,N_19784,N_19764);
and UO_2353 (O_2353,N_19686,N_19710);
nor UO_2354 (O_2354,N_19900,N_19951);
nor UO_2355 (O_2355,N_19847,N_19691);
or UO_2356 (O_2356,N_19958,N_19657);
or UO_2357 (O_2357,N_19897,N_19693);
nor UO_2358 (O_2358,N_19609,N_19667);
and UO_2359 (O_2359,N_19977,N_19981);
nor UO_2360 (O_2360,N_19857,N_19854);
xnor UO_2361 (O_2361,N_19990,N_19605);
nor UO_2362 (O_2362,N_19755,N_19694);
or UO_2363 (O_2363,N_19710,N_19953);
nand UO_2364 (O_2364,N_19624,N_19927);
xor UO_2365 (O_2365,N_19651,N_19790);
nand UO_2366 (O_2366,N_19757,N_19733);
xor UO_2367 (O_2367,N_19603,N_19857);
nand UO_2368 (O_2368,N_19723,N_19724);
or UO_2369 (O_2369,N_19623,N_19889);
nand UO_2370 (O_2370,N_19960,N_19835);
and UO_2371 (O_2371,N_19877,N_19984);
xor UO_2372 (O_2372,N_19999,N_19660);
and UO_2373 (O_2373,N_19616,N_19925);
nand UO_2374 (O_2374,N_19889,N_19709);
and UO_2375 (O_2375,N_19858,N_19702);
and UO_2376 (O_2376,N_19919,N_19654);
nor UO_2377 (O_2377,N_19824,N_19847);
nor UO_2378 (O_2378,N_19744,N_19635);
and UO_2379 (O_2379,N_19705,N_19874);
or UO_2380 (O_2380,N_19975,N_19652);
nor UO_2381 (O_2381,N_19844,N_19943);
and UO_2382 (O_2382,N_19839,N_19877);
and UO_2383 (O_2383,N_19761,N_19928);
and UO_2384 (O_2384,N_19834,N_19892);
or UO_2385 (O_2385,N_19838,N_19633);
nand UO_2386 (O_2386,N_19901,N_19810);
nand UO_2387 (O_2387,N_19932,N_19715);
or UO_2388 (O_2388,N_19685,N_19879);
xor UO_2389 (O_2389,N_19820,N_19849);
nor UO_2390 (O_2390,N_19714,N_19954);
or UO_2391 (O_2391,N_19981,N_19931);
or UO_2392 (O_2392,N_19930,N_19741);
nor UO_2393 (O_2393,N_19964,N_19681);
nand UO_2394 (O_2394,N_19633,N_19870);
nand UO_2395 (O_2395,N_19791,N_19979);
or UO_2396 (O_2396,N_19939,N_19703);
nand UO_2397 (O_2397,N_19676,N_19940);
or UO_2398 (O_2398,N_19669,N_19848);
or UO_2399 (O_2399,N_19964,N_19751);
nand UO_2400 (O_2400,N_19791,N_19619);
xor UO_2401 (O_2401,N_19909,N_19743);
and UO_2402 (O_2402,N_19730,N_19737);
or UO_2403 (O_2403,N_19630,N_19658);
and UO_2404 (O_2404,N_19706,N_19871);
nand UO_2405 (O_2405,N_19821,N_19926);
xor UO_2406 (O_2406,N_19984,N_19977);
and UO_2407 (O_2407,N_19638,N_19719);
or UO_2408 (O_2408,N_19770,N_19818);
xnor UO_2409 (O_2409,N_19688,N_19761);
nand UO_2410 (O_2410,N_19915,N_19837);
nand UO_2411 (O_2411,N_19739,N_19624);
and UO_2412 (O_2412,N_19871,N_19899);
and UO_2413 (O_2413,N_19697,N_19955);
or UO_2414 (O_2414,N_19829,N_19674);
nor UO_2415 (O_2415,N_19646,N_19804);
nand UO_2416 (O_2416,N_19773,N_19649);
and UO_2417 (O_2417,N_19668,N_19924);
nand UO_2418 (O_2418,N_19931,N_19812);
nor UO_2419 (O_2419,N_19699,N_19943);
nor UO_2420 (O_2420,N_19691,N_19888);
nor UO_2421 (O_2421,N_19636,N_19657);
and UO_2422 (O_2422,N_19869,N_19936);
nand UO_2423 (O_2423,N_19912,N_19957);
or UO_2424 (O_2424,N_19869,N_19884);
xnor UO_2425 (O_2425,N_19823,N_19859);
or UO_2426 (O_2426,N_19814,N_19904);
nand UO_2427 (O_2427,N_19625,N_19792);
nor UO_2428 (O_2428,N_19936,N_19609);
nor UO_2429 (O_2429,N_19696,N_19890);
nand UO_2430 (O_2430,N_19611,N_19787);
or UO_2431 (O_2431,N_19677,N_19895);
nand UO_2432 (O_2432,N_19926,N_19602);
or UO_2433 (O_2433,N_19763,N_19678);
nor UO_2434 (O_2434,N_19971,N_19920);
nand UO_2435 (O_2435,N_19857,N_19823);
and UO_2436 (O_2436,N_19892,N_19895);
nand UO_2437 (O_2437,N_19733,N_19994);
nor UO_2438 (O_2438,N_19653,N_19843);
nand UO_2439 (O_2439,N_19994,N_19879);
xnor UO_2440 (O_2440,N_19704,N_19755);
xor UO_2441 (O_2441,N_19716,N_19784);
or UO_2442 (O_2442,N_19762,N_19660);
nor UO_2443 (O_2443,N_19816,N_19962);
xor UO_2444 (O_2444,N_19633,N_19975);
and UO_2445 (O_2445,N_19796,N_19943);
nor UO_2446 (O_2446,N_19888,N_19904);
xor UO_2447 (O_2447,N_19705,N_19614);
or UO_2448 (O_2448,N_19852,N_19661);
nor UO_2449 (O_2449,N_19825,N_19856);
nor UO_2450 (O_2450,N_19662,N_19627);
nand UO_2451 (O_2451,N_19956,N_19754);
and UO_2452 (O_2452,N_19631,N_19975);
or UO_2453 (O_2453,N_19874,N_19724);
or UO_2454 (O_2454,N_19853,N_19864);
nor UO_2455 (O_2455,N_19622,N_19799);
xnor UO_2456 (O_2456,N_19771,N_19908);
and UO_2457 (O_2457,N_19729,N_19946);
xor UO_2458 (O_2458,N_19798,N_19622);
and UO_2459 (O_2459,N_19993,N_19614);
nor UO_2460 (O_2460,N_19972,N_19832);
nand UO_2461 (O_2461,N_19871,N_19698);
xnor UO_2462 (O_2462,N_19780,N_19734);
nor UO_2463 (O_2463,N_19800,N_19732);
and UO_2464 (O_2464,N_19909,N_19796);
nor UO_2465 (O_2465,N_19990,N_19682);
nor UO_2466 (O_2466,N_19803,N_19981);
xnor UO_2467 (O_2467,N_19828,N_19769);
and UO_2468 (O_2468,N_19840,N_19911);
xor UO_2469 (O_2469,N_19760,N_19618);
and UO_2470 (O_2470,N_19875,N_19846);
nand UO_2471 (O_2471,N_19912,N_19605);
or UO_2472 (O_2472,N_19676,N_19912);
or UO_2473 (O_2473,N_19976,N_19951);
nand UO_2474 (O_2474,N_19867,N_19762);
nand UO_2475 (O_2475,N_19798,N_19600);
nand UO_2476 (O_2476,N_19663,N_19668);
xnor UO_2477 (O_2477,N_19826,N_19978);
xnor UO_2478 (O_2478,N_19954,N_19774);
and UO_2479 (O_2479,N_19781,N_19620);
or UO_2480 (O_2480,N_19726,N_19940);
xor UO_2481 (O_2481,N_19623,N_19620);
or UO_2482 (O_2482,N_19602,N_19899);
nand UO_2483 (O_2483,N_19851,N_19633);
xor UO_2484 (O_2484,N_19883,N_19873);
nor UO_2485 (O_2485,N_19732,N_19791);
or UO_2486 (O_2486,N_19882,N_19952);
nand UO_2487 (O_2487,N_19730,N_19648);
nand UO_2488 (O_2488,N_19604,N_19981);
nand UO_2489 (O_2489,N_19867,N_19782);
xnor UO_2490 (O_2490,N_19818,N_19752);
and UO_2491 (O_2491,N_19740,N_19609);
xor UO_2492 (O_2492,N_19809,N_19935);
nand UO_2493 (O_2493,N_19889,N_19624);
and UO_2494 (O_2494,N_19620,N_19915);
nor UO_2495 (O_2495,N_19770,N_19663);
or UO_2496 (O_2496,N_19937,N_19660);
xor UO_2497 (O_2497,N_19652,N_19724);
nand UO_2498 (O_2498,N_19735,N_19882);
and UO_2499 (O_2499,N_19849,N_19722);
endmodule