module basic_2500_25000_3000_4_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19086,N_19087,N_19088,N_19089,N_19090,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19166,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19343,N_19344,N_19345,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19416,N_19417,N_19418,N_19419,N_19420,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19567,N_19568,N_19569,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19804,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19861,N_19862,N_19863,N_19864,N_19865,N_19867,N_19868,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20051,N_20052,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20462,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20610,N_20611,N_20612,N_20613,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20668,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20741,N_20742,N_20743,N_20744,N_20745,N_20747,N_20748,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21091,N_21092,N_21093,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21315,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21830,N_21833,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21863,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22346,N_22347,N_22348,N_22349,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23046,N_23047,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23078,N_23079,N_23080,N_23081,N_23082,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23369,N_23370,N_23371,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23613,N_23614,N_23615,N_23616,N_23618,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23689,N_23690,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23806,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24027,N_24028,N_24029,N_24030,N_24031,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24073,N_24074,N_24075,N_24076,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24190,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24445,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24533,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24565,N_24566,N_24567,N_24568,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24865,N_24866,N_24867,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24998,N_24999;
xor U0 (N_0,In_1810,In_1096);
or U1 (N_1,In_1275,In_9);
nand U2 (N_2,In_1066,In_446);
nor U3 (N_3,In_1381,In_1499);
and U4 (N_4,In_1815,In_89);
nor U5 (N_5,In_138,In_721);
nor U6 (N_6,In_1195,In_706);
and U7 (N_7,In_248,In_1765);
xnor U8 (N_8,In_1780,In_1332);
and U9 (N_9,In_2107,In_1553);
nand U10 (N_10,In_1512,In_1643);
or U11 (N_11,In_2018,In_1683);
nor U12 (N_12,In_389,In_2457);
or U13 (N_13,In_1985,In_1261);
nand U14 (N_14,In_2382,In_1049);
nand U15 (N_15,In_1216,In_2424);
or U16 (N_16,In_1540,In_2489);
or U17 (N_17,In_225,In_561);
xor U18 (N_18,In_1994,In_1671);
or U19 (N_19,In_1743,In_1874);
and U20 (N_20,In_278,In_117);
and U21 (N_21,In_2164,In_1483);
xnor U22 (N_22,In_2269,In_2182);
and U23 (N_23,In_101,In_321);
nand U24 (N_24,In_1674,In_130);
nand U25 (N_25,In_775,In_194);
nand U26 (N_26,In_429,In_370);
xor U27 (N_27,In_73,In_781);
or U28 (N_28,In_322,In_1284);
and U29 (N_29,In_1379,In_2290);
and U30 (N_30,In_2044,In_1238);
or U31 (N_31,In_50,In_2357);
nor U32 (N_32,In_2323,In_2300);
or U33 (N_33,In_590,In_943);
nand U34 (N_34,In_1117,In_698);
xnor U35 (N_35,In_908,In_1647);
and U36 (N_36,In_2062,In_1310);
and U37 (N_37,In_1201,In_1631);
nand U38 (N_38,In_113,In_1413);
nand U39 (N_39,In_399,In_1998);
nor U40 (N_40,In_1670,In_1484);
and U41 (N_41,In_806,In_1489);
nand U42 (N_42,In_975,In_715);
and U43 (N_43,In_1352,In_927);
nor U44 (N_44,In_1878,In_1684);
or U45 (N_45,In_425,In_2230);
and U46 (N_46,In_2003,In_653);
xnor U47 (N_47,In_1896,In_231);
or U48 (N_48,In_1894,In_739);
and U49 (N_49,In_1727,In_795);
nor U50 (N_50,In_944,In_2219);
nand U51 (N_51,In_1158,In_276);
or U52 (N_52,In_818,In_947);
nor U53 (N_53,In_1007,In_2498);
and U54 (N_54,In_286,In_722);
nor U55 (N_55,In_1939,In_1419);
or U56 (N_56,In_1470,In_801);
and U57 (N_57,In_723,In_2169);
nor U58 (N_58,In_1273,In_940);
or U59 (N_59,In_1079,In_666);
nor U60 (N_60,In_957,In_869);
and U61 (N_61,In_1526,In_651);
or U62 (N_62,In_1123,In_1708);
nand U63 (N_63,In_2244,In_346);
nor U64 (N_64,In_77,In_512);
nand U65 (N_65,In_2297,In_470);
nand U66 (N_66,In_240,In_1109);
and U67 (N_67,In_2209,In_137);
nor U68 (N_68,In_1370,In_99);
and U69 (N_69,In_1031,In_334);
nor U70 (N_70,In_1791,In_1229);
nor U71 (N_71,In_526,In_1294);
nor U72 (N_72,In_1303,In_1064);
or U73 (N_73,In_1562,In_308);
nor U74 (N_74,In_100,In_2017);
nand U75 (N_75,In_964,In_2070);
or U76 (N_76,In_1932,In_594);
or U77 (N_77,In_1783,In_931);
and U78 (N_78,In_2406,In_1384);
xnor U79 (N_79,In_491,In_1254);
xor U80 (N_80,In_424,In_1970);
xnor U81 (N_81,In_1607,In_1717);
nand U82 (N_82,In_1445,In_390);
nor U83 (N_83,In_1793,In_1407);
nor U84 (N_84,In_242,In_654);
nand U85 (N_85,In_513,In_460);
or U86 (N_86,In_352,In_1120);
nand U87 (N_87,In_788,In_1172);
nor U88 (N_88,In_1308,In_306);
and U89 (N_89,In_505,In_773);
nand U90 (N_90,In_1431,In_1668);
or U91 (N_91,In_333,In_112);
nand U92 (N_92,In_145,In_1113);
xnor U93 (N_93,In_2069,In_1068);
nand U94 (N_94,In_1637,In_1112);
nand U95 (N_95,In_93,In_216);
or U96 (N_96,In_2061,In_1231);
nand U97 (N_97,In_2354,In_2448);
and U98 (N_98,In_1129,In_391);
xor U99 (N_99,In_1974,In_320);
and U100 (N_100,In_1879,In_1888);
nand U101 (N_101,In_2478,In_1372);
nand U102 (N_102,In_1873,In_1619);
xor U103 (N_103,In_171,In_650);
nand U104 (N_104,In_1258,In_1301);
and U105 (N_105,In_1649,In_522);
and U106 (N_106,In_1136,In_1622);
nor U107 (N_107,In_2117,In_386);
nand U108 (N_108,In_1695,In_1111);
xnor U109 (N_109,In_1623,In_2040);
and U110 (N_110,In_400,In_2309);
or U111 (N_111,In_2405,In_1030);
nand U112 (N_112,In_790,In_1687);
xnor U113 (N_113,In_148,In_886);
and U114 (N_114,In_34,In_1421);
xnor U115 (N_115,In_392,In_374);
nand U116 (N_116,In_459,In_1106);
or U117 (N_117,In_15,In_408);
or U118 (N_118,In_1652,In_1346);
and U119 (N_119,In_335,In_1055);
nor U120 (N_120,In_945,In_1697);
nand U121 (N_121,In_2463,In_665);
nor U122 (N_122,In_1476,In_1980);
and U123 (N_123,In_829,In_1763);
or U124 (N_124,In_973,In_2023);
nand U125 (N_125,In_1130,In_376);
or U126 (N_126,In_246,In_147);
or U127 (N_127,In_398,In_1235);
or U128 (N_128,In_2370,In_1038);
nand U129 (N_129,In_1139,In_191);
or U130 (N_130,In_1203,In_1312);
xor U131 (N_131,In_1906,In_529);
xor U132 (N_132,In_625,In_342);
xor U133 (N_133,In_925,In_874);
nand U134 (N_134,In_1197,In_328);
nand U135 (N_135,In_480,In_559);
xnor U136 (N_136,In_444,In_803);
and U137 (N_137,In_2179,In_2221);
and U138 (N_138,In_903,In_2435);
nand U139 (N_139,In_1853,In_68);
and U140 (N_140,In_877,In_54);
or U141 (N_141,In_2291,In_555);
and U142 (N_142,In_1002,In_1253);
and U143 (N_143,In_208,In_827);
xnor U144 (N_144,In_1336,In_518);
and U145 (N_145,In_2301,In_1367);
nand U146 (N_146,In_1174,In_372);
or U147 (N_147,In_2490,In_1611);
nor U148 (N_148,In_865,In_179);
nor U149 (N_149,In_718,In_2051);
and U150 (N_150,In_441,In_1086);
xor U151 (N_151,In_2317,In_1550);
nand U152 (N_152,In_1321,In_1658);
nand U153 (N_153,In_1971,In_1114);
nor U154 (N_154,In_573,In_437);
xnor U155 (N_155,In_2304,In_2445);
or U156 (N_156,In_633,In_1324);
and U157 (N_157,In_2264,In_736);
or U158 (N_158,In_533,In_1358);
or U159 (N_159,In_2280,In_300);
xnor U160 (N_160,In_2008,In_679);
nor U161 (N_161,In_1406,In_546);
or U162 (N_162,In_747,In_115);
or U163 (N_163,In_1627,In_1462);
or U164 (N_164,In_678,In_1973);
nand U165 (N_165,In_2173,In_2094);
nand U166 (N_166,In_8,In_198);
nor U167 (N_167,In_493,In_65);
and U168 (N_168,In_2054,In_1961);
nor U169 (N_169,In_251,In_139);
and U170 (N_170,In_1916,In_144);
nor U171 (N_171,In_133,In_1871);
nand U172 (N_172,In_1731,In_2263);
nand U173 (N_173,In_1039,In_1048);
nand U174 (N_174,In_1849,In_898);
nand U175 (N_175,In_1983,In_2465);
nor U176 (N_176,In_1377,In_2254);
nor U177 (N_177,In_986,In_445);
and U178 (N_178,In_490,In_1065);
nand U179 (N_179,In_204,In_499);
and U180 (N_180,In_1897,In_2384);
and U181 (N_181,In_1278,In_1991);
nand U182 (N_182,In_1035,In_618);
or U183 (N_183,In_1325,In_929);
nand U184 (N_184,In_2377,In_2134);
and U185 (N_185,In_83,In_1295);
nor U186 (N_186,In_498,In_1778);
or U187 (N_187,In_1914,In_439);
and U188 (N_188,In_541,In_892);
or U189 (N_189,In_1075,In_1771);
nand U190 (N_190,In_2418,In_1577);
nor U191 (N_191,In_956,In_1601);
nor U192 (N_192,In_591,In_223);
or U193 (N_193,In_2315,In_212);
nor U194 (N_194,In_417,In_627);
or U195 (N_195,In_1350,In_2168);
nor U196 (N_196,In_1320,In_2245);
or U197 (N_197,In_2393,In_143);
nand U198 (N_198,In_1507,In_95);
xor U199 (N_199,In_2131,In_1245);
or U200 (N_200,In_2243,In_579);
nand U201 (N_201,In_1036,In_2319);
and U202 (N_202,In_188,In_861);
nand U203 (N_203,In_1584,In_1023);
nand U204 (N_204,In_1248,In_1669);
nor U205 (N_205,In_1576,In_712);
or U206 (N_206,In_2417,In_2242);
or U207 (N_207,In_692,In_1452);
and U208 (N_208,In_72,In_2082);
or U209 (N_209,In_1843,In_946);
and U210 (N_210,In_2262,In_582);
nor U211 (N_211,In_782,In_39);
nand U212 (N_212,In_135,In_291);
nor U213 (N_213,In_1144,In_707);
nor U214 (N_214,In_564,In_1207);
or U215 (N_215,In_2492,In_282);
nor U216 (N_216,In_46,In_482);
nor U217 (N_217,In_2128,In_277);
nor U218 (N_218,In_539,In_436);
nand U219 (N_219,In_1852,In_695);
nor U220 (N_220,In_40,In_1753);
or U221 (N_221,In_634,In_1221);
nand U222 (N_222,In_1872,In_2326);
nor U223 (N_223,In_1742,In_725);
and U224 (N_224,In_1063,In_1967);
nor U225 (N_225,In_911,In_507);
xor U226 (N_226,In_2027,In_1568);
nor U227 (N_227,In_1956,In_2089);
nand U228 (N_228,In_849,In_2225);
and U229 (N_229,In_932,In_870);
or U230 (N_230,In_624,In_1371);
or U231 (N_231,In_1761,In_1756);
or U232 (N_232,In_273,In_1796);
or U233 (N_233,In_2258,In_2096);
and U234 (N_234,In_1428,In_353);
and U235 (N_235,In_2006,In_2389);
nor U236 (N_236,In_2329,In_1861);
nand U237 (N_237,In_716,In_440);
nand U238 (N_238,In_2267,In_1600);
nand U239 (N_239,In_450,In_2476);
and U240 (N_240,In_2350,In_1903);
and U241 (N_241,In_1832,In_981);
nor U242 (N_242,In_2093,In_1713);
nor U243 (N_243,In_2193,In_1556);
nor U244 (N_244,In_2181,In_1001);
or U245 (N_245,In_2019,In_215);
and U246 (N_246,In_511,In_1881);
and U247 (N_247,In_2436,In_1091);
and U248 (N_248,In_2356,In_851);
nor U249 (N_249,In_868,In_14);
nor U250 (N_250,In_1214,In_1281);
or U251 (N_251,In_2004,In_1430);
nand U252 (N_252,In_1220,In_878);
or U253 (N_253,In_1645,In_1736);
or U254 (N_254,In_338,In_1792);
and U255 (N_255,In_686,In_2092);
or U256 (N_256,In_525,In_1538);
and U257 (N_257,In_2285,In_1095);
or U258 (N_258,In_2190,In_2105);
nor U259 (N_259,In_2143,In_833);
and U260 (N_260,In_1465,In_107);
nand U261 (N_261,In_348,In_548);
nand U262 (N_262,In_1898,In_819);
and U263 (N_263,In_1962,In_197);
nand U264 (N_264,In_2325,In_793);
nand U265 (N_265,In_2095,In_662);
or U266 (N_266,In_517,In_2126);
nand U267 (N_267,In_1058,In_1183);
nand U268 (N_268,In_1813,In_1453);
nor U269 (N_269,In_1493,In_70);
or U270 (N_270,In_454,In_229);
and U271 (N_271,In_266,In_2481);
nor U272 (N_272,In_97,In_2375);
nor U273 (N_273,In_356,In_1920);
nor U274 (N_274,In_1648,In_1630);
or U275 (N_275,In_2276,In_2340);
and U276 (N_276,In_1514,In_1348);
nand U277 (N_277,In_677,In_2265);
nor U278 (N_278,In_2125,In_1329);
or U279 (N_279,In_974,In_2238);
nor U280 (N_280,In_2078,In_1901);
nand U281 (N_281,In_1752,In_2239);
nand U282 (N_282,In_982,In_567);
and U283 (N_283,In_1770,In_2011);
nand U284 (N_284,In_2167,In_2275);
and U285 (N_285,In_794,In_1513);
xor U286 (N_286,In_1799,In_1676);
nand U287 (N_287,In_2480,In_1807);
nand U288 (N_288,In_999,In_1490);
xnor U289 (N_289,In_1046,In_2046);
and U290 (N_290,In_1839,In_2332);
nand U291 (N_291,In_1546,In_592);
nand U292 (N_292,In_1388,In_763);
nor U293 (N_293,In_318,In_2100);
nor U294 (N_294,In_2233,In_1076);
nor U295 (N_295,In_2189,In_280);
or U296 (N_296,In_131,In_1262);
nand U297 (N_297,In_2057,In_294);
or U298 (N_298,In_2270,In_655);
and U299 (N_299,In_2091,In_610);
or U300 (N_300,In_1899,In_1338);
and U301 (N_301,In_1527,In_743);
and U302 (N_302,In_1333,In_494);
or U303 (N_303,In_867,In_413);
nor U304 (N_304,In_2113,In_1104);
xnor U305 (N_305,In_2408,In_489);
nor U306 (N_306,In_2076,In_233);
and U307 (N_307,In_740,In_1184);
nand U308 (N_308,In_1167,In_2220);
or U309 (N_309,In_421,In_1252);
or U310 (N_310,In_411,In_1461);
nand U311 (N_311,In_501,In_1996);
nor U312 (N_312,In_1315,In_759);
or U313 (N_313,In_2154,In_761);
nand U314 (N_314,In_641,In_1525);
or U315 (N_315,In_585,In_1578);
nand U316 (N_316,In_1099,In_1927);
or U317 (N_317,In_2266,In_966);
nor U318 (N_318,In_896,In_2183);
nand U319 (N_319,In_1746,In_2240);
nand U320 (N_320,In_866,In_1755);
nand U321 (N_321,In_2009,In_2122);
and U322 (N_322,In_1260,In_405);
or U323 (N_323,In_367,In_1147);
xnor U324 (N_324,In_1784,In_700);
nand U325 (N_325,In_853,In_2344);
nand U326 (N_326,In_2289,In_1682);
nor U327 (N_327,In_2097,In_2214);
xor U328 (N_328,In_362,In_2376);
xnor U329 (N_329,In_2158,In_846);
nor U330 (N_330,In_119,In_1610);
nor U331 (N_331,In_186,In_427);
and U332 (N_332,In_1613,In_2074);
nor U333 (N_333,In_593,In_378);
nand U334 (N_334,In_1923,In_1298);
nor U335 (N_335,In_667,In_449);
or U336 (N_336,In_71,In_58);
or U337 (N_337,In_812,In_547);
nor U338 (N_338,In_735,In_811);
nand U339 (N_339,In_23,In_1467);
nor U340 (N_340,In_1053,In_1842);
or U341 (N_341,In_1660,In_52);
or U342 (N_342,In_176,In_642);
and U343 (N_343,In_1941,In_875);
nand U344 (N_344,In_1869,In_1100);
and U345 (N_345,In_953,In_422);
nor U346 (N_346,In_1327,In_1798);
and U347 (N_347,In_2216,In_1542);
nand U348 (N_348,In_1590,In_719);
nor U349 (N_349,In_871,In_910);
or U350 (N_350,In_1052,In_1171);
nand U351 (N_351,In_954,In_2058);
or U352 (N_352,In_1990,In_497);
and U353 (N_353,In_914,In_1311);
nor U354 (N_354,In_1522,In_2327);
and U355 (N_355,In_1558,In_1270);
nand U356 (N_356,In_2320,In_888);
or U357 (N_357,In_2075,In_1162);
and U358 (N_358,In_837,In_451);
nand U359 (N_359,In_1392,In_2438);
or U360 (N_360,In_1533,In_2161);
nand U361 (N_361,In_523,In_979);
or U362 (N_362,In_952,In_1191);
or U363 (N_363,In_1825,In_385);
xor U364 (N_364,In_1733,In_1767);
and U365 (N_365,In_473,In_984);
nand U366 (N_366,In_1827,In_469);
nand U367 (N_367,In_608,In_183);
xnor U368 (N_368,In_1418,In_2232);
nor U369 (N_369,In_557,In_502);
and U370 (N_370,In_1516,In_488);
nand U371 (N_371,In_521,In_281);
nand U372 (N_372,In_2055,In_1855);
nand U373 (N_373,In_121,In_1892);
and U374 (N_374,In_1887,In_272);
nand U375 (N_375,In_1455,In_2449);
nand U376 (N_376,In_1176,In_1760);
nand U377 (N_377,In_2380,In_174);
or U378 (N_378,In_478,In_160);
nand U379 (N_379,In_2460,In_688);
and U380 (N_380,In_2385,In_500);
or U381 (N_381,In_2403,In_2446);
and U382 (N_382,In_305,In_1164);
and U383 (N_383,In_1151,In_1279);
and U384 (N_384,In_492,In_1547);
nor U385 (N_385,In_1840,In_1360);
nor U386 (N_386,In_2369,In_1921);
nand U387 (N_387,In_2475,In_2022);
nand U388 (N_388,In_2303,In_2293);
nor U389 (N_389,In_855,In_2440);
and U390 (N_390,In_235,In_477);
or U391 (N_391,In_693,In_1933);
xnor U392 (N_392,In_2423,In_1858);
and U393 (N_393,In_433,In_1787);
nand U394 (N_394,In_1240,In_1126);
nor U395 (N_395,In_238,In_600);
nor U396 (N_396,In_638,In_2072);
xor U397 (N_397,In_1188,In_210);
or U398 (N_398,In_1532,In_967);
or U399 (N_399,In_506,In_2170);
or U400 (N_400,In_2390,In_993);
nand U401 (N_401,In_2483,In_339);
and U402 (N_402,In_2123,In_2349);
or U403 (N_403,In_689,In_37);
and U404 (N_404,In_2253,In_622);
nand U405 (N_405,In_456,In_1004);
nand U406 (N_406,In_1378,In_157);
or U407 (N_407,In_1585,In_1965);
nor U408 (N_408,In_2413,In_253);
or U409 (N_409,In_1101,In_181);
and U410 (N_410,In_2462,In_1937);
and U411 (N_411,In_1132,In_1);
nand U412 (N_412,In_1340,In_1276);
nor U413 (N_413,In_2260,In_1444);
and U414 (N_414,In_2016,In_1986);
and U415 (N_415,In_603,In_27);
or U416 (N_416,In_371,In_2177);
nand U417 (N_417,In_1369,In_261);
or U418 (N_418,In_2180,In_172);
nand U419 (N_419,In_122,In_968);
nor U420 (N_420,In_2261,In_2166);
nand U421 (N_421,In_1163,In_1154);
nand U422 (N_422,In_922,In_1434);
nor U423 (N_423,In_909,In_1560);
nor U424 (N_424,In_28,In_341);
nor U425 (N_425,In_336,In_103);
or U426 (N_426,In_1192,In_78);
xnor U427 (N_427,In_1472,In_2141);
or U428 (N_428,In_1289,In_2345);
nor U429 (N_429,In_1219,In_601);
or U430 (N_430,In_1441,In_207);
xor U431 (N_431,In_196,In_168);
and U432 (N_432,In_1711,In_770);
and U433 (N_433,In_1890,In_2295);
or U434 (N_434,In_792,In_1943);
and U435 (N_435,In_1847,In_598);
nand U436 (N_436,In_2336,In_161);
nand U437 (N_437,In_384,In_218);
and U438 (N_438,In_382,In_2084);
nand U439 (N_439,In_1306,In_1543);
or U440 (N_440,In_192,In_520);
nand U441 (N_441,In_2284,In_1387);
or U442 (N_442,In_232,In_76);
nor U443 (N_443,In_1213,In_349);
nor U444 (N_444,In_2472,In_1691);
or U445 (N_445,In_1042,In_1335);
nor U446 (N_446,In_1498,In_1339);
nor U447 (N_447,In_879,In_1215);
nor U448 (N_448,In_124,In_86);
and U449 (N_449,In_1729,In_535);
nand U450 (N_450,In_1963,In_508);
nor U451 (N_451,In_486,In_1644);
and U452 (N_452,In_2373,In_2104);
nand U453 (N_453,In_948,In_859);
or U454 (N_454,In_1491,In_504);
xnor U455 (N_455,In_2132,In_57);
or U456 (N_456,In_1835,In_2223);
or U457 (N_457,In_1605,In_1390);
nand U458 (N_458,In_753,In_1537);
nor U459 (N_459,In_1282,In_1433);
or U460 (N_460,In_1354,In_1364);
or U461 (N_461,In_631,In_1051);
or U462 (N_462,In_836,In_114);
nand U463 (N_463,In_1494,In_2434);
nor U464 (N_464,In_1715,In_1924);
or U465 (N_465,In_2185,In_1889);
or U466 (N_466,In_1698,In_120);
xnor U467 (N_467,In_1021,In_1280);
and U468 (N_468,In_140,In_809);
xnor U469 (N_469,In_2103,In_551);
nand U470 (N_470,In_1876,In_1745);
and U471 (N_471,In_2151,In_2334);
nor U472 (N_472,In_2012,In_1435);
or U473 (N_473,In_1628,In_891);
nand U474 (N_474,In_729,In_538);
nor U475 (N_475,In_2383,In_1447);
nand U476 (N_476,In_269,In_789);
nor U477 (N_477,In_1050,In_10);
xnor U478 (N_478,In_1409,In_767);
nor U479 (N_479,In_2414,In_2218);
nand U480 (N_480,In_862,In_2496);
or U481 (N_481,In_1766,In_1636);
nand U482 (N_482,In_1938,In_1088);
and U483 (N_483,In_1830,In_2030);
or U484 (N_484,In_1680,In_230);
or U485 (N_485,In_2200,In_2400);
and U486 (N_486,In_1081,In_1679);
nand U487 (N_487,In_1833,In_756);
nor U488 (N_488,In_110,In_2404);
or U489 (N_489,In_1177,In_314);
nand U490 (N_490,In_643,In_1383);
and U491 (N_491,In_438,In_2048);
nand U492 (N_492,In_562,In_1999);
and U493 (N_493,In_2355,In_2001);
nor U494 (N_494,In_2379,In_1246);
nor U495 (N_495,In_2176,In_2484);
and U496 (N_496,In_284,In_296);
and U497 (N_497,In_566,In_1561);
nand U498 (N_498,In_375,In_299);
nand U499 (N_499,In_1659,In_1529);
nor U500 (N_500,In_2307,In_2312);
or U501 (N_501,In_416,In_1194);
nor U502 (N_502,In_1015,In_1510);
and U503 (N_503,In_1313,In_193);
and U504 (N_504,In_918,In_2129);
nand U505 (N_505,In_1374,In_2471);
and U506 (N_506,In_254,In_2346);
nor U507 (N_507,In_249,In_381);
nand U508 (N_508,In_676,In_1119);
nor U509 (N_509,In_1653,In_363);
nor U510 (N_510,In_1115,In_1523);
or U511 (N_511,In_2495,In_640);
nor U512 (N_512,In_912,In_732);
nor U513 (N_513,In_1267,In_1782);
nand U514 (N_514,In_2083,In_597);
or U515 (N_515,In_913,In_304);
and U516 (N_516,In_754,In_1808);
xnor U517 (N_517,In_1323,In_1741);
nand U518 (N_518,In_1531,In_899);
nor U519 (N_519,In_1816,In_2066);
nand U520 (N_520,In_626,In_1426);
and U521 (N_521,In_823,In_2042);
xnor U522 (N_522,In_1316,In_1202);
nand U523 (N_523,In_1424,In_1964);
nand U524 (N_524,In_1272,In_158);
and U525 (N_525,In_2392,In_810);
nor U526 (N_526,In_1910,In_798);
nor U527 (N_527,In_2274,In_510);
nand U528 (N_528,In_1851,In_407);
or U529 (N_529,In_1460,In_1149);
or U530 (N_530,In_1632,In_900);
or U531 (N_531,In_466,In_220);
nand U532 (N_532,In_1629,In_487);
nand U533 (N_533,In_2337,In_1777);
and U534 (N_534,In_21,In_2124);
or U535 (N_535,In_1979,In_2228);
nor U536 (N_536,In_574,In_1138);
nor U537 (N_537,In_1210,In_727);
nand U538 (N_538,In_2443,In_1917);
and U539 (N_539,In_528,In_423);
nand U540 (N_540,In_1290,In_1902);
and U541 (N_541,In_2433,In_2045);
and U542 (N_542,In_902,In_1277);
xnor U543 (N_543,In_675,In_1477);
nand U544 (N_544,In_1509,In_2120);
nand U545 (N_545,In_2047,In_2175);
and U546 (N_546,In_1382,In_1948);
nand U547 (N_547,In_60,In_1028);
or U548 (N_548,In_609,In_519);
and U549 (N_549,In_228,In_1223);
and U550 (N_550,In_1580,In_2187);
or U551 (N_551,In_1730,In_1018);
or U552 (N_552,In_289,In_1029);
and U553 (N_553,In_2036,In_628);
nor U554 (N_554,In_1951,In_937);
nand U555 (N_555,In_1414,In_332);
and U556 (N_556,In_1408,In_2039);
nand U557 (N_557,In_1122,In_1738);
or U558 (N_558,In_1893,In_2364);
nand U559 (N_559,In_1818,In_184);
nor U560 (N_560,In_2281,In_1685);
nand U561 (N_561,In_369,In_0);
nand U562 (N_562,In_2116,In_1234);
or U563 (N_563,In_485,In_1694);
or U564 (N_564,In_1978,In_1618);
and U565 (N_565,In_1304,In_1166);
nor U566 (N_566,In_495,In_983);
and U567 (N_567,In_1700,In_1193);
or U568 (N_568,In_1182,In_1355);
nor U569 (N_569,In_1487,In_1451);
nand U570 (N_570,In_2279,In_1779);
or U571 (N_571,In_383,In_2425);
nor U572 (N_572,In_2178,In_558);
nand U573 (N_573,In_1400,In_2156);
or U574 (N_574,In_2049,In_224);
nand U575 (N_575,In_1972,In_1586);
nand U576 (N_576,In_2160,In_1740);
xor U577 (N_577,In_669,In_1161);
and U578 (N_578,In_2137,In_623);
and U579 (N_579,In_129,In_164);
nand U580 (N_580,In_1775,In_728);
nor U581 (N_581,In_1178,In_1581);
and U582 (N_582,In_2186,In_542);
and U583 (N_583,In_2399,In_1774);
xor U584 (N_584,In_1479,In_62);
xnor U585 (N_585,In_1639,In_1069);
or U586 (N_586,In_1721,In_1222);
nand U587 (N_587,In_720,In_1153);
nor U588 (N_588,In_1054,In_247);
or U589 (N_589,In_1094,In_1987);
nor U590 (N_590,In_757,In_1722);
and U591 (N_591,In_1809,In_569);
nand U592 (N_592,In_412,In_153);
nand U593 (N_593,In_1988,In_169);
nand U594 (N_594,In_1661,In_1506);
and U595 (N_595,In_319,In_784);
xor U596 (N_596,In_1877,In_302);
and U597 (N_597,In_167,In_257);
xor U598 (N_598,In_1173,In_1353);
nor U599 (N_599,In_962,In_315);
or U600 (N_600,In_831,In_1189);
nor U601 (N_601,In_361,In_1286);
xor U602 (N_602,In_344,In_2410);
nand U603 (N_603,In_704,In_572);
nor U604 (N_604,In_1573,In_347);
and U605 (N_605,In_2226,In_31);
or U606 (N_606,In_769,In_1398);
nor U607 (N_607,In_1909,In_617);
and U608 (N_608,In_2427,In_1087);
or U609 (N_609,In_1366,In_1198);
or U610 (N_610,In_324,In_2077);
or U611 (N_611,In_1781,In_1212);
or U612 (N_612,In_1226,In_2237);
and U613 (N_613,In_1084,In_20);
or U614 (N_614,In_1411,In_475);
or U615 (N_615,In_1067,In_1402);
nand U616 (N_616,In_1615,In_530);
nand U617 (N_617,In_1342,In_1690);
nor U618 (N_618,In_1891,In_2338);
or U619 (N_619,In_1157,In_2038);
nor U620 (N_620,In_2172,In_1912);
nand U621 (N_621,In_1635,In_1608);
or U622 (N_622,In_1218,In_1412);
or U623 (N_623,In_397,In_1922);
or U624 (N_624,In_990,In_1768);
nor U625 (N_625,In_1751,In_1875);
nand U626 (N_626,In_992,In_1341);
and U627 (N_627,In_2255,In_1846);
and U628 (N_628,In_1057,In_1656);
and U629 (N_629,In_1199,In_2318);
or U630 (N_630,In_209,In_7);
and U631 (N_631,In_1318,In_42);
and U632 (N_632,In_271,In_2060);
xnor U633 (N_633,In_1952,In_684);
and U634 (N_634,In_1061,In_1037);
or U635 (N_635,In_1145,In_2163);
and U636 (N_636,In_2155,In_1127);
or U637 (N_637,In_1307,In_1380);
or U638 (N_638,In_858,In_496);
nand U639 (N_639,In_2114,In_2111);
nor U640 (N_640,In_1592,In_1588);
nand U641 (N_641,In_2451,In_2374);
or U642 (N_642,In_942,In_1621);
nor U643 (N_643,In_1293,In_2468);
nand U644 (N_644,In_1720,In_796);
and U645 (N_645,In_2466,In_379);
xor U646 (N_646,In_47,In_1391);
and U647 (N_647,In_1975,In_1473);
nand U648 (N_648,In_2493,In_848);
and U649 (N_649,In_1299,In_1739);
nor U650 (N_650,In_1517,In_279);
nand U651 (N_651,In_2195,In_800);
nor U652 (N_652,In_738,In_649);
nor U653 (N_653,In_53,In_354);
nor U654 (N_654,In_1143,In_1397);
xor U655 (N_655,In_1232,In_1135);
or U656 (N_656,In_619,In_102);
xor U657 (N_657,In_18,In_199);
or U658 (N_658,In_467,In_1968);
and U659 (N_659,In_755,In_2294);
or U660 (N_660,In_2050,In_751);
and U661 (N_661,In_19,In_2333);
xor U662 (N_662,In_2442,In_663);
or U663 (N_663,In_1170,In_1884);
and U664 (N_664,In_2416,In_1326);
nor U665 (N_665,In_442,In_2347);
nand U666 (N_666,In_443,In_1440);
and U667 (N_667,In_1363,In_373);
or U668 (N_668,In_462,In_994);
nand U669 (N_669,In_1860,In_1425);
nand U670 (N_670,In_668,In_1822);
and U671 (N_671,In_163,In_1929);
nand U672 (N_672,In_2056,In_69);
nor U673 (N_673,In_1870,In_1757);
and U674 (N_674,In_465,In_1624);
or U675 (N_675,In_926,In_816);
or U676 (N_676,In_1569,In_1186);
and U677 (N_677,In_760,In_258);
nand U678 (N_678,In_2035,In_934);
nor U679 (N_679,In_1187,In_1505);
xor U680 (N_680,In_1105,In_856);
nand U681 (N_681,In_29,In_1257);
nand U682 (N_682,In_893,In_635);
and U683 (N_683,In_1150,In_1692);
and U684 (N_684,In_2272,In_394);
or U685 (N_685,In_2352,In_2079);
nor U686 (N_686,In_2415,In_845);
nand U687 (N_687,In_310,In_1142);
or U688 (N_688,In_1667,In_1657);
and U689 (N_689,In_758,In_1185);
nor U690 (N_690,In_2162,In_2247);
nor U691 (N_691,In_1895,In_1723);
and U692 (N_692,In_2296,In_1070);
nor U693 (N_693,In_1949,In_1155);
or U694 (N_694,In_1124,In_637);
and U695 (N_695,In_589,In_1609);
xnor U696 (N_696,In_2387,In_2007);
or U697 (N_697,In_772,In_629);
nand U698 (N_698,In_890,In_1944);
nand U699 (N_699,In_1675,In_415);
nor U700 (N_700,In_1982,In_997);
or U701 (N_701,In_67,In_1663);
nand U702 (N_702,In_435,In_345);
nand U703 (N_703,In_84,In_474);
nor U704 (N_704,In_537,In_1020);
or U705 (N_705,In_109,In_1626);
or U706 (N_706,In_2064,In_825);
or U707 (N_707,In_1131,In_998);
xnor U708 (N_708,In_881,In_1966);
xor U709 (N_709,In_1865,In_1828);
xor U710 (N_710,In_189,In_1528);
and U711 (N_711,In_1693,In_938);
or U712 (N_712,In_2488,In_578);
nor U713 (N_713,In_458,In_2429);
xor U714 (N_714,In_2395,In_1259);
and U715 (N_715,In_1612,In_1175);
and U716 (N_716,In_2106,In_1714);
nand U717 (N_717,In_1137,In_1848);
nand U718 (N_718,In_1217,In_985);
nand U719 (N_719,In_1249,In_1583);
xnor U720 (N_720,In_841,In_410);
xnor U721 (N_721,In_1373,In_1801);
nor U722 (N_722,In_1181,In_1469);
or U723 (N_723,In_1224,In_340);
nor U724 (N_724,In_1365,In_1134);
nand U725 (N_725,In_1314,In_1650);
nor U726 (N_726,In_190,In_141);
nor U727 (N_727,In_2014,In_690);
nor U728 (N_728,In_1032,In_1959);
and U729 (N_729,In_2299,In_1750);
nand U730 (N_730,In_916,In_2298);
nor U731 (N_731,In_1496,In_1417);
nor U732 (N_732,In_1518,In_2188);
nor U733 (N_733,In_309,In_13);
nand U734 (N_734,In_847,In_905);
and U735 (N_735,In_152,In_307);
xor U736 (N_736,In_2394,In_250);
nand U737 (N_737,In_2150,In_1376);
and U738 (N_738,In_1043,In_928);
nor U739 (N_739,In_2127,In_388);
nor U740 (N_740,In_1347,In_298);
nand U741 (N_741,In_214,In_481);
and U742 (N_742,In_901,In_1022);
nand U743 (N_743,In_1439,In_1749);
or U744 (N_744,In_431,In_1911);
nor U745 (N_745,In_1554,In_2165);
nand U746 (N_746,In_1786,In_1758);
or U747 (N_747,In_59,In_2198);
nand U748 (N_748,In_2447,In_419);
or U749 (N_749,In_2241,In_1570);
and U750 (N_750,In_155,In_750);
and U751 (N_751,In_56,In_705);
nand U752 (N_752,In_1803,In_1824);
nor U753 (N_753,In_1291,In_426);
nand U754 (N_754,In_2479,In_1640);
or U755 (N_755,In_1190,In_1389);
nand U756 (N_756,In_1090,In_4);
and U757 (N_757,In_857,In_1744);
and U758 (N_758,In_404,In_2053);
and U759 (N_759,In_1928,In_358);
and U760 (N_760,In_2494,In_696);
or U761 (N_761,In_1625,In_2184);
nor U762 (N_762,In_2130,In_387);
or U763 (N_763,In_2021,In_1501);
nand U764 (N_764,In_461,In_288);
xnor U765 (N_765,In_930,In_292);
or U766 (N_766,In_1934,In_660);
and U767 (N_767,In_515,In_907);
or U768 (N_768,In_2464,In_351);
or U769 (N_769,In_1458,In_1269);
nand U770 (N_770,In_2286,In_1977);
nand U771 (N_771,In_17,In_1169);
xor U772 (N_772,In_252,In_2153);
nor U773 (N_773,In_2,In_1776);
or U774 (N_774,In_1545,In_2353);
and U775 (N_775,In_98,In_553);
nand U776 (N_776,In_799,In_503);
nand U777 (N_777,In_1012,In_826);
and U778 (N_778,In_1854,In_1646);
nor U779 (N_779,In_2080,In_2453);
and U780 (N_780,In_749,In_989);
and U781 (N_781,In_51,In_726);
nand U782 (N_782,In_1593,In_2041);
and U783 (N_783,In_1200,In_2450);
and U784 (N_784,In_1908,In_2378);
nor U785 (N_785,In_1582,In_1802);
nand U786 (N_786,In_1283,In_2157);
nand U787 (N_787,In_1475,In_1571);
nor U788 (N_788,In_2013,In_920);
or U789 (N_789,In_1085,In_2217);
nor U790 (N_790,In_835,In_1534);
nor U791 (N_791,In_2068,In_434);
nand U792 (N_792,In_1880,In_1836);
nand U793 (N_793,In_1686,In_329);
nand U794 (N_794,In_917,In_1572);
and U795 (N_795,In_154,In_2135);
nor U796 (N_796,In_1337,In_1019);
nand U797 (N_797,In_1436,In_904);
and U798 (N_798,In_1204,In_2231);
nor U799 (N_799,In_2420,In_285);
or U800 (N_800,In_813,In_1797);
nand U801 (N_801,In_452,In_237);
nor U802 (N_802,In_1344,In_245);
and U803 (N_803,In_403,In_534);
nand U804 (N_804,In_1712,In_357);
nand U805 (N_805,In_2149,In_1551);
xor U806 (N_806,In_55,In_2331);
and U807 (N_807,In_1082,In_2205);
nand U808 (N_808,In_1850,In_85);
and U809 (N_809,In_312,In_1826);
and U810 (N_810,In_1319,In_822);
or U811 (N_811,In_1947,In_1602);
nand U812 (N_812,In_1255,In_1466);
and U813 (N_813,In_2419,In_2313);
or U814 (N_814,In_2067,In_1041);
and U815 (N_815,In_35,In_2222);
or U816 (N_816,In_303,In_766);
and U817 (N_817,In_648,In_804);
nor U818 (N_818,In_1225,In_2052);
and U819 (N_819,In_863,In_2441);
xor U820 (N_820,In_748,In_1829);
or U821 (N_821,In_1102,In_1432);
nand U822 (N_822,In_1287,In_1564);
or U823 (N_823,In_1256,In_268);
and U824 (N_824,In_2085,In_2234);
and U825 (N_825,In_1266,In_25);
and U826 (N_826,In_1343,In_1118);
or U827 (N_827,In_1415,In_1945);
nor U828 (N_828,In_1997,In_1396);
or U829 (N_829,In_325,In_2112);
nor U830 (N_830,In_2032,In_1958);
nand U831 (N_831,In_448,In_864);
or U832 (N_832,In_737,In_2409);
and U833 (N_833,In_808,In_694);
xnor U834 (N_834,In_2037,In_317);
or U835 (N_835,In_1709,In_1725);
and U836 (N_836,In_1841,In_1013);
or U837 (N_837,In_2063,In_187);
and U838 (N_838,In_996,In_1361);
nor U839 (N_839,In_1905,In_1005);
and U840 (N_840,In_1575,In_1056);
nand U841 (N_841,In_2371,In_1241);
and U842 (N_842,In_699,In_1940);
and U843 (N_843,In_418,In_1662);
and U844 (N_844,In_664,In_1764);
nor U845 (N_845,In_1014,In_1093);
nand U846 (N_846,In_1206,In_1699);
nand U847 (N_847,In_26,In_524);
xnor U848 (N_848,In_2366,In_2470);
or U849 (N_849,In_681,In_134);
nand U850 (N_850,In_1495,In_2236);
nor U851 (N_851,In_1008,In_1179);
nor U852 (N_852,In_746,In_12);
or U853 (N_853,In_1478,In_834);
and U854 (N_854,In_2196,In_2026);
and U855 (N_855,In_359,In_1817);
or U856 (N_856,In_393,In_1706);
nand U857 (N_857,In_1555,In_205);
and U858 (N_858,In_239,In_2381);
nor U859 (N_859,In_1500,In_396);
nand U860 (N_860,In_565,In_2020);
or U861 (N_861,In_1811,In_177);
and U862 (N_862,In_1953,In_36);
nand U863 (N_863,In_323,In_2499);
or U864 (N_864,In_2250,In_606);
nand U865 (N_865,In_1747,In_2043);
nor U866 (N_866,In_2454,In_283);
or U867 (N_867,In_2034,In_1665);
nor U868 (N_868,In_2439,In_6);
and U869 (N_869,In_1734,In_2401);
and U870 (N_870,In_1448,In_791);
xnor U871 (N_871,In_876,In_1482);
nand U872 (N_872,In_1485,In_1399);
nand U873 (N_873,In_621,In_1265);
nand U874 (N_874,In_1357,In_1579);
nor U875 (N_875,In_243,In_1394);
nand U876 (N_876,In_1773,In_1521);
and U877 (N_877,In_326,In_1559);
and U878 (N_878,In_939,In_43);
nand U879 (N_879,In_175,In_1140);
and U880 (N_880,In_1651,In_2287);
or U881 (N_881,In_1040,In_1160);
xor U882 (N_882,In_762,In_882);
nand U883 (N_883,In_2088,In_3);
nor U884 (N_884,In_104,In_1351);
and U885 (N_885,In_645,In_90);
or U886 (N_886,In_2306,In_2109);
or U887 (N_887,In_1420,In_1672);
or U888 (N_888,In_96,In_1450);
xnor U889 (N_889,In_2302,In_995);
nand U890 (N_890,In_195,In_2015);
and U891 (N_891,In_219,In_1930);
or U892 (N_892,In_1772,In_1401);
or U893 (N_893,In_1121,In_586);
nand U894 (N_894,In_1486,In_1196);
or U895 (N_895,In_2098,In_752);
or U896 (N_896,In_1634,In_568);
nor U897 (N_897,In_1103,In_105);
or U898 (N_898,In_527,In_543);
nand U899 (N_899,In_1474,In_267);
or U900 (N_900,In_588,In_976);
nor U901 (N_901,In_1960,In_24);
nand U902 (N_902,In_768,In_178);
nand U903 (N_903,In_264,In_647);
xnor U904 (N_904,In_2115,In_1574);
and U905 (N_905,In_1097,In_1606);
or U906 (N_906,In_1976,In_75);
or U907 (N_907,In_430,In_2486);
nand U908 (N_908,In_2108,In_1957);
nor U909 (N_909,In_406,In_646);
nor U910 (N_910,In_1702,In_670);
and U911 (N_911,In_48,In_2213);
nand U912 (N_912,In_343,In_575);
nand U913 (N_913,In_1701,In_1511);
nand U914 (N_914,In_1566,In_1003);
nand U915 (N_915,In_969,In_74);
xnor U916 (N_916,In_1904,In_2458);
and U917 (N_917,In_1011,In_2485);
and U918 (N_918,In_221,In_509);
and U919 (N_919,In_2133,In_1305);
and U920 (N_920,In_2421,In_965);
xnor U921 (N_921,In_2324,In_301);
nor U922 (N_922,In_2311,In_659);
nand U923 (N_923,In_532,In_1705);
nor U924 (N_924,In_1642,In_1823);
and U925 (N_925,In_889,In_1244);
and U926 (N_926,In_2292,In_1754);
nor U927 (N_927,In_2144,In_1589);
nand U928 (N_928,In_2206,In_797);
nand U929 (N_929,In_584,In_1268);
and U930 (N_930,In_1805,In_571);
and U931 (N_931,In_1520,In_1641);
or U932 (N_932,In_1393,In_612);
nand U933 (N_933,In_1769,In_1654);
and U934 (N_934,In_2073,In_1925);
and U935 (N_935,In_978,In_41);
xnor U936 (N_936,In_2199,In_839);
and U937 (N_937,In_364,In_1993);
and U938 (N_938,In_1356,In_81);
and U939 (N_939,In_1867,In_779);
nand U940 (N_940,In_457,In_873);
and U941 (N_941,In_265,In_2257);
nor U942 (N_942,In_1969,In_1302);
xnor U943 (N_943,In_1107,In_2487);
and U944 (N_944,In_1228,In_132);
and U945 (N_945,In_1604,In_1205);
xor U946 (N_946,In_843,In_1718);
or U947 (N_947,In_2467,In_1638);
nand U948 (N_948,In_1159,In_94);
nor U949 (N_949,In_1673,In_1616);
or U950 (N_950,In_1614,In_1541);
or U951 (N_951,In_2090,In_88);
and U952 (N_952,In_1116,In_1108);
nor U953 (N_953,In_1704,In_1557);
and U954 (N_954,In_2282,In_733);
nand U955 (N_955,In_1098,In_2372);
nor U956 (N_956,In_1696,In_685);
nand U957 (N_957,In_1735,In_297);
or U958 (N_958,In_2086,In_933);
xnor U959 (N_959,In_1524,In_958);
or U960 (N_960,In_2407,In_701);
and U961 (N_961,In_630,In_2339);
nand U962 (N_962,In_783,In_661);
nand U963 (N_963,In_2273,In_2396);
nand U964 (N_964,In_2367,In_2412);
nand U965 (N_965,In_2147,In_850);
and U966 (N_966,In_1395,In_126);
and U967 (N_967,In_1868,In_1535);
nand U968 (N_968,In_484,In_1863);
or U969 (N_969,In_1819,In_173);
nand U970 (N_970,In_2071,In_2469);
nand U971 (N_971,In_1587,In_977);
nand U972 (N_972,In_1033,In_516);
and U973 (N_973,In_1317,In_1732);
xnor U974 (N_974,In_2343,In_1125);
nor U975 (N_975,In_840,In_570);
nand U976 (N_976,In_1862,In_1942);
nor U977 (N_977,In_1918,In_146);
nand U978 (N_978,In_674,In_1502);
nand U979 (N_979,In_380,In_402);
or U980 (N_980,In_1328,In_786);
nand U981 (N_981,In_1236,In_514);
or U982 (N_982,In_1857,In_91);
and U983 (N_983,In_170,In_1285);
nor U984 (N_984,In_1247,In_79);
nand U985 (N_985,In_1047,In_936);
xnor U986 (N_986,In_1913,In_1530);
and U987 (N_987,In_832,In_2174);
nand U988 (N_988,In_709,In_852);
and U989 (N_989,In_2246,In_549);
or U990 (N_990,In_1504,In_2171);
nor U991 (N_991,In_1045,In_327);
and U992 (N_992,In_49,In_395);
or U993 (N_993,In_2251,In_2002);
nor U994 (N_994,In_365,In_1464);
and U995 (N_995,In_2335,In_1405);
nor U996 (N_996,In_531,In_1984);
and U997 (N_997,In_1885,In_1027);
xor U998 (N_998,In_2455,In_2087);
or U999 (N_999,In_1385,In_162);
and U1000 (N_1000,In_713,In_217);
nor U1001 (N_1001,In_2000,In_897);
nand U1002 (N_1002,In_180,In_652);
or U1003 (N_1003,In_293,In_360);
nand U1004 (N_1004,In_1955,In_256);
nand U1005 (N_1005,In_255,In_1026);
and U1006 (N_1006,In_259,In_2229);
xor U1007 (N_1007,In_596,In_780);
and U1008 (N_1008,In_1821,In_1233);
nand U1009 (N_1009,In_1790,In_1017);
nand U1010 (N_1010,In_1034,In_61);
nand U1011 (N_1011,In_724,In_1362);
or U1012 (N_1012,In_587,In_1762);
nor U1013 (N_1013,In_607,In_1438);
nor U1014 (N_1014,In_2191,In_2397);
xor U1015 (N_1015,In_2328,In_377);
nor U1016 (N_1016,In_2215,In_2031);
or U1017 (N_1017,In_200,In_1083);
nor U1018 (N_1018,In_1719,In_1156);
nor U1019 (N_1019,In_2033,In_1073);
nand U1020 (N_1020,In_1345,In_2025);
nand U1021 (N_1021,In_463,In_2314);
nor U1022 (N_1022,In_2146,In_1006);
nor U1023 (N_1023,In_1845,In_988);
nor U1024 (N_1024,In_540,In_2361);
nand U1025 (N_1025,In_1148,In_702);
nor U1026 (N_1026,In_577,In_1900);
nand U1027 (N_1027,In_602,In_1515);
or U1028 (N_1028,In_331,In_1292);
nor U1029 (N_1029,In_234,In_1443);
nand U1030 (N_1030,In_2431,In_1788);
nand U1031 (N_1031,In_714,In_1536);
and U1032 (N_1032,In_708,In_895);
nor U1033 (N_1033,In_906,In_1025);
nand U1034 (N_1034,In_149,In_764);
or U1035 (N_1035,In_2028,In_2152);
xor U1036 (N_1036,In_1071,In_151);
and U1037 (N_1037,In_2192,In_1812);
nor U1038 (N_1038,In_45,In_671);
xnor U1039 (N_1039,In_2010,In_1468);
nor U1040 (N_1040,In_884,In_1165);
and U1041 (N_1041,In_1503,In_872);
nand U1042 (N_1042,In_1565,In_2432);
xnor U1043 (N_1043,In_316,In_1681);
or U1044 (N_1044,In_1598,In_550);
nand U1045 (N_1045,In_260,In_1309);
nand U1046 (N_1046,In_1457,In_1263);
and U1047 (N_1047,In_711,In_745);
nand U1048 (N_1048,In_125,In_2391);
nand U1049 (N_1049,In_182,In_2248);
and U1050 (N_1050,In_915,In_128);
nand U1051 (N_1051,In_2308,In_468);
nor U1052 (N_1052,In_2101,In_1707);
xor U1053 (N_1053,In_2110,In_241);
nor U1054 (N_1054,In_2360,In_1010);
xnor U1055 (N_1055,In_805,In_1242);
nand U1056 (N_1056,In_1250,In_1331);
or U1057 (N_1057,In_1655,In_1080);
xnor U1058 (N_1058,In_1375,In_581);
nor U1059 (N_1059,In_778,In_2099);
nand U1060 (N_1060,In_453,In_595);
or U1061 (N_1061,In_1062,In_2477);
nor U1062 (N_1062,In_1954,In_330);
nand U1063 (N_1063,In_1322,In_2426);
and U1064 (N_1064,In_2197,In_580);
nor U1065 (N_1065,In_1989,In_949);
nor U1066 (N_1066,In_991,In_166);
nand U1067 (N_1067,In_1437,In_111);
nand U1068 (N_1068,In_82,In_142);
xnor U1069 (N_1069,In_2305,In_1422);
nand U1070 (N_1070,In_1992,In_1617);
and U1071 (N_1071,In_2388,In_2456);
xnor U1072 (N_1072,In_414,In_213);
or U1073 (N_1073,In_1678,In_854);
and U1074 (N_1074,In_1716,In_1243);
and U1075 (N_1075,In_2005,In_2411);
xnor U1076 (N_1076,In_1935,In_1508);
and U1077 (N_1077,In_2491,In_961);
nand U1078 (N_1078,In_366,In_1404);
nor U1079 (N_1079,In_552,In_1563);
nand U1080 (N_1080,In_1519,In_2252);
nor U1081 (N_1081,In_2227,In_1995);
nand U1082 (N_1082,In_771,In_1077);
or U1083 (N_1083,In_1146,In_118);
xnor U1084 (N_1084,In_1603,In_80);
xnor U1085 (N_1085,In_1427,In_1688);
nand U1086 (N_1086,In_1208,In_830);
and U1087 (N_1087,In_563,In_807);
nor U1088 (N_1088,In_355,In_313);
and U1089 (N_1089,In_1710,In_22);
and U1090 (N_1090,In_1794,In_203);
or U1091 (N_1091,In_222,In_1009);
nand U1092 (N_1092,In_262,In_2102);
nand U1093 (N_1093,In_63,In_1059);
xor U1094 (N_1094,In_2348,In_842);
and U1095 (N_1095,In_44,In_1806);
nand U1096 (N_1096,In_1737,In_290);
nor U1097 (N_1097,In_2459,In_2359);
nor U1098 (N_1098,In_287,In_644);
or U1099 (N_1099,In_656,In_741);
nand U1100 (N_1100,In_2208,In_476);
xnor U1101 (N_1101,In_1595,In_2422);
nor U1102 (N_1102,In_683,In_127);
nor U1103 (N_1103,In_821,In_1946);
xnor U1104 (N_1104,In_87,In_1463);
nand U1105 (N_1105,In_1981,In_824);
or U1106 (N_1106,In_1837,In_885);
and U1107 (N_1107,In_1168,In_1359);
and U1108 (N_1108,In_1591,In_2386);
and U1109 (N_1109,In_2139,In_447);
nand U1110 (N_1110,In_1844,In_1423);
or U1111 (N_1111,In_2368,In_464);
or U1112 (N_1112,In_1297,In_66);
and U1113 (N_1113,In_1831,In_2024);
and U1114 (N_1114,In_963,In_2118);
nor U1115 (N_1115,In_1368,In_2259);
or U1116 (N_1116,In_1789,In_2202);
and U1117 (N_1117,In_1481,In_64);
or U1118 (N_1118,In_2497,In_2310);
or U1119 (N_1119,In_894,In_2316);
nor U1120 (N_1120,In_1211,In_1859);
nand U1121 (N_1121,In_941,In_270);
nand U1122 (N_1122,In_632,In_202);
or U1123 (N_1123,In_2342,In_959);
nor U1124 (N_1124,In_2437,In_935);
and U1125 (N_1125,In_1677,In_1800);
and U1126 (N_1126,In_960,In_1334);
nor U1127 (N_1127,In_583,In_2119);
nor U1128 (N_1128,In_604,In_1548);
or U1129 (N_1129,In_672,In_883);
or U1130 (N_1130,In_923,In_2452);
or U1131 (N_1131,In_2428,In_2029);
nor U1132 (N_1132,In_2201,In_734);
or U1133 (N_1133,In_33,In_1024);
or U1134 (N_1134,In_1016,In_880);
and U1135 (N_1135,In_1931,In_2235);
and U1136 (N_1136,In_838,In_970);
and U1137 (N_1137,In_1386,In_2365);
or U1138 (N_1138,In_1666,In_2207);
and U1139 (N_1139,In_2362,In_951);
nand U1140 (N_1140,In_311,In_2398);
nor U1141 (N_1141,In_2277,In_150);
or U1142 (N_1142,In_401,In_1092);
or U1143 (N_1143,In_1748,In_1227);
nand U1144 (N_1144,In_2204,In_32);
xor U1145 (N_1145,In_1907,In_980);
or U1146 (N_1146,In_1230,In_185);
or U1147 (N_1147,In_2081,In_420);
nor U1148 (N_1148,In_1429,In_1544);
and U1149 (N_1149,In_201,In_1454);
xor U1150 (N_1150,In_658,In_1834);
nor U1151 (N_1151,In_2211,In_817);
nor U1152 (N_1152,In_2203,In_1403);
and U1153 (N_1153,In_1856,In_455);
nor U1154 (N_1154,In_244,In_776);
xor U1155 (N_1155,In_554,In_844);
xnor U1156 (N_1156,In_1000,In_673);
and U1157 (N_1157,In_16,In_350);
and U1158 (N_1158,In_1446,In_2363);
nand U1159 (N_1159,In_1795,In_1060);
nand U1160 (N_1160,In_2402,In_717);
or U1161 (N_1161,In_2474,In_2444);
nor U1162 (N_1162,In_2212,In_1209);
or U1163 (N_1163,In_814,In_1152);
and U1164 (N_1164,In_211,In_1724);
or U1165 (N_1165,In_1471,In_613);
or U1166 (N_1166,In_697,In_972);
nor U1167 (N_1167,In_615,In_815);
or U1168 (N_1168,In_1237,In_1620);
and U1169 (N_1169,In_1110,In_1689);
nor U1170 (N_1170,In_2142,In_1567);
and U1171 (N_1171,In_2283,In_1074);
nand U1172 (N_1172,In_2268,In_471);
and U1173 (N_1173,In_409,In_1497);
nor U1174 (N_1174,In_2322,In_1349);
nor U1175 (N_1175,In_616,In_576);
nand U1176 (N_1176,In_1883,In_5);
and U1177 (N_1177,In_1133,In_1814);
nand U1178 (N_1178,In_687,In_2159);
nand U1179 (N_1179,In_1330,In_1410);
or U1180 (N_1180,In_785,In_703);
or U1181 (N_1181,In_765,In_428);
and U1182 (N_1182,In_1596,In_368);
nor U1183 (N_1183,In_802,In_2194);
xnor U1184 (N_1184,In_2330,In_614);
and U1185 (N_1185,In_1759,In_2148);
and U1186 (N_1186,In_108,In_1726);
or U1187 (N_1187,In_1926,In_1180);
or U1188 (N_1188,In_2249,In_2065);
nor U1189 (N_1189,In_337,In_1239);
or U1190 (N_1190,In_657,In_987);
and U1191 (N_1191,In_38,In_1950);
or U1192 (N_1192,In_691,In_730);
nand U1193 (N_1193,In_1919,In_636);
and U1194 (N_1194,In_2210,In_2321);
or U1195 (N_1195,In_2136,In_1728);
xor U1196 (N_1196,In_1044,In_820);
or U1197 (N_1197,In_274,In_1936);
or U1198 (N_1198,In_227,In_1128);
or U1199 (N_1199,In_432,In_1599);
or U1200 (N_1200,In_921,In_1449);
nor U1201 (N_1201,In_159,In_1271);
nor U1202 (N_1202,In_919,In_955);
xnor U1203 (N_1203,In_1915,In_1089);
or U1204 (N_1204,In_275,In_1804);
and U1205 (N_1205,In_599,In_1480);
nand U1206 (N_1206,In_744,In_2138);
xor U1207 (N_1207,In_2358,In_1288);
nand U1208 (N_1208,In_680,In_2473);
or U1209 (N_1209,In_226,In_774);
and U1210 (N_1210,In_1882,In_639);
nor U1211 (N_1211,In_731,In_1594);
or U1212 (N_1212,In_924,In_206);
nor U1213 (N_1213,In_682,In_1552);
and U1214 (N_1214,In_1492,In_1264);
nor U1215 (N_1215,In_2256,In_2140);
and U1216 (N_1216,In_1785,In_544);
and U1217 (N_1217,In_2461,In_1141);
and U1218 (N_1218,In_92,In_742);
and U1219 (N_1219,In_556,In_483);
xor U1220 (N_1220,In_2145,In_236);
nor U1221 (N_1221,In_479,In_887);
nor U1222 (N_1222,In_106,In_2482);
nand U1223 (N_1223,In_2224,In_2351);
nand U1224 (N_1224,In_1549,In_1864);
xnor U1225 (N_1225,In_1703,In_1633);
and U1226 (N_1226,In_1597,In_1251);
nor U1227 (N_1227,In_30,In_611);
xnor U1228 (N_1228,In_971,In_710);
xnor U1229 (N_1229,In_1072,In_136);
nand U1230 (N_1230,In_1886,In_1456);
or U1231 (N_1231,In_2059,In_1488);
or U1232 (N_1232,In_2288,In_295);
or U1233 (N_1233,In_1866,In_123);
nand U1234 (N_1234,In_1300,In_777);
nor U1235 (N_1235,In_605,In_2121);
and U1236 (N_1236,In_2278,In_1416);
and U1237 (N_1237,In_545,In_950);
or U1238 (N_1238,In_116,In_263);
xor U1239 (N_1239,In_620,In_1078);
and U1240 (N_1240,In_860,In_2271);
and U1241 (N_1241,In_536,In_787);
nor U1242 (N_1242,In_1274,In_2430);
nand U1243 (N_1243,In_472,In_1459);
nor U1244 (N_1244,In_2341,In_1539);
nand U1245 (N_1245,In_828,In_560);
nor U1246 (N_1246,In_11,In_1296);
nand U1247 (N_1247,In_165,In_156);
nor U1248 (N_1248,In_1442,In_1838);
and U1249 (N_1249,In_1664,In_1820);
nand U1250 (N_1250,In_303,In_76);
xnor U1251 (N_1251,In_1305,In_288);
or U1252 (N_1252,In_1265,In_766);
and U1253 (N_1253,In_1417,In_2166);
nor U1254 (N_1254,In_1796,In_1852);
or U1255 (N_1255,In_592,In_1959);
xnor U1256 (N_1256,In_1637,In_1359);
and U1257 (N_1257,In_1612,In_321);
xor U1258 (N_1258,In_99,In_118);
nand U1259 (N_1259,In_2496,In_2117);
and U1260 (N_1260,In_934,In_2123);
nand U1261 (N_1261,In_1110,In_1657);
nand U1262 (N_1262,In_450,In_710);
and U1263 (N_1263,In_647,In_1772);
nor U1264 (N_1264,In_1594,In_421);
or U1265 (N_1265,In_2132,In_1576);
nand U1266 (N_1266,In_641,In_434);
nand U1267 (N_1267,In_491,In_835);
and U1268 (N_1268,In_1970,In_2144);
xnor U1269 (N_1269,In_21,In_355);
or U1270 (N_1270,In_1644,In_2103);
xor U1271 (N_1271,In_1277,In_2015);
nor U1272 (N_1272,In_2345,In_2142);
nor U1273 (N_1273,In_2375,In_1222);
nand U1274 (N_1274,In_1811,In_2076);
nor U1275 (N_1275,In_1855,In_786);
nand U1276 (N_1276,In_932,In_1573);
or U1277 (N_1277,In_175,In_1445);
or U1278 (N_1278,In_1576,In_2351);
or U1279 (N_1279,In_138,In_854);
or U1280 (N_1280,In_1497,In_789);
and U1281 (N_1281,In_815,In_2174);
or U1282 (N_1282,In_561,In_36);
or U1283 (N_1283,In_2037,In_2356);
nand U1284 (N_1284,In_954,In_159);
xnor U1285 (N_1285,In_624,In_1222);
and U1286 (N_1286,In_669,In_791);
and U1287 (N_1287,In_600,In_1430);
and U1288 (N_1288,In_2197,In_834);
nand U1289 (N_1289,In_2271,In_1162);
nand U1290 (N_1290,In_2303,In_252);
and U1291 (N_1291,In_1780,In_741);
nand U1292 (N_1292,In_716,In_903);
nor U1293 (N_1293,In_1927,In_915);
nand U1294 (N_1294,In_2495,In_2253);
nand U1295 (N_1295,In_1640,In_1106);
or U1296 (N_1296,In_363,In_163);
nand U1297 (N_1297,In_4,In_1036);
nor U1298 (N_1298,In_1321,In_1481);
nor U1299 (N_1299,In_476,In_29);
nor U1300 (N_1300,In_1297,In_2092);
or U1301 (N_1301,In_2166,In_297);
nand U1302 (N_1302,In_120,In_1403);
and U1303 (N_1303,In_17,In_1703);
and U1304 (N_1304,In_142,In_501);
or U1305 (N_1305,In_1666,In_1565);
and U1306 (N_1306,In_1701,In_704);
or U1307 (N_1307,In_982,In_1797);
or U1308 (N_1308,In_2377,In_1618);
or U1309 (N_1309,In_2327,In_813);
nand U1310 (N_1310,In_1024,In_659);
nand U1311 (N_1311,In_1167,In_1074);
and U1312 (N_1312,In_931,In_2270);
nand U1313 (N_1313,In_1473,In_167);
nor U1314 (N_1314,In_1209,In_391);
nand U1315 (N_1315,In_50,In_2306);
nor U1316 (N_1316,In_1334,In_59);
nand U1317 (N_1317,In_2387,In_417);
and U1318 (N_1318,In_1850,In_502);
xnor U1319 (N_1319,In_1581,In_1601);
xnor U1320 (N_1320,In_217,In_1953);
or U1321 (N_1321,In_862,In_1549);
or U1322 (N_1322,In_2426,In_1857);
nor U1323 (N_1323,In_1306,In_2098);
or U1324 (N_1324,In_111,In_855);
nor U1325 (N_1325,In_866,In_812);
and U1326 (N_1326,In_612,In_232);
nand U1327 (N_1327,In_599,In_1568);
xor U1328 (N_1328,In_2279,In_1809);
nor U1329 (N_1329,In_1604,In_1962);
xor U1330 (N_1330,In_875,In_548);
nor U1331 (N_1331,In_93,In_868);
and U1332 (N_1332,In_1414,In_1404);
or U1333 (N_1333,In_302,In_792);
and U1334 (N_1334,In_584,In_1231);
nand U1335 (N_1335,In_939,In_1791);
nor U1336 (N_1336,In_340,In_1005);
or U1337 (N_1337,In_1234,In_1414);
or U1338 (N_1338,In_403,In_820);
and U1339 (N_1339,In_1183,In_296);
or U1340 (N_1340,In_758,In_43);
nand U1341 (N_1341,In_793,In_1457);
nand U1342 (N_1342,In_1817,In_948);
xor U1343 (N_1343,In_476,In_32);
xnor U1344 (N_1344,In_1440,In_316);
nand U1345 (N_1345,In_933,In_1411);
or U1346 (N_1346,In_1424,In_141);
and U1347 (N_1347,In_54,In_1067);
or U1348 (N_1348,In_1272,In_1322);
xnor U1349 (N_1349,In_176,In_202);
nor U1350 (N_1350,In_784,In_1674);
xnor U1351 (N_1351,In_2209,In_1109);
xnor U1352 (N_1352,In_200,In_2218);
or U1353 (N_1353,In_785,In_2020);
or U1354 (N_1354,In_746,In_608);
or U1355 (N_1355,In_1127,In_1157);
xor U1356 (N_1356,In_150,In_769);
and U1357 (N_1357,In_1092,In_481);
or U1358 (N_1358,In_2181,In_1062);
nor U1359 (N_1359,In_2010,In_207);
nor U1360 (N_1360,In_1435,In_102);
nand U1361 (N_1361,In_1150,In_2387);
nand U1362 (N_1362,In_435,In_414);
nor U1363 (N_1363,In_1121,In_1637);
xor U1364 (N_1364,In_1868,In_1929);
nand U1365 (N_1365,In_988,In_767);
nand U1366 (N_1366,In_1716,In_624);
or U1367 (N_1367,In_2212,In_1506);
nor U1368 (N_1368,In_2350,In_410);
or U1369 (N_1369,In_81,In_2264);
nand U1370 (N_1370,In_2478,In_1682);
nor U1371 (N_1371,In_585,In_518);
or U1372 (N_1372,In_2205,In_1815);
and U1373 (N_1373,In_2435,In_1134);
or U1374 (N_1374,In_2487,In_912);
nor U1375 (N_1375,In_2243,In_1572);
and U1376 (N_1376,In_1670,In_1693);
nand U1377 (N_1377,In_1877,In_2419);
or U1378 (N_1378,In_512,In_2399);
xnor U1379 (N_1379,In_448,In_336);
nor U1380 (N_1380,In_2321,In_1434);
and U1381 (N_1381,In_847,In_1201);
and U1382 (N_1382,In_387,In_562);
or U1383 (N_1383,In_571,In_562);
and U1384 (N_1384,In_165,In_1);
nor U1385 (N_1385,In_1746,In_1572);
or U1386 (N_1386,In_2335,In_124);
and U1387 (N_1387,In_1329,In_1959);
or U1388 (N_1388,In_336,In_2126);
or U1389 (N_1389,In_190,In_195);
nor U1390 (N_1390,In_124,In_2489);
or U1391 (N_1391,In_1378,In_949);
nor U1392 (N_1392,In_1691,In_206);
and U1393 (N_1393,In_659,In_375);
nand U1394 (N_1394,In_2333,In_1554);
nand U1395 (N_1395,In_2304,In_123);
or U1396 (N_1396,In_1050,In_1746);
nor U1397 (N_1397,In_356,In_1204);
xor U1398 (N_1398,In_2106,In_1112);
and U1399 (N_1399,In_1529,In_741);
or U1400 (N_1400,In_1276,In_347);
and U1401 (N_1401,In_1626,In_14);
and U1402 (N_1402,In_1630,In_1177);
or U1403 (N_1403,In_1626,In_1019);
nand U1404 (N_1404,In_691,In_1727);
nor U1405 (N_1405,In_1831,In_308);
nor U1406 (N_1406,In_0,In_306);
nor U1407 (N_1407,In_1625,In_2243);
or U1408 (N_1408,In_139,In_2060);
nor U1409 (N_1409,In_2252,In_1780);
nor U1410 (N_1410,In_1798,In_1375);
or U1411 (N_1411,In_1871,In_858);
or U1412 (N_1412,In_1424,In_92);
and U1413 (N_1413,In_1599,In_368);
nor U1414 (N_1414,In_1409,In_1461);
and U1415 (N_1415,In_2447,In_2435);
and U1416 (N_1416,In_1866,In_1511);
and U1417 (N_1417,In_1953,In_760);
or U1418 (N_1418,In_257,In_1934);
or U1419 (N_1419,In_279,In_2474);
and U1420 (N_1420,In_2190,In_424);
nand U1421 (N_1421,In_1563,In_322);
nor U1422 (N_1422,In_1348,In_510);
nor U1423 (N_1423,In_313,In_724);
or U1424 (N_1424,In_45,In_286);
or U1425 (N_1425,In_1376,In_464);
or U1426 (N_1426,In_1862,In_1171);
nor U1427 (N_1427,In_1830,In_1783);
nand U1428 (N_1428,In_148,In_634);
xor U1429 (N_1429,In_858,In_2254);
nand U1430 (N_1430,In_1994,In_74);
and U1431 (N_1431,In_2046,In_1453);
nor U1432 (N_1432,In_557,In_1753);
or U1433 (N_1433,In_1968,In_1708);
nand U1434 (N_1434,In_1370,In_905);
nand U1435 (N_1435,In_1663,In_537);
xor U1436 (N_1436,In_1750,In_946);
or U1437 (N_1437,In_1471,In_1139);
nand U1438 (N_1438,In_1515,In_2184);
nand U1439 (N_1439,In_2445,In_812);
nor U1440 (N_1440,In_885,In_1336);
or U1441 (N_1441,In_2488,In_1935);
and U1442 (N_1442,In_551,In_990);
xor U1443 (N_1443,In_1565,In_2395);
or U1444 (N_1444,In_1782,In_1046);
nand U1445 (N_1445,In_2037,In_1341);
nor U1446 (N_1446,In_2473,In_2350);
xnor U1447 (N_1447,In_1458,In_1340);
nor U1448 (N_1448,In_460,In_1814);
nand U1449 (N_1449,In_1065,In_837);
nand U1450 (N_1450,In_1872,In_1447);
nand U1451 (N_1451,In_520,In_2156);
nor U1452 (N_1452,In_1550,In_389);
nor U1453 (N_1453,In_697,In_572);
or U1454 (N_1454,In_2123,In_1027);
and U1455 (N_1455,In_1259,In_1204);
nand U1456 (N_1456,In_1725,In_2283);
nand U1457 (N_1457,In_562,In_1669);
and U1458 (N_1458,In_2081,In_664);
nor U1459 (N_1459,In_1729,In_111);
nor U1460 (N_1460,In_713,In_198);
nor U1461 (N_1461,In_998,In_1424);
and U1462 (N_1462,In_296,In_1718);
or U1463 (N_1463,In_577,In_1891);
and U1464 (N_1464,In_1848,In_1278);
xor U1465 (N_1465,In_1649,In_1629);
nor U1466 (N_1466,In_205,In_858);
nor U1467 (N_1467,In_775,In_244);
nor U1468 (N_1468,In_539,In_666);
xnor U1469 (N_1469,In_579,In_98);
or U1470 (N_1470,In_1379,In_536);
or U1471 (N_1471,In_713,In_1418);
or U1472 (N_1472,In_1915,In_1925);
and U1473 (N_1473,In_1398,In_84);
nand U1474 (N_1474,In_1319,In_1671);
or U1475 (N_1475,In_66,In_2243);
and U1476 (N_1476,In_841,In_22);
and U1477 (N_1477,In_2396,In_1975);
or U1478 (N_1478,In_549,In_73);
nor U1479 (N_1479,In_1936,In_288);
and U1480 (N_1480,In_705,In_599);
or U1481 (N_1481,In_657,In_1278);
and U1482 (N_1482,In_1505,In_1313);
or U1483 (N_1483,In_1924,In_2017);
or U1484 (N_1484,In_854,In_986);
and U1485 (N_1485,In_83,In_1156);
nor U1486 (N_1486,In_1051,In_2048);
nor U1487 (N_1487,In_901,In_73);
and U1488 (N_1488,In_2235,In_1383);
or U1489 (N_1489,In_315,In_1599);
or U1490 (N_1490,In_657,In_2229);
and U1491 (N_1491,In_950,In_322);
nand U1492 (N_1492,In_1036,In_1114);
xor U1493 (N_1493,In_2462,In_486);
nand U1494 (N_1494,In_709,In_1696);
nand U1495 (N_1495,In_1298,In_1604);
xnor U1496 (N_1496,In_1308,In_1573);
nand U1497 (N_1497,In_2068,In_2120);
or U1498 (N_1498,In_2445,In_1550);
nor U1499 (N_1499,In_1280,In_128);
nand U1500 (N_1500,In_2370,In_1375);
and U1501 (N_1501,In_623,In_537);
xor U1502 (N_1502,In_1490,In_651);
nor U1503 (N_1503,In_1491,In_443);
and U1504 (N_1504,In_203,In_1472);
nor U1505 (N_1505,In_1871,In_1349);
nor U1506 (N_1506,In_1288,In_37);
nand U1507 (N_1507,In_1499,In_75);
or U1508 (N_1508,In_1367,In_1623);
and U1509 (N_1509,In_76,In_1805);
nor U1510 (N_1510,In_133,In_1429);
xor U1511 (N_1511,In_1636,In_1587);
nand U1512 (N_1512,In_2288,In_1413);
nor U1513 (N_1513,In_361,In_407);
xor U1514 (N_1514,In_1228,In_1082);
and U1515 (N_1515,In_1317,In_1627);
nand U1516 (N_1516,In_867,In_698);
or U1517 (N_1517,In_438,In_939);
and U1518 (N_1518,In_2131,In_83);
xor U1519 (N_1519,In_1664,In_1450);
nand U1520 (N_1520,In_1968,In_750);
nor U1521 (N_1521,In_53,In_954);
nand U1522 (N_1522,In_362,In_887);
or U1523 (N_1523,In_339,In_2095);
nor U1524 (N_1524,In_1123,In_2313);
nand U1525 (N_1525,In_1790,In_1016);
or U1526 (N_1526,In_773,In_2046);
and U1527 (N_1527,In_2091,In_1564);
nor U1528 (N_1528,In_1065,In_981);
nand U1529 (N_1529,In_1067,In_1833);
nor U1530 (N_1530,In_337,In_1157);
or U1531 (N_1531,In_202,In_1313);
xnor U1532 (N_1532,In_1268,In_1490);
nor U1533 (N_1533,In_527,In_1637);
or U1534 (N_1534,In_410,In_448);
nand U1535 (N_1535,In_1853,In_1896);
and U1536 (N_1536,In_2334,In_1186);
or U1537 (N_1537,In_610,In_2188);
or U1538 (N_1538,In_201,In_1673);
nor U1539 (N_1539,In_2323,In_1455);
or U1540 (N_1540,In_1142,In_1885);
nor U1541 (N_1541,In_147,In_1653);
xor U1542 (N_1542,In_728,In_2109);
nand U1543 (N_1543,In_1525,In_703);
and U1544 (N_1544,In_438,In_275);
or U1545 (N_1545,In_448,In_1798);
nor U1546 (N_1546,In_2223,In_7);
or U1547 (N_1547,In_1017,In_2119);
nand U1548 (N_1548,In_1304,In_714);
nand U1549 (N_1549,In_1967,In_250);
or U1550 (N_1550,In_2072,In_704);
nand U1551 (N_1551,In_641,In_2328);
nand U1552 (N_1552,In_430,In_2437);
nand U1553 (N_1553,In_2405,In_90);
nand U1554 (N_1554,In_2044,In_758);
or U1555 (N_1555,In_1849,In_1654);
nand U1556 (N_1556,In_848,In_1541);
xnor U1557 (N_1557,In_442,In_790);
and U1558 (N_1558,In_1201,In_2488);
xnor U1559 (N_1559,In_62,In_483);
nor U1560 (N_1560,In_1819,In_2020);
or U1561 (N_1561,In_1257,In_708);
nor U1562 (N_1562,In_1577,In_1167);
nor U1563 (N_1563,In_592,In_1583);
or U1564 (N_1564,In_2069,In_1941);
and U1565 (N_1565,In_1185,In_1604);
nand U1566 (N_1566,In_1074,In_831);
nor U1567 (N_1567,In_954,In_2419);
nor U1568 (N_1568,In_2085,In_2024);
nor U1569 (N_1569,In_1663,In_2410);
or U1570 (N_1570,In_1660,In_1859);
nor U1571 (N_1571,In_2444,In_784);
nand U1572 (N_1572,In_1034,In_1280);
and U1573 (N_1573,In_333,In_2174);
nor U1574 (N_1574,In_352,In_1032);
nand U1575 (N_1575,In_404,In_96);
nor U1576 (N_1576,In_1494,In_1545);
nor U1577 (N_1577,In_1851,In_1769);
and U1578 (N_1578,In_912,In_689);
nand U1579 (N_1579,In_1189,In_1532);
nor U1580 (N_1580,In_2491,In_785);
and U1581 (N_1581,In_514,In_2101);
nor U1582 (N_1582,In_1448,In_1983);
or U1583 (N_1583,In_1808,In_1228);
nand U1584 (N_1584,In_1811,In_1159);
nand U1585 (N_1585,In_223,In_1449);
nand U1586 (N_1586,In_119,In_296);
nor U1587 (N_1587,In_700,In_2402);
nand U1588 (N_1588,In_565,In_2310);
or U1589 (N_1589,In_1285,In_1548);
and U1590 (N_1590,In_749,In_2108);
or U1591 (N_1591,In_1937,In_2);
and U1592 (N_1592,In_2373,In_1685);
nor U1593 (N_1593,In_209,In_286);
nor U1594 (N_1594,In_2106,In_2313);
and U1595 (N_1595,In_18,In_1068);
or U1596 (N_1596,In_1759,In_2179);
nor U1597 (N_1597,In_780,In_2271);
nor U1598 (N_1598,In_1097,In_1536);
nor U1599 (N_1599,In_678,In_2478);
or U1600 (N_1600,In_1043,In_1830);
nand U1601 (N_1601,In_1094,In_2301);
nor U1602 (N_1602,In_2363,In_941);
or U1603 (N_1603,In_1698,In_2102);
and U1604 (N_1604,In_1986,In_1999);
nand U1605 (N_1605,In_856,In_550);
nand U1606 (N_1606,In_1380,In_54);
and U1607 (N_1607,In_56,In_1452);
nand U1608 (N_1608,In_1773,In_242);
or U1609 (N_1609,In_2,In_1177);
and U1610 (N_1610,In_2341,In_2071);
nand U1611 (N_1611,In_1688,In_939);
or U1612 (N_1612,In_421,In_1916);
nor U1613 (N_1613,In_1476,In_813);
or U1614 (N_1614,In_1112,In_2249);
nand U1615 (N_1615,In_282,In_2281);
nand U1616 (N_1616,In_1072,In_2190);
or U1617 (N_1617,In_1068,In_1625);
nor U1618 (N_1618,In_1332,In_1176);
nor U1619 (N_1619,In_587,In_2366);
or U1620 (N_1620,In_2497,In_2093);
and U1621 (N_1621,In_1627,In_80);
nand U1622 (N_1622,In_708,In_1388);
nor U1623 (N_1623,In_481,In_2148);
or U1624 (N_1624,In_566,In_1690);
nor U1625 (N_1625,In_1541,In_1640);
nor U1626 (N_1626,In_1671,In_831);
nor U1627 (N_1627,In_1171,In_366);
nor U1628 (N_1628,In_1604,In_1558);
nor U1629 (N_1629,In_646,In_1217);
nor U1630 (N_1630,In_2171,In_1431);
xor U1631 (N_1631,In_351,In_1173);
or U1632 (N_1632,In_2191,In_2208);
nor U1633 (N_1633,In_1553,In_664);
nand U1634 (N_1634,In_442,In_311);
nor U1635 (N_1635,In_2099,In_1931);
and U1636 (N_1636,In_336,In_2098);
nor U1637 (N_1637,In_1843,In_1382);
or U1638 (N_1638,In_2332,In_1572);
and U1639 (N_1639,In_2248,In_2056);
nand U1640 (N_1640,In_886,In_303);
nor U1641 (N_1641,In_274,In_988);
xnor U1642 (N_1642,In_2003,In_1269);
and U1643 (N_1643,In_873,In_1632);
xor U1644 (N_1644,In_2340,In_1095);
or U1645 (N_1645,In_1280,In_2010);
nor U1646 (N_1646,In_1057,In_377);
nor U1647 (N_1647,In_179,In_638);
nand U1648 (N_1648,In_1675,In_738);
or U1649 (N_1649,In_939,In_1802);
xnor U1650 (N_1650,In_441,In_2264);
nor U1651 (N_1651,In_930,In_377);
and U1652 (N_1652,In_167,In_884);
and U1653 (N_1653,In_2498,In_670);
and U1654 (N_1654,In_86,In_625);
and U1655 (N_1655,In_1915,In_981);
nand U1656 (N_1656,In_1324,In_882);
nand U1657 (N_1657,In_933,In_1581);
xor U1658 (N_1658,In_1986,In_791);
or U1659 (N_1659,In_90,In_1167);
nor U1660 (N_1660,In_1232,In_2197);
xor U1661 (N_1661,In_212,In_981);
and U1662 (N_1662,In_437,In_188);
nand U1663 (N_1663,In_1432,In_2484);
and U1664 (N_1664,In_878,In_518);
or U1665 (N_1665,In_1551,In_742);
or U1666 (N_1666,In_1823,In_2452);
or U1667 (N_1667,In_573,In_510);
xnor U1668 (N_1668,In_2470,In_1907);
nand U1669 (N_1669,In_540,In_2438);
or U1670 (N_1670,In_2296,In_1093);
and U1671 (N_1671,In_673,In_1127);
nor U1672 (N_1672,In_737,In_590);
or U1673 (N_1673,In_1880,In_2355);
or U1674 (N_1674,In_1417,In_168);
nand U1675 (N_1675,In_1241,In_1333);
nand U1676 (N_1676,In_539,In_2326);
nor U1677 (N_1677,In_497,In_1916);
nand U1678 (N_1678,In_2082,In_1407);
nand U1679 (N_1679,In_1877,In_2130);
or U1680 (N_1680,In_2433,In_2051);
xnor U1681 (N_1681,In_1017,In_1068);
or U1682 (N_1682,In_511,In_1194);
nand U1683 (N_1683,In_885,In_579);
or U1684 (N_1684,In_1366,In_718);
nand U1685 (N_1685,In_608,In_2388);
nor U1686 (N_1686,In_482,In_2100);
and U1687 (N_1687,In_1116,In_1302);
or U1688 (N_1688,In_2232,In_805);
and U1689 (N_1689,In_913,In_2269);
nor U1690 (N_1690,In_1796,In_1532);
or U1691 (N_1691,In_338,In_479);
and U1692 (N_1692,In_1129,In_2316);
and U1693 (N_1693,In_2305,In_1449);
and U1694 (N_1694,In_885,In_1618);
or U1695 (N_1695,In_483,In_1579);
or U1696 (N_1696,In_2476,In_1712);
nand U1697 (N_1697,In_1646,In_424);
and U1698 (N_1698,In_1726,In_2383);
or U1699 (N_1699,In_1734,In_1093);
and U1700 (N_1700,In_1483,In_634);
and U1701 (N_1701,In_124,In_1963);
nor U1702 (N_1702,In_1520,In_1222);
and U1703 (N_1703,In_1208,In_886);
and U1704 (N_1704,In_852,In_704);
xnor U1705 (N_1705,In_1262,In_2037);
nor U1706 (N_1706,In_1120,In_1997);
nand U1707 (N_1707,In_787,In_747);
and U1708 (N_1708,In_1471,In_1778);
or U1709 (N_1709,In_1142,In_792);
xnor U1710 (N_1710,In_1214,In_1726);
xor U1711 (N_1711,In_1609,In_884);
nand U1712 (N_1712,In_926,In_460);
xnor U1713 (N_1713,In_1744,In_2368);
nand U1714 (N_1714,In_389,In_310);
nand U1715 (N_1715,In_1160,In_1862);
nand U1716 (N_1716,In_2106,In_818);
or U1717 (N_1717,In_1265,In_1688);
xor U1718 (N_1718,In_1893,In_387);
nand U1719 (N_1719,In_823,In_1574);
and U1720 (N_1720,In_1377,In_1135);
nand U1721 (N_1721,In_1571,In_1466);
nand U1722 (N_1722,In_1222,In_485);
and U1723 (N_1723,In_388,In_1982);
and U1724 (N_1724,In_2204,In_511);
nor U1725 (N_1725,In_1486,In_696);
nand U1726 (N_1726,In_2468,In_858);
nand U1727 (N_1727,In_2497,In_696);
and U1728 (N_1728,In_378,In_2415);
nor U1729 (N_1729,In_87,In_2325);
nor U1730 (N_1730,In_493,In_1942);
nand U1731 (N_1731,In_1542,In_244);
and U1732 (N_1732,In_1457,In_1488);
and U1733 (N_1733,In_996,In_1202);
xor U1734 (N_1734,In_1970,In_677);
xnor U1735 (N_1735,In_1561,In_266);
nand U1736 (N_1736,In_1127,In_1250);
or U1737 (N_1737,In_1669,In_806);
nor U1738 (N_1738,In_778,In_2323);
or U1739 (N_1739,In_2442,In_672);
or U1740 (N_1740,In_302,In_570);
and U1741 (N_1741,In_970,In_2299);
and U1742 (N_1742,In_298,In_1149);
nor U1743 (N_1743,In_1293,In_1309);
nor U1744 (N_1744,In_1253,In_2100);
nand U1745 (N_1745,In_1347,In_1601);
nor U1746 (N_1746,In_753,In_1743);
nor U1747 (N_1747,In_244,In_1975);
or U1748 (N_1748,In_1907,In_2103);
nor U1749 (N_1749,In_816,In_2031);
or U1750 (N_1750,In_2054,In_1543);
nand U1751 (N_1751,In_1800,In_1013);
nand U1752 (N_1752,In_1468,In_725);
or U1753 (N_1753,In_1039,In_1388);
and U1754 (N_1754,In_1247,In_2010);
nor U1755 (N_1755,In_862,In_2359);
or U1756 (N_1756,In_1147,In_1703);
or U1757 (N_1757,In_742,In_2414);
nand U1758 (N_1758,In_10,In_1186);
or U1759 (N_1759,In_1392,In_392);
xnor U1760 (N_1760,In_935,In_355);
and U1761 (N_1761,In_608,In_1860);
xnor U1762 (N_1762,In_2121,In_297);
and U1763 (N_1763,In_556,In_679);
nand U1764 (N_1764,In_171,In_620);
and U1765 (N_1765,In_754,In_1690);
xor U1766 (N_1766,In_955,In_1064);
nand U1767 (N_1767,In_265,In_357);
and U1768 (N_1768,In_1648,In_2061);
nor U1769 (N_1769,In_1246,In_87);
nor U1770 (N_1770,In_2274,In_1169);
nor U1771 (N_1771,In_717,In_10);
nand U1772 (N_1772,In_1654,In_2096);
nand U1773 (N_1773,In_2226,In_815);
xnor U1774 (N_1774,In_1449,In_1294);
nor U1775 (N_1775,In_1232,In_1041);
nand U1776 (N_1776,In_1155,In_1875);
nand U1777 (N_1777,In_831,In_2295);
or U1778 (N_1778,In_715,In_1748);
nor U1779 (N_1779,In_1164,In_383);
nor U1780 (N_1780,In_801,In_1616);
nor U1781 (N_1781,In_577,In_636);
nand U1782 (N_1782,In_909,In_1892);
or U1783 (N_1783,In_1201,In_2333);
nand U1784 (N_1784,In_2046,In_2272);
nand U1785 (N_1785,In_1096,In_1489);
nand U1786 (N_1786,In_1567,In_2439);
nor U1787 (N_1787,In_44,In_1019);
or U1788 (N_1788,In_2396,In_930);
and U1789 (N_1789,In_998,In_2040);
nand U1790 (N_1790,In_541,In_437);
nor U1791 (N_1791,In_308,In_2495);
nor U1792 (N_1792,In_244,In_662);
or U1793 (N_1793,In_2208,In_1204);
nor U1794 (N_1794,In_2289,In_1537);
xor U1795 (N_1795,In_486,In_814);
or U1796 (N_1796,In_2161,In_774);
nand U1797 (N_1797,In_2242,In_1203);
nand U1798 (N_1798,In_726,In_2481);
nand U1799 (N_1799,In_2372,In_815);
and U1800 (N_1800,In_818,In_2435);
nand U1801 (N_1801,In_306,In_1420);
nand U1802 (N_1802,In_994,In_973);
nor U1803 (N_1803,In_2088,In_191);
or U1804 (N_1804,In_1752,In_1638);
nand U1805 (N_1805,In_2,In_1038);
nand U1806 (N_1806,In_2134,In_1630);
nor U1807 (N_1807,In_634,In_1410);
xor U1808 (N_1808,In_1530,In_2002);
nor U1809 (N_1809,In_2067,In_867);
nand U1810 (N_1810,In_11,In_2369);
nand U1811 (N_1811,In_2380,In_667);
xnor U1812 (N_1812,In_2036,In_975);
or U1813 (N_1813,In_788,In_2056);
and U1814 (N_1814,In_513,In_1665);
and U1815 (N_1815,In_1583,In_759);
nor U1816 (N_1816,In_498,In_2125);
or U1817 (N_1817,In_1062,In_430);
and U1818 (N_1818,In_1997,In_2409);
or U1819 (N_1819,In_1751,In_1022);
nand U1820 (N_1820,In_2152,In_1464);
or U1821 (N_1821,In_2349,In_437);
or U1822 (N_1822,In_2087,In_1298);
xnor U1823 (N_1823,In_1523,In_693);
nand U1824 (N_1824,In_257,In_1495);
nand U1825 (N_1825,In_699,In_2282);
xnor U1826 (N_1826,In_1063,In_664);
or U1827 (N_1827,In_1510,In_170);
nor U1828 (N_1828,In_38,In_1721);
nor U1829 (N_1829,In_992,In_298);
nand U1830 (N_1830,In_1692,In_628);
or U1831 (N_1831,In_821,In_355);
or U1832 (N_1832,In_289,In_381);
or U1833 (N_1833,In_1750,In_2251);
nand U1834 (N_1834,In_1644,In_529);
nand U1835 (N_1835,In_1334,In_2232);
or U1836 (N_1836,In_1129,In_2318);
and U1837 (N_1837,In_1543,In_1024);
and U1838 (N_1838,In_363,In_33);
or U1839 (N_1839,In_2040,In_1276);
xor U1840 (N_1840,In_2091,In_1748);
nand U1841 (N_1841,In_1426,In_319);
and U1842 (N_1842,In_1033,In_440);
or U1843 (N_1843,In_2222,In_2418);
or U1844 (N_1844,In_225,In_1042);
or U1845 (N_1845,In_608,In_410);
and U1846 (N_1846,In_1765,In_208);
nand U1847 (N_1847,In_1910,In_2379);
and U1848 (N_1848,In_2223,In_1638);
nor U1849 (N_1849,In_2482,In_1299);
and U1850 (N_1850,In_513,In_80);
xnor U1851 (N_1851,In_1470,In_22);
and U1852 (N_1852,In_2199,In_152);
and U1853 (N_1853,In_842,In_1639);
nand U1854 (N_1854,In_554,In_1383);
or U1855 (N_1855,In_467,In_2317);
nor U1856 (N_1856,In_1921,In_2405);
or U1857 (N_1857,In_2097,In_376);
and U1858 (N_1858,In_820,In_2138);
nand U1859 (N_1859,In_1688,In_2174);
and U1860 (N_1860,In_1274,In_724);
nand U1861 (N_1861,In_1503,In_1897);
and U1862 (N_1862,In_804,In_1737);
and U1863 (N_1863,In_1540,In_716);
or U1864 (N_1864,In_2388,In_1656);
nor U1865 (N_1865,In_1113,In_339);
nand U1866 (N_1866,In_697,In_2300);
nand U1867 (N_1867,In_863,In_1344);
and U1868 (N_1868,In_665,In_972);
and U1869 (N_1869,In_897,In_1346);
or U1870 (N_1870,In_949,In_1453);
and U1871 (N_1871,In_914,In_1029);
and U1872 (N_1872,In_193,In_1884);
and U1873 (N_1873,In_1955,In_711);
xor U1874 (N_1874,In_1380,In_28);
nor U1875 (N_1875,In_1464,In_1181);
nand U1876 (N_1876,In_2425,In_1257);
nor U1877 (N_1877,In_56,In_616);
nor U1878 (N_1878,In_2071,In_785);
nor U1879 (N_1879,In_30,In_1013);
nand U1880 (N_1880,In_1213,In_2307);
or U1881 (N_1881,In_1413,In_2421);
nor U1882 (N_1882,In_218,In_1507);
nor U1883 (N_1883,In_424,In_670);
nand U1884 (N_1884,In_280,In_1450);
or U1885 (N_1885,In_268,In_2477);
and U1886 (N_1886,In_772,In_1062);
nor U1887 (N_1887,In_2358,In_1545);
nor U1888 (N_1888,In_901,In_2461);
or U1889 (N_1889,In_2001,In_1144);
and U1890 (N_1890,In_434,In_88);
nor U1891 (N_1891,In_12,In_1709);
and U1892 (N_1892,In_1365,In_1861);
nand U1893 (N_1893,In_2031,In_1983);
or U1894 (N_1894,In_726,In_143);
and U1895 (N_1895,In_999,In_2335);
and U1896 (N_1896,In_2314,In_616);
or U1897 (N_1897,In_809,In_1922);
or U1898 (N_1898,In_211,In_494);
and U1899 (N_1899,In_1629,In_1155);
or U1900 (N_1900,In_2189,In_127);
nor U1901 (N_1901,In_609,In_1501);
nand U1902 (N_1902,In_2195,In_2492);
xnor U1903 (N_1903,In_1906,In_768);
or U1904 (N_1904,In_2227,In_366);
or U1905 (N_1905,In_1577,In_321);
or U1906 (N_1906,In_1241,In_1019);
nor U1907 (N_1907,In_573,In_2233);
and U1908 (N_1908,In_15,In_520);
and U1909 (N_1909,In_1234,In_1817);
and U1910 (N_1910,In_1650,In_1662);
nor U1911 (N_1911,In_222,In_1033);
nor U1912 (N_1912,In_2198,In_972);
or U1913 (N_1913,In_733,In_2165);
or U1914 (N_1914,In_2334,In_1838);
nand U1915 (N_1915,In_1355,In_931);
and U1916 (N_1916,In_1196,In_1567);
nor U1917 (N_1917,In_973,In_260);
nor U1918 (N_1918,In_2244,In_1281);
or U1919 (N_1919,In_2469,In_893);
nand U1920 (N_1920,In_2499,In_1972);
or U1921 (N_1921,In_1049,In_572);
and U1922 (N_1922,In_71,In_1348);
and U1923 (N_1923,In_314,In_1487);
or U1924 (N_1924,In_379,In_1362);
xnor U1925 (N_1925,In_28,In_594);
and U1926 (N_1926,In_670,In_1510);
nand U1927 (N_1927,In_849,In_2279);
nor U1928 (N_1928,In_161,In_1143);
or U1929 (N_1929,In_2068,In_2002);
and U1930 (N_1930,In_1767,In_1236);
nor U1931 (N_1931,In_566,In_74);
nor U1932 (N_1932,In_1184,In_1433);
and U1933 (N_1933,In_1197,In_2260);
or U1934 (N_1934,In_2118,In_367);
nor U1935 (N_1935,In_242,In_2476);
nand U1936 (N_1936,In_729,In_1897);
nand U1937 (N_1937,In_840,In_271);
and U1938 (N_1938,In_477,In_348);
or U1939 (N_1939,In_1504,In_1780);
xor U1940 (N_1940,In_2213,In_1837);
nand U1941 (N_1941,In_1870,In_1246);
nor U1942 (N_1942,In_1998,In_324);
or U1943 (N_1943,In_916,In_2171);
or U1944 (N_1944,In_1815,In_1508);
or U1945 (N_1945,In_249,In_2184);
and U1946 (N_1946,In_2215,In_1236);
xor U1947 (N_1947,In_886,In_2361);
nand U1948 (N_1948,In_71,In_2286);
or U1949 (N_1949,In_436,In_1897);
or U1950 (N_1950,In_1354,In_1470);
nand U1951 (N_1951,In_28,In_4);
or U1952 (N_1952,In_1079,In_1085);
nand U1953 (N_1953,In_2085,In_1200);
and U1954 (N_1954,In_1537,In_712);
or U1955 (N_1955,In_829,In_176);
or U1956 (N_1956,In_2337,In_891);
nand U1957 (N_1957,In_1120,In_500);
nand U1958 (N_1958,In_275,In_2149);
and U1959 (N_1959,In_972,In_319);
and U1960 (N_1960,In_1347,In_1687);
nor U1961 (N_1961,In_2389,In_117);
xor U1962 (N_1962,In_2360,In_2411);
nand U1963 (N_1963,In_688,In_1314);
xor U1964 (N_1964,In_903,In_1008);
or U1965 (N_1965,In_2485,In_1246);
or U1966 (N_1966,In_787,In_1503);
xnor U1967 (N_1967,In_1140,In_1987);
or U1968 (N_1968,In_1358,In_146);
or U1969 (N_1969,In_843,In_2116);
nand U1970 (N_1970,In_861,In_60);
or U1971 (N_1971,In_20,In_2231);
nor U1972 (N_1972,In_847,In_519);
and U1973 (N_1973,In_1442,In_177);
and U1974 (N_1974,In_210,In_2106);
xor U1975 (N_1975,In_389,In_502);
or U1976 (N_1976,In_887,In_988);
and U1977 (N_1977,In_1670,In_1618);
and U1978 (N_1978,In_1367,In_2099);
nand U1979 (N_1979,In_1750,In_2231);
and U1980 (N_1980,In_1529,In_263);
or U1981 (N_1981,In_1783,In_960);
nor U1982 (N_1982,In_1435,In_635);
nand U1983 (N_1983,In_2468,In_2220);
or U1984 (N_1984,In_1206,In_551);
nand U1985 (N_1985,In_2168,In_644);
or U1986 (N_1986,In_1810,In_2144);
or U1987 (N_1987,In_1219,In_1355);
or U1988 (N_1988,In_636,In_126);
and U1989 (N_1989,In_1204,In_2264);
nor U1990 (N_1990,In_1070,In_1830);
xnor U1991 (N_1991,In_503,In_1805);
and U1992 (N_1992,In_1186,In_1130);
or U1993 (N_1993,In_349,In_674);
xor U1994 (N_1994,In_3,In_2029);
or U1995 (N_1995,In_224,In_2137);
and U1996 (N_1996,In_2470,In_2174);
nor U1997 (N_1997,In_2219,In_1250);
and U1998 (N_1998,In_1506,In_1757);
nand U1999 (N_1999,In_881,In_688);
and U2000 (N_2000,In_612,In_1005);
nand U2001 (N_2001,In_1209,In_1371);
and U2002 (N_2002,In_46,In_2356);
nand U2003 (N_2003,In_1439,In_1108);
or U2004 (N_2004,In_1077,In_1522);
and U2005 (N_2005,In_2186,In_1081);
nand U2006 (N_2006,In_76,In_342);
and U2007 (N_2007,In_830,In_1377);
and U2008 (N_2008,In_809,In_191);
or U2009 (N_2009,In_588,In_1053);
nor U2010 (N_2010,In_612,In_1012);
and U2011 (N_2011,In_1167,In_1808);
nand U2012 (N_2012,In_1319,In_1004);
xor U2013 (N_2013,In_363,In_2383);
or U2014 (N_2014,In_2495,In_727);
xnor U2015 (N_2015,In_359,In_224);
and U2016 (N_2016,In_2359,In_2296);
nor U2017 (N_2017,In_2207,In_398);
or U2018 (N_2018,In_1977,In_1020);
or U2019 (N_2019,In_2316,In_1986);
or U2020 (N_2020,In_631,In_1904);
nor U2021 (N_2021,In_1201,In_1581);
xor U2022 (N_2022,In_1618,In_1087);
nor U2023 (N_2023,In_1663,In_1057);
nor U2024 (N_2024,In_780,In_664);
or U2025 (N_2025,In_484,In_1011);
nand U2026 (N_2026,In_152,In_556);
xor U2027 (N_2027,In_137,In_1622);
nor U2028 (N_2028,In_506,In_138);
and U2029 (N_2029,In_2312,In_42);
or U2030 (N_2030,In_740,In_1707);
and U2031 (N_2031,In_335,In_2248);
or U2032 (N_2032,In_648,In_1323);
xnor U2033 (N_2033,In_391,In_1562);
xor U2034 (N_2034,In_2222,In_976);
nand U2035 (N_2035,In_1615,In_2183);
or U2036 (N_2036,In_780,In_1780);
nor U2037 (N_2037,In_448,In_460);
nor U2038 (N_2038,In_2005,In_1605);
and U2039 (N_2039,In_104,In_908);
or U2040 (N_2040,In_1186,In_659);
and U2041 (N_2041,In_206,In_95);
and U2042 (N_2042,In_989,In_2399);
nand U2043 (N_2043,In_1792,In_1205);
nand U2044 (N_2044,In_1053,In_193);
nand U2045 (N_2045,In_640,In_1545);
xnor U2046 (N_2046,In_1943,In_1745);
or U2047 (N_2047,In_1913,In_1206);
and U2048 (N_2048,In_961,In_269);
nand U2049 (N_2049,In_1313,In_1406);
nand U2050 (N_2050,In_2120,In_1674);
xnor U2051 (N_2051,In_1906,In_2460);
nand U2052 (N_2052,In_2373,In_573);
and U2053 (N_2053,In_1677,In_1381);
nand U2054 (N_2054,In_2181,In_1002);
or U2055 (N_2055,In_1831,In_1376);
and U2056 (N_2056,In_1722,In_648);
or U2057 (N_2057,In_126,In_916);
xnor U2058 (N_2058,In_787,In_824);
nor U2059 (N_2059,In_1075,In_824);
xnor U2060 (N_2060,In_209,In_2078);
or U2061 (N_2061,In_185,In_2391);
nor U2062 (N_2062,In_1409,In_1337);
xnor U2063 (N_2063,In_2491,In_1950);
nor U2064 (N_2064,In_1308,In_106);
nor U2065 (N_2065,In_1417,In_558);
and U2066 (N_2066,In_655,In_920);
nand U2067 (N_2067,In_582,In_1452);
nor U2068 (N_2068,In_2467,In_422);
xnor U2069 (N_2069,In_2084,In_1387);
nor U2070 (N_2070,In_502,In_1351);
xnor U2071 (N_2071,In_1868,In_239);
or U2072 (N_2072,In_2071,In_1580);
or U2073 (N_2073,In_305,In_1019);
xor U2074 (N_2074,In_2106,In_2296);
nor U2075 (N_2075,In_5,In_2289);
and U2076 (N_2076,In_837,In_1867);
xnor U2077 (N_2077,In_173,In_1104);
or U2078 (N_2078,In_1040,In_809);
and U2079 (N_2079,In_43,In_226);
nor U2080 (N_2080,In_618,In_1020);
and U2081 (N_2081,In_1128,In_1949);
or U2082 (N_2082,In_1077,In_1267);
xnor U2083 (N_2083,In_34,In_2032);
nand U2084 (N_2084,In_2482,In_1995);
nand U2085 (N_2085,In_712,In_1029);
xor U2086 (N_2086,In_1418,In_2222);
and U2087 (N_2087,In_967,In_732);
or U2088 (N_2088,In_24,In_1399);
nor U2089 (N_2089,In_237,In_1985);
nor U2090 (N_2090,In_866,In_883);
and U2091 (N_2091,In_0,In_1642);
or U2092 (N_2092,In_1300,In_1092);
nor U2093 (N_2093,In_1774,In_2108);
nor U2094 (N_2094,In_1942,In_1437);
xor U2095 (N_2095,In_697,In_1437);
or U2096 (N_2096,In_1609,In_1170);
nor U2097 (N_2097,In_1041,In_187);
nand U2098 (N_2098,In_2292,In_2495);
or U2099 (N_2099,In_1827,In_634);
nand U2100 (N_2100,In_180,In_959);
and U2101 (N_2101,In_990,In_1687);
nor U2102 (N_2102,In_424,In_1827);
xor U2103 (N_2103,In_693,In_794);
or U2104 (N_2104,In_960,In_1479);
and U2105 (N_2105,In_779,In_941);
nand U2106 (N_2106,In_952,In_889);
nand U2107 (N_2107,In_67,In_1799);
and U2108 (N_2108,In_502,In_1521);
nand U2109 (N_2109,In_1391,In_2484);
or U2110 (N_2110,In_1709,In_1198);
and U2111 (N_2111,In_2169,In_2308);
nor U2112 (N_2112,In_1293,In_2480);
nand U2113 (N_2113,In_1473,In_313);
nor U2114 (N_2114,In_1649,In_914);
nor U2115 (N_2115,In_2292,In_695);
or U2116 (N_2116,In_1309,In_2139);
nor U2117 (N_2117,In_732,In_1904);
or U2118 (N_2118,In_2351,In_503);
nor U2119 (N_2119,In_1695,In_2025);
or U2120 (N_2120,In_2087,In_2347);
nand U2121 (N_2121,In_936,In_1512);
xor U2122 (N_2122,In_1138,In_430);
and U2123 (N_2123,In_159,In_891);
xnor U2124 (N_2124,In_676,In_170);
nor U2125 (N_2125,In_208,In_1527);
nor U2126 (N_2126,In_1012,In_1983);
xnor U2127 (N_2127,In_1149,In_1724);
nor U2128 (N_2128,In_1130,In_896);
and U2129 (N_2129,In_1835,In_625);
nor U2130 (N_2130,In_497,In_607);
or U2131 (N_2131,In_363,In_1738);
or U2132 (N_2132,In_2020,In_1897);
and U2133 (N_2133,In_2081,In_1408);
or U2134 (N_2134,In_455,In_2202);
nand U2135 (N_2135,In_464,In_363);
nor U2136 (N_2136,In_1901,In_2275);
xnor U2137 (N_2137,In_2142,In_121);
or U2138 (N_2138,In_153,In_2470);
nor U2139 (N_2139,In_1595,In_1529);
and U2140 (N_2140,In_458,In_1787);
nand U2141 (N_2141,In_1912,In_343);
and U2142 (N_2142,In_1097,In_1317);
or U2143 (N_2143,In_981,In_1321);
and U2144 (N_2144,In_2392,In_1897);
and U2145 (N_2145,In_1302,In_1196);
or U2146 (N_2146,In_2319,In_2392);
nor U2147 (N_2147,In_126,In_1654);
and U2148 (N_2148,In_447,In_553);
nand U2149 (N_2149,In_352,In_1398);
and U2150 (N_2150,In_1584,In_1399);
nand U2151 (N_2151,In_1043,In_1804);
nand U2152 (N_2152,In_1901,In_342);
or U2153 (N_2153,In_2064,In_470);
or U2154 (N_2154,In_1125,In_664);
nand U2155 (N_2155,In_557,In_1714);
or U2156 (N_2156,In_2297,In_2427);
nand U2157 (N_2157,In_1871,In_545);
and U2158 (N_2158,In_2055,In_555);
nor U2159 (N_2159,In_1257,In_21);
or U2160 (N_2160,In_987,In_49);
nand U2161 (N_2161,In_2380,In_598);
and U2162 (N_2162,In_583,In_707);
and U2163 (N_2163,In_858,In_414);
nand U2164 (N_2164,In_166,In_715);
nor U2165 (N_2165,In_359,In_2465);
xnor U2166 (N_2166,In_1799,In_1698);
and U2167 (N_2167,In_2198,In_2228);
nand U2168 (N_2168,In_1998,In_2229);
and U2169 (N_2169,In_2282,In_314);
nand U2170 (N_2170,In_1517,In_1983);
nor U2171 (N_2171,In_284,In_1340);
or U2172 (N_2172,In_2231,In_290);
and U2173 (N_2173,In_2084,In_1242);
nor U2174 (N_2174,In_121,In_1503);
nand U2175 (N_2175,In_1352,In_2224);
nor U2176 (N_2176,In_1329,In_292);
nand U2177 (N_2177,In_1868,In_2168);
nor U2178 (N_2178,In_601,In_971);
nand U2179 (N_2179,In_1273,In_142);
nand U2180 (N_2180,In_68,In_680);
or U2181 (N_2181,In_1419,In_2133);
or U2182 (N_2182,In_406,In_297);
nand U2183 (N_2183,In_90,In_626);
or U2184 (N_2184,In_2227,In_1484);
nand U2185 (N_2185,In_822,In_916);
nand U2186 (N_2186,In_2109,In_897);
nor U2187 (N_2187,In_648,In_746);
nor U2188 (N_2188,In_2153,In_1576);
and U2189 (N_2189,In_525,In_441);
and U2190 (N_2190,In_1628,In_736);
nor U2191 (N_2191,In_447,In_1559);
nand U2192 (N_2192,In_2356,In_1839);
nand U2193 (N_2193,In_1488,In_868);
nor U2194 (N_2194,In_1008,In_157);
and U2195 (N_2195,In_527,In_1464);
or U2196 (N_2196,In_1717,In_554);
nor U2197 (N_2197,In_594,In_775);
or U2198 (N_2198,In_2281,In_1140);
or U2199 (N_2199,In_264,In_26);
nand U2200 (N_2200,In_1748,In_954);
nand U2201 (N_2201,In_2439,In_2247);
nand U2202 (N_2202,In_443,In_1748);
and U2203 (N_2203,In_265,In_1833);
and U2204 (N_2204,In_1580,In_2048);
or U2205 (N_2205,In_2489,In_1845);
and U2206 (N_2206,In_2105,In_2139);
or U2207 (N_2207,In_2308,In_2090);
and U2208 (N_2208,In_2435,In_341);
nor U2209 (N_2209,In_2440,In_751);
or U2210 (N_2210,In_1505,In_574);
nand U2211 (N_2211,In_1270,In_1240);
and U2212 (N_2212,In_1548,In_1489);
nand U2213 (N_2213,In_1232,In_2171);
nand U2214 (N_2214,In_322,In_1451);
nor U2215 (N_2215,In_2291,In_963);
nand U2216 (N_2216,In_1244,In_94);
nand U2217 (N_2217,In_321,In_840);
nand U2218 (N_2218,In_408,In_578);
nand U2219 (N_2219,In_72,In_110);
nor U2220 (N_2220,In_321,In_299);
nor U2221 (N_2221,In_2345,In_1348);
nor U2222 (N_2222,In_478,In_1388);
xor U2223 (N_2223,In_1698,In_1056);
and U2224 (N_2224,In_127,In_1373);
nor U2225 (N_2225,In_1849,In_1739);
nor U2226 (N_2226,In_2186,In_470);
and U2227 (N_2227,In_107,In_1491);
nand U2228 (N_2228,In_976,In_1053);
xor U2229 (N_2229,In_1954,In_2339);
nand U2230 (N_2230,In_1412,In_1299);
or U2231 (N_2231,In_1480,In_1458);
nor U2232 (N_2232,In_1788,In_224);
nor U2233 (N_2233,In_1190,In_523);
xnor U2234 (N_2234,In_1598,In_2098);
xnor U2235 (N_2235,In_1589,In_1045);
or U2236 (N_2236,In_505,In_1546);
and U2237 (N_2237,In_1356,In_2475);
nand U2238 (N_2238,In_1206,In_2178);
and U2239 (N_2239,In_2384,In_977);
and U2240 (N_2240,In_2425,In_427);
or U2241 (N_2241,In_186,In_566);
or U2242 (N_2242,In_627,In_2125);
or U2243 (N_2243,In_1268,In_1303);
or U2244 (N_2244,In_2233,In_191);
nand U2245 (N_2245,In_315,In_2468);
and U2246 (N_2246,In_263,In_1037);
xor U2247 (N_2247,In_853,In_205);
or U2248 (N_2248,In_524,In_865);
nor U2249 (N_2249,In_1381,In_952);
nor U2250 (N_2250,In_2131,In_1743);
and U2251 (N_2251,In_372,In_821);
and U2252 (N_2252,In_1882,In_1397);
nand U2253 (N_2253,In_1298,In_2332);
nand U2254 (N_2254,In_187,In_1238);
nor U2255 (N_2255,In_1884,In_1937);
xnor U2256 (N_2256,In_1509,In_2381);
nand U2257 (N_2257,In_608,In_1148);
or U2258 (N_2258,In_2284,In_2499);
and U2259 (N_2259,In_1587,In_1088);
nand U2260 (N_2260,In_1483,In_1666);
and U2261 (N_2261,In_2334,In_2379);
and U2262 (N_2262,In_1267,In_2455);
and U2263 (N_2263,In_1136,In_826);
or U2264 (N_2264,In_1957,In_739);
nor U2265 (N_2265,In_707,In_2225);
and U2266 (N_2266,In_286,In_1895);
or U2267 (N_2267,In_1668,In_911);
and U2268 (N_2268,In_622,In_1441);
xor U2269 (N_2269,In_2169,In_2259);
nand U2270 (N_2270,In_633,In_1117);
and U2271 (N_2271,In_451,In_550);
or U2272 (N_2272,In_2178,In_1269);
nor U2273 (N_2273,In_101,In_2026);
nor U2274 (N_2274,In_405,In_119);
or U2275 (N_2275,In_2202,In_79);
and U2276 (N_2276,In_128,In_1952);
or U2277 (N_2277,In_2073,In_388);
or U2278 (N_2278,In_1584,In_1254);
and U2279 (N_2279,In_452,In_1449);
nand U2280 (N_2280,In_2462,In_1184);
nor U2281 (N_2281,In_272,In_1392);
or U2282 (N_2282,In_588,In_172);
nor U2283 (N_2283,In_1730,In_2349);
nor U2284 (N_2284,In_2032,In_2031);
xor U2285 (N_2285,In_610,In_1464);
nand U2286 (N_2286,In_839,In_2005);
and U2287 (N_2287,In_1073,In_1776);
nand U2288 (N_2288,In_422,In_1584);
and U2289 (N_2289,In_1700,In_308);
or U2290 (N_2290,In_2279,In_2375);
and U2291 (N_2291,In_476,In_1513);
nand U2292 (N_2292,In_689,In_2332);
xnor U2293 (N_2293,In_1385,In_2066);
nand U2294 (N_2294,In_234,In_1777);
and U2295 (N_2295,In_858,In_2153);
and U2296 (N_2296,In_2074,In_1729);
and U2297 (N_2297,In_1513,In_524);
and U2298 (N_2298,In_2198,In_763);
nor U2299 (N_2299,In_2024,In_445);
nor U2300 (N_2300,In_367,In_1073);
nand U2301 (N_2301,In_1450,In_499);
nor U2302 (N_2302,In_777,In_2003);
or U2303 (N_2303,In_9,In_1068);
and U2304 (N_2304,In_1771,In_2445);
nand U2305 (N_2305,In_1217,In_1602);
xnor U2306 (N_2306,In_1718,In_1904);
or U2307 (N_2307,In_1845,In_2272);
xor U2308 (N_2308,In_1340,In_2173);
or U2309 (N_2309,In_595,In_393);
and U2310 (N_2310,In_1689,In_1226);
or U2311 (N_2311,In_596,In_1363);
or U2312 (N_2312,In_24,In_1941);
nor U2313 (N_2313,In_1496,In_621);
nand U2314 (N_2314,In_305,In_1244);
and U2315 (N_2315,In_1162,In_1694);
and U2316 (N_2316,In_2417,In_1354);
or U2317 (N_2317,In_2062,In_737);
nor U2318 (N_2318,In_2182,In_1522);
or U2319 (N_2319,In_979,In_2194);
and U2320 (N_2320,In_199,In_778);
or U2321 (N_2321,In_922,In_1233);
or U2322 (N_2322,In_163,In_823);
xnor U2323 (N_2323,In_1765,In_2312);
nor U2324 (N_2324,In_1073,In_404);
xor U2325 (N_2325,In_673,In_995);
nor U2326 (N_2326,In_0,In_921);
nor U2327 (N_2327,In_573,In_2229);
and U2328 (N_2328,In_190,In_789);
nor U2329 (N_2329,In_1111,In_1441);
and U2330 (N_2330,In_615,In_1204);
xnor U2331 (N_2331,In_1351,In_396);
nand U2332 (N_2332,In_1567,In_247);
nor U2333 (N_2333,In_1437,In_1672);
nor U2334 (N_2334,In_487,In_1530);
or U2335 (N_2335,In_2014,In_798);
or U2336 (N_2336,In_2244,In_1693);
nor U2337 (N_2337,In_884,In_1346);
nor U2338 (N_2338,In_2411,In_1008);
and U2339 (N_2339,In_2349,In_1443);
xnor U2340 (N_2340,In_2348,In_2069);
or U2341 (N_2341,In_1898,In_269);
and U2342 (N_2342,In_1581,In_1617);
xor U2343 (N_2343,In_1661,In_1908);
nand U2344 (N_2344,In_1574,In_184);
nor U2345 (N_2345,In_1302,In_722);
nor U2346 (N_2346,In_722,In_1947);
and U2347 (N_2347,In_329,In_1226);
nand U2348 (N_2348,In_1426,In_1005);
nand U2349 (N_2349,In_2380,In_837);
nor U2350 (N_2350,In_572,In_1029);
nor U2351 (N_2351,In_1953,In_1648);
or U2352 (N_2352,In_2249,In_2153);
nand U2353 (N_2353,In_1280,In_1664);
or U2354 (N_2354,In_356,In_696);
nor U2355 (N_2355,In_1160,In_1759);
nor U2356 (N_2356,In_2303,In_553);
nand U2357 (N_2357,In_1845,In_1311);
and U2358 (N_2358,In_97,In_704);
nand U2359 (N_2359,In_1379,In_712);
nand U2360 (N_2360,In_1098,In_1396);
nand U2361 (N_2361,In_427,In_1969);
and U2362 (N_2362,In_1133,In_884);
nand U2363 (N_2363,In_1279,In_2431);
and U2364 (N_2364,In_1731,In_726);
or U2365 (N_2365,In_2249,In_257);
nand U2366 (N_2366,In_2246,In_1101);
or U2367 (N_2367,In_1479,In_1183);
or U2368 (N_2368,In_2246,In_596);
nor U2369 (N_2369,In_1902,In_2201);
and U2370 (N_2370,In_896,In_10);
and U2371 (N_2371,In_78,In_1318);
or U2372 (N_2372,In_389,In_2455);
and U2373 (N_2373,In_2102,In_833);
nand U2374 (N_2374,In_1567,In_2424);
or U2375 (N_2375,In_1186,In_2415);
or U2376 (N_2376,In_1330,In_1287);
or U2377 (N_2377,In_1757,In_2085);
nor U2378 (N_2378,In_2479,In_1570);
and U2379 (N_2379,In_368,In_233);
xnor U2380 (N_2380,In_2478,In_75);
xor U2381 (N_2381,In_2023,In_1121);
xor U2382 (N_2382,In_2339,In_1904);
and U2383 (N_2383,In_1684,In_2457);
and U2384 (N_2384,In_1494,In_709);
nor U2385 (N_2385,In_2060,In_2098);
nor U2386 (N_2386,In_2254,In_1822);
nand U2387 (N_2387,In_826,In_885);
and U2388 (N_2388,In_1797,In_2237);
or U2389 (N_2389,In_1158,In_2160);
or U2390 (N_2390,In_2261,In_117);
nor U2391 (N_2391,In_1189,In_717);
xnor U2392 (N_2392,In_2151,In_315);
nor U2393 (N_2393,In_1218,In_497);
or U2394 (N_2394,In_1120,In_2444);
or U2395 (N_2395,In_1943,In_818);
and U2396 (N_2396,In_563,In_2405);
and U2397 (N_2397,In_1374,In_1166);
xor U2398 (N_2398,In_1828,In_186);
xnor U2399 (N_2399,In_403,In_247);
and U2400 (N_2400,In_356,In_2035);
nand U2401 (N_2401,In_1992,In_251);
and U2402 (N_2402,In_1916,In_1471);
xor U2403 (N_2403,In_2399,In_1934);
nor U2404 (N_2404,In_1610,In_166);
nand U2405 (N_2405,In_1973,In_581);
nor U2406 (N_2406,In_1805,In_1240);
or U2407 (N_2407,In_161,In_1698);
or U2408 (N_2408,In_1257,In_2252);
or U2409 (N_2409,In_454,In_1685);
nor U2410 (N_2410,In_1125,In_1473);
and U2411 (N_2411,In_1138,In_1270);
xnor U2412 (N_2412,In_1891,In_1060);
nand U2413 (N_2413,In_2061,In_1375);
nand U2414 (N_2414,In_1486,In_840);
nand U2415 (N_2415,In_46,In_1371);
or U2416 (N_2416,In_1885,In_2087);
xnor U2417 (N_2417,In_2457,In_543);
xor U2418 (N_2418,In_2229,In_546);
nor U2419 (N_2419,In_603,In_2246);
and U2420 (N_2420,In_1737,In_261);
and U2421 (N_2421,In_695,In_2413);
xor U2422 (N_2422,In_62,In_1775);
nor U2423 (N_2423,In_1013,In_533);
or U2424 (N_2424,In_870,In_886);
nor U2425 (N_2425,In_1434,In_21);
or U2426 (N_2426,In_113,In_2031);
nor U2427 (N_2427,In_1915,In_344);
and U2428 (N_2428,In_67,In_130);
and U2429 (N_2429,In_419,In_1408);
and U2430 (N_2430,In_1885,In_634);
or U2431 (N_2431,In_384,In_429);
or U2432 (N_2432,In_2253,In_1251);
or U2433 (N_2433,In_2264,In_987);
and U2434 (N_2434,In_2052,In_2142);
and U2435 (N_2435,In_956,In_412);
and U2436 (N_2436,In_193,In_1716);
nand U2437 (N_2437,In_371,In_2028);
or U2438 (N_2438,In_683,In_2082);
nand U2439 (N_2439,In_131,In_1191);
or U2440 (N_2440,In_926,In_1591);
and U2441 (N_2441,In_1658,In_815);
nand U2442 (N_2442,In_529,In_711);
nor U2443 (N_2443,In_675,In_800);
or U2444 (N_2444,In_606,In_438);
xor U2445 (N_2445,In_1407,In_1529);
or U2446 (N_2446,In_1989,In_1211);
nor U2447 (N_2447,In_1263,In_805);
nand U2448 (N_2448,In_1662,In_288);
nand U2449 (N_2449,In_344,In_1158);
nor U2450 (N_2450,In_2160,In_1261);
nand U2451 (N_2451,In_851,In_1117);
nor U2452 (N_2452,In_300,In_675);
nand U2453 (N_2453,In_1773,In_1772);
and U2454 (N_2454,In_159,In_274);
xnor U2455 (N_2455,In_525,In_57);
nor U2456 (N_2456,In_202,In_2136);
and U2457 (N_2457,In_1793,In_850);
nor U2458 (N_2458,In_2151,In_1539);
and U2459 (N_2459,In_2143,In_1898);
or U2460 (N_2460,In_2485,In_835);
and U2461 (N_2461,In_22,In_769);
or U2462 (N_2462,In_2458,In_212);
or U2463 (N_2463,In_460,In_1619);
or U2464 (N_2464,In_315,In_1913);
nand U2465 (N_2465,In_156,In_144);
or U2466 (N_2466,In_288,In_1730);
nand U2467 (N_2467,In_711,In_1890);
nand U2468 (N_2468,In_1820,In_2460);
nor U2469 (N_2469,In_1171,In_1406);
or U2470 (N_2470,In_1803,In_1490);
nor U2471 (N_2471,In_2013,In_341);
nand U2472 (N_2472,In_2382,In_667);
and U2473 (N_2473,In_543,In_1254);
and U2474 (N_2474,In_529,In_621);
or U2475 (N_2475,In_1513,In_123);
xnor U2476 (N_2476,In_397,In_174);
nor U2477 (N_2477,In_1309,In_1468);
xor U2478 (N_2478,In_1847,In_2285);
nand U2479 (N_2479,In_609,In_1987);
nor U2480 (N_2480,In_2179,In_717);
nand U2481 (N_2481,In_609,In_1484);
nor U2482 (N_2482,In_395,In_294);
nor U2483 (N_2483,In_1108,In_1047);
and U2484 (N_2484,In_2453,In_549);
nor U2485 (N_2485,In_1833,In_2103);
or U2486 (N_2486,In_710,In_2029);
and U2487 (N_2487,In_1126,In_2223);
nand U2488 (N_2488,In_1675,In_1202);
and U2489 (N_2489,In_441,In_2128);
xor U2490 (N_2490,In_2379,In_2315);
nor U2491 (N_2491,In_248,In_629);
nor U2492 (N_2492,In_179,In_833);
xnor U2493 (N_2493,In_1155,In_2433);
or U2494 (N_2494,In_404,In_736);
or U2495 (N_2495,In_1265,In_14);
xnor U2496 (N_2496,In_1293,In_1419);
nand U2497 (N_2497,In_799,In_419);
nand U2498 (N_2498,In_1683,In_1424);
and U2499 (N_2499,In_2408,In_334);
nand U2500 (N_2500,In_2407,In_1304);
nand U2501 (N_2501,In_2184,In_822);
or U2502 (N_2502,In_2100,In_612);
nand U2503 (N_2503,In_1813,In_499);
xnor U2504 (N_2504,In_1815,In_136);
nor U2505 (N_2505,In_390,In_1340);
nand U2506 (N_2506,In_1938,In_119);
and U2507 (N_2507,In_2043,In_578);
nand U2508 (N_2508,In_161,In_227);
or U2509 (N_2509,In_328,In_1073);
or U2510 (N_2510,In_277,In_2429);
and U2511 (N_2511,In_1980,In_1477);
and U2512 (N_2512,In_492,In_2381);
nor U2513 (N_2513,In_315,In_1927);
or U2514 (N_2514,In_2255,In_1757);
nor U2515 (N_2515,In_1863,In_1755);
xor U2516 (N_2516,In_217,In_1600);
nand U2517 (N_2517,In_340,In_1288);
or U2518 (N_2518,In_2046,In_1621);
nor U2519 (N_2519,In_1540,In_1098);
or U2520 (N_2520,In_1948,In_2331);
nor U2521 (N_2521,In_82,In_1266);
or U2522 (N_2522,In_1696,In_1228);
or U2523 (N_2523,In_1233,In_174);
nor U2524 (N_2524,In_1265,In_1548);
xnor U2525 (N_2525,In_245,In_338);
or U2526 (N_2526,In_2481,In_384);
or U2527 (N_2527,In_1972,In_117);
nor U2528 (N_2528,In_2379,In_1199);
and U2529 (N_2529,In_1257,In_1330);
nand U2530 (N_2530,In_415,In_1029);
nor U2531 (N_2531,In_1754,In_555);
or U2532 (N_2532,In_46,In_1816);
or U2533 (N_2533,In_356,In_1651);
and U2534 (N_2534,In_286,In_1250);
and U2535 (N_2535,In_1264,In_1140);
nor U2536 (N_2536,In_909,In_181);
nand U2537 (N_2537,In_1959,In_2176);
or U2538 (N_2538,In_2137,In_2152);
or U2539 (N_2539,In_2232,In_1310);
nor U2540 (N_2540,In_1631,In_1502);
nand U2541 (N_2541,In_2234,In_1785);
nand U2542 (N_2542,In_1297,In_190);
nor U2543 (N_2543,In_1430,In_615);
nand U2544 (N_2544,In_46,In_1349);
nand U2545 (N_2545,In_1762,In_2366);
or U2546 (N_2546,In_144,In_955);
nand U2547 (N_2547,In_1613,In_246);
xor U2548 (N_2548,In_254,In_916);
xnor U2549 (N_2549,In_885,In_1940);
and U2550 (N_2550,In_920,In_1895);
nor U2551 (N_2551,In_1272,In_175);
xor U2552 (N_2552,In_253,In_440);
or U2553 (N_2553,In_1062,In_1496);
nor U2554 (N_2554,In_1766,In_607);
xnor U2555 (N_2555,In_1399,In_1752);
nor U2556 (N_2556,In_1446,In_1456);
and U2557 (N_2557,In_1600,In_1921);
nor U2558 (N_2558,In_1477,In_1007);
nor U2559 (N_2559,In_756,In_557);
or U2560 (N_2560,In_1050,In_276);
or U2561 (N_2561,In_188,In_1504);
and U2562 (N_2562,In_945,In_1797);
xnor U2563 (N_2563,In_2070,In_1264);
nor U2564 (N_2564,In_1534,In_2268);
nor U2565 (N_2565,In_1629,In_216);
and U2566 (N_2566,In_792,In_1183);
or U2567 (N_2567,In_2056,In_1239);
or U2568 (N_2568,In_988,In_259);
nor U2569 (N_2569,In_26,In_597);
nor U2570 (N_2570,In_848,In_2384);
nand U2571 (N_2571,In_1912,In_1277);
nor U2572 (N_2572,In_655,In_880);
xor U2573 (N_2573,In_2105,In_1491);
nand U2574 (N_2574,In_1335,In_12);
nor U2575 (N_2575,In_2416,In_1056);
nand U2576 (N_2576,In_1055,In_105);
or U2577 (N_2577,In_1092,In_174);
or U2578 (N_2578,In_1268,In_133);
nor U2579 (N_2579,In_169,In_618);
or U2580 (N_2580,In_1839,In_942);
and U2581 (N_2581,In_1426,In_2404);
nor U2582 (N_2582,In_1853,In_826);
nand U2583 (N_2583,In_1877,In_258);
nand U2584 (N_2584,In_1771,In_149);
nand U2585 (N_2585,In_1647,In_2411);
and U2586 (N_2586,In_1915,In_433);
nand U2587 (N_2587,In_1791,In_2382);
or U2588 (N_2588,In_620,In_2391);
nand U2589 (N_2589,In_2332,In_1792);
nand U2590 (N_2590,In_2177,In_1075);
and U2591 (N_2591,In_593,In_1388);
nand U2592 (N_2592,In_412,In_565);
nand U2593 (N_2593,In_471,In_1630);
or U2594 (N_2594,In_1695,In_2411);
nand U2595 (N_2595,In_1306,In_969);
nor U2596 (N_2596,In_855,In_1166);
and U2597 (N_2597,In_795,In_1241);
nor U2598 (N_2598,In_608,In_1561);
nor U2599 (N_2599,In_1217,In_1642);
or U2600 (N_2600,In_89,In_2366);
nand U2601 (N_2601,In_1823,In_2365);
or U2602 (N_2602,In_548,In_1078);
nor U2603 (N_2603,In_1098,In_428);
xor U2604 (N_2604,In_515,In_2046);
nor U2605 (N_2605,In_1618,In_1568);
nor U2606 (N_2606,In_903,In_673);
nor U2607 (N_2607,In_1987,In_1759);
and U2608 (N_2608,In_1635,In_494);
and U2609 (N_2609,In_1315,In_2269);
and U2610 (N_2610,In_590,In_1564);
nor U2611 (N_2611,In_1991,In_1106);
and U2612 (N_2612,In_2431,In_58);
nand U2613 (N_2613,In_1740,In_216);
nand U2614 (N_2614,In_668,In_2217);
nor U2615 (N_2615,In_1052,In_2163);
nor U2616 (N_2616,In_2149,In_1758);
or U2617 (N_2617,In_1745,In_2474);
nand U2618 (N_2618,In_2081,In_2390);
nand U2619 (N_2619,In_1615,In_831);
nor U2620 (N_2620,In_2424,In_79);
nand U2621 (N_2621,In_1304,In_185);
or U2622 (N_2622,In_1261,In_2325);
or U2623 (N_2623,In_323,In_901);
nand U2624 (N_2624,In_1320,In_1538);
nand U2625 (N_2625,In_280,In_2330);
nand U2626 (N_2626,In_1207,In_1674);
nor U2627 (N_2627,In_1939,In_2294);
and U2628 (N_2628,In_1585,In_914);
and U2629 (N_2629,In_78,In_2178);
or U2630 (N_2630,In_835,In_1255);
and U2631 (N_2631,In_2171,In_875);
and U2632 (N_2632,In_941,In_1715);
nand U2633 (N_2633,In_331,In_1531);
nor U2634 (N_2634,In_1653,In_2183);
and U2635 (N_2635,In_235,In_791);
and U2636 (N_2636,In_1946,In_140);
nor U2637 (N_2637,In_10,In_1288);
xor U2638 (N_2638,In_751,In_1445);
nand U2639 (N_2639,In_1755,In_1225);
nand U2640 (N_2640,In_780,In_2379);
and U2641 (N_2641,In_1533,In_548);
or U2642 (N_2642,In_720,In_908);
nor U2643 (N_2643,In_1815,In_1855);
xnor U2644 (N_2644,In_277,In_716);
nor U2645 (N_2645,In_622,In_221);
and U2646 (N_2646,In_510,In_768);
nor U2647 (N_2647,In_126,In_1760);
and U2648 (N_2648,In_148,In_1750);
or U2649 (N_2649,In_1666,In_637);
xnor U2650 (N_2650,In_1617,In_1201);
and U2651 (N_2651,In_1054,In_1483);
nand U2652 (N_2652,In_1721,In_2118);
and U2653 (N_2653,In_1497,In_1587);
xor U2654 (N_2654,In_381,In_972);
or U2655 (N_2655,In_784,In_726);
and U2656 (N_2656,In_2357,In_516);
nand U2657 (N_2657,In_1054,In_913);
nor U2658 (N_2658,In_252,In_1247);
or U2659 (N_2659,In_1171,In_1674);
or U2660 (N_2660,In_187,In_1135);
and U2661 (N_2661,In_795,In_974);
xor U2662 (N_2662,In_957,In_1841);
and U2663 (N_2663,In_1866,In_43);
nor U2664 (N_2664,In_2167,In_1437);
nand U2665 (N_2665,In_1226,In_450);
and U2666 (N_2666,In_530,In_1849);
or U2667 (N_2667,In_796,In_497);
xor U2668 (N_2668,In_1130,In_2055);
nor U2669 (N_2669,In_1587,In_792);
and U2670 (N_2670,In_1487,In_2278);
nor U2671 (N_2671,In_684,In_1968);
nor U2672 (N_2672,In_1846,In_1728);
nor U2673 (N_2673,In_848,In_2170);
nor U2674 (N_2674,In_2496,In_2285);
or U2675 (N_2675,In_502,In_2193);
xor U2676 (N_2676,In_666,In_599);
or U2677 (N_2677,In_7,In_2496);
or U2678 (N_2678,In_952,In_1489);
and U2679 (N_2679,In_2225,In_869);
or U2680 (N_2680,In_2202,In_66);
nor U2681 (N_2681,In_1985,In_1807);
xor U2682 (N_2682,In_81,In_1194);
nand U2683 (N_2683,In_2397,In_1311);
xor U2684 (N_2684,In_17,In_1964);
and U2685 (N_2685,In_2017,In_165);
or U2686 (N_2686,In_1527,In_733);
xnor U2687 (N_2687,In_1918,In_937);
nand U2688 (N_2688,In_1740,In_2100);
nand U2689 (N_2689,In_213,In_1282);
and U2690 (N_2690,In_2315,In_1817);
nor U2691 (N_2691,In_90,In_1357);
or U2692 (N_2692,In_709,In_976);
or U2693 (N_2693,In_1602,In_2412);
and U2694 (N_2694,In_1387,In_1123);
and U2695 (N_2695,In_1179,In_530);
nor U2696 (N_2696,In_1872,In_1819);
nand U2697 (N_2697,In_1218,In_2383);
or U2698 (N_2698,In_217,In_1206);
nor U2699 (N_2699,In_1280,In_2417);
nor U2700 (N_2700,In_881,In_66);
or U2701 (N_2701,In_332,In_921);
and U2702 (N_2702,In_695,In_584);
and U2703 (N_2703,In_788,In_1196);
or U2704 (N_2704,In_2420,In_368);
and U2705 (N_2705,In_1425,In_1403);
nor U2706 (N_2706,In_296,In_805);
nand U2707 (N_2707,In_789,In_2265);
nor U2708 (N_2708,In_7,In_395);
and U2709 (N_2709,In_2132,In_1490);
and U2710 (N_2710,In_1995,In_427);
and U2711 (N_2711,In_1919,In_33);
and U2712 (N_2712,In_965,In_2043);
or U2713 (N_2713,In_420,In_807);
or U2714 (N_2714,In_440,In_1160);
nor U2715 (N_2715,In_1934,In_407);
or U2716 (N_2716,In_438,In_541);
nand U2717 (N_2717,In_1169,In_807);
or U2718 (N_2718,In_1307,In_1323);
nand U2719 (N_2719,In_1413,In_1214);
nand U2720 (N_2720,In_1708,In_1355);
and U2721 (N_2721,In_1314,In_1905);
nor U2722 (N_2722,In_2161,In_1567);
nand U2723 (N_2723,In_1792,In_26);
nand U2724 (N_2724,In_180,In_28);
and U2725 (N_2725,In_1603,In_429);
and U2726 (N_2726,In_30,In_1839);
or U2727 (N_2727,In_2,In_1112);
nand U2728 (N_2728,In_2065,In_1869);
or U2729 (N_2729,In_287,In_1794);
xor U2730 (N_2730,In_1090,In_21);
or U2731 (N_2731,In_2203,In_2143);
nor U2732 (N_2732,In_2338,In_2375);
xor U2733 (N_2733,In_100,In_520);
or U2734 (N_2734,In_133,In_2033);
and U2735 (N_2735,In_20,In_1207);
and U2736 (N_2736,In_405,In_533);
and U2737 (N_2737,In_2154,In_242);
and U2738 (N_2738,In_2002,In_314);
nand U2739 (N_2739,In_1749,In_942);
nor U2740 (N_2740,In_1012,In_603);
or U2741 (N_2741,In_2019,In_2323);
nor U2742 (N_2742,In_822,In_1484);
nor U2743 (N_2743,In_283,In_675);
or U2744 (N_2744,In_201,In_2321);
and U2745 (N_2745,In_741,In_195);
or U2746 (N_2746,In_351,In_825);
xnor U2747 (N_2747,In_655,In_835);
nand U2748 (N_2748,In_1535,In_1069);
nor U2749 (N_2749,In_762,In_1529);
nand U2750 (N_2750,In_2446,In_2086);
nor U2751 (N_2751,In_1250,In_1045);
nor U2752 (N_2752,In_2077,In_1150);
or U2753 (N_2753,In_1626,In_994);
or U2754 (N_2754,In_322,In_577);
nor U2755 (N_2755,In_1132,In_1042);
nor U2756 (N_2756,In_1728,In_974);
nor U2757 (N_2757,In_2401,In_125);
xnor U2758 (N_2758,In_1880,In_786);
or U2759 (N_2759,In_1403,In_1003);
and U2760 (N_2760,In_321,In_2333);
or U2761 (N_2761,In_105,In_1996);
or U2762 (N_2762,In_1000,In_1969);
nand U2763 (N_2763,In_2143,In_1495);
and U2764 (N_2764,In_948,In_1609);
and U2765 (N_2765,In_2061,In_594);
nor U2766 (N_2766,In_2134,In_360);
nand U2767 (N_2767,In_1706,In_1572);
nand U2768 (N_2768,In_1594,In_1739);
nor U2769 (N_2769,In_241,In_699);
nand U2770 (N_2770,In_354,In_1287);
nor U2771 (N_2771,In_1396,In_1317);
or U2772 (N_2772,In_331,In_2324);
and U2773 (N_2773,In_472,In_1332);
and U2774 (N_2774,In_166,In_385);
and U2775 (N_2775,In_2418,In_1042);
or U2776 (N_2776,In_1291,In_32);
xor U2777 (N_2777,In_1417,In_1638);
or U2778 (N_2778,In_2095,In_537);
nand U2779 (N_2779,In_493,In_1856);
or U2780 (N_2780,In_1645,In_25);
and U2781 (N_2781,In_2345,In_261);
xor U2782 (N_2782,In_2472,In_320);
xor U2783 (N_2783,In_409,In_433);
nor U2784 (N_2784,In_1070,In_417);
and U2785 (N_2785,In_366,In_1255);
or U2786 (N_2786,In_1632,In_411);
nand U2787 (N_2787,In_75,In_215);
and U2788 (N_2788,In_1791,In_1650);
or U2789 (N_2789,In_1964,In_106);
nand U2790 (N_2790,In_1441,In_1395);
xor U2791 (N_2791,In_2306,In_2302);
and U2792 (N_2792,In_1982,In_427);
nand U2793 (N_2793,In_1582,In_1810);
xor U2794 (N_2794,In_1296,In_2422);
nor U2795 (N_2795,In_697,In_746);
or U2796 (N_2796,In_350,In_2314);
nor U2797 (N_2797,In_560,In_1292);
nor U2798 (N_2798,In_41,In_2130);
nand U2799 (N_2799,In_967,In_914);
and U2800 (N_2800,In_266,In_373);
nand U2801 (N_2801,In_658,In_124);
and U2802 (N_2802,In_359,In_1391);
or U2803 (N_2803,In_2416,In_683);
and U2804 (N_2804,In_1335,In_2309);
nor U2805 (N_2805,In_740,In_505);
and U2806 (N_2806,In_1499,In_2330);
xnor U2807 (N_2807,In_413,In_339);
nand U2808 (N_2808,In_1208,In_209);
nand U2809 (N_2809,In_1494,In_590);
xnor U2810 (N_2810,In_1578,In_2339);
or U2811 (N_2811,In_2288,In_890);
and U2812 (N_2812,In_1603,In_1026);
and U2813 (N_2813,In_2034,In_1456);
nor U2814 (N_2814,In_890,In_51);
nor U2815 (N_2815,In_1929,In_1638);
nand U2816 (N_2816,In_167,In_36);
xor U2817 (N_2817,In_58,In_2107);
nor U2818 (N_2818,In_73,In_2099);
nand U2819 (N_2819,In_537,In_1056);
xor U2820 (N_2820,In_2354,In_1755);
nand U2821 (N_2821,In_1961,In_221);
nor U2822 (N_2822,In_618,In_1801);
and U2823 (N_2823,In_173,In_776);
nand U2824 (N_2824,In_1265,In_529);
or U2825 (N_2825,In_1943,In_1066);
nor U2826 (N_2826,In_2126,In_811);
and U2827 (N_2827,In_331,In_2216);
nand U2828 (N_2828,In_2093,In_1847);
nor U2829 (N_2829,In_1586,In_2394);
xnor U2830 (N_2830,In_1757,In_46);
xor U2831 (N_2831,In_1279,In_1886);
nor U2832 (N_2832,In_2303,In_1514);
and U2833 (N_2833,In_557,In_1289);
nor U2834 (N_2834,In_546,In_845);
and U2835 (N_2835,In_2438,In_1070);
nor U2836 (N_2836,In_895,In_1215);
nand U2837 (N_2837,In_2221,In_1678);
nor U2838 (N_2838,In_2372,In_615);
or U2839 (N_2839,In_258,In_2320);
xor U2840 (N_2840,In_1649,In_794);
nand U2841 (N_2841,In_2336,In_2130);
nor U2842 (N_2842,In_1981,In_1574);
nand U2843 (N_2843,In_1736,In_2167);
and U2844 (N_2844,In_1964,In_2495);
or U2845 (N_2845,In_2481,In_1338);
nor U2846 (N_2846,In_740,In_2469);
nor U2847 (N_2847,In_539,In_791);
nand U2848 (N_2848,In_778,In_61);
and U2849 (N_2849,In_1600,In_1798);
and U2850 (N_2850,In_864,In_1757);
and U2851 (N_2851,In_2319,In_965);
and U2852 (N_2852,In_1575,In_2254);
xor U2853 (N_2853,In_1018,In_331);
xor U2854 (N_2854,In_1895,In_951);
nor U2855 (N_2855,In_1516,In_1416);
nor U2856 (N_2856,In_1949,In_1391);
nand U2857 (N_2857,In_196,In_1981);
or U2858 (N_2858,In_2265,In_2268);
xor U2859 (N_2859,In_349,In_1241);
or U2860 (N_2860,In_1286,In_2111);
or U2861 (N_2861,In_1423,In_507);
or U2862 (N_2862,In_2380,In_988);
nand U2863 (N_2863,In_2444,In_1833);
and U2864 (N_2864,In_216,In_1239);
nor U2865 (N_2865,In_359,In_2253);
or U2866 (N_2866,In_2169,In_1595);
nor U2867 (N_2867,In_1587,In_1629);
nand U2868 (N_2868,In_2072,In_1759);
and U2869 (N_2869,In_1595,In_1929);
and U2870 (N_2870,In_1649,In_1952);
or U2871 (N_2871,In_303,In_1059);
xnor U2872 (N_2872,In_1455,In_2123);
or U2873 (N_2873,In_499,In_2483);
nor U2874 (N_2874,In_2364,In_816);
nor U2875 (N_2875,In_1773,In_591);
xnor U2876 (N_2876,In_394,In_1027);
and U2877 (N_2877,In_1499,In_86);
nor U2878 (N_2878,In_123,In_1230);
nor U2879 (N_2879,In_473,In_1607);
xor U2880 (N_2880,In_2339,In_1055);
or U2881 (N_2881,In_1058,In_2471);
nand U2882 (N_2882,In_2221,In_881);
nor U2883 (N_2883,In_996,In_1844);
nor U2884 (N_2884,In_1599,In_1425);
xnor U2885 (N_2885,In_2350,In_2248);
nor U2886 (N_2886,In_1700,In_2131);
nand U2887 (N_2887,In_1059,In_1340);
and U2888 (N_2888,In_11,In_2041);
nor U2889 (N_2889,In_593,In_313);
nor U2890 (N_2890,In_592,In_1947);
nor U2891 (N_2891,In_1527,In_1482);
nor U2892 (N_2892,In_2318,In_2092);
nor U2893 (N_2893,In_786,In_287);
nor U2894 (N_2894,In_2449,In_1833);
xor U2895 (N_2895,In_689,In_2189);
nand U2896 (N_2896,In_859,In_2379);
xor U2897 (N_2897,In_1398,In_617);
nor U2898 (N_2898,In_490,In_1737);
or U2899 (N_2899,In_91,In_1029);
and U2900 (N_2900,In_568,In_2444);
and U2901 (N_2901,In_1732,In_371);
or U2902 (N_2902,In_69,In_1022);
nand U2903 (N_2903,In_1490,In_2126);
or U2904 (N_2904,In_2162,In_307);
nor U2905 (N_2905,In_1544,In_2474);
or U2906 (N_2906,In_94,In_2245);
nor U2907 (N_2907,In_1095,In_1422);
nor U2908 (N_2908,In_347,In_619);
nor U2909 (N_2909,In_1476,In_694);
or U2910 (N_2910,In_1081,In_156);
nor U2911 (N_2911,In_1568,In_771);
and U2912 (N_2912,In_1841,In_1625);
nor U2913 (N_2913,In_2293,In_1138);
nand U2914 (N_2914,In_230,In_2106);
and U2915 (N_2915,In_1570,In_247);
nor U2916 (N_2916,In_2334,In_309);
nand U2917 (N_2917,In_245,In_1216);
nand U2918 (N_2918,In_881,In_1102);
and U2919 (N_2919,In_277,In_2470);
nand U2920 (N_2920,In_2083,In_2408);
or U2921 (N_2921,In_889,In_1540);
nor U2922 (N_2922,In_1833,In_980);
xnor U2923 (N_2923,In_1959,In_1217);
or U2924 (N_2924,In_1634,In_841);
xnor U2925 (N_2925,In_2177,In_1474);
nor U2926 (N_2926,In_629,In_978);
or U2927 (N_2927,In_1064,In_2255);
or U2928 (N_2928,In_1396,In_2224);
nand U2929 (N_2929,In_1407,In_188);
or U2930 (N_2930,In_2233,In_1151);
or U2931 (N_2931,In_815,In_1325);
nor U2932 (N_2932,In_506,In_2149);
nand U2933 (N_2933,In_83,In_2064);
xor U2934 (N_2934,In_1628,In_153);
and U2935 (N_2935,In_1112,In_1422);
nor U2936 (N_2936,In_2292,In_1242);
nand U2937 (N_2937,In_1623,In_744);
and U2938 (N_2938,In_1828,In_1469);
xnor U2939 (N_2939,In_214,In_401);
nor U2940 (N_2940,In_580,In_2262);
or U2941 (N_2941,In_1474,In_90);
nor U2942 (N_2942,In_785,In_973);
and U2943 (N_2943,In_1738,In_337);
or U2944 (N_2944,In_1676,In_694);
nand U2945 (N_2945,In_742,In_256);
or U2946 (N_2946,In_1558,In_1759);
nand U2947 (N_2947,In_1026,In_590);
nand U2948 (N_2948,In_63,In_369);
nor U2949 (N_2949,In_1526,In_1497);
xor U2950 (N_2950,In_1387,In_1808);
nor U2951 (N_2951,In_1746,In_1096);
and U2952 (N_2952,In_272,In_400);
or U2953 (N_2953,In_263,In_64);
nand U2954 (N_2954,In_1250,In_902);
xor U2955 (N_2955,In_699,In_1176);
nand U2956 (N_2956,In_1888,In_2250);
nand U2957 (N_2957,In_765,In_1749);
and U2958 (N_2958,In_576,In_1830);
nor U2959 (N_2959,In_2136,In_1404);
and U2960 (N_2960,In_1978,In_1250);
nand U2961 (N_2961,In_2088,In_524);
and U2962 (N_2962,In_2438,In_819);
or U2963 (N_2963,In_385,In_843);
or U2964 (N_2964,In_2442,In_875);
xnor U2965 (N_2965,In_1223,In_1550);
or U2966 (N_2966,In_2327,In_2238);
xor U2967 (N_2967,In_2394,In_1321);
or U2968 (N_2968,In_1888,In_1339);
nor U2969 (N_2969,In_1844,In_881);
nand U2970 (N_2970,In_1446,In_1357);
and U2971 (N_2971,In_683,In_373);
and U2972 (N_2972,In_2046,In_1840);
and U2973 (N_2973,In_2305,In_2262);
nor U2974 (N_2974,In_1129,In_1321);
and U2975 (N_2975,In_2047,In_2497);
and U2976 (N_2976,In_711,In_919);
and U2977 (N_2977,In_184,In_826);
or U2978 (N_2978,In_1117,In_2309);
nand U2979 (N_2979,In_1834,In_2456);
nand U2980 (N_2980,In_2114,In_1104);
and U2981 (N_2981,In_829,In_2465);
nor U2982 (N_2982,In_1426,In_750);
or U2983 (N_2983,In_929,In_720);
or U2984 (N_2984,In_1584,In_2363);
or U2985 (N_2985,In_2222,In_2151);
and U2986 (N_2986,In_2077,In_742);
nor U2987 (N_2987,In_1311,In_1484);
and U2988 (N_2988,In_1067,In_1400);
and U2989 (N_2989,In_2133,In_854);
or U2990 (N_2990,In_834,In_1079);
or U2991 (N_2991,In_1493,In_1155);
or U2992 (N_2992,In_863,In_1394);
nand U2993 (N_2993,In_763,In_1746);
and U2994 (N_2994,In_1659,In_1643);
and U2995 (N_2995,In_1229,In_623);
nor U2996 (N_2996,In_2283,In_1276);
nand U2997 (N_2997,In_824,In_174);
nor U2998 (N_2998,In_433,In_1538);
and U2999 (N_2999,In_2120,In_499);
and U3000 (N_3000,In_712,In_2309);
or U3001 (N_3001,In_924,In_1215);
nand U3002 (N_3002,In_1243,In_2125);
and U3003 (N_3003,In_805,In_217);
nand U3004 (N_3004,In_1622,In_1712);
and U3005 (N_3005,In_1381,In_1605);
nand U3006 (N_3006,In_2157,In_1374);
nand U3007 (N_3007,In_1523,In_1294);
xnor U3008 (N_3008,In_367,In_644);
nor U3009 (N_3009,In_1789,In_145);
nand U3010 (N_3010,In_2122,In_283);
or U3011 (N_3011,In_343,In_2019);
nor U3012 (N_3012,In_2316,In_2214);
and U3013 (N_3013,In_2346,In_1590);
or U3014 (N_3014,In_1017,In_2464);
nand U3015 (N_3015,In_1419,In_427);
nand U3016 (N_3016,In_1243,In_1601);
and U3017 (N_3017,In_1356,In_1271);
or U3018 (N_3018,In_516,In_812);
and U3019 (N_3019,In_2278,In_1605);
and U3020 (N_3020,In_768,In_490);
nand U3021 (N_3021,In_962,In_1275);
nand U3022 (N_3022,In_175,In_33);
nor U3023 (N_3023,In_2472,In_914);
or U3024 (N_3024,In_85,In_271);
nand U3025 (N_3025,In_329,In_998);
and U3026 (N_3026,In_2308,In_1922);
xor U3027 (N_3027,In_1122,In_1572);
and U3028 (N_3028,In_89,In_1445);
and U3029 (N_3029,In_1319,In_1367);
nand U3030 (N_3030,In_2164,In_1830);
nand U3031 (N_3031,In_724,In_78);
xor U3032 (N_3032,In_689,In_1622);
nand U3033 (N_3033,In_1725,In_2439);
nand U3034 (N_3034,In_1852,In_1637);
nor U3035 (N_3035,In_179,In_1797);
or U3036 (N_3036,In_1594,In_2437);
or U3037 (N_3037,In_2471,In_243);
nor U3038 (N_3038,In_698,In_1700);
xor U3039 (N_3039,In_19,In_1597);
nand U3040 (N_3040,In_2007,In_2016);
nor U3041 (N_3041,In_750,In_148);
or U3042 (N_3042,In_172,In_2415);
or U3043 (N_3043,In_251,In_2255);
or U3044 (N_3044,In_2078,In_1372);
xnor U3045 (N_3045,In_1937,In_935);
xnor U3046 (N_3046,In_1709,In_1935);
nand U3047 (N_3047,In_2312,In_976);
nand U3048 (N_3048,In_2178,In_1074);
and U3049 (N_3049,In_2493,In_1740);
and U3050 (N_3050,In_199,In_1398);
or U3051 (N_3051,In_2000,In_1661);
or U3052 (N_3052,In_415,In_1087);
nand U3053 (N_3053,In_1691,In_945);
xnor U3054 (N_3054,In_936,In_1331);
xnor U3055 (N_3055,In_1040,In_313);
nor U3056 (N_3056,In_1288,In_2210);
and U3057 (N_3057,In_914,In_955);
and U3058 (N_3058,In_536,In_2453);
and U3059 (N_3059,In_1654,In_1506);
or U3060 (N_3060,In_981,In_1931);
and U3061 (N_3061,In_1270,In_1343);
or U3062 (N_3062,In_210,In_882);
or U3063 (N_3063,In_2399,In_1534);
nand U3064 (N_3064,In_872,In_2077);
nor U3065 (N_3065,In_1281,In_2479);
or U3066 (N_3066,In_2316,In_1590);
or U3067 (N_3067,In_1678,In_2241);
or U3068 (N_3068,In_390,In_810);
or U3069 (N_3069,In_2020,In_401);
xnor U3070 (N_3070,In_813,In_115);
nand U3071 (N_3071,In_1178,In_2437);
or U3072 (N_3072,In_2068,In_2456);
nor U3073 (N_3073,In_31,In_271);
or U3074 (N_3074,In_1493,In_1112);
or U3075 (N_3075,In_1385,In_1506);
nor U3076 (N_3076,In_380,In_2421);
or U3077 (N_3077,In_112,In_1853);
and U3078 (N_3078,In_2492,In_1327);
nand U3079 (N_3079,In_1086,In_1522);
nor U3080 (N_3080,In_1387,In_2047);
and U3081 (N_3081,In_1638,In_1380);
and U3082 (N_3082,In_398,In_1690);
or U3083 (N_3083,In_24,In_601);
nor U3084 (N_3084,In_1952,In_1262);
xnor U3085 (N_3085,In_1134,In_1622);
or U3086 (N_3086,In_1838,In_1173);
and U3087 (N_3087,In_2452,In_793);
and U3088 (N_3088,In_1814,In_171);
and U3089 (N_3089,In_2128,In_452);
or U3090 (N_3090,In_1057,In_1643);
nand U3091 (N_3091,In_2160,In_170);
xnor U3092 (N_3092,In_504,In_2248);
nand U3093 (N_3093,In_945,In_1694);
and U3094 (N_3094,In_1380,In_1605);
nor U3095 (N_3095,In_166,In_581);
nor U3096 (N_3096,In_552,In_878);
or U3097 (N_3097,In_581,In_2087);
and U3098 (N_3098,In_367,In_1338);
nor U3099 (N_3099,In_2091,In_1141);
nand U3100 (N_3100,In_1430,In_1193);
and U3101 (N_3101,In_289,In_2285);
or U3102 (N_3102,In_886,In_1809);
nand U3103 (N_3103,In_1979,In_1732);
nand U3104 (N_3104,In_2243,In_477);
or U3105 (N_3105,In_405,In_1342);
nand U3106 (N_3106,In_599,In_1615);
or U3107 (N_3107,In_516,In_653);
nor U3108 (N_3108,In_791,In_2222);
and U3109 (N_3109,In_2135,In_2436);
nor U3110 (N_3110,In_2263,In_534);
and U3111 (N_3111,In_1444,In_1045);
xnor U3112 (N_3112,In_148,In_2095);
xnor U3113 (N_3113,In_1617,In_88);
and U3114 (N_3114,In_169,In_1633);
and U3115 (N_3115,In_874,In_1270);
nand U3116 (N_3116,In_1551,In_1625);
and U3117 (N_3117,In_1008,In_332);
nor U3118 (N_3118,In_2015,In_140);
and U3119 (N_3119,In_2165,In_2395);
nand U3120 (N_3120,In_1335,In_1196);
nor U3121 (N_3121,In_978,In_749);
xor U3122 (N_3122,In_2437,In_1352);
and U3123 (N_3123,In_455,In_1374);
nand U3124 (N_3124,In_1746,In_1264);
nand U3125 (N_3125,In_1652,In_734);
and U3126 (N_3126,In_1313,In_2427);
nand U3127 (N_3127,In_2426,In_78);
and U3128 (N_3128,In_1163,In_385);
nand U3129 (N_3129,In_950,In_1321);
or U3130 (N_3130,In_401,In_118);
and U3131 (N_3131,In_2497,In_916);
nor U3132 (N_3132,In_1479,In_470);
nor U3133 (N_3133,In_1104,In_109);
nand U3134 (N_3134,In_1987,In_2107);
and U3135 (N_3135,In_560,In_1966);
nand U3136 (N_3136,In_1991,In_2126);
nor U3137 (N_3137,In_1417,In_1312);
nand U3138 (N_3138,In_537,In_9);
and U3139 (N_3139,In_823,In_1872);
nor U3140 (N_3140,In_889,In_2127);
or U3141 (N_3141,In_1928,In_2104);
nor U3142 (N_3142,In_917,In_724);
and U3143 (N_3143,In_1650,In_349);
nor U3144 (N_3144,In_1362,In_1240);
nor U3145 (N_3145,In_2470,In_1699);
or U3146 (N_3146,In_1080,In_1671);
nand U3147 (N_3147,In_425,In_1465);
nor U3148 (N_3148,In_2451,In_2453);
and U3149 (N_3149,In_2067,In_1905);
nor U3150 (N_3150,In_870,In_896);
nand U3151 (N_3151,In_309,In_261);
nor U3152 (N_3152,In_1505,In_1547);
nand U3153 (N_3153,In_1827,In_1464);
nand U3154 (N_3154,In_397,In_260);
nand U3155 (N_3155,In_2150,In_177);
nand U3156 (N_3156,In_1274,In_45);
and U3157 (N_3157,In_1291,In_390);
or U3158 (N_3158,In_456,In_1090);
and U3159 (N_3159,In_283,In_1167);
nor U3160 (N_3160,In_448,In_524);
nor U3161 (N_3161,In_291,In_1627);
and U3162 (N_3162,In_1899,In_2432);
nor U3163 (N_3163,In_2232,In_413);
or U3164 (N_3164,In_1177,In_516);
or U3165 (N_3165,In_1622,In_954);
nor U3166 (N_3166,In_1288,In_184);
or U3167 (N_3167,In_1339,In_2000);
nor U3168 (N_3168,In_1102,In_1923);
nand U3169 (N_3169,In_605,In_13);
nor U3170 (N_3170,In_2291,In_2130);
nand U3171 (N_3171,In_2062,In_701);
nor U3172 (N_3172,In_2334,In_1868);
nor U3173 (N_3173,In_1982,In_892);
nor U3174 (N_3174,In_593,In_2077);
nor U3175 (N_3175,In_753,In_1040);
nand U3176 (N_3176,In_1511,In_1093);
nand U3177 (N_3177,In_1111,In_1976);
xnor U3178 (N_3178,In_984,In_623);
nand U3179 (N_3179,In_1138,In_594);
nand U3180 (N_3180,In_353,In_1409);
xor U3181 (N_3181,In_478,In_1101);
or U3182 (N_3182,In_406,In_1252);
or U3183 (N_3183,In_63,In_1474);
nand U3184 (N_3184,In_1872,In_219);
or U3185 (N_3185,In_1346,In_1909);
nor U3186 (N_3186,In_2349,In_1746);
nand U3187 (N_3187,In_1691,In_526);
nor U3188 (N_3188,In_1630,In_1975);
and U3189 (N_3189,In_756,In_1357);
and U3190 (N_3190,In_2464,In_820);
nor U3191 (N_3191,In_2424,In_195);
nor U3192 (N_3192,In_2341,In_1394);
nand U3193 (N_3193,In_1252,In_1267);
nand U3194 (N_3194,In_316,In_1668);
or U3195 (N_3195,In_1230,In_752);
nor U3196 (N_3196,In_1100,In_211);
and U3197 (N_3197,In_1655,In_1589);
and U3198 (N_3198,In_1648,In_1998);
nand U3199 (N_3199,In_1703,In_2301);
nor U3200 (N_3200,In_946,In_2041);
and U3201 (N_3201,In_454,In_1008);
xnor U3202 (N_3202,In_2171,In_775);
xnor U3203 (N_3203,In_1928,In_483);
nor U3204 (N_3204,In_1485,In_1014);
or U3205 (N_3205,In_1362,In_760);
and U3206 (N_3206,In_31,In_740);
nor U3207 (N_3207,In_149,In_947);
nor U3208 (N_3208,In_2059,In_1536);
and U3209 (N_3209,In_619,In_139);
or U3210 (N_3210,In_594,In_323);
xnor U3211 (N_3211,In_2215,In_249);
nand U3212 (N_3212,In_1596,In_591);
or U3213 (N_3213,In_2138,In_2192);
or U3214 (N_3214,In_1310,In_306);
or U3215 (N_3215,In_1846,In_512);
and U3216 (N_3216,In_873,In_907);
nand U3217 (N_3217,In_1006,In_220);
or U3218 (N_3218,In_1688,In_745);
xor U3219 (N_3219,In_2094,In_940);
or U3220 (N_3220,In_1365,In_1546);
and U3221 (N_3221,In_552,In_2046);
and U3222 (N_3222,In_247,In_1690);
nand U3223 (N_3223,In_1660,In_1956);
and U3224 (N_3224,In_711,In_1503);
nand U3225 (N_3225,In_388,In_1580);
and U3226 (N_3226,In_396,In_2243);
or U3227 (N_3227,In_1079,In_460);
nand U3228 (N_3228,In_429,In_574);
or U3229 (N_3229,In_1728,In_1682);
nor U3230 (N_3230,In_106,In_1199);
and U3231 (N_3231,In_573,In_2302);
nand U3232 (N_3232,In_1561,In_2420);
or U3233 (N_3233,In_2126,In_2412);
nand U3234 (N_3234,In_1382,In_2182);
and U3235 (N_3235,In_87,In_2386);
nand U3236 (N_3236,In_1261,In_989);
and U3237 (N_3237,In_1957,In_1445);
nor U3238 (N_3238,In_822,In_2269);
nor U3239 (N_3239,In_2038,In_1372);
or U3240 (N_3240,In_22,In_1712);
xor U3241 (N_3241,In_1637,In_1027);
nand U3242 (N_3242,In_1459,In_1236);
xor U3243 (N_3243,In_727,In_2486);
nor U3244 (N_3244,In_463,In_1655);
nand U3245 (N_3245,In_2029,In_1293);
and U3246 (N_3246,In_1752,In_462);
xor U3247 (N_3247,In_1630,In_563);
nor U3248 (N_3248,In_31,In_321);
and U3249 (N_3249,In_909,In_872);
or U3250 (N_3250,In_626,In_1584);
or U3251 (N_3251,In_463,In_403);
and U3252 (N_3252,In_1177,In_2143);
or U3253 (N_3253,In_498,In_118);
or U3254 (N_3254,In_1918,In_698);
nand U3255 (N_3255,In_1090,In_475);
or U3256 (N_3256,In_1708,In_421);
or U3257 (N_3257,In_2004,In_1629);
or U3258 (N_3258,In_1601,In_1462);
or U3259 (N_3259,In_615,In_1404);
nand U3260 (N_3260,In_1342,In_2162);
nand U3261 (N_3261,In_587,In_11);
nand U3262 (N_3262,In_634,In_79);
nor U3263 (N_3263,In_276,In_1378);
and U3264 (N_3264,In_510,In_1366);
nand U3265 (N_3265,In_1442,In_1086);
nand U3266 (N_3266,In_2085,In_134);
or U3267 (N_3267,In_1890,In_762);
nor U3268 (N_3268,In_744,In_2030);
and U3269 (N_3269,In_472,In_608);
nand U3270 (N_3270,In_2080,In_865);
nand U3271 (N_3271,In_1480,In_102);
nor U3272 (N_3272,In_1576,In_969);
or U3273 (N_3273,In_1138,In_784);
nor U3274 (N_3274,In_21,In_1726);
or U3275 (N_3275,In_2251,In_1369);
and U3276 (N_3276,In_1772,In_583);
or U3277 (N_3277,In_1302,In_1380);
and U3278 (N_3278,In_1189,In_1762);
and U3279 (N_3279,In_1630,In_1132);
xnor U3280 (N_3280,In_1001,In_2141);
or U3281 (N_3281,In_159,In_136);
and U3282 (N_3282,In_2112,In_795);
nor U3283 (N_3283,In_1869,In_543);
nand U3284 (N_3284,In_960,In_1276);
nand U3285 (N_3285,In_2071,In_1469);
or U3286 (N_3286,In_190,In_40);
nor U3287 (N_3287,In_1672,In_662);
and U3288 (N_3288,In_76,In_731);
or U3289 (N_3289,In_1703,In_691);
nand U3290 (N_3290,In_1898,In_2034);
or U3291 (N_3291,In_859,In_2453);
or U3292 (N_3292,In_1347,In_1927);
or U3293 (N_3293,In_370,In_928);
nand U3294 (N_3294,In_601,In_985);
nand U3295 (N_3295,In_819,In_1991);
nor U3296 (N_3296,In_1590,In_1776);
and U3297 (N_3297,In_787,In_48);
nor U3298 (N_3298,In_1254,In_457);
nand U3299 (N_3299,In_2253,In_2041);
nand U3300 (N_3300,In_1945,In_1511);
nor U3301 (N_3301,In_1471,In_768);
nor U3302 (N_3302,In_449,In_582);
or U3303 (N_3303,In_1333,In_1433);
xnor U3304 (N_3304,In_1773,In_2180);
and U3305 (N_3305,In_1739,In_2421);
and U3306 (N_3306,In_722,In_1863);
nor U3307 (N_3307,In_56,In_225);
or U3308 (N_3308,In_1183,In_1677);
and U3309 (N_3309,In_1423,In_1929);
or U3310 (N_3310,In_1210,In_900);
or U3311 (N_3311,In_281,In_87);
nand U3312 (N_3312,In_1241,In_447);
and U3313 (N_3313,In_1112,In_2399);
and U3314 (N_3314,In_1513,In_1415);
nand U3315 (N_3315,In_813,In_1592);
and U3316 (N_3316,In_1466,In_1741);
or U3317 (N_3317,In_1855,In_1556);
nor U3318 (N_3318,In_767,In_203);
nand U3319 (N_3319,In_742,In_1714);
nand U3320 (N_3320,In_1266,In_627);
nand U3321 (N_3321,In_2345,In_2224);
nor U3322 (N_3322,In_2251,In_1757);
nand U3323 (N_3323,In_1921,In_1661);
xor U3324 (N_3324,In_217,In_1321);
nor U3325 (N_3325,In_1588,In_2427);
or U3326 (N_3326,In_234,In_1408);
nor U3327 (N_3327,In_2411,In_283);
and U3328 (N_3328,In_474,In_1515);
and U3329 (N_3329,In_436,In_2155);
xnor U3330 (N_3330,In_1202,In_2279);
or U3331 (N_3331,In_677,In_954);
nand U3332 (N_3332,In_839,In_869);
and U3333 (N_3333,In_1388,In_1205);
or U3334 (N_3334,In_6,In_565);
nor U3335 (N_3335,In_1713,In_1150);
nand U3336 (N_3336,In_981,In_669);
or U3337 (N_3337,In_928,In_1230);
and U3338 (N_3338,In_1245,In_2203);
nand U3339 (N_3339,In_1514,In_518);
nor U3340 (N_3340,In_698,In_1964);
nand U3341 (N_3341,In_1763,In_2009);
or U3342 (N_3342,In_2049,In_756);
and U3343 (N_3343,In_2337,In_1675);
nand U3344 (N_3344,In_2364,In_2277);
nand U3345 (N_3345,In_1893,In_1444);
nand U3346 (N_3346,In_1787,In_5);
or U3347 (N_3347,In_2497,In_2361);
and U3348 (N_3348,In_1834,In_609);
nor U3349 (N_3349,In_14,In_477);
or U3350 (N_3350,In_1416,In_690);
and U3351 (N_3351,In_1804,In_244);
nor U3352 (N_3352,In_1435,In_1035);
and U3353 (N_3353,In_2446,In_725);
nand U3354 (N_3354,In_1309,In_132);
nor U3355 (N_3355,In_1276,In_271);
nand U3356 (N_3356,In_1028,In_2025);
or U3357 (N_3357,In_794,In_2050);
or U3358 (N_3358,In_1361,In_1773);
nand U3359 (N_3359,In_1758,In_1949);
and U3360 (N_3360,In_2390,In_1518);
nor U3361 (N_3361,In_1690,In_1090);
and U3362 (N_3362,In_1539,In_2292);
nor U3363 (N_3363,In_1429,In_1099);
xor U3364 (N_3364,In_2462,In_1914);
nor U3365 (N_3365,In_2448,In_31);
and U3366 (N_3366,In_459,In_1163);
and U3367 (N_3367,In_2251,In_1672);
nand U3368 (N_3368,In_813,In_1704);
or U3369 (N_3369,In_1982,In_2119);
nand U3370 (N_3370,In_1761,In_2345);
or U3371 (N_3371,In_833,In_2153);
nand U3372 (N_3372,In_2230,In_1592);
or U3373 (N_3373,In_1869,In_380);
or U3374 (N_3374,In_1070,In_553);
xor U3375 (N_3375,In_1731,In_1845);
xor U3376 (N_3376,In_1897,In_1907);
nand U3377 (N_3377,In_1115,In_730);
xnor U3378 (N_3378,In_183,In_1376);
nor U3379 (N_3379,In_1155,In_820);
nand U3380 (N_3380,In_495,In_1098);
nor U3381 (N_3381,In_1221,In_1470);
nor U3382 (N_3382,In_1136,In_852);
or U3383 (N_3383,In_1857,In_1283);
nand U3384 (N_3384,In_1270,In_210);
nand U3385 (N_3385,In_151,In_1334);
nand U3386 (N_3386,In_1968,In_462);
nor U3387 (N_3387,In_1410,In_1568);
nand U3388 (N_3388,In_203,In_871);
nor U3389 (N_3389,In_1951,In_882);
or U3390 (N_3390,In_1884,In_1287);
nor U3391 (N_3391,In_1997,In_410);
and U3392 (N_3392,In_577,In_1132);
nor U3393 (N_3393,In_1912,In_203);
and U3394 (N_3394,In_1765,In_274);
or U3395 (N_3395,In_470,In_101);
or U3396 (N_3396,In_1886,In_257);
nor U3397 (N_3397,In_827,In_178);
nor U3398 (N_3398,In_389,In_2302);
nand U3399 (N_3399,In_1941,In_1803);
or U3400 (N_3400,In_2300,In_1949);
nor U3401 (N_3401,In_609,In_292);
nor U3402 (N_3402,In_1189,In_766);
and U3403 (N_3403,In_1688,In_1647);
or U3404 (N_3404,In_679,In_328);
or U3405 (N_3405,In_1858,In_2354);
nand U3406 (N_3406,In_192,In_1202);
nor U3407 (N_3407,In_2395,In_2374);
and U3408 (N_3408,In_2371,In_202);
and U3409 (N_3409,In_1534,In_1300);
or U3410 (N_3410,In_1838,In_1746);
nor U3411 (N_3411,In_1041,In_1918);
xor U3412 (N_3412,In_1668,In_1878);
nand U3413 (N_3413,In_1806,In_393);
nand U3414 (N_3414,In_1572,In_1823);
or U3415 (N_3415,In_1921,In_1650);
nand U3416 (N_3416,In_221,In_2005);
nor U3417 (N_3417,In_311,In_2167);
nor U3418 (N_3418,In_1341,In_1411);
and U3419 (N_3419,In_1352,In_1562);
nor U3420 (N_3420,In_1510,In_1603);
nand U3421 (N_3421,In_1906,In_287);
nand U3422 (N_3422,In_1436,In_1698);
and U3423 (N_3423,In_1311,In_1562);
and U3424 (N_3424,In_502,In_535);
nor U3425 (N_3425,In_2202,In_405);
or U3426 (N_3426,In_611,In_1999);
nor U3427 (N_3427,In_604,In_1851);
nand U3428 (N_3428,In_1525,In_1929);
and U3429 (N_3429,In_1930,In_1788);
nand U3430 (N_3430,In_145,In_1207);
or U3431 (N_3431,In_500,In_2392);
nor U3432 (N_3432,In_10,In_513);
or U3433 (N_3433,In_1615,In_846);
or U3434 (N_3434,In_2468,In_1928);
and U3435 (N_3435,In_629,In_380);
nor U3436 (N_3436,In_1933,In_161);
xnor U3437 (N_3437,In_1498,In_1218);
and U3438 (N_3438,In_504,In_1981);
or U3439 (N_3439,In_1322,In_567);
or U3440 (N_3440,In_990,In_2239);
nand U3441 (N_3441,In_23,In_797);
nor U3442 (N_3442,In_861,In_975);
or U3443 (N_3443,In_39,In_302);
nand U3444 (N_3444,In_2315,In_79);
xor U3445 (N_3445,In_31,In_1451);
or U3446 (N_3446,In_1657,In_387);
xor U3447 (N_3447,In_2174,In_1925);
nand U3448 (N_3448,In_1375,In_1935);
or U3449 (N_3449,In_863,In_1970);
nor U3450 (N_3450,In_945,In_543);
nand U3451 (N_3451,In_2200,In_1423);
xnor U3452 (N_3452,In_330,In_54);
or U3453 (N_3453,In_1810,In_2234);
nor U3454 (N_3454,In_1189,In_1348);
and U3455 (N_3455,In_2020,In_97);
and U3456 (N_3456,In_953,In_2420);
or U3457 (N_3457,In_1287,In_2291);
or U3458 (N_3458,In_203,In_1350);
or U3459 (N_3459,In_372,In_458);
nor U3460 (N_3460,In_1608,In_939);
xor U3461 (N_3461,In_2053,In_2083);
and U3462 (N_3462,In_2009,In_1341);
or U3463 (N_3463,In_1519,In_462);
nand U3464 (N_3464,In_2422,In_2266);
xor U3465 (N_3465,In_1970,In_707);
nand U3466 (N_3466,In_2057,In_964);
nor U3467 (N_3467,In_1577,In_989);
and U3468 (N_3468,In_1969,In_157);
nor U3469 (N_3469,In_2120,In_2478);
and U3470 (N_3470,In_1941,In_1279);
and U3471 (N_3471,In_850,In_865);
and U3472 (N_3472,In_931,In_1416);
nand U3473 (N_3473,In_1806,In_415);
and U3474 (N_3474,In_2166,In_251);
or U3475 (N_3475,In_961,In_425);
nand U3476 (N_3476,In_92,In_2362);
nor U3477 (N_3477,In_104,In_146);
nand U3478 (N_3478,In_388,In_317);
nor U3479 (N_3479,In_1699,In_1875);
or U3480 (N_3480,In_342,In_1005);
or U3481 (N_3481,In_311,In_790);
and U3482 (N_3482,In_676,In_1499);
or U3483 (N_3483,In_2016,In_2067);
and U3484 (N_3484,In_1866,In_749);
and U3485 (N_3485,In_429,In_1511);
nor U3486 (N_3486,In_1055,In_453);
nor U3487 (N_3487,In_1998,In_1132);
and U3488 (N_3488,In_954,In_1854);
or U3489 (N_3489,In_306,In_442);
nor U3490 (N_3490,In_2038,In_2103);
xor U3491 (N_3491,In_45,In_2304);
nand U3492 (N_3492,In_853,In_2296);
or U3493 (N_3493,In_641,In_1615);
nand U3494 (N_3494,In_1490,In_2354);
and U3495 (N_3495,In_2118,In_618);
nor U3496 (N_3496,In_882,In_201);
nand U3497 (N_3497,In_535,In_465);
and U3498 (N_3498,In_814,In_1786);
or U3499 (N_3499,In_2088,In_1319);
nor U3500 (N_3500,In_1616,In_1183);
or U3501 (N_3501,In_1147,In_1171);
nand U3502 (N_3502,In_1564,In_249);
or U3503 (N_3503,In_1062,In_1423);
nand U3504 (N_3504,In_288,In_2312);
or U3505 (N_3505,In_2192,In_1457);
nor U3506 (N_3506,In_280,In_143);
or U3507 (N_3507,In_1993,In_982);
and U3508 (N_3508,In_2071,In_1064);
nand U3509 (N_3509,In_912,In_1180);
xor U3510 (N_3510,In_1937,In_1932);
and U3511 (N_3511,In_1484,In_1089);
and U3512 (N_3512,In_2239,In_1157);
nand U3513 (N_3513,In_1302,In_735);
and U3514 (N_3514,In_1011,In_2001);
nand U3515 (N_3515,In_560,In_148);
xnor U3516 (N_3516,In_391,In_1411);
nor U3517 (N_3517,In_979,In_91);
nand U3518 (N_3518,In_1371,In_165);
nand U3519 (N_3519,In_2466,In_217);
and U3520 (N_3520,In_2205,In_996);
or U3521 (N_3521,In_972,In_1770);
or U3522 (N_3522,In_1153,In_273);
and U3523 (N_3523,In_500,In_1702);
or U3524 (N_3524,In_192,In_2456);
or U3525 (N_3525,In_1262,In_621);
nor U3526 (N_3526,In_2357,In_1551);
and U3527 (N_3527,In_109,In_611);
nand U3528 (N_3528,In_1634,In_3);
nor U3529 (N_3529,In_864,In_2213);
and U3530 (N_3530,In_1498,In_1471);
nand U3531 (N_3531,In_674,In_416);
xor U3532 (N_3532,In_1352,In_524);
xor U3533 (N_3533,In_2313,In_1956);
or U3534 (N_3534,In_467,In_818);
nand U3535 (N_3535,In_1327,In_1678);
and U3536 (N_3536,In_1644,In_277);
nor U3537 (N_3537,In_1441,In_1776);
and U3538 (N_3538,In_1323,In_2350);
nand U3539 (N_3539,In_1439,In_2176);
nor U3540 (N_3540,In_2038,In_2232);
nand U3541 (N_3541,In_903,In_1281);
xor U3542 (N_3542,In_734,In_2010);
nor U3543 (N_3543,In_245,In_1830);
nor U3544 (N_3544,In_1160,In_466);
nand U3545 (N_3545,In_2443,In_407);
or U3546 (N_3546,In_485,In_2417);
nor U3547 (N_3547,In_2369,In_172);
and U3548 (N_3548,In_2259,In_908);
or U3549 (N_3549,In_1458,In_982);
and U3550 (N_3550,In_1899,In_494);
and U3551 (N_3551,In_673,In_1079);
or U3552 (N_3552,In_418,In_1016);
nor U3553 (N_3553,In_244,In_1685);
and U3554 (N_3554,In_484,In_154);
and U3555 (N_3555,In_2128,In_590);
or U3556 (N_3556,In_570,In_1641);
nor U3557 (N_3557,In_1271,In_1253);
nand U3558 (N_3558,In_1821,In_849);
and U3559 (N_3559,In_2496,In_1110);
nand U3560 (N_3560,In_830,In_341);
and U3561 (N_3561,In_181,In_182);
nand U3562 (N_3562,In_457,In_2177);
xor U3563 (N_3563,In_960,In_2);
nand U3564 (N_3564,In_2096,In_850);
nand U3565 (N_3565,In_725,In_939);
nand U3566 (N_3566,In_1561,In_1410);
or U3567 (N_3567,In_1361,In_598);
nor U3568 (N_3568,In_2049,In_1857);
nor U3569 (N_3569,In_2257,In_1670);
nand U3570 (N_3570,In_1171,In_2493);
xnor U3571 (N_3571,In_2086,In_2035);
nor U3572 (N_3572,In_150,In_1317);
nand U3573 (N_3573,In_1144,In_1528);
or U3574 (N_3574,In_1404,In_1861);
or U3575 (N_3575,In_2235,In_1670);
nor U3576 (N_3576,In_2341,In_656);
nor U3577 (N_3577,In_1326,In_2011);
nand U3578 (N_3578,In_1206,In_554);
nand U3579 (N_3579,In_987,In_1497);
xor U3580 (N_3580,In_1054,In_1426);
nand U3581 (N_3581,In_244,In_633);
and U3582 (N_3582,In_1773,In_248);
nand U3583 (N_3583,In_984,In_1060);
nor U3584 (N_3584,In_2156,In_1672);
or U3585 (N_3585,In_2407,In_2066);
xnor U3586 (N_3586,In_1787,In_2257);
or U3587 (N_3587,In_2023,In_951);
nor U3588 (N_3588,In_1521,In_148);
and U3589 (N_3589,In_1087,In_1579);
or U3590 (N_3590,In_738,In_505);
and U3591 (N_3591,In_2429,In_630);
or U3592 (N_3592,In_1669,In_1581);
or U3593 (N_3593,In_775,In_273);
or U3594 (N_3594,In_1150,In_729);
xnor U3595 (N_3595,In_2144,In_1415);
nand U3596 (N_3596,In_1229,In_1305);
or U3597 (N_3597,In_396,In_1073);
or U3598 (N_3598,In_2379,In_390);
nor U3599 (N_3599,In_1538,In_1794);
or U3600 (N_3600,In_1473,In_412);
or U3601 (N_3601,In_1202,In_1848);
nand U3602 (N_3602,In_2104,In_774);
and U3603 (N_3603,In_1763,In_327);
or U3604 (N_3604,In_1183,In_732);
or U3605 (N_3605,In_80,In_1496);
nand U3606 (N_3606,In_2355,In_1901);
nand U3607 (N_3607,In_2279,In_1418);
xor U3608 (N_3608,In_117,In_483);
nor U3609 (N_3609,In_1495,In_99);
nand U3610 (N_3610,In_702,In_6);
nor U3611 (N_3611,In_50,In_1463);
nor U3612 (N_3612,In_162,In_408);
xnor U3613 (N_3613,In_2479,In_2035);
xnor U3614 (N_3614,In_1084,In_320);
nor U3615 (N_3615,In_775,In_605);
or U3616 (N_3616,In_66,In_311);
or U3617 (N_3617,In_1499,In_663);
xor U3618 (N_3618,In_1562,In_1684);
xnor U3619 (N_3619,In_277,In_2036);
nor U3620 (N_3620,In_2184,In_1838);
or U3621 (N_3621,In_2157,In_2199);
nor U3622 (N_3622,In_2403,In_1855);
nand U3623 (N_3623,In_2150,In_1969);
and U3624 (N_3624,In_2230,In_1493);
or U3625 (N_3625,In_2465,In_1756);
nand U3626 (N_3626,In_2094,In_1068);
nor U3627 (N_3627,In_319,In_1847);
nor U3628 (N_3628,In_2252,In_312);
nor U3629 (N_3629,In_2225,In_804);
nand U3630 (N_3630,In_875,In_1178);
nor U3631 (N_3631,In_1495,In_702);
nand U3632 (N_3632,In_491,In_1908);
nand U3633 (N_3633,In_2275,In_1113);
nor U3634 (N_3634,In_853,In_315);
nand U3635 (N_3635,In_2311,In_1648);
nand U3636 (N_3636,In_1850,In_397);
or U3637 (N_3637,In_1946,In_1885);
and U3638 (N_3638,In_1750,In_1620);
nand U3639 (N_3639,In_166,In_2468);
nor U3640 (N_3640,In_435,In_1223);
and U3641 (N_3641,In_1416,In_2023);
or U3642 (N_3642,In_1767,In_1622);
nand U3643 (N_3643,In_1158,In_1681);
nor U3644 (N_3644,In_1,In_1537);
nor U3645 (N_3645,In_2347,In_1515);
or U3646 (N_3646,In_69,In_1425);
nand U3647 (N_3647,In_932,In_664);
and U3648 (N_3648,In_1717,In_1466);
or U3649 (N_3649,In_527,In_2061);
nand U3650 (N_3650,In_855,In_1487);
and U3651 (N_3651,In_1888,In_2413);
nand U3652 (N_3652,In_15,In_83);
nand U3653 (N_3653,In_411,In_2001);
and U3654 (N_3654,In_2099,In_1330);
and U3655 (N_3655,In_1910,In_74);
nand U3656 (N_3656,In_1263,In_518);
nor U3657 (N_3657,In_1262,In_718);
nand U3658 (N_3658,In_2328,In_555);
xnor U3659 (N_3659,In_1156,In_1552);
nor U3660 (N_3660,In_1474,In_2466);
xnor U3661 (N_3661,In_2345,In_468);
or U3662 (N_3662,In_1311,In_2442);
nor U3663 (N_3663,In_523,In_1674);
nand U3664 (N_3664,In_925,In_2260);
or U3665 (N_3665,In_1447,In_1893);
nor U3666 (N_3666,In_1290,In_817);
nand U3667 (N_3667,In_1033,In_857);
and U3668 (N_3668,In_1846,In_1968);
or U3669 (N_3669,In_1151,In_817);
or U3670 (N_3670,In_1585,In_167);
and U3671 (N_3671,In_2394,In_2010);
nor U3672 (N_3672,In_495,In_2446);
and U3673 (N_3673,In_2389,In_1729);
and U3674 (N_3674,In_401,In_120);
xor U3675 (N_3675,In_828,In_959);
nor U3676 (N_3676,In_349,In_1296);
nand U3677 (N_3677,In_2103,In_1822);
nor U3678 (N_3678,In_1898,In_1741);
nor U3679 (N_3679,In_945,In_1259);
and U3680 (N_3680,In_2330,In_1302);
nand U3681 (N_3681,In_271,In_1140);
and U3682 (N_3682,In_371,In_366);
and U3683 (N_3683,In_1348,In_884);
nor U3684 (N_3684,In_1251,In_842);
nand U3685 (N_3685,In_806,In_1404);
nor U3686 (N_3686,In_1677,In_422);
or U3687 (N_3687,In_121,In_2065);
and U3688 (N_3688,In_833,In_2085);
and U3689 (N_3689,In_681,In_2370);
nand U3690 (N_3690,In_2499,In_1825);
and U3691 (N_3691,In_134,In_781);
or U3692 (N_3692,In_434,In_1818);
nand U3693 (N_3693,In_1386,In_2167);
nor U3694 (N_3694,In_420,In_404);
xor U3695 (N_3695,In_905,In_1238);
nand U3696 (N_3696,In_1719,In_492);
or U3697 (N_3697,In_341,In_1007);
nand U3698 (N_3698,In_105,In_1727);
nor U3699 (N_3699,In_335,In_466);
or U3700 (N_3700,In_1128,In_2174);
or U3701 (N_3701,In_2121,In_2291);
nor U3702 (N_3702,In_1245,In_411);
and U3703 (N_3703,In_1306,In_154);
xor U3704 (N_3704,In_2311,In_1915);
and U3705 (N_3705,In_1340,In_1014);
nor U3706 (N_3706,In_1798,In_246);
or U3707 (N_3707,In_257,In_696);
nand U3708 (N_3708,In_821,In_928);
and U3709 (N_3709,In_582,In_1854);
nor U3710 (N_3710,In_2189,In_1717);
nor U3711 (N_3711,In_1984,In_396);
nor U3712 (N_3712,In_1053,In_1227);
and U3713 (N_3713,In_1652,In_2046);
and U3714 (N_3714,In_352,In_1066);
or U3715 (N_3715,In_2178,In_706);
nand U3716 (N_3716,In_1395,In_2139);
nor U3717 (N_3717,In_107,In_807);
or U3718 (N_3718,In_251,In_1256);
nand U3719 (N_3719,In_1201,In_2291);
and U3720 (N_3720,In_226,In_300);
and U3721 (N_3721,In_1397,In_717);
nor U3722 (N_3722,In_1374,In_1713);
xnor U3723 (N_3723,In_716,In_1968);
and U3724 (N_3724,In_729,In_1466);
xor U3725 (N_3725,In_880,In_1177);
xnor U3726 (N_3726,In_559,In_1653);
nor U3727 (N_3727,In_106,In_2018);
and U3728 (N_3728,In_1421,In_1493);
nand U3729 (N_3729,In_847,In_2203);
and U3730 (N_3730,In_1027,In_1092);
or U3731 (N_3731,In_943,In_1671);
nand U3732 (N_3732,In_1613,In_2263);
nor U3733 (N_3733,In_805,In_638);
and U3734 (N_3734,In_2261,In_2003);
nor U3735 (N_3735,In_1773,In_938);
or U3736 (N_3736,In_1611,In_1391);
or U3737 (N_3737,In_620,In_348);
or U3738 (N_3738,In_1838,In_1883);
nor U3739 (N_3739,In_2408,In_823);
nand U3740 (N_3740,In_2112,In_2097);
nand U3741 (N_3741,In_1257,In_1759);
or U3742 (N_3742,In_2284,In_2201);
and U3743 (N_3743,In_1042,In_1322);
nand U3744 (N_3744,In_1299,In_344);
xnor U3745 (N_3745,In_903,In_424);
nand U3746 (N_3746,In_1417,In_2086);
nand U3747 (N_3747,In_1206,In_2303);
or U3748 (N_3748,In_775,In_2309);
or U3749 (N_3749,In_1540,In_582);
and U3750 (N_3750,In_1947,In_34);
or U3751 (N_3751,In_345,In_1497);
nand U3752 (N_3752,In_1543,In_1150);
nand U3753 (N_3753,In_2008,In_1518);
or U3754 (N_3754,In_405,In_1112);
and U3755 (N_3755,In_834,In_2091);
and U3756 (N_3756,In_1251,In_805);
or U3757 (N_3757,In_1759,In_217);
nor U3758 (N_3758,In_1344,In_1468);
or U3759 (N_3759,In_441,In_968);
or U3760 (N_3760,In_26,In_3);
nand U3761 (N_3761,In_345,In_979);
nand U3762 (N_3762,In_841,In_148);
and U3763 (N_3763,In_1316,In_112);
nand U3764 (N_3764,In_1174,In_461);
xor U3765 (N_3765,In_480,In_2042);
or U3766 (N_3766,In_2276,In_962);
or U3767 (N_3767,In_1065,In_677);
nor U3768 (N_3768,In_2135,In_1192);
nor U3769 (N_3769,In_778,In_1448);
or U3770 (N_3770,In_1891,In_1961);
or U3771 (N_3771,In_2355,In_1597);
or U3772 (N_3772,In_2171,In_1584);
or U3773 (N_3773,In_1366,In_377);
and U3774 (N_3774,In_754,In_1095);
nand U3775 (N_3775,In_691,In_1693);
or U3776 (N_3776,In_121,In_1021);
nand U3777 (N_3777,In_1119,In_580);
nand U3778 (N_3778,In_150,In_229);
or U3779 (N_3779,In_1833,In_2383);
nor U3780 (N_3780,In_835,In_1044);
xnor U3781 (N_3781,In_746,In_250);
xor U3782 (N_3782,In_953,In_72);
nor U3783 (N_3783,In_1451,In_2276);
nand U3784 (N_3784,In_2190,In_784);
and U3785 (N_3785,In_1788,In_896);
or U3786 (N_3786,In_640,In_1071);
nor U3787 (N_3787,In_292,In_1904);
nor U3788 (N_3788,In_697,In_2195);
nand U3789 (N_3789,In_2012,In_1858);
nand U3790 (N_3790,In_1843,In_249);
nor U3791 (N_3791,In_1548,In_148);
and U3792 (N_3792,In_919,In_2214);
nor U3793 (N_3793,In_2249,In_1226);
nor U3794 (N_3794,In_1121,In_488);
or U3795 (N_3795,In_840,In_2496);
or U3796 (N_3796,In_891,In_188);
nor U3797 (N_3797,In_2467,In_633);
or U3798 (N_3798,In_1602,In_1845);
nand U3799 (N_3799,In_1782,In_201);
nand U3800 (N_3800,In_1541,In_906);
xnor U3801 (N_3801,In_1697,In_9);
xnor U3802 (N_3802,In_1252,In_2193);
or U3803 (N_3803,In_1711,In_1841);
nand U3804 (N_3804,In_951,In_1420);
and U3805 (N_3805,In_1174,In_1255);
or U3806 (N_3806,In_2345,In_774);
and U3807 (N_3807,In_1020,In_1136);
and U3808 (N_3808,In_383,In_302);
or U3809 (N_3809,In_2130,In_2182);
nand U3810 (N_3810,In_1861,In_665);
nand U3811 (N_3811,In_1477,In_1760);
nor U3812 (N_3812,In_357,In_1185);
and U3813 (N_3813,In_1761,In_1793);
and U3814 (N_3814,In_110,In_2183);
or U3815 (N_3815,In_1348,In_2328);
xnor U3816 (N_3816,In_1944,In_498);
nand U3817 (N_3817,In_1172,In_356);
xnor U3818 (N_3818,In_604,In_929);
and U3819 (N_3819,In_1330,In_1871);
nand U3820 (N_3820,In_1544,In_1865);
nor U3821 (N_3821,In_2316,In_350);
nand U3822 (N_3822,In_640,In_1623);
nand U3823 (N_3823,In_623,In_1093);
nand U3824 (N_3824,In_1929,In_434);
and U3825 (N_3825,In_841,In_1088);
xor U3826 (N_3826,In_1205,In_2117);
nor U3827 (N_3827,In_307,In_833);
nand U3828 (N_3828,In_782,In_892);
or U3829 (N_3829,In_913,In_50);
and U3830 (N_3830,In_710,In_1087);
xor U3831 (N_3831,In_343,In_845);
or U3832 (N_3832,In_1806,In_725);
or U3833 (N_3833,In_1491,In_1505);
or U3834 (N_3834,In_1947,In_507);
xnor U3835 (N_3835,In_1624,In_1259);
and U3836 (N_3836,In_1985,In_1822);
nor U3837 (N_3837,In_935,In_997);
xor U3838 (N_3838,In_1276,In_435);
nand U3839 (N_3839,In_851,In_2401);
or U3840 (N_3840,In_1857,In_1234);
nor U3841 (N_3841,In_1396,In_488);
nor U3842 (N_3842,In_1547,In_1484);
xor U3843 (N_3843,In_78,In_596);
or U3844 (N_3844,In_2292,In_639);
nand U3845 (N_3845,In_1455,In_2256);
or U3846 (N_3846,In_2454,In_1125);
xor U3847 (N_3847,In_384,In_254);
and U3848 (N_3848,In_178,In_842);
and U3849 (N_3849,In_2108,In_2220);
nand U3850 (N_3850,In_1659,In_1954);
nand U3851 (N_3851,In_696,In_31);
and U3852 (N_3852,In_1562,In_1372);
nor U3853 (N_3853,In_1108,In_1203);
nand U3854 (N_3854,In_1732,In_1642);
nand U3855 (N_3855,In_399,In_201);
nand U3856 (N_3856,In_1636,In_1767);
or U3857 (N_3857,In_2459,In_301);
nand U3858 (N_3858,In_1048,In_574);
or U3859 (N_3859,In_2382,In_569);
or U3860 (N_3860,In_141,In_217);
nor U3861 (N_3861,In_2406,In_594);
and U3862 (N_3862,In_219,In_1867);
nor U3863 (N_3863,In_1036,In_1730);
and U3864 (N_3864,In_904,In_572);
or U3865 (N_3865,In_1033,In_1836);
nand U3866 (N_3866,In_938,In_2441);
nand U3867 (N_3867,In_357,In_923);
or U3868 (N_3868,In_1419,In_1701);
nor U3869 (N_3869,In_2111,In_1723);
nand U3870 (N_3870,In_1167,In_1807);
and U3871 (N_3871,In_338,In_2220);
nand U3872 (N_3872,In_2252,In_664);
nand U3873 (N_3873,In_2014,In_329);
nand U3874 (N_3874,In_19,In_2174);
nand U3875 (N_3875,In_1570,In_1646);
xor U3876 (N_3876,In_1824,In_597);
xor U3877 (N_3877,In_2117,In_2204);
xnor U3878 (N_3878,In_904,In_181);
nand U3879 (N_3879,In_1488,In_40);
nand U3880 (N_3880,In_2281,In_129);
nor U3881 (N_3881,In_501,In_517);
xor U3882 (N_3882,In_2374,In_555);
nand U3883 (N_3883,In_1491,In_60);
nand U3884 (N_3884,In_1414,In_2250);
nor U3885 (N_3885,In_450,In_588);
nand U3886 (N_3886,In_2071,In_404);
nand U3887 (N_3887,In_1144,In_2496);
nand U3888 (N_3888,In_1461,In_1894);
or U3889 (N_3889,In_887,In_2145);
and U3890 (N_3890,In_1725,In_1378);
and U3891 (N_3891,In_2071,In_1109);
or U3892 (N_3892,In_1244,In_1024);
nand U3893 (N_3893,In_2344,In_2311);
or U3894 (N_3894,In_1214,In_615);
xnor U3895 (N_3895,In_2027,In_2430);
nand U3896 (N_3896,In_482,In_1507);
nand U3897 (N_3897,In_1153,In_982);
nand U3898 (N_3898,In_315,In_585);
nand U3899 (N_3899,In_1671,In_2007);
or U3900 (N_3900,In_596,In_2203);
nand U3901 (N_3901,In_808,In_2357);
nand U3902 (N_3902,In_1016,In_1987);
nand U3903 (N_3903,In_1936,In_1791);
xnor U3904 (N_3904,In_536,In_795);
nor U3905 (N_3905,In_1302,In_730);
nand U3906 (N_3906,In_169,In_790);
nor U3907 (N_3907,In_1937,In_646);
and U3908 (N_3908,In_641,In_271);
and U3909 (N_3909,In_447,In_130);
xnor U3910 (N_3910,In_2086,In_496);
nor U3911 (N_3911,In_1204,In_1342);
nor U3912 (N_3912,In_1284,In_1405);
or U3913 (N_3913,In_1194,In_1486);
or U3914 (N_3914,In_2163,In_2415);
and U3915 (N_3915,In_1320,In_1078);
nand U3916 (N_3916,In_1050,In_172);
and U3917 (N_3917,In_2209,In_1352);
or U3918 (N_3918,In_1788,In_2361);
xnor U3919 (N_3919,In_1594,In_651);
nor U3920 (N_3920,In_904,In_558);
or U3921 (N_3921,In_1837,In_528);
or U3922 (N_3922,In_2338,In_2255);
nand U3923 (N_3923,In_1763,In_117);
nor U3924 (N_3924,In_453,In_27);
nand U3925 (N_3925,In_1865,In_373);
and U3926 (N_3926,In_1118,In_1283);
nor U3927 (N_3927,In_1260,In_2424);
or U3928 (N_3928,In_370,In_1340);
nor U3929 (N_3929,In_925,In_1091);
nor U3930 (N_3930,In_2271,In_1844);
or U3931 (N_3931,In_818,In_709);
and U3932 (N_3932,In_2122,In_1479);
or U3933 (N_3933,In_606,In_177);
and U3934 (N_3934,In_2019,In_173);
nand U3935 (N_3935,In_115,In_657);
or U3936 (N_3936,In_1179,In_2328);
and U3937 (N_3937,In_1100,In_2376);
or U3938 (N_3938,In_104,In_222);
nand U3939 (N_3939,In_1211,In_1865);
nand U3940 (N_3940,In_931,In_2249);
and U3941 (N_3941,In_2310,In_628);
and U3942 (N_3942,In_1920,In_2437);
nor U3943 (N_3943,In_1579,In_764);
and U3944 (N_3944,In_1964,In_1090);
nor U3945 (N_3945,In_1192,In_2461);
nor U3946 (N_3946,In_1132,In_557);
or U3947 (N_3947,In_1863,In_1739);
and U3948 (N_3948,In_1865,In_1149);
xnor U3949 (N_3949,In_780,In_173);
nor U3950 (N_3950,In_754,In_1223);
nor U3951 (N_3951,In_701,In_685);
and U3952 (N_3952,In_895,In_392);
or U3953 (N_3953,In_1950,In_1631);
nand U3954 (N_3954,In_222,In_1876);
or U3955 (N_3955,In_1975,In_1897);
or U3956 (N_3956,In_384,In_853);
or U3957 (N_3957,In_1957,In_1684);
nor U3958 (N_3958,In_2111,In_1766);
or U3959 (N_3959,In_1279,In_2392);
and U3960 (N_3960,In_2463,In_856);
and U3961 (N_3961,In_1720,In_98);
and U3962 (N_3962,In_1879,In_1058);
or U3963 (N_3963,In_139,In_983);
nor U3964 (N_3964,In_187,In_890);
and U3965 (N_3965,In_2187,In_349);
and U3966 (N_3966,In_694,In_1960);
or U3967 (N_3967,In_103,In_957);
nand U3968 (N_3968,In_911,In_617);
nor U3969 (N_3969,In_905,In_765);
nand U3970 (N_3970,In_1930,In_940);
nor U3971 (N_3971,In_1749,In_2064);
nor U3972 (N_3972,In_1360,In_1386);
and U3973 (N_3973,In_2384,In_2300);
and U3974 (N_3974,In_2396,In_258);
nor U3975 (N_3975,In_1755,In_2488);
nor U3976 (N_3976,In_1547,In_772);
and U3977 (N_3977,In_945,In_1067);
or U3978 (N_3978,In_367,In_323);
or U3979 (N_3979,In_1438,In_1275);
and U3980 (N_3980,In_1513,In_32);
nor U3981 (N_3981,In_121,In_2000);
nor U3982 (N_3982,In_819,In_2432);
and U3983 (N_3983,In_1199,In_711);
and U3984 (N_3984,In_556,In_1083);
and U3985 (N_3985,In_1627,In_2205);
and U3986 (N_3986,In_400,In_1797);
nand U3987 (N_3987,In_1620,In_1932);
and U3988 (N_3988,In_1638,In_2330);
xnor U3989 (N_3989,In_1132,In_154);
nor U3990 (N_3990,In_2436,In_508);
nor U3991 (N_3991,In_820,In_605);
or U3992 (N_3992,In_274,In_2158);
nand U3993 (N_3993,In_1842,In_1369);
or U3994 (N_3994,In_109,In_1761);
and U3995 (N_3995,In_264,In_1448);
or U3996 (N_3996,In_1293,In_762);
and U3997 (N_3997,In_737,In_7);
or U3998 (N_3998,In_1526,In_917);
xor U3999 (N_3999,In_1098,In_957);
nand U4000 (N_4000,In_1942,In_1462);
xnor U4001 (N_4001,In_2087,In_1833);
nand U4002 (N_4002,In_2262,In_965);
and U4003 (N_4003,In_846,In_167);
or U4004 (N_4004,In_1527,In_2325);
nor U4005 (N_4005,In_152,In_2290);
nand U4006 (N_4006,In_1990,In_1212);
and U4007 (N_4007,In_1644,In_1496);
xor U4008 (N_4008,In_1506,In_1829);
or U4009 (N_4009,In_2029,In_162);
nor U4010 (N_4010,In_1971,In_258);
nor U4011 (N_4011,In_62,In_1208);
nand U4012 (N_4012,In_1150,In_1680);
xor U4013 (N_4013,In_2251,In_1379);
nor U4014 (N_4014,In_2006,In_1946);
nor U4015 (N_4015,In_240,In_1005);
nor U4016 (N_4016,In_421,In_610);
and U4017 (N_4017,In_340,In_315);
and U4018 (N_4018,In_1595,In_1179);
nor U4019 (N_4019,In_463,In_2171);
nor U4020 (N_4020,In_1314,In_517);
or U4021 (N_4021,In_2344,In_2362);
and U4022 (N_4022,In_1371,In_1099);
xor U4023 (N_4023,In_1171,In_1248);
nand U4024 (N_4024,In_1100,In_2402);
nor U4025 (N_4025,In_2116,In_2084);
xor U4026 (N_4026,In_2255,In_1615);
nor U4027 (N_4027,In_1340,In_1386);
and U4028 (N_4028,In_501,In_1271);
or U4029 (N_4029,In_1451,In_754);
nor U4030 (N_4030,In_1084,In_635);
nand U4031 (N_4031,In_856,In_1719);
xnor U4032 (N_4032,In_344,In_325);
xnor U4033 (N_4033,In_564,In_1981);
or U4034 (N_4034,In_1944,In_2409);
or U4035 (N_4035,In_683,In_93);
nand U4036 (N_4036,In_1389,In_358);
and U4037 (N_4037,In_1078,In_2230);
or U4038 (N_4038,In_16,In_933);
and U4039 (N_4039,In_1510,In_2412);
nor U4040 (N_4040,In_2285,In_1103);
nand U4041 (N_4041,In_2138,In_2130);
or U4042 (N_4042,In_2176,In_507);
and U4043 (N_4043,In_1314,In_2034);
or U4044 (N_4044,In_2439,In_24);
nor U4045 (N_4045,In_1017,In_2057);
and U4046 (N_4046,In_220,In_2439);
xnor U4047 (N_4047,In_358,In_841);
and U4048 (N_4048,In_24,In_657);
and U4049 (N_4049,In_2254,In_2352);
nand U4050 (N_4050,In_589,In_2107);
or U4051 (N_4051,In_1419,In_2441);
and U4052 (N_4052,In_181,In_2366);
nand U4053 (N_4053,In_1888,In_1622);
nand U4054 (N_4054,In_6,In_281);
nand U4055 (N_4055,In_529,In_2071);
and U4056 (N_4056,In_1204,In_273);
nor U4057 (N_4057,In_1582,In_1569);
xnor U4058 (N_4058,In_667,In_841);
nand U4059 (N_4059,In_1421,In_1964);
nand U4060 (N_4060,In_1025,In_1033);
or U4061 (N_4061,In_1598,In_2456);
and U4062 (N_4062,In_1222,In_680);
or U4063 (N_4063,In_757,In_1597);
or U4064 (N_4064,In_320,In_2236);
or U4065 (N_4065,In_1131,In_1049);
xnor U4066 (N_4066,In_831,In_516);
xnor U4067 (N_4067,In_817,In_1302);
or U4068 (N_4068,In_868,In_2228);
nand U4069 (N_4069,In_34,In_2469);
xor U4070 (N_4070,In_1310,In_30);
nand U4071 (N_4071,In_17,In_1604);
and U4072 (N_4072,In_1166,In_1114);
nor U4073 (N_4073,In_2007,In_2410);
and U4074 (N_4074,In_741,In_1809);
nand U4075 (N_4075,In_420,In_2152);
or U4076 (N_4076,In_1385,In_726);
and U4077 (N_4077,In_2491,In_433);
nor U4078 (N_4078,In_1918,In_2096);
or U4079 (N_4079,In_1572,In_1293);
and U4080 (N_4080,In_1656,In_1686);
nor U4081 (N_4081,In_44,In_2046);
nand U4082 (N_4082,In_1563,In_1236);
or U4083 (N_4083,In_2047,In_1570);
nor U4084 (N_4084,In_1068,In_2374);
and U4085 (N_4085,In_1570,In_2455);
and U4086 (N_4086,In_1880,In_589);
and U4087 (N_4087,In_2128,In_1045);
or U4088 (N_4088,In_1853,In_422);
xor U4089 (N_4089,In_661,In_913);
and U4090 (N_4090,In_85,In_1958);
or U4091 (N_4091,In_2100,In_813);
and U4092 (N_4092,In_2321,In_133);
or U4093 (N_4093,In_1959,In_1533);
and U4094 (N_4094,In_1579,In_1920);
nor U4095 (N_4095,In_621,In_3);
and U4096 (N_4096,In_1201,In_194);
or U4097 (N_4097,In_1663,In_2341);
nor U4098 (N_4098,In_2375,In_554);
or U4099 (N_4099,In_1523,In_1742);
nand U4100 (N_4100,In_2402,In_343);
or U4101 (N_4101,In_1035,In_1190);
or U4102 (N_4102,In_1475,In_1927);
nand U4103 (N_4103,In_1721,In_1585);
nand U4104 (N_4104,In_472,In_2225);
nor U4105 (N_4105,In_11,In_1743);
nor U4106 (N_4106,In_1187,In_1575);
nand U4107 (N_4107,In_1112,In_2163);
nand U4108 (N_4108,In_609,In_2042);
or U4109 (N_4109,In_2082,In_1563);
or U4110 (N_4110,In_134,In_425);
nand U4111 (N_4111,In_1104,In_2019);
and U4112 (N_4112,In_590,In_104);
nor U4113 (N_4113,In_636,In_655);
nor U4114 (N_4114,In_374,In_1593);
or U4115 (N_4115,In_1844,In_1561);
nor U4116 (N_4116,In_565,In_1481);
nand U4117 (N_4117,In_1025,In_1507);
and U4118 (N_4118,In_2082,In_2104);
nand U4119 (N_4119,In_1253,In_996);
and U4120 (N_4120,In_1665,In_1754);
nand U4121 (N_4121,In_1989,In_2146);
and U4122 (N_4122,In_1532,In_2226);
or U4123 (N_4123,In_1803,In_703);
and U4124 (N_4124,In_2254,In_177);
nand U4125 (N_4125,In_157,In_1465);
nor U4126 (N_4126,In_2022,In_1731);
nand U4127 (N_4127,In_261,In_282);
nand U4128 (N_4128,In_855,In_2411);
and U4129 (N_4129,In_505,In_1458);
or U4130 (N_4130,In_1651,In_1913);
nand U4131 (N_4131,In_2019,In_1532);
and U4132 (N_4132,In_1788,In_1493);
nor U4133 (N_4133,In_179,In_1965);
or U4134 (N_4134,In_1177,In_1452);
nor U4135 (N_4135,In_489,In_2291);
or U4136 (N_4136,In_1122,In_803);
and U4137 (N_4137,In_705,In_1515);
nor U4138 (N_4138,In_2180,In_2206);
nor U4139 (N_4139,In_1255,In_1497);
xor U4140 (N_4140,In_370,In_1202);
or U4141 (N_4141,In_2164,In_1597);
or U4142 (N_4142,In_2200,In_795);
nor U4143 (N_4143,In_1880,In_632);
nor U4144 (N_4144,In_907,In_1936);
or U4145 (N_4145,In_698,In_1703);
xor U4146 (N_4146,In_1315,In_665);
nand U4147 (N_4147,In_116,In_1966);
and U4148 (N_4148,In_1477,In_1673);
nand U4149 (N_4149,In_2198,In_2489);
nand U4150 (N_4150,In_1663,In_1912);
and U4151 (N_4151,In_1916,In_298);
nor U4152 (N_4152,In_44,In_1352);
and U4153 (N_4153,In_32,In_2028);
or U4154 (N_4154,In_1536,In_1339);
or U4155 (N_4155,In_2428,In_1132);
and U4156 (N_4156,In_393,In_87);
or U4157 (N_4157,In_592,In_1812);
and U4158 (N_4158,In_482,In_1210);
nand U4159 (N_4159,In_2087,In_960);
or U4160 (N_4160,In_1135,In_191);
and U4161 (N_4161,In_2046,In_208);
nand U4162 (N_4162,In_2087,In_2290);
and U4163 (N_4163,In_22,In_1687);
nor U4164 (N_4164,In_699,In_2384);
nor U4165 (N_4165,In_2478,In_1435);
nor U4166 (N_4166,In_1881,In_2012);
nand U4167 (N_4167,In_1859,In_1145);
and U4168 (N_4168,In_1393,In_1757);
and U4169 (N_4169,In_337,In_1167);
or U4170 (N_4170,In_762,In_94);
or U4171 (N_4171,In_1942,In_802);
or U4172 (N_4172,In_1322,In_462);
nor U4173 (N_4173,In_1496,In_1457);
or U4174 (N_4174,In_1883,In_424);
nor U4175 (N_4175,In_1325,In_800);
or U4176 (N_4176,In_1356,In_939);
nor U4177 (N_4177,In_1926,In_1843);
nand U4178 (N_4178,In_1641,In_2142);
nand U4179 (N_4179,In_261,In_1229);
nor U4180 (N_4180,In_986,In_2317);
nor U4181 (N_4181,In_2369,In_2214);
nor U4182 (N_4182,In_1460,In_2125);
nand U4183 (N_4183,In_2041,In_154);
nand U4184 (N_4184,In_1832,In_676);
nand U4185 (N_4185,In_1065,In_2094);
nor U4186 (N_4186,In_396,In_890);
or U4187 (N_4187,In_540,In_371);
nor U4188 (N_4188,In_959,In_503);
nand U4189 (N_4189,In_476,In_93);
nand U4190 (N_4190,In_1689,In_890);
nor U4191 (N_4191,In_1469,In_1717);
xor U4192 (N_4192,In_1106,In_1100);
or U4193 (N_4193,In_288,In_725);
nor U4194 (N_4194,In_114,In_1057);
nand U4195 (N_4195,In_2197,In_216);
xnor U4196 (N_4196,In_941,In_1844);
nor U4197 (N_4197,In_2420,In_1166);
and U4198 (N_4198,In_2001,In_2436);
and U4199 (N_4199,In_905,In_1347);
nand U4200 (N_4200,In_50,In_583);
nand U4201 (N_4201,In_476,In_227);
nor U4202 (N_4202,In_2405,In_2407);
and U4203 (N_4203,In_2358,In_504);
nand U4204 (N_4204,In_567,In_2306);
xor U4205 (N_4205,In_1677,In_1078);
nand U4206 (N_4206,In_920,In_598);
or U4207 (N_4207,In_2241,In_64);
and U4208 (N_4208,In_713,In_1989);
nand U4209 (N_4209,In_2271,In_403);
and U4210 (N_4210,In_1484,In_1511);
nand U4211 (N_4211,In_1972,In_535);
nor U4212 (N_4212,In_157,In_1281);
nor U4213 (N_4213,In_520,In_0);
nand U4214 (N_4214,In_279,In_797);
xnor U4215 (N_4215,In_1023,In_1186);
and U4216 (N_4216,In_1027,In_2216);
nand U4217 (N_4217,In_670,In_1259);
and U4218 (N_4218,In_1403,In_1450);
and U4219 (N_4219,In_1902,In_762);
nand U4220 (N_4220,In_2308,In_2270);
nor U4221 (N_4221,In_994,In_2009);
nand U4222 (N_4222,In_428,In_579);
nor U4223 (N_4223,In_847,In_1908);
nor U4224 (N_4224,In_1460,In_1951);
or U4225 (N_4225,In_288,In_1054);
xnor U4226 (N_4226,In_1773,In_536);
nand U4227 (N_4227,In_1038,In_1031);
or U4228 (N_4228,In_332,In_1762);
nor U4229 (N_4229,In_64,In_509);
or U4230 (N_4230,In_167,In_1018);
and U4231 (N_4231,In_746,In_171);
or U4232 (N_4232,In_1436,In_2252);
or U4233 (N_4233,In_1019,In_595);
nand U4234 (N_4234,In_735,In_1825);
nand U4235 (N_4235,In_2004,In_391);
nor U4236 (N_4236,In_358,In_2211);
or U4237 (N_4237,In_1700,In_56);
nand U4238 (N_4238,In_740,In_2223);
nor U4239 (N_4239,In_1561,In_666);
nor U4240 (N_4240,In_2112,In_580);
nand U4241 (N_4241,In_2152,In_1875);
and U4242 (N_4242,In_2119,In_1230);
nand U4243 (N_4243,In_2260,In_402);
nor U4244 (N_4244,In_744,In_400);
or U4245 (N_4245,In_1268,In_426);
nor U4246 (N_4246,In_1074,In_705);
nor U4247 (N_4247,In_347,In_1140);
nor U4248 (N_4248,In_1428,In_2268);
nand U4249 (N_4249,In_1168,In_1612);
and U4250 (N_4250,In_2125,In_2126);
or U4251 (N_4251,In_1344,In_318);
nand U4252 (N_4252,In_918,In_1313);
nand U4253 (N_4253,In_1830,In_1751);
and U4254 (N_4254,In_682,In_2054);
and U4255 (N_4255,In_1954,In_370);
or U4256 (N_4256,In_803,In_2367);
xnor U4257 (N_4257,In_2244,In_1669);
or U4258 (N_4258,In_101,In_783);
nand U4259 (N_4259,In_1273,In_1103);
and U4260 (N_4260,In_1500,In_2208);
nor U4261 (N_4261,In_952,In_2005);
and U4262 (N_4262,In_617,In_366);
and U4263 (N_4263,In_594,In_1964);
nor U4264 (N_4264,In_445,In_2238);
and U4265 (N_4265,In_495,In_1360);
nor U4266 (N_4266,In_1214,In_118);
or U4267 (N_4267,In_1540,In_363);
xnor U4268 (N_4268,In_1194,In_1803);
nor U4269 (N_4269,In_2171,In_94);
and U4270 (N_4270,In_2046,In_720);
nand U4271 (N_4271,In_1055,In_1477);
nor U4272 (N_4272,In_639,In_1723);
and U4273 (N_4273,In_1619,In_2267);
nand U4274 (N_4274,In_2180,In_465);
nand U4275 (N_4275,In_1164,In_1379);
or U4276 (N_4276,In_69,In_2024);
nand U4277 (N_4277,In_2127,In_952);
or U4278 (N_4278,In_788,In_796);
nor U4279 (N_4279,In_73,In_570);
and U4280 (N_4280,In_34,In_1443);
nand U4281 (N_4281,In_855,In_2069);
nand U4282 (N_4282,In_1216,In_1154);
nand U4283 (N_4283,In_1056,In_530);
nor U4284 (N_4284,In_1603,In_2367);
xnor U4285 (N_4285,In_83,In_815);
nor U4286 (N_4286,In_585,In_1288);
nand U4287 (N_4287,In_2340,In_1656);
nor U4288 (N_4288,In_1685,In_1267);
nand U4289 (N_4289,In_300,In_1235);
nor U4290 (N_4290,In_1813,In_240);
and U4291 (N_4291,In_200,In_1578);
and U4292 (N_4292,In_1080,In_1339);
and U4293 (N_4293,In_2087,In_1250);
nand U4294 (N_4294,In_2024,In_2345);
nor U4295 (N_4295,In_1557,In_1062);
nor U4296 (N_4296,In_131,In_695);
nor U4297 (N_4297,In_2104,In_973);
nor U4298 (N_4298,In_193,In_842);
nor U4299 (N_4299,In_1428,In_903);
or U4300 (N_4300,In_1956,In_723);
nand U4301 (N_4301,In_1153,In_1133);
or U4302 (N_4302,In_919,In_1745);
nand U4303 (N_4303,In_1500,In_1338);
and U4304 (N_4304,In_1627,In_822);
xor U4305 (N_4305,In_1805,In_647);
nand U4306 (N_4306,In_392,In_792);
xor U4307 (N_4307,In_49,In_1435);
and U4308 (N_4308,In_1356,In_812);
nor U4309 (N_4309,In_766,In_100);
nand U4310 (N_4310,In_1970,In_1703);
or U4311 (N_4311,In_407,In_2410);
and U4312 (N_4312,In_196,In_818);
nand U4313 (N_4313,In_322,In_2347);
nand U4314 (N_4314,In_2106,In_307);
or U4315 (N_4315,In_107,In_2131);
and U4316 (N_4316,In_2182,In_1828);
nand U4317 (N_4317,In_1487,In_1573);
nor U4318 (N_4318,In_1361,In_310);
xnor U4319 (N_4319,In_222,In_2424);
nand U4320 (N_4320,In_1631,In_414);
or U4321 (N_4321,In_235,In_139);
and U4322 (N_4322,In_1928,In_1605);
nand U4323 (N_4323,In_887,In_813);
nand U4324 (N_4324,In_298,In_1982);
nand U4325 (N_4325,In_332,In_439);
nor U4326 (N_4326,In_2379,In_1749);
or U4327 (N_4327,In_1928,In_513);
and U4328 (N_4328,In_1271,In_1964);
or U4329 (N_4329,In_653,In_1800);
nand U4330 (N_4330,In_939,In_392);
nor U4331 (N_4331,In_762,In_344);
and U4332 (N_4332,In_213,In_2225);
or U4333 (N_4333,In_2087,In_1185);
xor U4334 (N_4334,In_1365,In_223);
xnor U4335 (N_4335,In_2004,In_2282);
xnor U4336 (N_4336,In_1909,In_1969);
xnor U4337 (N_4337,In_1114,In_1137);
and U4338 (N_4338,In_762,In_748);
and U4339 (N_4339,In_1569,In_1665);
nor U4340 (N_4340,In_995,In_1886);
nand U4341 (N_4341,In_2250,In_1691);
nor U4342 (N_4342,In_61,In_463);
nor U4343 (N_4343,In_1079,In_618);
nand U4344 (N_4344,In_1805,In_625);
nand U4345 (N_4345,In_1587,In_1393);
nor U4346 (N_4346,In_167,In_943);
or U4347 (N_4347,In_181,In_180);
nor U4348 (N_4348,In_131,In_2018);
nand U4349 (N_4349,In_1825,In_1846);
nor U4350 (N_4350,In_1961,In_2492);
nor U4351 (N_4351,In_291,In_855);
nor U4352 (N_4352,In_981,In_534);
and U4353 (N_4353,In_1359,In_1938);
nor U4354 (N_4354,In_1303,In_733);
or U4355 (N_4355,In_1864,In_536);
nor U4356 (N_4356,In_2032,In_862);
xnor U4357 (N_4357,In_1811,In_817);
or U4358 (N_4358,In_24,In_1889);
nand U4359 (N_4359,In_503,In_1113);
or U4360 (N_4360,In_1308,In_1643);
nand U4361 (N_4361,In_542,In_2098);
and U4362 (N_4362,In_2321,In_1351);
or U4363 (N_4363,In_1703,In_303);
nor U4364 (N_4364,In_719,In_1279);
nor U4365 (N_4365,In_914,In_1881);
and U4366 (N_4366,In_2040,In_1107);
and U4367 (N_4367,In_1738,In_1991);
nor U4368 (N_4368,In_1984,In_2251);
nor U4369 (N_4369,In_1117,In_672);
nor U4370 (N_4370,In_709,In_2138);
and U4371 (N_4371,In_2344,In_1013);
nor U4372 (N_4372,In_1147,In_1938);
nand U4373 (N_4373,In_1185,In_2290);
nand U4374 (N_4374,In_1810,In_529);
or U4375 (N_4375,In_314,In_1030);
nor U4376 (N_4376,In_1023,In_581);
or U4377 (N_4377,In_1981,In_2470);
and U4378 (N_4378,In_2078,In_1692);
nand U4379 (N_4379,In_1396,In_1522);
and U4380 (N_4380,In_1128,In_2255);
nor U4381 (N_4381,In_544,In_697);
xor U4382 (N_4382,In_201,In_1232);
xnor U4383 (N_4383,In_297,In_1788);
nand U4384 (N_4384,In_626,In_2082);
nand U4385 (N_4385,In_869,In_1797);
and U4386 (N_4386,In_1535,In_1441);
or U4387 (N_4387,In_1260,In_1672);
and U4388 (N_4388,In_1400,In_500);
nor U4389 (N_4389,In_381,In_151);
and U4390 (N_4390,In_1322,In_2398);
or U4391 (N_4391,In_1794,In_275);
xnor U4392 (N_4392,In_799,In_1059);
nand U4393 (N_4393,In_938,In_275);
or U4394 (N_4394,In_937,In_1433);
and U4395 (N_4395,In_1970,In_745);
nor U4396 (N_4396,In_2482,In_1578);
and U4397 (N_4397,In_1988,In_2092);
and U4398 (N_4398,In_1678,In_2461);
nand U4399 (N_4399,In_2379,In_1253);
nand U4400 (N_4400,In_2047,In_952);
nand U4401 (N_4401,In_430,In_2304);
nor U4402 (N_4402,In_1291,In_2442);
nor U4403 (N_4403,In_527,In_812);
nand U4404 (N_4404,In_1408,In_241);
xnor U4405 (N_4405,In_1278,In_1525);
or U4406 (N_4406,In_1413,In_1031);
xor U4407 (N_4407,In_714,In_1127);
nor U4408 (N_4408,In_1379,In_101);
nand U4409 (N_4409,In_2461,In_1915);
and U4410 (N_4410,In_689,In_326);
and U4411 (N_4411,In_369,In_98);
xnor U4412 (N_4412,In_1354,In_1817);
nand U4413 (N_4413,In_430,In_1645);
nand U4414 (N_4414,In_1995,In_2026);
and U4415 (N_4415,In_2202,In_392);
nand U4416 (N_4416,In_1100,In_272);
or U4417 (N_4417,In_983,In_1631);
xnor U4418 (N_4418,In_2359,In_1093);
and U4419 (N_4419,In_471,In_1928);
or U4420 (N_4420,In_2294,In_50);
nor U4421 (N_4421,In_1564,In_512);
or U4422 (N_4422,In_2233,In_882);
or U4423 (N_4423,In_2265,In_2241);
nor U4424 (N_4424,In_2179,In_217);
nand U4425 (N_4425,In_422,In_1990);
nand U4426 (N_4426,In_902,In_2118);
nand U4427 (N_4427,In_902,In_1471);
nand U4428 (N_4428,In_2171,In_2353);
or U4429 (N_4429,In_23,In_2222);
and U4430 (N_4430,In_1752,In_18);
nor U4431 (N_4431,In_1154,In_1841);
or U4432 (N_4432,In_1933,In_2292);
nand U4433 (N_4433,In_590,In_316);
nor U4434 (N_4434,In_2186,In_723);
nor U4435 (N_4435,In_991,In_2369);
and U4436 (N_4436,In_659,In_2);
or U4437 (N_4437,In_1833,In_772);
nor U4438 (N_4438,In_1130,In_1432);
or U4439 (N_4439,In_1237,In_1514);
or U4440 (N_4440,In_1543,In_120);
nand U4441 (N_4441,In_324,In_1881);
nand U4442 (N_4442,In_1177,In_1219);
and U4443 (N_4443,In_2,In_1014);
nor U4444 (N_4444,In_1484,In_106);
or U4445 (N_4445,In_998,In_1839);
and U4446 (N_4446,In_1378,In_1044);
and U4447 (N_4447,In_2395,In_2233);
nor U4448 (N_4448,In_1963,In_291);
xor U4449 (N_4449,In_1997,In_744);
or U4450 (N_4450,In_1243,In_1202);
and U4451 (N_4451,In_1598,In_581);
xnor U4452 (N_4452,In_786,In_1157);
nand U4453 (N_4453,In_1360,In_2136);
or U4454 (N_4454,In_2039,In_687);
nand U4455 (N_4455,In_1599,In_11);
nor U4456 (N_4456,In_1655,In_2280);
or U4457 (N_4457,In_1047,In_327);
or U4458 (N_4458,In_691,In_2479);
nand U4459 (N_4459,In_2411,In_1180);
xor U4460 (N_4460,In_345,In_1897);
or U4461 (N_4461,In_535,In_1748);
or U4462 (N_4462,In_170,In_997);
and U4463 (N_4463,In_1314,In_59);
or U4464 (N_4464,In_1814,In_558);
nor U4465 (N_4465,In_1127,In_1553);
xor U4466 (N_4466,In_289,In_2048);
xor U4467 (N_4467,In_864,In_1842);
nand U4468 (N_4468,In_345,In_1381);
nor U4469 (N_4469,In_1191,In_1032);
or U4470 (N_4470,In_514,In_578);
or U4471 (N_4471,In_481,In_1250);
or U4472 (N_4472,In_171,In_2373);
or U4473 (N_4473,In_1915,In_1446);
nor U4474 (N_4474,In_1958,In_561);
and U4475 (N_4475,In_206,In_1290);
nand U4476 (N_4476,In_2304,In_813);
nor U4477 (N_4477,In_1767,In_1490);
or U4478 (N_4478,In_1781,In_1630);
nor U4479 (N_4479,In_2365,In_1323);
and U4480 (N_4480,In_1066,In_362);
or U4481 (N_4481,In_470,In_1727);
nor U4482 (N_4482,In_1626,In_1745);
nand U4483 (N_4483,In_383,In_485);
or U4484 (N_4484,In_1635,In_2255);
or U4485 (N_4485,In_1881,In_171);
nor U4486 (N_4486,In_751,In_1285);
and U4487 (N_4487,In_867,In_2237);
or U4488 (N_4488,In_2234,In_594);
nor U4489 (N_4489,In_979,In_1325);
nor U4490 (N_4490,In_2148,In_1085);
or U4491 (N_4491,In_944,In_1503);
or U4492 (N_4492,In_451,In_1281);
nor U4493 (N_4493,In_1091,In_1549);
or U4494 (N_4494,In_2075,In_483);
nand U4495 (N_4495,In_1253,In_2084);
nand U4496 (N_4496,In_1254,In_1175);
nor U4497 (N_4497,In_1503,In_1452);
or U4498 (N_4498,In_670,In_1582);
and U4499 (N_4499,In_1752,In_2408);
or U4500 (N_4500,In_2330,In_711);
nor U4501 (N_4501,In_491,In_1474);
and U4502 (N_4502,In_863,In_369);
or U4503 (N_4503,In_277,In_647);
nand U4504 (N_4504,In_249,In_370);
or U4505 (N_4505,In_711,In_2376);
nor U4506 (N_4506,In_1915,In_2134);
nand U4507 (N_4507,In_978,In_367);
and U4508 (N_4508,In_1909,In_1988);
nand U4509 (N_4509,In_176,In_606);
and U4510 (N_4510,In_2266,In_515);
or U4511 (N_4511,In_2073,In_313);
or U4512 (N_4512,In_1095,In_816);
and U4513 (N_4513,In_2055,In_296);
nor U4514 (N_4514,In_553,In_940);
and U4515 (N_4515,In_786,In_1355);
and U4516 (N_4516,In_285,In_1882);
or U4517 (N_4517,In_1530,In_1976);
xnor U4518 (N_4518,In_265,In_110);
nand U4519 (N_4519,In_1529,In_765);
or U4520 (N_4520,In_1904,In_365);
nor U4521 (N_4521,In_172,In_81);
or U4522 (N_4522,In_1367,In_2458);
nor U4523 (N_4523,In_955,In_1586);
and U4524 (N_4524,In_930,In_2398);
nor U4525 (N_4525,In_2096,In_1515);
nand U4526 (N_4526,In_218,In_1845);
and U4527 (N_4527,In_2011,In_1635);
xnor U4528 (N_4528,In_2236,In_235);
nand U4529 (N_4529,In_419,In_1572);
nand U4530 (N_4530,In_1581,In_286);
nor U4531 (N_4531,In_1924,In_381);
nand U4532 (N_4532,In_621,In_868);
and U4533 (N_4533,In_2177,In_1884);
nor U4534 (N_4534,In_165,In_546);
or U4535 (N_4535,In_382,In_606);
and U4536 (N_4536,In_1014,In_2384);
nor U4537 (N_4537,In_2328,In_1585);
or U4538 (N_4538,In_2423,In_1677);
or U4539 (N_4539,In_1407,In_2044);
and U4540 (N_4540,In_171,In_29);
nor U4541 (N_4541,In_1281,In_1974);
xnor U4542 (N_4542,In_795,In_1674);
or U4543 (N_4543,In_1032,In_511);
and U4544 (N_4544,In_695,In_2253);
xor U4545 (N_4545,In_2083,In_1145);
or U4546 (N_4546,In_60,In_1794);
nand U4547 (N_4547,In_789,In_1469);
and U4548 (N_4548,In_126,In_455);
and U4549 (N_4549,In_1527,In_1152);
or U4550 (N_4550,In_481,In_2265);
xor U4551 (N_4551,In_416,In_171);
nor U4552 (N_4552,In_987,In_978);
and U4553 (N_4553,In_755,In_766);
and U4554 (N_4554,In_198,In_481);
and U4555 (N_4555,In_807,In_1457);
nor U4556 (N_4556,In_2039,In_1952);
or U4557 (N_4557,In_1266,In_1770);
nand U4558 (N_4558,In_752,In_677);
nand U4559 (N_4559,In_2174,In_1757);
nand U4560 (N_4560,In_1263,In_1295);
nand U4561 (N_4561,In_240,In_696);
nor U4562 (N_4562,In_1854,In_597);
or U4563 (N_4563,In_1719,In_1204);
nand U4564 (N_4564,In_1936,In_85);
nor U4565 (N_4565,In_1826,In_750);
and U4566 (N_4566,In_68,In_789);
or U4567 (N_4567,In_1186,In_1036);
nor U4568 (N_4568,In_1258,In_169);
nand U4569 (N_4569,In_1694,In_873);
and U4570 (N_4570,In_1002,In_454);
nand U4571 (N_4571,In_1824,In_562);
or U4572 (N_4572,In_1851,In_45);
nor U4573 (N_4573,In_1950,In_850);
nor U4574 (N_4574,In_577,In_1399);
nor U4575 (N_4575,In_2499,In_1131);
nor U4576 (N_4576,In_1612,In_406);
and U4577 (N_4577,In_1036,In_320);
and U4578 (N_4578,In_469,In_235);
xnor U4579 (N_4579,In_315,In_2382);
nor U4580 (N_4580,In_1707,In_1039);
nand U4581 (N_4581,In_721,In_1432);
or U4582 (N_4582,In_395,In_593);
nand U4583 (N_4583,In_1296,In_2182);
nor U4584 (N_4584,In_689,In_924);
or U4585 (N_4585,In_1771,In_933);
nor U4586 (N_4586,In_659,In_1789);
nand U4587 (N_4587,In_1859,In_1705);
nor U4588 (N_4588,In_1389,In_589);
and U4589 (N_4589,In_107,In_1082);
nor U4590 (N_4590,In_1961,In_2258);
nor U4591 (N_4591,In_1405,In_2453);
or U4592 (N_4592,In_723,In_336);
or U4593 (N_4593,In_1320,In_1890);
nor U4594 (N_4594,In_2300,In_956);
or U4595 (N_4595,In_2477,In_2232);
or U4596 (N_4596,In_442,In_632);
xor U4597 (N_4597,In_655,In_2438);
nand U4598 (N_4598,In_474,In_856);
and U4599 (N_4599,In_914,In_2414);
and U4600 (N_4600,In_322,In_1099);
xnor U4601 (N_4601,In_621,In_211);
or U4602 (N_4602,In_1745,In_284);
nor U4603 (N_4603,In_747,In_2465);
nor U4604 (N_4604,In_336,In_1131);
nor U4605 (N_4605,In_746,In_2067);
nand U4606 (N_4606,In_2216,In_1477);
nor U4607 (N_4607,In_1476,In_1707);
xnor U4608 (N_4608,In_1227,In_2130);
and U4609 (N_4609,In_1609,In_6);
nand U4610 (N_4610,In_2147,In_1085);
and U4611 (N_4611,In_2080,In_1754);
or U4612 (N_4612,In_1320,In_1365);
or U4613 (N_4613,In_2241,In_535);
nand U4614 (N_4614,In_852,In_181);
nor U4615 (N_4615,In_519,In_1354);
nand U4616 (N_4616,In_1123,In_1923);
and U4617 (N_4617,In_301,In_128);
nand U4618 (N_4618,In_0,In_405);
and U4619 (N_4619,In_1681,In_532);
xor U4620 (N_4620,In_528,In_2024);
or U4621 (N_4621,In_1993,In_2151);
or U4622 (N_4622,In_1447,In_1821);
or U4623 (N_4623,In_479,In_2111);
and U4624 (N_4624,In_1802,In_2381);
or U4625 (N_4625,In_2424,In_378);
nand U4626 (N_4626,In_1883,In_1329);
nand U4627 (N_4627,In_1101,In_345);
xor U4628 (N_4628,In_2051,In_1096);
nand U4629 (N_4629,In_231,In_1075);
nand U4630 (N_4630,In_1645,In_1092);
nand U4631 (N_4631,In_1229,In_1660);
nand U4632 (N_4632,In_1689,In_863);
nand U4633 (N_4633,In_519,In_1213);
nand U4634 (N_4634,In_91,In_683);
nand U4635 (N_4635,In_820,In_1735);
or U4636 (N_4636,In_1069,In_1053);
nand U4637 (N_4637,In_976,In_2285);
or U4638 (N_4638,In_177,In_2385);
nor U4639 (N_4639,In_1712,In_709);
or U4640 (N_4640,In_1089,In_2416);
and U4641 (N_4641,In_498,In_1694);
nand U4642 (N_4642,In_179,In_1879);
nor U4643 (N_4643,In_1501,In_981);
or U4644 (N_4644,In_2496,In_2251);
and U4645 (N_4645,In_959,In_766);
nand U4646 (N_4646,In_363,In_1053);
and U4647 (N_4647,In_2104,In_1647);
nand U4648 (N_4648,In_1287,In_1779);
or U4649 (N_4649,In_1220,In_1945);
or U4650 (N_4650,In_1574,In_66);
and U4651 (N_4651,In_1215,In_1945);
and U4652 (N_4652,In_335,In_2047);
and U4653 (N_4653,In_882,In_786);
nand U4654 (N_4654,In_682,In_1334);
or U4655 (N_4655,In_2451,In_2158);
and U4656 (N_4656,In_273,In_1570);
or U4657 (N_4657,In_496,In_2490);
and U4658 (N_4658,In_2042,In_2161);
or U4659 (N_4659,In_2070,In_1127);
and U4660 (N_4660,In_1599,In_1804);
nand U4661 (N_4661,In_550,In_1891);
xor U4662 (N_4662,In_1845,In_1003);
or U4663 (N_4663,In_2139,In_2007);
and U4664 (N_4664,In_1344,In_1653);
nand U4665 (N_4665,In_289,In_3);
nand U4666 (N_4666,In_1220,In_2064);
nand U4667 (N_4667,In_898,In_285);
nor U4668 (N_4668,In_1518,In_2078);
nand U4669 (N_4669,In_849,In_1612);
nand U4670 (N_4670,In_2123,In_2419);
nand U4671 (N_4671,In_38,In_1906);
nand U4672 (N_4672,In_682,In_272);
nor U4673 (N_4673,In_1829,In_1503);
and U4674 (N_4674,In_1496,In_1939);
and U4675 (N_4675,In_987,In_140);
and U4676 (N_4676,In_1177,In_1288);
nor U4677 (N_4677,In_1135,In_1653);
and U4678 (N_4678,In_335,In_1982);
or U4679 (N_4679,In_587,In_949);
nand U4680 (N_4680,In_1239,In_533);
xnor U4681 (N_4681,In_534,In_1066);
and U4682 (N_4682,In_929,In_1091);
nor U4683 (N_4683,In_960,In_2028);
nor U4684 (N_4684,In_2238,In_1150);
nand U4685 (N_4685,In_1510,In_1815);
xor U4686 (N_4686,In_1169,In_238);
or U4687 (N_4687,In_2319,In_1342);
and U4688 (N_4688,In_851,In_1349);
or U4689 (N_4689,In_160,In_1845);
nor U4690 (N_4690,In_2173,In_810);
nor U4691 (N_4691,In_637,In_1921);
or U4692 (N_4692,In_1788,In_1054);
or U4693 (N_4693,In_1428,In_1423);
xor U4694 (N_4694,In_1628,In_567);
nand U4695 (N_4695,In_1751,In_264);
nor U4696 (N_4696,In_322,In_2219);
nand U4697 (N_4697,In_627,In_1560);
and U4698 (N_4698,In_434,In_159);
nor U4699 (N_4699,In_815,In_1009);
and U4700 (N_4700,In_1694,In_418);
and U4701 (N_4701,In_1361,In_2045);
xnor U4702 (N_4702,In_1288,In_1894);
nand U4703 (N_4703,In_1511,In_1714);
nor U4704 (N_4704,In_2173,In_1403);
or U4705 (N_4705,In_2245,In_1154);
nand U4706 (N_4706,In_226,In_1285);
and U4707 (N_4707,In_185,In_2279);
and U4708 (N_4708,In_2169,In_2418);
and U4709 (N_4709,In_1541,In_151);
and U4710 (N_4710,In_1322,In_1459);
xnor U4711 (N_4711,In_1110,In_1038);
nand U4712 (N_4712,In_1578,In_582);
and U4713 (N_4713,In_1522,In_1455);
or U4714 (N_4714,In_2304,In_629);
nor U4715 (N_4715,In_1272,In_1789);
and U4716 (N_4716,In_1339,In_1611);
or U4717 (N_4717,In_1939,In_1953);
nor U4718 (N_4718,In_60,In_1946);
nor U4719 (N_4719,In_388,In_372);
or U4720 (N_4720,In_612,In_2465);
nand U4721 (N_4721,In_1849,In_1878);
and U4722 (N_4722,In_238,In_2027);
xor U4723 (N_4723,In_1736,In_335);
or U4724 (N_4724,In_1037,In_1912);
nor U4725 (N_4725,In_2400,In_855);
nand U4726 (N_4726,In_2435,In_1271);
and U4727 (N_4727,In_283,In_1101);
xnor U4728 (N_4728,In_1172,In_587);
nand U4729 (N_4729,In_2300,In_945);
nor U4730 (N_4730,In_2341,In_796);
and U4731 (N_4731,In_2074,In_2440);
nor U4732 (N_4732,In_32,In_1531);
or U4733 (N_4733,In_2146,In_1103);
or U4734 (N_4734,In_946,In_1679);
or U4735 (N_4735,In_1304,In_557);
nand U4736 (N_4736,In_1635,In_1238);
and U4737 (N_4737,In_1713,In_56);
and U4738 (N_4738,In_1987,In_2450);
nor U4739 (N_4739,In_1994,In_2199);
nand U4740 (N_4740,In_101,In_1191);
or U4741 (N_4741,In_993,In_628);
nor U4742 (N_4742,In_244,In_2229);
and U4743 (N_4743,In_1617,In_2084);
and U4744 (N_4744,In_345,In_285);
and U4745 (N_4745,In_1652,In_564);
and U4746 (N_4746,In_2421,In_2009);
and U4747 (N_4747,In_1122,In_1119);
and U4748 (N_4748,In_903,In_1944);
nor U4749 (N_4749,In_1401,In_2207);
nand U4750 (N_4750,In_168,In_120);
xnor U4751 (N_4751,In_956,In_1501);
or U4752 (N_4752,In_380,In_2380);
nand U4753 (N_4753,In_1327,In_2006);
nor U4754 (N_4754,In_2263,In_2356);
xor U4755 (N_4755,In_952,In_1915);
nand U4756 (N_4756,In_901,In_884);
nor U4757 (N_4757,In_2380,In_679);
or U4758 (N_4758,In_1262,In_862);
or U4759 (N_4759,In_1749,In_1424);
xnor U4760 (N_4760,In_1975,In_348);
and U4761 (N_4761,In_1676,In_230);
xor U4762 (N_4762,In_598,In_885);
nand U4763 (N_4763,In_2224,In_931);
and U4764 (N_4764,In_2145,In_208);
and U4765 (N_4765,In_1978,In_1224);
nor U4766 (N_4766,In_2227,In_1069);
nor U4767 (N_4767,In_2353,In_623);
and U4768 (N_4768,In_149,In_2024);
nand U4769 (N_4769,In_1678,In_120);
nor U4770 (N_4770,In_1332,In_137);
and U4771 (N_4771,In_347,In_556);
xnor U4772 (N_4772,In_216,In_645);
nand U4773 (N_4773,In_1412,In_534);
or U4774 (N_4774,In_2088,In_2347);
nand U4775 (N_4775,In_844,In_1704);
or U4776 (N_4776,In_1713,In_1805);
and U4777 (N_4777,In_2359,In_2066);
and U4778 (N_4778,In_2491,In_734);
or U4779 (N_4779,In_719,In_439);
and U4780 (N_4780,In_741,In_183);
nand U4781 (N_4781,In_1360,In_1395);
and U4782 (N_4782,In_2342,In_1167);
nand U4783 (N_4783,In_1518,In_1033);
and U4784 (N_4784,In_1747,In_24);
and U4785 (N_4785,In_2160,In_1844);
nand U4786 (N_4786,In_1501,In_1469);
xnor U4787 (N_4787,In_1839,In_975);
and U4788 (N_4788,In_984,In_293);
or U4789 (N_4789,In_212,In_296);
and U4790 (N_4790,In_597,In_772);
and U4791 (N_4791,In_2473,In_1530);
and U4792 (N_4792,In_2184,In_596);
nand U4793 (N_4793,In_2372,In_169);
xor U4794 (N_4794,In_2375,In_530);
or U4795 (N_4795,In_1296,In_1867);
xor U4796 (N_4796,In_280,In_2102);
and U4797 (N_4797,In_948,In_827);
nand U4798 (N_4798,In_453,In_2289);
nor U4799 (N_4799,In_502,In_641);
nor U4800 (N_4800,In_760,In_186);
or U4801 (N_4801,In_2307,In_1184);
nand U4802 (N_4802,In_482,In_319);
or U4803 (N_4803,In_1479,In_117);
and U4804 (N_4804,In_1075,In_1955);
nand U4805 (N_4805,In_1363,In_1605);
xnor U4806 (N_4806,In_800,In_1675);
and U4807 (N_4807,In_2495,In_422);
nor U4808 (N_4808,In_1575,In_1018);
and U4809 (N_4809,In_2277,In_100);
or U4810 (N_4810,In_542,In_1818);
nor U4811 (N_4811,In_1250,In_525);
nor U4812 (N_4812,In_1408,In_365);
and U4813 (N_4813,In_1412,In_2438);
nor U4814 (N_4814,In_2142,In_422);
nor U4815 (N_4815,In_2235,In_1544);
or U4816 (N_4816,In_1904,In_2152);
nand U4817 (N_4817,In_428,In_241);
xnor U4818 (N_4818,In_510,In_1143);
or U4819 (N_4819,In_1691,In_229);
or U4820 (N_4820,In_1587,In_587);
xor U4821 (N_4821,In_1009,In_2082);
nand U4822 (N_4822,In_1494,In_1700);
xnor U4823 (N_4823,In_77,In_695);
nand U4824 (N_4824,In_269,In_1177);
nor U4825 (N_4825,In_1684,In_768);
nand U4826 (N_4826,In_2322,In_2221);
and U4827 (N_4827,In_764,In_194);
nor U4828 (N_4828,In_1991,In_564);
and U4829 (N_4829,In_874,In_1659);
or U4830 (N_4830,In_2408,In_894);
and U4831 (N_4831,In_271,In_2279);
nor U4832 (N_4832,In_1307,In_442);
nand U4833 (N_4833,In_1436,In_583);
or U4834 (N_4834,In_1333,In_1999);
or U4835 (N_4835,In_519,In_2);
or U4836 (N_4836,In_2017,In_1366);
and U4837 (N_4837,In_1569,In_2157);
nor U4838 (N_4838,In_2222,In_2201);
or U4839 (N_4839,In_2366,In_106);
or U4840 (N_4840,In_1527,In_955);
or U4841 (N_4841,In_2491,In_992);
or U4842 (N_4842,In_1178,In_322);
nor U4843 (N_4843,In_1757,In_226);
xnor U4844 (N_4844,In_1785,In_827);
or U4845 (N_4845,In_1615,In_883);
nand U4846 (N_4846,In_1989,In_1901);
or U4847 (N_4847,In_610,In_265);
xnor U4848 (N_4848,In_1446,In_1931);
nand U4849 (N_4849,In_2367,In_669);
nor U4850 (N_4850,In_2216,In_2342);
xor U4851 (N_4851,In_1191,In_1795);
nand U4852 (N_4852,In_1345,In_2375);
and U4853 (N_4853,In_2065,In_1142);
and U4854 (N_4854,In_1137,In_1478);
or U4855 (N_4855,In_708,In_1567);
and U4856 (N_4856,In_1433,In_1940);
xor U4857 (N_4857,In_310,In_137);
or U4858 (N_4858,In_1729,In_984);
or U4859 (N_4859,In_125,In_2494);
nand U4860 (N_4860,In_1120,In_1850);
nor U4861 (N_4861,In_533,In_2396);
and U4862 (N_4862,In_433,In_838);
nand U4863 (N_4863,In_1993,In_520);
nand U4864 (N_4864,In_212,In_117);
xor U4865 (N_4865,In_1370,In_2415);
xnor U4866 (N_4866,In_335,In_136);
or U4867 (N_4867,In_107,In_482);
xnor U4868 (N_4868,In_1574,In_1000);
nand U4869 (N_4869,In_549,In_119);
nand U4870 (N_4870,In_201,In_2093);
nor U4871 (N_4871,In_2153,In_2098);
and U4872 (N_4872,In_282,In_272);
nand U4873 (N_4873,In_514,In_11);
nor U4874 (N_4874,In_2183,In_1289);
nor U4875 (N_4875,In_638,In_1233);
nand U4876 (N_4876,In_2474,In_1111);
and U4877 (N_4877,In_717,In_973);
nand U4878 (N_4878,In_1400,In_1646);
or U4879 (N_4879,In_2220,In_1303);
and U4880 (N_4880,In_2063,In_64);
or U4881 (N_4881,In_1906,In_1325);
nand U4882 (N_4882,In_1188,In_890);
or U4883 (N_4883,In_1290,In_2147);
or U4884 (N_4884,In_1546,In_1075);
nand U4885 (N_4885,In_492,In_834);
nand U4886 (N_4886,In_855,In_1359);
and U4887 (N_4887,In_857,In_393);
nor U4888 (N_4888,In_2479,In_1880);
nand U4889 (N_4889,In_2079,In_2452);
nor U4890 (N_4890,In_2264,In_1320);
nand U4891 (N_4891,In_1030,In_655);
nor U4892 (N_4892,In_1286,In_708);
nand U4893 (N_4893,In_1792,In_1057);
or U4894 (N_4894,In_1536,In_2249);
nand U4895 (N_4895,In_1256,In_1204);
nor U4896 (N_4896,In_80,In_1328);
or U4897 (N_4897,In_2453,In_1236);
nand U4898 (N_4898,In_387,In_1160);
nor U4899 (N_4899,In_1569,In_1936);
or U4900 (N_4900,In_219,In_1109);
and U4901 (N_4901,In_555,In_1831);
nor U4902 (N_4902,In_380,In_290);
and U4903 (N_4903,In_1968,In_1085);
nand U4904 (N_4904,In_615,In_1941);
and U4905 (N_4905,In_466,In_442);
nand U4906 (N_4906,In_1569,In_477);
nand U4907 (N_4907,In_758,In_24);
nor U4908 (N_4908,In_700,In_2485);
or U4909 (N_4909,In_749,In_1071);
nor U4910 (N_4910,In_484,In_2058);
or U4911 (N_4911,In_929,In_128);
nand U4912 (N_4912,In_2270,In_698);
xnor U4913 (N_4913,In_352,In_1445);
xor U4914 (N_4914,In_459,In_2080);
or U4915 (N_4915,In_1267,In_305);
nand U4916 (N_4916,In_1138,In_1429);
and U4917 (N_4917,In_950,In_27);
and U4918 (N_4918,In_571,In_252);
and U4919 (N_4919,In_2338,In_2298);
and U4920 (N_4920,In_726,In_2247);
and U4921 (N_4921,In_565,In_2263);
and U4922 (N_4922,In_2469,In_2189);
nor U4923 (N_4923,In_981,In_1096);
nor U4924 (N_4924,In_89,In_298);
or U4925 (N_4925,In_1472,In_2494);
and U4926 (N_4926,In_291,In_1205);
nor U4927 (N_4927,In_2067,In_1786);
nor U4928 (N_4928,In_381,In_674);
and U4929 (N_4929,In_139,In_1885);
nor U4930 (N_4930,In_273,In_1143);
xor U4931 (N_4931,In_1454,In_2139);
or U4932 (N_4932,In_167,In_450);
or U4933 (N_4933,In_1463,In_1897);
and U4934 (N_4934,In_1176,In_1516);
and U4935 (N_4935,In_46,In_1386);
or U4936 (N_4936,In_1742,In_1764);
or U4937 (N_4937,In_311,In_2037);
nand U4938 (N_4938,In_1674,In_1826);
or U4939 (N_4939,In_1875,In_1342);
nor U4940 (N_4940,In_1336,In_735);
or U4941 (N_4941,In_1098,In_513);
nor U4942 (N_4942,In_1605,In_2065);
and U4943 (N_4943,In_505,In_76);
and U4944 (N_4944,In_1731,In_1701);
and U4945 (N_4945,In_1145,In_352);
nor U4946 (N_4946,In_1669,In_1892);
or U4947 (N_4947,In_247,In_140);
xnor U4948 (N_4948,In_2083,In_2022);
nand U4949 (N_4949,In_1314,In_1678);
xor U4950 (N_4950,In_2458,In_439);
nor U4951 (N_4951,In_530,In_1840);
nor U4952 (N_4952,In_44,In_1219);
or U4953 (N_4953,In_1254,In_132);
and U4954 (N_4954,In_1611,In_761);
nor U4955 (N_4955,In_729,In_587);
xor U4956 (N_4956,In_1155,In_1369);
nor U4957 (N_4957,In_2206,In_419);
and U4958 (N_4958,In_472,In_995);
nand U4959 (N_4959,In_1491,In_2397);
nand U4960 (N_4960,In_207,In_918);
nor U4961 (N_4961,In_664,In_577);
nor U4962 (N_4962,In_2380,In_415);
nand U4963 (N_4963,In_818,In_1383);
or U4964 (N_4964,In_918,In_2449);
and U4965 (N_4965,In_1250,In_2443);
nand U4966 (N_4966,In_2206,In_139);
and U4967 (N_4967,In_1157,In_26);
xor U4968 (N_4968,In_1009,In_1613);
nand U4969 (N_4969,In_2138,In_894);
and U4970 (N_4970,In_1759,In_1100);
and U4971 (N_4971,In_201,In_341);
nor U4972 (N_4972,In_1640,In_927);
or U4973 (N_4973,In_754,In_620);
xor U4974 (N_4974,In_278,In_1157);
nor U4975 (N_4975,In_987,In_2309);
and U4976 (N_4976,In_2196,In_1624);
nor U4977 (N_4977,In_2374,In_1040);
nor U4978 (N_4978,In_1614,In_1896);
or U4979 (N_4979,In_960,In_19);
nor U4980 (N_4980,In_157,In_1812);
or U4981 (N_4981,In_957,In_1832);
or U4982 (N_4982,In_592,In_184);
or U4983 (N_4983,In_1028,In_544);
nor U4984 (N_4984,In_1151,In_276);
nand U4985 (N_4985,In_2398,In_1682);
xnor U4986 (N_4986,In_168,In_1941);
and U4987 (N_4987,In_250,In_2323);
nor U4988 (N_4988,In_2340,In_951);
and U4989 (N_4989,In_2215,In_379);
xnor U4990 (N_4990,In_292,In_58);
and U4991 (N_4991,In_261,In_1636);
xnor U4992 (N_4992,In_1890,In_2334);
nand U4993 (N_4993,In_394,In_275);
nand U4994 (N_4994,In_306,In_80);
nor U4995 (N_4995,In_2211,In_1996);
nand U4996 (N_4996,In_667,In_2260);
nand U4997 (N_4997,In_1307,In_1138);
nor U4998 (N_4998,In_622,In_2451);
nor U4999 (N_4999,In_159,In_1559);
and U5000 (N_5000,In_2205,In_2050);
nand U5001 (N_5001,In_1917,In_1203);
nand U5002 (N_5002,In_1608,In_205);
nand U5003 (N_5003,In_1314,In_658);
and U5004 (N_5004,In_1664,In_1170);
nor U5005 (N_5005,In_1730,In_987);
nor U5006 (N_5006,In_2061,In_1645);
nand U5007 (N_5007,In_1455,In_2408);
xnor U5008 (N_5008,In_1084,In_255);
or U5009 (N_5009,In_418,In_749);
nand U5010 (N_5010,In_1018,In_816);
and U5011 (N_5011,In_123,In_789);
nand U5012 (N_5012,In_54,In_2216);
or U5013 (N_5013,In_1491,In_824);
nor U5014 (N_5014,In_1518,In_855);
nand U5015 (N_5015,In_2147,In_1947);
nand U5016 (N_5016,In_2367,In_660);
nand U5017 (N_5017,In_1030,In_1595);
and U5018 (N_5018,In_654,In_1884);
nor U5019 (N_5019,In_2457,In_538);
and U5020 (N_5020,In_7,In_1245);
nand U5021 (N_5021,In_1033,In_1666);
and U5022 (N_5022,In_2423,In_2288);
and U5023 (N_5023,In_390,In_2063);
nand U5024 (N_5024,In_527,In_1247);
and U5025 (N_5025,In_2498,In_346);
or U5026 (N_5026,In_2258,In_47);
and U5027 (N_5027,In_1051,In_529);
nand U5028 (N_5028,In_773,In_2405);
nand U5029 (N_5029,In_2410,In_1275);
nor U5030 (N_5030,In_1310,In_2367);
xnor U5031 (N_5031,In_1801,In_1938);
nand U5032 (N_5032,In_134,In_1004);
or U5033 (N_5033,In_526,In_1747);
nor U5034 (N_5034,In_563,In_2233);
and U5035 (N_5035,In_2043,In_2297);
xnor U5036 (N_5036,In_136,In_67);
or U5037 (N_5037,In_1988,In_2392);
nor U5038 (N_5038,In_2363,In_1880);
or U5039 (N_5039,In_2433,In_2275);
nand U5040 (N_5040,In_1824,In_79);
or U5041 (N_5041,In_1276,In_878);
nor U5042 (N_5042,In_1944,In_1742);
or U5043 (N_5043,In_893,In_807);
nand U5044 (N_5044,In_1060,In_403);
xor U5045 (N_5045,In_2047,In_1093);
nor U5046 (N_5046,In_1867,In_1184);
nor U5047 (N_5047,In_2008,In_653);
or U5048 (N_5048,In_527,In_174);
nor U5049 (N_5049,In_802,In_1778);
or U5050 (N_5050,In_1798,In_110);
and U5051 (N_5051,In_2463,In_2177);
nor U5052 (N_5052,In_423,In_697);
or U5053 (N_5053,In_777,In_683);
and U5054 (N_5054,In_178,In_1952);
and U5055 (N_5055,In_1085,In_608);
and U5056 (N_5056,In_576,In_367);
nand U5057 (N_5057,In_2336,In_820);
and U5058 (N_5058,In_2385,In_2395);
or U5059 (N_5059,In_2068,In_1244);
and U5060 (N_5060,In_1616,In_13);
nor U5061 (N_5061,In_2362,In_827);
or U5062 (N_5062,In_1479,In_1843);
nor U5063 (N_5063,In_1773,In_1523);
nor U5064 (N_5064,In_1563,In_1745);
xor U5065 (N_5065,In_930,In_2249);
nand U5066 (N_5066,In_2064,In_97);
or U5067 (N_5067,In_2359,In_187);
nor U5068 (N_5068,In_954,In_623);
or U5069 (N_5069,In_630,In_2280);
or U5070 (N_5070,In_1763,In_1024);
or U5071 (N_5071,In_2236,In_52);
or U5072 (N_5072,In_1889,In_929);
xnor U5073 (N_5073,In_1729,In_435);
or U5074 (N_5074,In_2081,In_562);
nand U5075 (N_5075,In_300,In_1811);
nor U5076 (N_5076,In_724,In_1987);
nor U5077 (N_5077,In_2083,In_137);
or U5078 (N_5078,In_1291,In_744);
nand U5079 (N_5079,In_228,In_1760);
or U5080 (N_5080,In_2296,In_828);
and U5081 (N_5081,In_1978,In_286);
or U5082 (N_5082,In_1273,In_2424);
nand U5083 (N_5083,In_2036,In_2069);
and U5084 (N_5084,In_453,In_637);
nor U5085 (N_5085,In_1974,In_2121);
or U5086 (N_5086,In_989,In_921);
or U5087 (N_5087,In_675,In_1012);
nand U5088 (N_5088,In_1982,In_1282);
nor U5089 (N_5089,In_1928,In_2124);
or U5090 (N_5090,In_1045,In_637);
nand U5091 (N_5091,In_319,In_938);
nor U5092 (N_5092,In_864,In_200);
and U5093 (N_5093,In_1846,In_1047);
nor U5094 (N_5094,In_2263,In_1735);
or U5095 (N_5095,In_1,In_1352);
nor U5096 (N_5096,In_492,In_737);
or U5097 (N_5097,In_594,In_1551);
xnor U5098 (N_5098,In_492,In_2066);
xnor U5099 (N_5099,In_980,In_1028);
nand U5100 (N_5100,In_1545,In_1426);
nand U5101 (N_5101,In_1986,In_473);
and U5102 (N_5102,In_1744,In_2311);
nand U5103 (N_5103,In_1499,In_1589);
and U5104 (N_5104,In_756,In_2451);
or U5105 (N_5105,In_96,In_2087);
or U5106 (N_5106,In_211,In_1958);
and U5107 (N_5107,In_636,In_527);
and U5108 (N_5108,In_240,In_1588);
nor U5109 (N_5109,In_1507,In_731);
nor U5110 (N_5110,In_348,In_2153);
and U5111 (N_5111,In_1049,In_1825);
nand U5112 (N_5112,In_1538,In_808);
nand U5113 (N_5113,In_2225,In_769);
xnor U5114 (N_5114,In_377,In_956);
and U5115 (N_5115,In_177,In_668);
nand U5116 (N_5116,In_613,In_1523);
and U5117 (N_5117,In_464,In_570);
and U5118 (N_5118,In_1300,In_1671);
nor U5119 (N_5119,In_1194,In_673);
xnor U5120 (N_5120,In_550,In_521);
and U5121 (N_5121,In_789,In_684);
nand U5122 (N_5122,In_2160,In_1214);
nand U5123 (N_5123,In_21,In_898);
nand U5124 (N_5124,In_911,In_1905);
xor U5125 (N_5125,In_354,In_1455);
and U5126 (N_5126,In_1871,In_139);
or U5127 (N_5127,In_1718,In_1565);
or U5128 (N_5128,In_2082,In_582);
or U5129 (N_5129,In_488,In_1618);
and U5130 (N_5130,In_1454,In_139);
nor U5131 (N_5131,In_1381,In_1956);
and U5132 (N_5132,In_480,In_897);
and U5133 (N_5133,In_1766,In_1223);
nor U5134 (N_5134,In_2377,In_1788);
xnor U5135 (N_5135,In_1845,In_1806);
nor U5136 (N_5136,In_1329,In_641);
and U5137 (N_5137,In_15,In_279);
nand U5138 (N_5138,In_1905,In_1621);
nand U5139 (N_5139,In_2408,In_804);
nor U5140 (N_5140,In_478,In_2081);
or U5141 (N_5141,In_2202,In_1947);
xnor U5142 (N_5142,In_1130,In_1675);
and U5143 (N_5143,In_1511,In_502);
nor U5144 (N_5144,In_2360,In_2167);
and U5145 (N_5145,In_642,In_2422);
and U5146 (N_5146,In_2304,In_2471);
nor U5147 (N_5147,In_1442,In_1333);
nor U5148 (N_5148,In_1539,In_1800);
nand U5149 (N_5149,In_1847,In_1196);
nor U5150 (N_5150,In_1300,In_1172);
or U5151 (N_5151,In_1887,In_2499);
nand U5152 (N_5152,In_67,In_97);
nor U5153 (N_5153,In_1526,In_53);
and U5154 (N_5154,In_1226,In_940);
and U5155 (N_5155,In_1380,In_1192);
or U5156 (N_5156,In_2209,In_1922);
nand U5157 (N_5157,In_559,In_1169);
and U5158 (N_5158,In_1614,In_1216);
or U5159 (N_5159,In_24,In_901);
xnor U5160 (N_5160,In_845,In_2409);
xor U5161 (N_5161,In_2254,In_415);
or U5162 (N_5162,In_312,In_2313);
or U5163 (N_5163,In_393,In_750);
nand U5164 (N_5164,In_1057,In_2445);
xor U5165 (N_5165,In_1199,In_1569);
or U5166 (N_5166,In_1671,In_1673);
nand U5167 (N_5167,In_442,In_479);
nor U5168 (N_5168,In_166,In_780);
nand U5169 (N_5169,In_1971,In_1223);
or U5170 (N_5170,In_2420,In_2340);
xor U5171 (N_5171,In_492,In_1808);
nand U5172 (N_5172,In_1810,In_2202);
nor U5173 (N_5173,In_1080,In_1144);
xor U5174 (N_5174,In_431,In_916);
nand U5175 (N_5175,In_38,In_2272);
nor U5176 (N_5176,In_304,In_1021);
nand U5177 (N_5177,In_2175,In_1058);
and U5178 (N_5178,In_2328,In_382);
or U5179 (N_5179,In_922,In_11);
and U5180 (N_5180,In_2162,In_1496);
and U5181 (N_5181,In_2073,In_1950);
nor U5182 (N_5182,In_1212,In_1870);
or U5183 (N_5183,In_2225,In_1279);
and U5184 (N_5184,In_1448,In_1590);
nor U5185 (N_5185,In_1353,In_501);
nor U5186 (N_5186,In_145,In_1145);
nand U5187 (N_5187,In_1810,In_1482);
or U5188 (N_5188,In_2365,In_969);
nand U5189 (N_5189,In_1730,In_704);
xnor U5190 (N_5190,In_856,In_2216);
xnor U5191 (N_5191,In_1938,In_1572);
or U5192 (N_5192,In_1423,In_236);
or U5193 (N_5193,In_1971,In_1142);
or U5194 (N_5194,In_885,In_1650);
or U5195 (N_5195,In_2468,In_692);
and U5196 (N_5196,In_394,In_119);
or U5197 (N_5197,In_1339,In_783);
nor U5198 (N_5198,In_1209,In_2475);
and U5199 (N_5199,In_2101,In_1841);
and U5200 (N_5200,In_767,In_601);
nand U5201 (N_5201,In_580,In_2390);
and U5202 (N_5202,In_2174,In_1242);
or U5203 (N_5203,In_441,In_87);
and U5204 (N_5204,In_1995,In_1683);
nand U5205 (N_5205,In_2469,In_2000);
and U5206 (N_5206,In_698,In_264);
nand U5207 (N_5207,In_2212,In_761);
or U5208 (N_5208,In_1087,In_1785);
nand U5209 (N_5209,In_562,In_2292);
nor U5210 (N_5210,In_155,In_1307);
nand U5211 (N_5211,In_1278,In_1308);
nor U5212 (N_5212,In_1157,In_461);
and U5213 (N_5213,In_2451,In_2234);
or U5214 (N_5214,In_2492,In_2376);
or U5215 (N_5215,In_1845,In_32);
nor U5216 (N_5216,In_154,In_2255);
and U5217 (N_5217,In_1525,In_975);
and U5218 (N_5218,In_1851,In_374);
xnor U5219 (N_5219,In_1370,In_404);
and U5220 (N_5220,In_1848,In_920);
or U5221 (N_5221,In_2011,In_873);
nor U5222 (N_5222,In_1913,In_1727);
nand U5223 (N_5223,In_2075,In_331);
and U5224 (N_5224,In_1313,In_2076);
or U5225 (N_5225,In_673,In_2403);
nand U5226 (N_5226,In_2072,In_1742);
nand U5227 (N_5227,In_2468,In_2203);
nand U5228 (N_5228,In_2455,In_762);
nor U5229 (N_5229,In_329,In_715);
or U5230 (N_5230,In_1320,In_965);
xor U5231 (N_5231,In_2464,In_1960);
or U5232 (N_5232,In_1736,In_1248);
or U5233 (N_5233,In_2426,In_62);
and U5234 (N_5234,In_620,In_1968);
nand U5235 (N_5235,In_775,In_431);
nand U5236 (N_5236,In_243,In_159);
or U5237 (N_5237,In_1011,In_710);
nand U5238 (N_5238,In_1032,In_121);
nand U5239 (N_5239,In_374,In_857);
nor U5240 (N_5240,In_587,In_2024);
xnor U5241 (N_5241,In_2498,In_906);
xor U5242 (N_5242,In_2495,In_1950);
nand U5243 (N_5243,In_209,In_1602);
nor U5244 (N_5244,In_1661,In_848);
nand U5245 (N_5245,In_103,In_1590);
nor U5246 (N_5246,In_133,In_1474);
or U5247 (N_5247,In_146,In_1297);
nor U5248 (N_5248,In_666,In_2415);
and U5249 (N_5249,In_258,In_979);
and U5250 (N_5250,In_1709,In_1507);
nand U5251 (N_5251,In_1513,In_175);
or U5252 (N_5252,In_1059,In_1228);
or U5253 (N_5253,In_459,In_1947);
and U5254 (N_5254,In_485,In_14);
and U5255 (N_5255,In_1406,In_1162);
or U5256 (N_5256,In_27,In_2089);
nand U5257 (N_5257,In_1,In_1761);
or U5258 (N_5258,In_1069,In_612);
or U5259 (N_5259,In_1450,In_2448);
nor U5260 (N_5260,In_1224,In_109);
nor U5261 (N_5261,In_2129,In_1543);
nor U5262 (N_5262,In_1462,In_312);
and U5263 (N_5263,In_2038,In_710);
nand U5264 (N_5264,In_1407,In_132);
nor U5265 (N_5265,In_1295,In_1482);
nor U5266 (N_5266,In_672,In_1604);
or U5267 (N_5267,In_2240,In_13);
or U5268 (N_5268,In_1363,In_934);
or U5269 (N_5269,In_1454,In_893);
nand U5270 (N_5270,In_1491,In_1723);
xor U5271 (N_5271,In_421,In_328);
and U5272 (N_5272,In_454,In_876);
nand U5273 (N_5273,In_1643,In_270);
nand U5274 (N_5274,In_99,In_989);
and U5275 (N_5275,In_520,In_1136);
nor U5276 (N_5276,In_1026,In_392);
nand U5277 (N_5277,In_2310,In_1410);
nand U5278 (N_5278,In_41,In_1106);
or U5279 (N_5279,In_1638,In_2173);
xor U5280 (N_5280,In_1618,In_2311);
or U5281 (N_5281,In_1984,In_1450);
or U5282 (N_5282,In_516,In_1258);
or U5283 (N_5283,In_1620,In_1915);
or U5284 (N_5284,In_161,In_346);
and U5285 (N_5285,In_2409,In_1267);
nand U5286 (N_5286,In_1378,In_395);
or U5287 (N_5287,In_1274,In_1767);
nor U5288 (N_5288,In_281,In_755);
nand U5289 (N_5289,In_1988,In_754);
nor U5290 (N_5290,In_1950,In_2338);
or U5291 (N_5291,In_1613,In_73);
and U5292 (N_5292,In_2130,In_1966);
and U5293 (N_5293,In_2041,In_2014);
nor U5294 (N_5294,In_2104,In_278);
and U5295 (N_5295,In_18,In_2431);
and U5296 (N_5296,In_186,In_855);
or U5297 (N_5297,In_660,In_947);
and U5298 (N_5298,In_442,In_423);
and U5299 (N_5299,In_328,In_124);
or U5300 (N_5300,In_1395,In_1217);
nor U5301 (N_5301,In_1157,In_2264);
nand U5302 (N_5302,In_824,In_1070);
and U5303 (N_5303,In_1431,In_527);
or U5304 (N_5304,In_1336,In_1122);
or U5305 (N_5305,In_1017,In_2345);
and U5306 (N_5306,In_2105,In_1206);
or U5307 (N_5307,In_240,In_1675);
nand U5308 (N_5308,In_2394,In_2070);
nor U5309 (N_5309,In_1693,In_1871);
or U5310 (N_5310,In_1147,In_2389);
nand U5311 (N_5311,In_770,In_873);
and U5312 (N_5312,In_1492,In_992);
and U5313 (N_5313,In_1966,In_2129);
and U5314 (N_5314,In_1031,In_239);
nor U5315 (N_5315,In_871,In_2218);
xnor U5316 (N_5316,In_681,In_1926);
nor U5317 (N_5317,In_877,In_953);
or U5318 (N_5318,In_1233,In_489);
nand U5319 (N_5319,In_2293,In_983);
and U5320 (N_5320,In_2262,In_760);
nand U5321 (N_5321,In_1627,In_711);
nor U5322 (N_5322,In_398,In_740);
or U5323 (N_5323,In_1954,In_1275);
nor U5324 (N_5324,In_576,In_231);
or U5325 (N_5325,In_2298,In_723);
and U5326 (N_5326,In_638,In_1198);
and U5327 (N_5327,In_2290,In_1587);
and U5328 (N_5328,In_1893,In_25);
xor U5329 (N_5329,In_1252,In_2464);
and U5330 (N_5330,In_378,In_595);
and U5331 (N_5331,In_2361,In_1848);
or U5332 (N_5332,In_1397,In_1900);
or U5333 (N_5333,In_252,In_1831);
and U5334 (N_5334,In_1573,In_1548);
or U5335 (N_5335,In_988,In_859);
and U5336 (N_5336,In_2266,In_993);
nand U5337 (N_5337,In_572,In_999);
nand U5338 (N_5338,In_88,In_1394);
nand U5339 (N_5339,In_278,In_828);
nand U5340 (N_5340,In_2396,In_717);
or U5341 (N_5341,In_1898,In_2221);
or U5342 (N_5342,In_638,In_1153);
nand U5343 (N_5343,In_1946,In_1650);
nor U5344 (N_5344,In_1102,In_2413);
nand U5345 (N_5345,In_251,In_888);
and U5346 (N_5346,In_695,In_645);
xor U5347 (N_5347,In_1302,In_1897);
nor U5348 (N_5348,In_2052,In_1901);
nand U5349 (N_5349,In_2232,In_1205);
or U5350 (N_5350,In_635,In_680);
or U5351 (N_5351,In_359,In_668);
nor U5352 (N_5352,In_2488,In_1367);
or U5353 (N_5353,In_198,In_1420);
and U5354 (N_5354,In_1835,In_1305);
and U5355 (N_5355,In_763,In_1027);
or U5356 (N_5356,In_1130,In_2096);
and U5357 (N_5357,In_2284,In_1440);
or U5358 (N_5358,In_1610,In_228);
nor U5359 (N_5359,In_530,In_1288);
or U5360 (N_5360,In_2375,In_1200);
nand U5361 (N_5361,In_864,In_1817);
nor U5362 (N_5362,In_591,In_428);
xnor U5363 (N_5363,In_896,In_740);
nand U5364 (N_5364,In_1843,In_2435);
nand U5365 (N_5365,In_912,In_1435);
and U5366 (N_5366,In_448,In_975);
xor U5367 (N_5367,In_1242,In_1572);
and U5368 (N_5368,In_1284,In_1319);
or U5369 (N_5369,In_1448,In_476);
nor U5370 (N_5370,In_731,In_43);
xnor U5371 (N_5371,In_1558,In_416);
nor U5372 (N_5372,In_2156,In_2189);
nor U5373 (N_5373,In_62,In_2237);
nor U5374 (N_5374,In_2455,In_2230);
nand U5375 (N_5375,In_604,In_1994);
nand U5376 (N_5376,In_2306,In_412);
nor U5377 (N_5377,In_2164,In_698);
xor U5378 (N_5378,In_2037,In_2468);
and U5379 (N_5379,In_2413,In_90);
nand U5380 (N_5380,In_1476,In_428);
nor U5381 (N_5381,In_2208,In_1797);
or U5382 (N_5382,In_1030,In_2496);
and U5383 (N_5383,In_2280,In_247);
nand U5384 (N_5384,In_1340,In_2335);
or U5385 (N_5385,In_1741,In_26);
and U5386 (N_5386,In_3,In_2350);
nand U5387 (N_5387,In_367,In_1738);
or U5388 (N_5388,In_2179,In_202);
nand U5389 (N_5389,In_1077,In_1600);
and U5390 (N_5390,In_150,In_1985);
xor U5391 (N_5391,In_1183,In_393);
xor U5392 (N_5392,In_2090,In_427);
and U5393 (N_5393,In_595,In_1229);
nand U5394 (N_5394,In_1204,In_594);
and U5395 (N_5395,In_1640,In_2059);
nand U5396 (N_5396,In_259,In_391);
nand U5397 (N_5397,In_1825,In_2067);
or U5398 (N_5398,In_2239,In_585);
xnor U5399 (N_5399,In_1949,In_1922);
or U5400 (N_5400,In_1214,In_1876);
nor U5401 (N_5401,In_771,In_1850);
or U5402 (N_5402,In_1332,In_1367);
nand U5403 (N_5403,In_395,In_1479);
or U5404 (N_5404,In_599,In_940);
nand U5405 (N_5405,In_1968,In_484);
or U5406 (N_5406,In_518,In_305);
nand U5407 (N_5407,In_1995,In_2437);
nand U5408 (N_5408,In_1876,In_715);
nor U5409 (N_5409,In_1758,In_1880);
or U5410 (N_5410,In_696,In_2222);
nand U5411 (N_5411,In_984,In_806);
nand U5412 (N_5412,In_287,In_1069);
nand U5413 (N_5413,In_289,In_2221);
nand U5414 (N_5414,In_19,In_744);
nor U5415 (N_5415,In_1727,In_2456);
and U5416 (N_5416,In_1445,In_1782);
or U5417 (N_5417,In_1819,In_676);
or U5418 (N_5418,In_1588,In_684);
xor U5419 (N_5419,In_494,In_2164);
or U5420 (N_5420,In_1256,In_257);
and U5421 (N_5421,In_1409,In_2370);
and U5422 (N_5422,In_2195,In_1064);
or U5423 (N_5423,In_728,In_814);
nand U5424 (N_5424,In_902,In_2429);
nor U5425 (N_5425,In_1404,In_1154);
or U5426 (N_5426,In_621,In_1413);
nor U5427 (N_5427,In_1024,In_260);
nand U5428 (N_5428,In_1430,In_1401);
nor U5429 (N_5429,In_77,In_727);
and U5430 (N_5430,In_1272,In_1888);
and U5431 (N_5431,In_754,In_1415);
nand U5432 (N_5432,In_2281,In_944);
or U5433 (N_5433,In_2007,In_1526);
nor U5434 (N_5434,In_548,In_907);
nor U5435 (N_5435,In_1440,In_2465);
and U5436 (N_5436,In_992,In_1428);
nor U5437 (N_5437,In_343,In_381);
nand U5438 (N_5438,In_606,In_720);
xor U5439 (N_5439,In_2022,In_2021);
nand U5440 (N_5440,In_2241,In_978);
or U5441 (N_5441,In_906,In_2216);
nand U5442 (N_5442,In_1404,In_582);
and U5443 (N_5443,In_496,In_2352);
and U5444 (N_5444,In_755,In_1179);
and U5445 (N_5445,In_342,In_352);
and U5446 (N_5446,In_654,In_2302);
xnor U5447 (N_5447,In_1258,In_2001);
nor U5448 (N_5448,In_2226,In_1933);
or U5449 (N_5449,In_2124,In_2154);
nor U5450 (N_5450,In_732,In_1139);
and U5451 (N_5451,In_388,In_2392);
or U5452 (N_5452,In_1179,In_1965);
or U5453 (N_5453,In_1124,In_1203);
xor U5454 (N_5454,In_931,In_1968);
nor U5455 (N_5455,In_681,In_838);
or U5456 (N_5456,In_2302,In_2219);
nor U5457 (N_5457,In_114,In_1854);
or U5458 (N_5458,In_1152,In_1812);
nor U5459 (N_5459,In_30,In_678);
xnor U5460 (N_5460,In_1293,In_861);
nand U5461 (N_5461,In_1024,In_1206);
or U5462 (N_5462,In_2095,In_940);
nor U5463 (N_5463,In_1310,In_567);
nor U5464 (N_5464,In_2490,In_1917);
or U5465 (N_5465,In_2457,In_1254);
nor U5466 (N_5466,In_162,In_1591);
nand U5467 (N_5467,In_271,In_125);
xnor U5468 (N_5468,In_1231,In_845);
nand U5469 (N_5469,In_1766,In_2083);
nor U5470 (N_5470,In_941,In_2214);
or U5471 (N_5471,In_235,In_2392);
nand U5472 (N_5472,In_1366,In_1595);
or U5473 (N_5473,In_2227,In_1657);
nand U5474 (N_5474,In_852,In_1312);
nand U5475 (N_5475,In_942,In_1362);
xnor U5476 (N_5476,In_2200,In_1205);
or U5477 (N_5477,In_1769,In_845);
nor U5478 (N_5478,In_1053,In_361);
nand U5479 (N_5479,In_2167,In_83);
nor U5480 (N_5480,In_62,In_2381);
and U5481 (N_5481,In_2338,In_632);
nor U5482 (N_5482,In_1912,In_843);
xor U5483 (N_5483,In_419,In_838);
nor U5484 (N_5484,In_1475,In_2053);
or U5485 (N_5485,In_395,In_847);
nor U5486 (N_5486,In_1603,In_43);
and U5487 (N_5487,In_2482,In_532);
or U5488 (N_5488,In_1514,In_1626);
or U5489 (N_5489,In_1249,In_2226);
and U5490 (N_5490,In_476,In_603);
nand U5491 (N_5491,In_1185,In_654);
nand U5492 (N_5492,In_714,In_2010);
nand U5493 (N_5493,In_1000,In_636);
nor U5494 (N_5494,In_2180,In_1789);
xnor U5495 (N_5495,In_1814,In_2058);
nor U5496 (N_5496,In_2200,In_193);
nand U5497 (N_5497,In_2027,In_2140);
or U5498 (N_5498,In_1221,In_1927);
nor U5499 (N_5499,In_47,In_355);
nand U5500 (N_5500,In_581,In_1097);
and U5501 (N_5501,In_905,In_415);
nand U5502 (N_5502,In_1535,In_414);
or U5503 (N_5503,In_1629,In_2293);
nand U5504 (N_5504,In_95,In_2080);
nor U5505 (N_5505,In_1464,In_861);
xnor U5506 (N_5506,In_690,In_5);
or U5507 (N_5507,In_1636,In_1309);
nor U5508 (N_5508,In_1652,In_1187);
xnor U5509 (N_5509,In_861,In_1975);
nor U5510 (N_5510,In_191,In_780);
and U5511 (N_5511,In_844,In_2027);
or U5512 (N_5512,In_982,In_658);
and U5513 (N_5513,In_2458,In_285);
and U5514 (N_5514,In_2142,In_2128);
and U5515 (N_5515,In_1538,In_283);
or U5516 (N_5516,In_50,In_1423);
and U5517 (N_5517,In_2258,In_324);
nand U5518 (N_5518,In_1588,In_185);
nor U5519 (N_5519,In_449,In_1792);
nand U5520 (N_5520,In_241,In_761);
or U5521 (N_5521,In_716,In_2085);
and U5522 (N_5522,In_1132,In_363);
nand U5523 (N_5523,In_1317,In_2347);
nor U5524 (N_5524,In_1054,In_2228);
and U5525 (N_5525,In_2151,In_66);
and U5526 (N_5526,In_1790,In_1197);
and U5527 (N_5527,In_1904,In_2491);
or U5528 (N_5528,In_1206,In_2110);
and U5529 (N_5529,In_2164,In_215);
or U5530 (N_5530,In_1907,In_1876);
and U5531 (N_5531,In_1115,In_1784);
xor U5532 (N_5532,In_74,In_369);
nand U5533 (N_5533,In_1165,In_333);
nand U5534 (N_5534,In_1914,In_2003);
or U5535 (N_5535,In_981,In_289);
and U5536 (N_5536,In_931,In_292);
or U5537 (N_5537,In_2459,In_2370);
nor U5538 (N_5538,In_840,In_1712);
xor U5539 (N_5539,In_46,In_2463);
nor U5540 (N_5540,In_18,In_1616);
and U5541 (N_5541,In_1544,In_2277);
or U5542 (N_5542,In_1608,In_1886);
nand U5543 (N_5543,In_1937,In_740);
and U5544 (N_5544,In_577,In_1661);
or U5545 (N_5545,In_829,In_411);
or U5546 (N_5546,In_32,In_1994);
nand U5547 (N_5547,In_2479,In_671);
xnor U5548 (N_5548,In_905,In_1826);
nand U5549 (N_5549,In_1614,In_1447);
nor U5550 (N_5550,In_659,In_1330);
nor U5551 (N_5551,In_2053,In_1084);
nand U5552 (N_5552,In_177,In_1370);
or U5553 (N_5553,In_1582,In_1065);
xnor U5554 (N_5554,In_1738,In_608);
nand U5555 (N_5555,In_2141,In_276);
or U5556 (N_5556,In_830,In_731);
and U5557 (N_5557,In_641,In_1250);
nor U5558 (N_5558,In_703,In_2310);
and U5559 (N_5559,In_974,In_1753);
nor U5560 (N_5560,In_147,In_2046);
or U5561 (N_5561,In_612,In_769);
xnor U5562 (N_5562,In_15,In_1819);
or U5563 (N_5563,In_1848,In_1979);
nand U5564 (N_5564,In_569,In_1972);
nor U5565 (N_5565,In_1476,In_1214);
nand U5566 (N_5566,In_1388,In_637);
xnor U5567 (N_5567,In_1835,In_2024);
or U5568 (N_5568,In_2499,In_2488);
and U5569 (N_5569,In_878,In_608);
and U5570 (N_5570,In_1495,In_1020);
xnor U5571 (N_5571,In_1534,In_2369);
nand U5572 (N_5572,In_486,In_751);
nand U5573 (N_5573,In_2080,In_2161);
and U5574 (N_5574,In_1001,In_1626);
and U5575 (N_5575,In_612,In_379);
or U5576 (N_5576,In_2122,In_1557);
xor U5577 (N_5577,In_2043,In_2344);
or U5578 (N_5578,In_928,In_64);
nand U5579 (N_5579,In_1546,In_1572);
and U5580 (N_5580,In_1413,In_1507);
or U5581 (N_5581,In_2444,In_451);
or U5582 (N_5582,In_705,In_1735);
nor U5583 (N_5583,In_2018,In_1916);
nand U5584 (N_5584,In_2040,In_799);
and U5585 (N_5585,In_225,In_1083);
nor U5586 (N_5586,In_2305,In_2034);
nand U5587 (N_5587,In_201,In_1431);
and U5588 (N_5588,In_701,In_1106);
and U5589 (N_5589,In_1956,In_785);
nor U5590 (N_5590,In_904,In_346);
and U5591 (N_5591,In_498,In_1286);
and U5592 (N_5592,In_1724,In_1405);
and U5593 (N_5593,In_1864,In_1648);
nand U5594 (N_5594,In_974,In_688);
or U5595 (N_5595,In_795,In_1272);
or U5596 (N_5596,In_215,In_1149);
and U5597 (N_5597,In_720,In_2326);
nor U5598 (N_5598,In_2257,In_2386);
xor U5599 (N_5599,In_326,In_1252);
and U5600 (N_5600,In_1168,In_981);
and U5601 (N_5601,In_1203,In_245);
nor U5602 (N_5602,In_1513,In_760);
or U5603 (N_5603,In_262,In_2265);
and U5604 (N_5604,In_961,In_1817);
or U5605 (N_5605,In_410,In_1211);
or U5606 (N_5606,In_1454,In_1755);
nor U5607 (N_5607,In_2281,In_1005);
and U5608 (N_5608,In_321,In_1125);
nand U5609 (N_5609,In_238,In_637);
nand U5610 (N_5610,In_1179,In_1650);
and U5611 (N_5611,In_270,In_1662);
or U5612 (N_5612,In_1748,In_343);
nor U5613 (N_5613,In_110,In_570);
or U5614 (N_5614,In_2136,In_1888);
nor U5615 (N_5615,In_1476,In_659);
nor U5616 (N_5616,In_1285,In_1099);
nand U5617 (N_5617,In_1671,In_1614);
nor U5618 (N_5618,In_2191,In_272);
nor U5619 (N_5619,In_2414,In_1963);
xor U5620 (N_5620,In_21,In_509);
nor U5621 (N_5621,In_1819,In_1689);
or U5622 (N_5622,In_827,In_2356);
nor U5623 (N_5623,In_2324,In_1486);
or U5624 (N_5624,In_1238,In_1843);
and U5625 (N_5625,In_2431,In_690);
or U5626 (N_5626,In_1108,In_411);
or U5627 (N_5627,In_1576,In_2370);
and U5628 (N_5628,In_978,In_1502);
nor U5629 (N_5629,In_1729,In_2496);
xnor U5630 (N_5630,In_1516,In_1495);
or U5631 (N_5631,In_819,In_453);
and U5632 (N_5632,In_2472,In_456);
or U5633 (N_5633,In_1045,In_532);
xnor U5634 (N_5634,In_2137,In_252);
nor U5635 (N_5635,In_372,In_10);
nand U5636 (N_5636,In_2003,In_1678);
or U5637 (N_5637,In_1287,In_1406);
or U5638 (N_5638,In_2021,In_977);
and U5639 (N_5639,In_2054,In_819);
xnor U5640 (N_5640,In_476,In_1276);
nand U5641 (N_5641,In_2464,In_921);
nand U5642 (N_5642,In_134,In_1995);
or U5643 (N_5643,In_491,In_1723);
nand U5644 (N_5644,In_981,In_1901);
or U5645 (N_5645,In_1696,In_1232);
nand U5646 (N_5646,In_1300,In_111);
or U5647 (N_5647,In_138,In_2237);
nor U5648 (N_5648,In_1325,In_1263);
nor U5649 (N_5649,In_811,In_2422);
nand U5650 (N_5650,In_1666,In_1506);
xnor U5651 (N_5651,In_1871,In_671);
or U5652 (N_5652,In_562,In_1502);
or U5653 (N_5653,In_1355,In_2126);
nand U5654 (N_5654,In_2096,In_1934);
nor U5655 (N_5655,In_333,In_168);
and U5656 (N_5656,In_1166,In_996);
and U5657 (N_5657,In_901,In_1681);
nand U5658 (N_5658,In_1974,In_1614);
nand U5659 (N_5659,In_969,In_633);
or U5660 (N_5660,In_1264,In_1905);
nand U5661 (N_5661,In_437,In_2218);
or U5662 (N_5662,In_2125,In_1867);
xor U5663 (N_5663,In_558,In_2037);
and U5664 (N_5664,In_1625,In_1648);
and U5665 (N_5665,In_650,In_491);
nand U5666 (N_5666,In_1554,In_964);
and U5667 (N_5667,In_1289,In_288);
or U5668 (N_5668,In_2109,In_16);
nor U5669 (N_5669,In_1790,In_134);
nor U5670 (N_5670,In_2,In_175);
nor U5671 (N_5671,In_1726,In_299);
xor U5672 (N_5672,In_1529,In_751);
nand U5673 (N_5673,In_48,In_1082);
nand U5674 (N_5674,In_1323,In_1155);
nand U5675 (N_5675,In_1235,In_2410);
nor U5676 (N_5676,In_2178,In_410);
nor U5677 (N_5677,In_1042,In_2389);
or U5678 (N_5678,In_2205,In_1283);
and U5679 (N_5679,In_104,In_774);
and U5680 (N_5680,In_1741,In_1073);
nor U5681 (N_5681,In_1568,In_67);
or U5682 (N_5682,In_2259,In_790);
or U5683 (N_5683,In_1614,In_93);
nor U5684 (N_5684,In_2077,In_1629);
or U5685 (N_5685,In_403,In_524);
or U5686 (N_5686,In_1589,In_2107);
or U5687 (N_5687,In_667,In_912);
xnor U5688 (N_5688,In_193,In_1952);
and U5689 (N_5689,In_1258,In_1100);
or U5690 (N_5690,In_535,In_365);
nand U5691 (N_5691,In_24,In_2206);
nand U5692 (N_5692,In_780,In_1865);
nand U5693 (N_5693,In_1730,In_1744);
and U5694 (N_5694,In_91,In_1323);
and U5695 (N_5695,In_771,In_1885);
or U5696 (N_5696,In_899,In_1987);
nand U5697 (N_5697,In_635,In_1313);
nor U5698 (N_5698,In_2154,In_406);
and U5699 (N_5699,In_1550,In_1032);
nand U5700 (N_5700,In_622,In_1532);
nor U5701 (N_5701,In_664,In_653);
nand U5702 (N_5702,In_2246,In_2482);
nand U5703 (N_5703,In_1539,In_1398);
nor U5704 (N_5704,In_1629,In_2475);
xnor U5705 (N_5705,In_1039,In_757);
nand U5706 (N_5706,In_1397,In_990);
nand U5707 (N_5707,In_365,In_953);
or U5708 (N_5708,In_1152,In_1027);
and U5709 (N_5709,In_1708,In_659);
nor U5710 (N_5710,In_1998,In_186);
nor U5711 (N_5711,In_74,In_1419);
or U5712 (N_5712,In_1191,In_1955);
nand U5713 (N_5713,In_475,In_1441);
or U5714 (N_5714,In_935,In_1959);
nor U5715 (N_5715,In_1133,In_833);
nor U5716 (N_5716,In_2147,In_1330);
nand U5717 (N_5717,In_1468,In_193);
nor U5718 (N_5718,In_958,In_1340);
and U5719 (N_5719,In_1926,In_1270);
xor U5720 (N_5720,In_2334,In_1276);
nand U5721 (N_5721,In_1488,In_522);
or U5722 (N_5722,In_1995,In_1483);
or U5723 (N_5723,In_1236,In_1363);
nor U5724 (N_5724,In_200,In_979);
nand U5725 (N_5725,In_2276,In_1850);
or U5726 (N_5726,In_1542,In_2434);
and U5727 (N_5727,In_1066,In_174);
and U5728 (N_5728,In_55,In_2089);
or U5729 (N_5729,In_636,In_105);
or U5730 (N_5730,In_347,In_696);
nand U5731 (N_5731,In_404,In_2043);
or U5732 (N_5732,In_984,In_19);
xor U5733 (N_5733,In_200,In_437);
or U5734 (N_5734,In_2032,In_125);
and U5735 (N_5735,In_1404,In_1503);
nand U5736 (N_5736,In_2365,In_408);
nor U5737 (N_5737,In_287,In_1549);
or U5738 (N_5738,In_241,In_123);
xor U5739 (N_5739,In_788,In_1935);
or U5740 (N_5740,In_2358,In_1460);
or U5741 (N_5741,In_1903,In_2067);
nand U5742 (N_5742,In_2391,In_304);
or U5743 (N_5743,In_523,In_2320);
or U5744 (N_5744,In_1436,In_1880);
or U5745 (N_5745,In_1707,In_599);
nor U5746 (N_5746,In_392,In_572);
xnor U5747 (N_5747,In_1698,In_966);
nand U5748 (N_5748,In_332,In_1127);
or U5749 (N_5749,In_1784,In_1609);
or U5750 (N_5750,In_136,In_1019);
xnor U5751 (N_5751,In_2225,In_160);
xnor U5752 (N_5752,In_1657,In_882);
nor U5753 (N_5753,In_1889,In_2168);
or U5754 (N_5754,In_2050,In_545);
and U5755 (N_5755,In_1136,In_1163);
and U5756 (N_5756,In_403,In_2208);
nand U5757 (N_5757,In_1198,In_1929);
and U5758 (N_5758,In_2267,In_673);
and U5759 (N_5759,In_1682,In_1277);
nand U5760 (N_5760,In_264,In_425);
nor U5761 (N_5761,In_1768,In_1600);
nor U5762 (N_5762,In_320,In_981);
or U5763 (N_5763,In_982,In_2485);
and U5764 (N_5764,In_607,In_82);
or U5765 (N_5765,In_1062,In_1442);
nor U5766 (N_5766,In_1684,In_1406);
and U5767 (N_5767,In_1839,In_1393);
and U5768 (N_5768,In_1704,In_287);
or U5769 (N_5769,In_1986,In_1195);
and U5770 (N_5770,In_454,In_2196);
or U5771 (N_5771,In_638,In_2120);
nor U5772 (N_5772,In_648,In_253);
xnor U5773 (N_5773,In_1910,In_787);
and U5774 (N_5774,In_861,In_740);
and U5775 (N_5775,In_307,In_1468);
nor U5776 (N_5776,In_184,In_1202);
nor U5777 (N_5777,In_945,In_1998);
nor U5778 (N_5778,In_2379,In_2071);
and U5779 (N_5779,In_573,In_1585);
and U5780 (N_5780,In_770,In_629);
or U5781 (N_5781,In_799,In_1277);
nand U5782 (N_5782,In_852,In_1692);
or U5783 (N_5783,In_1667,In_1963);
nor U5784 (N_5784,In_988,In_342);
and U5785 (N_5785,In_1795,In_1289);
or U5786 (N_5786,In_45,In_1984);
xor U5787 (N_5787,In_544,In_824);
and U5788 (N_5788,In_897,In_986);
nor U5789 (N_5789,In_1366,In_1958);
or U5790 (N_5790,In_1991,In_2106);
or U5791 (N_5791,In_131,In_729);
nand U5792 (N_5792,In_1947,In_176);
nor U5793 (N_5793,In_537,In_2289);
nand U5794 (N_5794,In_388,In_1933);
nand U5795 (N_5795,In_2153,In_713);
nand U5796 (N_5796,In_14,In_590);
nor U5797 (N_5797,In_344,In_1317);
and U5798 (N_5798,In_1019,In_924);
nor U5799 (N_5799,In_1008,In_225);
or U5800 (N_5800,In_2104,In_2088);
or U5801 (N_5801,In_48,In_1307);
nor U5802 (N_5802,In_373,In_1047);
or U5803 (N_5803,In_820,In_545);
nor U5804 (N_5804,In_1865,In_2424);
nor U5805 (N_5805,In_2240,In_2219);
nor U5806 (N_5806,In_1085,In_2372);
or U5807 (N_5807,In_826,In_1228);
and U5808 (N_5808,In_1638,In_1693);
or U5809 (N_5809,In_1425,In_404);
nand U5810 (N_5810,In_718,In_374);
nor U5811 (N_5811,In_451,In_1494);
nor U5812 (N_5812,In_1559,In_940);
or U5813 (N_5813,In_1715,In_1766);
nand U5814 (N_5814,In_1036,In_1374);
and U5815 (N_5815,In_181,In_757);
nor U5816 (N_5816,In_1477,In_2278);
and U5817 (N_5817,In_258,In_1347);
xnor U5818 (N_5818,In_1450,In_2381);
nor U5819 (N_5819,In_842,In_1362);
or U5820 (N_5820,In_1460,In_2192);
and U5821 (N_5821,In_1201,In_2192);
and U5822 (N_5822,In_2169,In_2212);
nor U5823 (N_5823,In_78,In_201);
nor U5824 (N_5824,In_945,In_1948);
nor U5825 (N_5825,In_392,In_2409);
or U5826 (N_5826,In_2122,In_958);
and U5827 (N_5827,In_396,In_1858);
or U5828 (N_5828,In_1731,In_283);
or U5829 (N_5829,In_138,In_2211);
nand U5830 (N_5830,In_1432,In_1134);
and U5831 (N_5831,In_1877,In_2193);
nor U5832 (N_5832,In_177,In_2413);
nor U5833 (N_5833,In_814,In_1405);
xor U5834 (N_5834,In_1754,In_1003);
xnor U5835 (N_5835,In_1916,In_1487);
nand U5836 (N_5836,In_1468,In_2430);
nand U5837 (N_5837,In_2136,In_1890);
and U5838 (N_5838,In_819,In_185);
nor U5839 (N_5839,In_1119,In_986);
and U5840 (N_5840,In_224,In_1478);
nor U5841 (N_5841,In_492,In_892);
or U5842 (N_5842,In_2313,In_921);
nor U5843 (N_5843,In_1916,In_778);
and U5844 (N_5844,In_1414,In_1881);
nand U5845 (N_5845,In_1235,In_723);
and U5846 (N_5846,In_2128,In_1373);
nor U5847 (N_5847,In_1948,In_1139);
or U5848 (N_5848,In_165,In_1377);
nor U5849 (N_5849,In_22,In_1597);
and U5850 (N_5850,In_205,In_2460);
xor U5851 (N_5851,In_1540,In_1532);
and U5852 (N_5852,In_1438,In_639);
nor U5853 (N_5853,In_1937,In_2423);
or U5854 (N_5854,In_926,In_2295);
nor U5855 (N_5855,In_1346,In_852);
nand U5856 (N_5856,In_580,In_1757);
nor U5857 (N_5857,In_2256,In_2440);
xor U5858 (N_5858,In_2296,In_1841);
nor U5859 (N_5859,In_971,In_1366);
or U5860 (N_5860,In_855,In_2161);
nand U5861 (N_5861,In_677,In_1041);
nor U5862 (N_5862,In_1927,In_1366);
nor U5863 (N_5863,In_1243,In_889);
nand U5864 (N_5864,In_1308,In_1499);
and U5865 (N_5865,In_500,In_571);
or U5866 (N_5866,In_58,In_1366);
nand U5867 (N_5867,In_2238,In_1735);
and U5868 (N_5868,In_1803,In_1622);
nor U5869 (N_5869,In_1271,In_720);
nor U5870 (N_5870,In_1534,In_2476);
nand U5871 (N_5871,In_2317,In_810);
nor U5872 (N_5872,In_177,In_1647);
or U5873 (N_5873,In_1560,In_1052);
nand U5874 (N_5874,In_758,In_2311);
nand U5875 (N_5875,In_447,In_91);
and U5876 (N_5876,In_1758,In_291);
nand U5877 (N_5877,In_1369,In_2234);
nor U5878 (N_5878,In_152,In_1340);
or U5879 (N_5879,In_1798,In_1794);
nand U5880 (N_5880,In_1712,In_1581);
or U5881 (N_5881,In_766,In_476);
or U5882 (N_5882,In_1820,In_2311);
nor U5883 (N_5883,In_1076,In_383);
nor U5884 (N_5884,In_1437,In_2338);
and U5885 (N_5885,In_1704,In_1787);
nand U5886 (N_5886,In_1227,In_1629);
nor U5887 (N_5887,In_615,In_376);
and U5888 (N_5888,In_145,In_1234);
nor U5889 (N_5889,In_151,In_2275);
or U5890 (N_5890,In_1157,In_522);
or U5891 (N_5891,In_977,In_345);
and U5892 (N_5892,In_952,In_2185);
nor U5893 (N_5893,In_1074,In_144);
and U5894 (N_5894,In_1724,In_355);
or U5895 (N_5895,In_2440,In_2023);
nand U5896 (N_5896,In_1790,In_1458);
or U5897 (N_5897,In_2213,In_370);
nand U5898 (N_5898,In_1962,In_96);
or U5899 (N_5899,In_921,In_1263);
nor U5900 (N_5900,In_2049,In_2333);
nand U5901 (N_5901,In_2489,In_2309);
or U5902 (N_5902,In_2458,In_2283);
and U5903 (N_5903,In_2397,In_938);
or U5904 (N_5904,In_1594,In_1188);
or U5905 (N_5905,In_36,In_291);
nor U5906 (N_5906,In_1445,In_309);
and U5907 (N_5907,In_2042,In_1662);
and U5908 (N_5908,In_857,In_883);
or U5909 (N_5909,In_1748,In_1313);
or U5910 (N_5910,In_1690,In_2458);
nand U5911 (N_5911,In_427,In_742);
xor U5912 (N_5912,In_1180,In_1735);
or U5913 (N_5913,In_1721,In_1201);
nor U5914 (N_5914,In_1368,In_1844);
nand U5915 (N_5915,In_1726,In_2264);
nor U5916 (N_5916,In_257,In_2310);
nor U5917 (N_5917,In_1504,In_453);
nand U5918 (N_5918,In_1565,In_1295);
nand U5919 (N_5919,In_174,In_769);
or U5920 (N_5920,In_1453,In_593);
nor U5921 (N_5921,In_1253,In_1923);
nor U5922 (N_5922,In_1337,In_1360);
and U5923 (N_5923,In_1084,In_769);
nor U5924 (N_5924,In_1933,In_1246);
xor U5925 (N_5925,In_820,In_1761);
xnor U5926 (N_5926,In_509,In_218);
or U5927 (N_5927,In_888,In_2178);
and U5928 (N_5928,In_2111,In_39);
and U5929 (N_5929,In_1423,In_1127);
nand U5930 (N_5930,In_1472,In_1730);
xnor U5931 (N_5931,In_2203,In_1989);
or U5932 (N_5932,In_1575,In_329);
or U5933 (N_5933,In_382,In_938);
nor U5934 (N_5934,In_703,In_339);
nand U5935 (N_5935,In_1722,In_714);
nor U5936 (N_5936,In_1191,In_167);
and U5937 (N_5937,In_589,In_63);
nor U5938 (N_5938,In_875,In_2044);
or U5939 (N_5939,In_1571,In_260);
nand U5940 (N_5940,In_1780,In_1591);
nand U5941 (N_5941,In_1708,In_920);
nand U5942 (N_5942,In_2255,In_2428);
nor U5943 (N_5943,In_492,In_1820);
nand U5944 (N_5944,In_1890,In_61);
nor U5945 (N_5945,In_1029,In_1201);
and U5946 (N_5946,In_1080,In_1948);
and U5947 (N_5947,In_83,In_2497);
and U5948 (N_5948,In_1136,In_2288);
nor U5949 (N_5949,In_1568,In_1338);
nand U5950 (N_5950,In_1806,In_960);
xnor U5951 (N_5951,In_1945,In_1195);
nand U5952 (N_5952,In_650,In_70);
and U5953 (N_5953,In_1440,In_1634);
nand U5954 (N_5954,In_2339,In_1461);
nand U5955 (N_5955,In_1233,In_305);
nand U5956 (N_5956,In_2291,In_779);
nor U5957 (N_5957,In_1745,In_1445);
nor U5958 (N_5958,In_1995,In_323);
nor U5959 (N_5959,In_505,In_1565);
and U5960 (N_5960,In_14,In_2059);
and U5961 (N_5961,In_1366,In_959);
xnor U5962 (N_5962,In_677,In_1532);
nor U5963 (N_5963,In_2286,In_1850);
xor U5964 (N_5964,In_282,In_1976);
or U5965 (N_5965,In_1296,In_1117);
nor U5966 (N_5966,In_2197,In_673);
or U5967 (N_5967,In_2035,In_1144);
or U5968 (N_5968,In_1631,In_1116);
nand U5969 (N_5969,In_1073,In_1018);
or U5970 (N_5970,In_1276,In_1337);
nand U5971 (N_5971,In_2239,In_654);
nand U5972 (N_5972,In_44,In_908);
nand U5973 (N_5973,In_229,In_515);
and U5974 (N_5974,In_1221,In_1943);
xnor U5975 (N_5975,In_1942,In_528);
and U5976 (N_5976,In_572,In_2353);
nand U5977 (N_5977,In_1373,In_1055);
xor U5978 (N_5978,In_966,In_214);
nor U5979 (N_5979,In_1996,In_1204);
nand U5980 (N_5980,In_833,In_165);
nor U5981 (N_5981,In_2195,In_1322);
or U5982 (N_5982,In_1531,In_284);
nand U5983 (N_5983,In_1087,In_19);
nand U5984 (N_5984,In_820,In_913);
or U5985 (N_5985,In_1674,In_1014);
nand U5986 (N_5986,In_1606,In_1981);
and U5987 (N_5987,In_855,In_270);
nand U5988 (N_5988,In_659,In_1604);
nand U5989 (N_5989,In_2430,In_584);
or U5990 (N_5990,In_1517,In_2054);
xnor U5991 (N_5991,In_2257,In_1256);
and U5992 (N_5992,In_862,In_1864);
or U5993 (N_5993,In_1243,In_1635);
xnor U5994 (N_5994,In_844,In_721);
xor U5995 (N_5995,In_1696,In_272);
nand U5996 (N_5996,In_847,In_2018);
nor U5997 (N_5997,In_1589,In_2335);
and U5998 (N_5998,In_356,In_797);
nand U5999 (N_5999,In_1571,In_1651);
nand U6000 (N_6000,In_2271,In_1186);
nor U6001 (N_6001,In_1880,In_1886);
nor U6002 (N_6002,In_2038,In_394);
and U6003 (N_6003,In_1894,In_266);
nor U6004 (N_6004,In_2410,In_593);
nor U6005 (N_6005,In_1884,In_2017);
nor U6006 (N_6006,In_505,In_1301);
nand U6007 (N_6007,In_611,In_2214);
and U6008 (N_6008,In_964,In_1186);
nor U6009 (N_6009,In_687,In_1205);
or U6010 (N_6010,In_1607,In_2059);
nand U6011 (N_6011,In_494,In_468);
nor U6012 (N_6012,In_1944,In_1685);
or U6013 (N_6013,In_1068,In_708);
nor U6014 (N_6014,In_1911,In_1342);
or U6015 (N_6015,In_2497,In_77);
or U6016 (N_6016,In_1360,In_2093);
nand U6017 (N_6017,In_2082,In_66);
nand U6018 (N_6018,In_2489,In_636);
and U6019 (N_6019,In_1529,In_119);
and U6020 (N_6020,In_1718,In_1927);
and U6021 (N_6021,In_1239,In_790);
or U6022 (N_6022,In_1146,In_2151);
nor U6023 (N_6023,In_2430,In_177);
nand U6024 (N_6024,In_1080,In_576);
nor U6025 (N_6025,In_962,In_451);
or U6026 (N_6026,In_1637,In_1625);
and U6027 (N_6027,In_2393,In_431);
nor U6028 (N_6028,In_748,In_2362);
nor U6029 (N_6029,In_233,In_1910);
or U6030 (N_6030,In_728,In_2407);
nand U6031 (N_6031,In_921,In_248);
or U6032 (N_6032,In_1789,In_2135);
nand U6033 (N_6033,In_1724,In_587);
or U6034 (N_6034,In_2447,In_1795);
or U6035 (N_6035,In_1909,In_2078);
nand U6036 (N_6036,In_1019,In_139);
and U6037 (N_6037,In_1440,In_1466);
nor U6038 (N_6038,In_1529,In_1374);
and U6039 (N_6039,In_257,In_1892);
xor U6040 (N_6040,In_329,In_1318);
and U6041 (N_6041,In_180,In_2312);
nand U6042 (N_6042,In_2316,In_2088);
nand U6043 (N_6043,In_1911,In_1857);
or U6044 (N_6044,In_882,In_542);
or U6045 (N_6045,In_684,In_697);
nand U6046 (N_6046,In_1913,In_1712);
and U6047 (N_6047,In_1534,In_2278);
or U6048 (N_6048,In_1042,In_672);
nand U6049 (N_6049,In_2294,In_5);
nand U6050 (N_6050,In_1476,In_907);
nand U6051 (N_6051,In_795,In_1108);
nand U6052 (N_6052,In_1320,In_10);
nor U6053 (N_6053,In_1035,In_2081);
nand U6054 (N_6054,In_860,In_806);
and U6055 (N_6055,In_717,In_2154);
and U6056 (N_6056,In_748,In_1973);
nand U6057 (N_6057,In_1026,In_2247);
nor U6058 (N_6058,In_294,In_1919);
nand U6059 (N_6059,In_1703,In_2208);
nand U6060 (N_6060,In_1314,In_361);
nand U6061 (N_6061,In_2443,In_820);
xor U6062 (N_6062,In_2190,In_599);
and U6063 (N_6063,In_821,In_930);
xor U6064 (N_6064,In_2315,In_472);
nand U6065 (N_6065,In_214,In_79);
or U6066 (N_6066,In_102,In_2077);
xnor U6067 (N_6067,In_639,In_433);
nand U6068 (N_6068,In_1183,In_972);
or U6069 (N_6069,In_1072,In_2470);
nor U6070 (N_6070,In_1935,In_2349);
nand U6071 (N_6071,In_1621,In_2222);
xor U6072 (N_6072,In_1201,In_961);
nand U6073 (N_6073,In_398,In_1712);
nor U6074 (N_6074,In_1301,In_2374);
or U6075 (N_6075,In_1725,In_972);
and U6076 (N_6076,In_1681,In_1669);
or U6077 (N_6077,In_2484,In_1556);
or U6078 (N_6078,In_322,In_2228);
or U6079 (N_6079,In_27,In_1402);
and U6080 (N_6080,In_1173,In_491);
and U6081 (N_6081,In_2074,In_1176);
or U6082 (N_6082,In_1051,In_1213);
nor U6083 (N_6083,In_46,In_544);
nand U6084 (N_6084,In_1815,In_611);
or U6085 (N_6085,In_927,In_1404);
and U6086 (N_6086,In_636,In_51);
and U6087 (N_6087,In_1123,In_892);
and U6088 (N_6088,In_615,In_1573);
and U6089 (N_6089,In_1309,In_977);
nor U6090 (N_6090,In_2415,In_636);
nor U6091 (N_6091,In_1716,In_378);
or U6092 (N_6092,In_531,In_915);
nor U6093 (N_6093,In_2293,In_1509);
or U6094 (N_6094,In_1096,In_2249);
nand U6095 (N_6095,In_1215,In_215);
nor U6096 (N_6096,In_1257,In_1181);
nand U6097 (N_6097,In_327,In_1676);
nor U6098 (N_6098,In_2045,In_68);
nor U6099 (N_6099,In_714,In_666);
and U6100 (N_6100,In_1626,In_1143);
nand U6101 (N_6101,In_1358,In_2379);
nor U6102 (N_6102,In_1395,In_2439);
or U6103 (N_6103,In_1861,In_1932);
xor U6104 (N_6104,In_282,In_1712);
nor U6105 (N_6105,In_2231,In_1714);
nand U6106 (N_6106,In_2279,In_1905);
nor U6107 (N_6107,In_273,In_2152);
xor U6108 (N_6108,In_624,In_1384);
xnor U6109 (N_6109,In_1494,In_1275);
nor U6110 (N_6110,In_2160,In_1847);
and U6111 (N_6111,In_1850,In_1368);
or U6112 (N_6112,In_837,In_890);
nand U6113 (N_6113,In_2344,In_1208);
and U6114 (N_6114,In_170,In_464);
nor U6115 (N_6115,In_433,In_1307);
or U6116 (N_6116,In_1174,In_424);
and U6117 (N_6117,In_1509,In_44);
and U6118 (N_6118,In_875,In_676);
nand U6119 (N_6119,In_1602,In_2264);
or U6120 (N_6120,In_1018,In_143);
xnor U6121 (N_6121,In_1086,In_1548);
nand U6122 (N_6122,In_1227,In_2090);
nand U6123 (N_6123,In_2370,In_1652);
nand U6124 (N_6124,In_2111,In_2033);
or U6125 (N_6125,In_1416,In_1705);
nor U6126 (N_6126,In_251,In_1728);
or U6127 (N_6127,In_1340,In_1685);
nand U6128 (N_6128,In_17,In_403);
and U6129 (N_6129,In_2079,In_2336);
nand U6130 (N_6130,In_764,In_318);
nand U6131 (N_6131,In_2462,In_702);
xnor U6132 (N_6132,In_1760,In_961);
nor U6133 (N_6133,In_1816,In_1516);
nor U6134 (N_6134,In_596,In_1975);
nor U6135 (N_6135,In_100,In_1669);
and U6136 (N_6136,In_91,In_1777);
nand U6137 (N_6137,In_2274,In_467);
nor U6138 (N_6138,In_1516,In_1915);
or U6139 (N_6139,In_258,In_1410);
nand U6140 (N_6140,In_2024,In_1938);
nand U6141 (N_6141,In_2142,In_893);
nor U6142 (N_6142,In_1478,In_2112);
or U6143 (N_6143,In_1877,In_531);
nor U6144 (N_6144,In_1929,In_1339);
nor U6145 (N_6145,In_554,In_1095);
nand U6146 (N_6146,In_1399,In_777);
nor U6147 (N_6147,In_247,In_890);
nor U6148 (N_6148,In_287,In_2138);
nor U6149 (N_6149,In_727,In_956);
nand U6150 (N_6150,In_309,In_2053);
or U6151 (N_6151,In_1302,In_46);
or U6152 (N_6152,In_320,In_1919);
or U6153 (N_6153,In_2423,In_469);
or U6154 (N_6154,In_1607,In_141);
or U6155 (N_6155,In_800,In_2287);
or U6156 (N_6156,In_900,In_1044);
nor U6157 (N_6157,In_1925,In_869);
and U6158 (N_6158,In_90,In_658);
or U6159 (N_6159,In_1487,In_1361);
nand U6160 (N_6160,In_1539,In_2232);
xor U6161 (N_6161,In_1250,In_1442);
or U6162 (N_6162,In_1288,In_2196);
and U6163 (N_6163,In_489,In_664);
and U6164 (N_6164,In_595,In_633);
nand U6165 (N_6165,In_800,In_2073);
or U6166 (N_6166,In_2466,In_1879);
nand U6167 (N_6167,In_2110,In_0);
nand U6168 (N_6168,In_776,In_2376);
nand U6169 (N_6169,In_1712,In_513);
nor U6170 (N_6170,In_1813,In_1999);
nor U6171 (N_6171,In_945,In_2384);
or U6172 (N_6172,In_519,In_2096);
nor U6173 (N_6173,In_2352,In_551);
nor U6174 (N_6174,In_1906,In_1509);
or U6175 (N_6175,In_2356,In_1664);
and U6176 (N_6176,In_814,In_494);
and U6177 (N_6177,In_1038,In_1265);
or U6178 (N_6178,In_526,In_2302);
and U6179 (N_6179,In_541,In_1303);
or U6180 (N_6180,In_531,In_1520);
and U6181 (N_6181,In_1094,In_2346);
xor U6182 (N_6182,In_568,In_504);
nand U6183 (N_6183,In_1319,In_1873);
nor U6184 (N_6184,In_252,In_2373);
nor U6185 (N_6185,In_1860,In_109);
xor U6186 (N_6186,In_1038,In_159);
nor U6187 (N_6187,In_1284,In_1383);
and U6188 (N_6188,In_1294,In_2454);
nor U6189 (N_6189,In_2410,In_2449);
or U6190 (N_6190,In_406,In_1958);
nand U6191 (N_6191,In_119,In_1261);
and U6192 (N_6192,In_2408,In_1981);
nand U6193 (N_6193,In_1935,In_259);
and U6194 (N_6194,In_1116,In_231);
nand U6195 (N_6195,In_1776,In_2380);
and U6196 (N_6196,In_2124,In_616);
or U6197 (N_6197,In_2411,In_903);
nand U6198 (N_6198,In_1817,In_1263);
and U6199 (N_6199,In_1347,In_320);
and U6200 (N_6200,In_950,In_1141);
and U6201 (N_6201,In_2381,In_1130);
nor U6202 (N_6202,In_1787,In_2176);
nand U6203 (N_6203,In_954,In_506);
nand U6204 (N_6204,In_1666,In_309);
and U6205 (N_6205,In_2301,In_756);
or U6206 (N_6206,In_328,In_1749);
xnor U6207 (N_6207,In_411,In_526);
nor U6208 (N_6208,In_299,In_1172);
nor U6209 (N_6209,In_2417,In_184);
and U6210 (N_6210,In_1695,In_550);
and U6211 (N_6211,In_772,In_657);
xor U6212 (N_6212,In_427,In_1967);
nor U6213 (N_6213,In_1774,In_57);
or U6214 (N_6214,In_304,In_2161);
or U6215 (N_6215,In_1502,In_282);
or U6216 (N_6216,In_2076,In_2293);
nor U6217 (N_6217,In_856,In_465);
or U6218 (N_6218,In_2033,In_1530);
and U6219 (N_6219,In_972,In_617);
and U6220 (N_6220,In_2182,In_415);
or U6221 (N_6221,In_1182,In_1035);
and U6222 (N_6222,In_180,In_84);
nand U6223 (N_6223,In_140,In_1719);
nor U6224 (N_6224,In_1612,In_1676);
and U6225 (N_6225,In_2294,In_1514);
or U6226 (N_6226,In_400,In_750);
xor U6227 (N_6227,In_92,In_2235);
nor U6228 (N_6228,In_2458,In_1837);
nor U6229 (N_6229,In_2092,In_1953);
xnor U6230 (N_6230,In_1166,In_534);
nor U6231 (N_6231,In_1324,In_959);
nor U6232 (N_6232,In_1334,In_1470);
and U6233 (N_6233,In_1865,In_1147);
and U6234 (N_6234,In_2020,In_2154);
and U6235 (N_6235,In_708,In_2101);
nand U6236 (N_6236,In_1304,In_2486);
or U6237 (N_6237,In_392,In_847);
or U6238 (N_6238,In_1075,In_706);
or U6239 (N_6239,In_1335,In_1215);
xor U6240 (N_6240,In_1470,In_1183);
or U6241 (N_6241,In_466,In_410);
xor U6242 (N_6242,In_2179,In_1135);
and U6243 (N_6243,In_1459,In_174);
or U6244 (N_6244,In_1784,In_1847);
and U6245 (N_6245,In_301,In_2341);
and U6246 (N_6246,In_1853,In_901);
xor U6247 (N_6247,In_1698,In_565);
and U6248 (N_6248,In_576,In_1615);
or U6249 (N_6249,In_585,In_1412);
nor U6250 (N_6250,N_3333,N_1632);
and U6251 (N_6251,N_3357,N_419);
and U6252 (N_6252,N_4570,N_246);
nand U6253 (N_6253,N_3563,N_2942);
nand U6254 (N_6254,N_4874,N_3525);
or U6255 (N_6255,N_4562,N_4516);
and U6256 (N_6256,N_1024,N_5074);
and U6257 (N_6257,N_3721,N_2989);
nor U6258 (N_6258,N_5340,N_3531);
and U6259 (N_6259,N_5,N_3875);
or U6260 (N_6260,N_230,N_2781);
xor U6261 (N_6261,N_64,N_2537);
and U6262 (N_6262,N_1289,N_3025);
xor U6263 (N_6263,N_259,N_291);
and U6264 (N_6264,N_956,N_1190);
nor U6265 (N_6265,N_3626,N_1777);
and U6266 (N_6266,N_5754,N_5815);
and U6267 (N_6267,N_616,N_2292);
and U6268 (N_6268,N_5579,N_3271);
nor U6269 (N_6269,N_4277,N_5686);
and U6270 (N_6270,N_3782,N_2107);
nand U6271 (N_6271,N_2055,N_1172);
nor U6272 (N_6272,N_2843,N_2608);
nor U6273 (N_6273,N_1713,N_3887);
nor U6274 (N_6274,N_2098,N_2409);
nand U6275 (N_6275,N_1443,N_1905);
and U6276 (N_6276,N_3308,N_312);
nor U6277 (N_6277,N_2952,N_382);
and U6278 (N_6278,N_3767,N_3809);
nor U6279 (N_6279,N_100,N_617);
and U6280 (N_6280,N_3344,N_2842);
and U6281 (N_6281,N_5491,N_2184);
and U6282 (N_6282,N_2158,N_5442);
nand U6283 (N_6283,N_5293,N_5228);
nand U6284 (N_6284,N_86,N_592);
and U6285 (N_6285,N_354,N_5605);
nand U6286 (N_6286,N_6239,N_5114);
and U6287 (N_6287,N_1245,N_1394);
nor U6288 (N_6288,N_1376,N_1506);
or U6289 (N_6289,N_547,N_4717);
and U6290 (N_6290,N_5997,N_334);
and U6291 (N_6291,N_137,N_3494);
or U6292 (N_6292,N_4532,N_3734);
and U6293 (N_6293,N_2466,N_5709);
and U6294 (N_6294,N_448,N_4306);
nor U6295 (N_6295,N_5985,N_2762);
nor U6296 (N_6296,N_1765,N_646);
nand U6297 (N_6297,N_987,N_5351);
nor U6298 (N_6298,N_871,N_5971);
nor U6299 (N_6299,N_872,N_2848);
nor U6300 (N_6300,N_2511,N_1247);
nand U6301 (N_6301,N_2986,N_5071);
nor U6302 (N_6302,N_5708,N_5390);
nor U6303 (N_6303,N_2396,N_953);
and U6304 (N_6304,N_4037,N_4703);
and U6305 (N_6305,N_633,N_2565);
xnor U6306 (N_6306,N_1988,N_2063);
nor U6307 (N_6307,N_4273,N_55);
nor U6308 (N_6308,N_974,N_301);
or U6309 (N_6309,N_895,N_545);
nand U6310 (N_6310,N_1037,N_1234);
nor U6311 (N_6311,N_6136,N_356);
or U6312 (N_6312,N_5669,N_5067);
nor U6313 (N_6313,N_1427,N_5732);
nor U6314 (N_6314,N_695,N_5848);
nand U6315 (N_6315,N_94,N_3003);
nand U6316 (N_6316,N_5799,N_1388);
and U6317 (N_6317,N_2241,N_368);
xor U6318 (N_6318,N_1865,N_1271);
nor U6319 (N_6319,N_5559,N_5464);
nand U6320 (N_6320,N_1815,N_3437);
nor U6321 (N_6321,N_2891,N_4585);
nand U6322 (N_6322,N_1498,N_846);
nand U6323 (N_6323,N_4375,N_1950);
nand U6324 (N_6324,N_3099,N_1744);
or U6325 (N_6325,N_4961,N_387);
nand U6326 (N_6326,N_3665,N_5952);
nand U6327 (N_6327,N_1346,N_6161);
and U6328 (N_6328,N_1739,N_6044);
xor U6329 (N_6329,N_4088,N_4328);
xor U6330 (N_6330,N_188,N_678);
nor U6331 (N_6331,N_1682,N_6);
or U6332 (N_6332,N_3805,N_3114);
and U6333 (N_6333,N_1468,N_2317);
nand U6334 (N_6334,N_746,N_3222);
and U6335 (N_6335,N_5253,N_4108);
xor U6336 (N_6336,N_4063,N_1099);
and U6337 (N_6337,N_2517,N_1292);
nor U6338 (N_6338,N_2044,N_4225);
or U6339 (N_6339,N_3266,N_4429);
nor U6340 (N_6340,N_1729,N_5950);
nand U6341 (N_6341,N_4545,N_797);
and U6342 (N_6342,N_2138,N_5480);
or U6343 (N_6343,N_1614,N_823);
and U6344 (N_6344,N_763,N_5958);
or U6345 (N_6345,N_2878,N_3218);
and U6346 (N_6346,N_5587,N_5783);
and U6347 (N_6347,N_287,N_3162);
and U6348 (N_6348,N_2926,N_5531);
nand U6349 (N_6349,N_3440,N_5793);
and U6350 (N_6350,N_4718,N_1731);
and U6351 (N_6351,N_3658,N_4907);
and U6352 (N_6352,N_3815,N_299);
nand U6353 (N_6353,N_1568,N_3368);
nor U6354 (N_6354,N_4269,N_1360);
or U6355 (N_6355,N_4126,N_5303);
and U6356 (N_6356,N_2935,N_3459);
or U6357 (N_6357,N_4606,N_3486);
xor U6358 (N_6358,N_3965,N_4481);
nand U6359 (N_6359,N_3178,N_4136);
nand U6360 (N_6360,N_6120,N_6143);
or U6361 (N_6361,N_3256,N_572);
and U6362 (N_6362,N_5688,N_5248);
nand U6363 (N_6363,N_4480,N_6058);
nor U6364 (N_6364,N_6125,N_3108);
or U6365 (N_6365,N_4355,N_3462);
nor U6366 (N_6366,N_2258,N_983);
or U6367 (N_6367,N_5513,N_3680);
and U6368 (N_6368,N_4927,N_2687);
or U6369 (N_6369,N_2563,N_5737);
or U6370 (N_6370,N_4503,N_2137);
and U6371 (N_6371,N_812,N_3435);
and U6372 (N_6372,N_5924,N_5244);
or U6373 (N_6373,N_3781,N_4173);
and U6374 (N_6374,N_3931,N_3628);
nand U6375 (N_6375,N_5199,N_1470);
nor U6376 (N_6376,N_6153,N_1314);
nand U6377 (N_6377,N_2615,N_4471);
or U6378 (N_6378,N_5837,N_5250);
nor U6379 (N_6379,N_1939,N_5112);
nand U6380 (N_6380,N_4762,N_526);
nor U6381 (N_6381,N_6211,N_3766);
xnor U6382 (N_6382,N_6027,N_4816);
nor U6383 (N_6383,N_4864,N_1983);
and U6384 (N_6384,N_566,N_3436);
nand U6385 (N_6385,N_3501,N_3712);
nand U6386 (N_6386,N_1123,N_5054);
nor U6387 (N_6387,N_5213,N_691);
and U6388 (N_6388,N_4695,N_2057);
nand U6389 (N_6389,N_6182,N_2358);
nor U6390 (N_6390,N_5653,N_1280);
or U6391 (N_6391,N_6004,N_4906);
nand U6392 (N_6392,N_1871,N_2080);
and U6393 (N_6393,N_3950,N_5400);
xnor U6394 (N_6394,N_1011,N_5164);
nand U6395 (N_6395,N_370,N_2304);
and U6396 (N_6396,N_194,N_5595);
nand U6397 (N_6397,N_3112,N_5874);
or U6398 (N_6398,N_11,N_2778);
and U6399 (N_6399,N_2232,N_3465);
or U6400 (N_6400,N_5887,N_1825);
nor U6401 (N_6401,N_4497,N_4008);
nand U6402 (N_6402,N_2357,N_1134);
xor U6403 (N_6403,N_5841,N_5329);
nand U6404 (N_6404,N_5052,N_5994);
or U6405 (N_6405,N_2974,N_2593);
and U6406 (N_6406,N_935,N_2779);
nand U6407 (N_6407,N_6199,N_151);
nand U6408 (N_6408,N_982,N_5109);
or U6409 (N_6409,N_4604,N_4148);
and U6410 (N_6410,N_1358,N_508);
nand U6411 (N_6411,N_3239,N_331);
nor U6412 (N_6412,N_770,N_4209);
xor U6413 (N_6413,N_568,N_4401);
or U6414 (N_6414,N_3879,N_320);
or U6415 (N_6415,N_5483,N_965);
nor U6416 (N_6416,N_5201,N_283);
xnor U6417 (N_6417,N_4383,N_1081);
and U6418 (N_6418,N_5909,N_5530);
nor U6419 (N_6419,N_1406,N_3954);
nor U6420 (N_6420,N_1933,N_1879);
nor U6421 (N_6421,N_5714,N_5585);
nand U6422 (N_6422,N_3476,N_1993);
and U6423 (N_6423,N_5582,N_5586);
nor U6424 (N_6424,N_4094,N_5945);
xnor U6425 (N_6425,N_3483,N_1956);
xnor U6426 (N_6426,N_3696,N_1778);
and U6427 (N_6427,N_2909,N_2074);
and U6428 (N_6428,N_4915,N_2718);
and U6429 (N_6429,N_5078,N_1447);
nand U6430 (N_6430,N_4826,N_1162);
or U6431 (N_6431,N_2135,N_5493);
and U6432 (N_6432,N_1251,N_1603);
xnor U6433 (N_6433,N_3659,N_2210);
and U6434 (N_6434,N_4664,N_3104);
nor U6435 (N_6435,N_5238,N_2289);
nor U6436 (N_6436,N_2908,N_2649);
xor U6437 (N_6437,N_5743,N_1429);
nor U6438 (N_6438,N_4655,N_648);
and U6439 (N_6439,N_4614,N_2716);
or U6440 (N_6440,N_5193,N_5439);
nor U6441 (N_6441,N_3754,N_4992);
nand U6442 (N_6442,N_5929,N_4246);
nor U6443 (N_6443,N_5728,N_1357);
nand U6444 (N_6444,N_4200,N_5296);
nor U6445 (N_6445,N_5256,N_2523);
and U6446 (N_6446,N_2420,N_4395);
and U6447 (N_6447,N_3513,N_3845);
nand U6448 (N_6448,N_4778,N_4680);
xor U6449 (N_6449,N_3516,N_4847);
xnor U6450 (N_6450,N_5580,N_2798);
and U6451 (N_6451,N_3229,N_1003);
or U6452 (N_6452,N_5227,N_6001);
nand U6453 (N_6453,N_4476,N_4607);
and U6454 (N_6454,N_3923,N_6207);
xnor U6455 (N_6455,N_1069,N_1296);
xor U6456 (N_6456,N_4842,N_4353);
nor U6457 (N_6457,N_1093,N_950);
nor U6458 (N_6458,N_3894,N_2949);
nor U6459 (N_6459,N_5086,N_4956);
nor U6460 (N_6460,N_2859,N_2225);
or U6461 (N_6461,N_5735,N_3038);
and U6462 (N_6462,N_4917,N_681);
nand U6463 (N_6463,N_1244,N_2309);
nand U6464 (N_6464,N_1350,N_1593);
nand U6465 (N_6465,N_4160,N_2215);
xor U6466 (N_6466,N_1555,N_6247);
nand U6467 (N_6467,N_5640,N_1638);
nand U6468 (N_6468,N_4899,N_3360);
or U6469 (N_6469,N_1091,N_2657);
nand U6470 (N_6470,N_1088,N_4810);
nor U6471 (N_6471,N_3846,N_3370);
or U6472 (N_6472,N_1762,N_4560);
or U6473 (N_6473,N_6010,N_3936);
nand U6474 (N_6474,N_3687,N_225);
nand U6475 (N_6475,N_3913,N_2922);
or U6476 (N_6476,N_3461,N_5385);
or U6477 (N_6477,N_4467,N_1868);
nor U6478 (N_6478,N_655,N_3005);
nor U6479 (N_6479,N_3996,N_3136);
and U6480 (N_6480,N_3132,N_4449);
nor U6481 (N_6481,N_6138,N_3568);
and U6482 (N_6482,N_4393,N_2693);
and U6483 (N_6483,N_3532,N_2482);
or U6484 (N_6484,N_2012,N_4100);
nand U6485 (N_6485,N_1587,N_5477);
and U6486 (N_6486,N_3201,N_1471);
and U6487 (N_6487,N_3185,N_3830);
or U6488 (N_6488,N_3241,N_1813);
xor U6489 (N_6489,N_70,N_5875);
nand U6490 (N_6490,N_89,N_517);
or U6491 (N_6491,N_3240,N_2016);
nor U6492 (N_6492,N_3983,N_3883);
nor U6493 (N_6493,N_5853,N_5654);
nand U6494 (N_6494,N_4642,N_4775);
nand U6495 (N_6495,N_1742,N_2486);
or U6496 (N_6496,N_1161,N_5687);
nor U6497 (N_6497,N_2576,N_2653);
and U6498 (N_6498,N_4889,N_1237);
or U6499 (N_6499,N_2103,N_3200);
and U6500 (N_6500,N_338,N_604);
nor U6501 (N_6501,N_5149,N_5287);
and U6502 (N_6502,N_5167,N_281);
nand U6503 (N_6503,N_2515,N_3834);
or U6504 (N_6504,N_2220,N_5581);
nor U6505 (N_6505,N_3073,N_2166);
xor U6506 (N_6506,N_415,N_1521);
nand U6507 (N_6507,N_5346,N_5890);
nor U6508 (N_6508,N_4167,N_5065);
nor U6509 (N_6509,N_832,N_5902);
or U6510 (N_6510,N_538,N_2586);
and U6511 (N_6511,N_4682,N_6062);
nor U6512 (N_6512,N_5370,N_6180);
nand U6513 (N_6513,N_4065,N_1979);
or U6514 (N_6514,N_2129,N_1628);
or U6515 (N_6515,N_1483,N_3219);
and U6516 (N_6516,N_1408,N_6146);
xnor U6517 (N_6517,N_63,N_1030);
nor U6518 (N_6518,N_3036,N_4032);
nand U6519 (N_6519,N_584,N_6039);
nand U6520 (N_6520,N_4257,N_4519);
or U6521 (N_6521,N_5048,N_3943);
or U6522 (N_6522,N_1610,N_927);
and U6523 (N_6523,N_4352,N_3776);
nand U6524 (N_6524,N_5174,N_2697);
or U6525 (N_6525,N_1583,N_4153);
or U6526 (N_6526,N_979,N_5658);
xnor U6527 (N_6527,N_4568,N_3994);
and U6528 (N_6528,N_4112,N_2816);
xnor U6529 (N_6529,N_2690,N_3796);
xor U6530 (N_6530,N_4530,N_5805);
or U6531 (N_6531,N_5214,N_2282);
or U6532 (N_6532,N_2709,N_6244);
or U6533 (N_6533,N_469,N_454);
nand U6534 (N_6534,N_1757,N_4948);
nand U6535 (N_6535,N_2679,N_2964);
or U6536 (N_6536,N_571,N_4182);
nor U6537 (N_6537,N_5009,N_790);
and U6538 (N_6538,N_1195,N_2046);
nor U6539 (N_6539,N_436,N_1362);
nor U6540 (N_6540,N_6158,N_565);
and U6541 (N_6541,N_4223,N_3473);
or U6542 (N_6542,N_625,N_4806);
nand U6543 (N_6543,N_4260,N_2068);
or U6544 (N_6544,N_4749,N_837);
and U6545 (N_6545,N_5018,N_424);
nand U6546 (N_6546,N_736,N_2400);
and U6547 (N_6547,N_4598,N_643);
or U6548 (N_6548,N_1936,N_29);
xor U6549 (N_6549,N_4990,N_3422);
nand U6550 (N_6550,N_3737,N_6059);
or U6551 (N_6551,N_208,N_980);
or U6552 (N_6552,N_1708,N_4211);
nor U6553 (N_6553,N_3300,N_975);
or U6554 (N_6554,N_6097,N_4483);
or U6555 (N_6555,N_2815,N_4374);
xor U6556 (N_6556,N_4969,N_4567);
xor U6557 (N_6557,N_4207,N_561);
or U6558 (N_6558,N_4895,N_730);
or U6559 (N_6559,N_1964,N_205);
or U6560 (N_6560,N_1163,N_1320);
nand U6561 (N_6561,N_4397,N_1110);
nand U6562 (N_6562,N_1844,N_5484);
nor U6563 (N_6563,N_674,N_4796);
nand U6564 (N_6564,N_5552,N_986);
nor U6565 (N_6565,N_1927,N_5755);
and U6566 (N_6566,N_2316,N_5410);
or U6567 (N_6567,N_343,N_5964);
or U6568 (N_6568,N_3210,N_2619);
nor U6569 (N_6569,N_1353,N_1820);
nand U6570 (N_6570,N_2665,N_108);
and U6571 (N_6571,N_1399,N_5892);
nand U6572 (N_6572,N_2470,N_1229);
and U6573 (N_6573,N_3281,N_1496);
or U6574 (N_6574,N_6238,N_4671);
and U6575 (N_6575,N_6155,N_1106);
nor U6576 (N_6576,N_2950,N_1193);
nand U6577 (N_6577,N_4880,N_1938);
and U6578 (N_6578,N_1660,N_3111);
nand U6579 (N_6579,N_1442,N_1227);
nor U6580 (N_6580,N_5272,N_6071);
nor U6581 (N_6581,N_756,N_1196);
xor U6582 (N_6582,N_4600,N_3230);
and U6583 (N_6583,N_5431,N_3928);
nand U6584 (N_6584,N_4785,N_5547);
or U6585 (N_6585,N_5839,N_5759);
and U6586 (N_6586,N_641,N_5860);
nand U6587 (N_6587,N_2946,N_1248);
nor U6588 (N_6588,N_3014,N_5497);
and U6589 (N_6589,N_704,N_2799);
or U6590 (N_6590,N_391,N_4364);
nor U6591 (N_6591,N_4935,N_1788);
xor U6592 (N_6592,N_3352,N_5621);
nor U6593 (N_6593,N_731,N_969);
or U6594 (N_6594,N_866,N_4168);
and U6595 (N_6595,N_1896,N_236);
and U6596 (N_6596,N_3867,N_585);
xor U6597 (N_6597,N_1543,N_803);
nand U6598 (N_6598,N_4085,N_4723);
xnor U6599 (N_6599,N_5515,N_1410);
and U6600 (N_6600,N_3481,N_4737);
nor U6601 (N_6601,N_2100,N_5498);
and U6602 (N_6602,N_810,N_4406);
or U6603 (N_6603,N_819,N_1274);
and U6604 (N_6604,N_2978,N_1662);
nor U6605 (N_6605,N_3706,N_420);
nand U6606 (N_6606,N_3749,N_2027);
and U6607 (N_6607,N_2469,N_1434);
nor U6608 (N_6608,N_6241,N_5844);
and U6609 (N_6609,N_6085,N_4314);
nor U6610 (N_6610,N_680,N_2948);
nor U6611 (N_6611,N_1335,N_3000);
nor U6612 (N_6612,N_2505,N_4287);
or U6613 (N_6613,N_773,N_180);
xor U6614 (N_6614,N_3446,N_2992);
nand U6615 (N_6615,N_712,N_2773);
nand U6616 (N_6616,N_5539,N_3947);
or U6617 (N_6617,N_5867,N_2402);
and U6618 (N_6618,N_5866,N_3068);
and U6619 (N_6619,N_1887,N_5718);
nor U6620 (N_6620,N_2536,N_2668);
and U6621 (N_6621,N_5251,N_2095);
nand U6622 (N_6622,N_3748,N_5151);
nand U6623 (N_6623,N_166,N_2895);
nand U6624 (N_6624,N_2970,N_1535);
nand U6625 (N_6625,N_1685,N_906);
or U6626 (N_6626,N_2390,N_3756);
and U6627 (N_6627,N_1574,N_4934);
or U6628 (N_6628,N_1317,N_6178);
and U6629 (N_6629,N_1854,N_3052);
and U6630 (N_6630,N_2460,N_562);
xor U6631 (N_6631,N_1822,N_6185);
and U6632 (N_6632,N_4902,N_5494);
nand U6633 (N_6633,N_2367,N_1942);
nor U6634 (N_6634,N_3499,N_239);
or U6635 (N_6635,N_1281,N_4981);
nor U6636 (N_6636,N_5241,N_824);
and U6637 (N_6637,N_181,N_335);
nor U6638 (N_6638,N_2056,N_3678);
nand U6639 (N_6639,N_5594,N_4028);
xor U6640 (N_6640,N_4804,N_3306);
nand U6641 (N_6641,N_1780,N_4477);
and U6642 (N_6642,N_5341,N_4676);
nor U6643 (N_6643,N_711,N_4311);
and U6644 (N_6644,N_4665,N_3);
nor U6645 (N_6645,N_5936,N_1425);
nor U6646 (N_6646,N_5758,N_1381);
and U6647 (N_6647,N_2202,N_3179);
or U6648 (N_6648,N_6056,N_1990);
nor U6649 (N_6649,N_4910,N_5920);
and U6650 (N_6650,N_2194,N_5116);
nand U6651 (N_6651,N_1035,N_2876);
and U6652 (N_6652,N_1748,N_5673);
nand U6653 (N_6653,N_2928,N_1803);
nand U6654 (N_6654,N_5624,N_3282);
and U6655 (N_6655,N_1930,N_5428);
nor U6656 (N_6656,N_2575,N_5968);
nor U6657 (N_6657,N_2662,N_2719);
and U6658 (N_6658,N_1667,N_5292);
nor U6659 (N_6659,N_5268,N_4528);
and U6660 (N_6660,N_4978,N_1456);
and U6661 (N_6661,N_2589,N_5571);
nand U6662 (N_6662,N_3757,N_3371);
xor U6663 (N_6663,N_3438,N_4115);
or U6664 (N_6664,N_3597,N_2967);
or U6665 (N_6665,N_1951,N_4904);
nor U6666 (N_6666,N_2113,N_3668);
or U6667 (N_6667,N_3021,N_4840);
or U6668 (N_6668,N_2875,N_3193);
and U6669 (N_6669,N_4292,N_595);
xor U6670 (N_6670,N_3810,N_1111);
nand U6671 (N_6671,N_6160,N_3573);
nor U6672 (N_6672,N_388,N_2899);
nor U6673 (N_6673,N_5795,N_1678);
and U6674 (N_6674,N_3558,N_802);
and U6675 (N_6675,N_6157,N_556);
and U6676 (N_6676,N_4959,N_3471);
and U6677 (N_6677,N_397,N_5443);
or U6678 (N_6678,N_2483,N_5265);
or U6679 (N_6679,N_3751,N_2014);
nor U6680 (N_6680,N_613,N_978);
nand U6681 (N_6681,N_541,N_3492);
or U6682 (N_6682,N_4815,N_5807);
or U6683 (N_6683,N_332,N_2097);
or U6684 (N_6684,N_2297,N_4356);
or U6685 (N_6685,N_411,N_549);
and U6686 (N_6686,N_3414,N_4463);
and U6687 (N_6687,N_2213,N_2578);
xor U6688 (N_6688,N_4290,N_3470);
and U6689 (N_6689,N_5257,N_2508);
nand U6690 (N_6690,N_2939,N_3528);
nand U6691 (N_6691,N_3717,N_1795);
nand U6692 (N_6692,N_37,N_1634);
nor U6693 (N_6693,N_6137,N_6204);
or U6694 (N_6694,N_2287,N_2963);
nor U6695 (N_6695,N_5118,N_2509);
or U6696 (N_6696,N_1857,N_23);
xnor U6697 (N_6697,N_3321,N_6017);
and U6698 (N_6698,N_3944,N_2853);
nand U6699 (N_6699,N_3130,N_3017);
or U6700 (N_6700,N_5229,N_3889);
nand U6701 (N_6701,N_631,N_5925);
nand U6702 (N_6702,N_536,N_3263);
or U6703 (N_6703,N_1580,N_5589);
xor U6704 (N_6704,N_2245,N_2273);
and U6705 (N_6705,N_203,N_190);
nand U6706 (N_6706,N_1031,N_1570);
and U6707 (N_6707,N_818,N_1530);
xor U6708 (N_6708,N_2330,N_2994);
and U6709 (N_6709,N_4087,N_3579);
or U6710 (N_6710,N_1351,N_1596);
or U6711 (N_6711,N_3366,N_1661);
and U6712 (N_6712,N_4145,N_5665);
and U6713 (N_6713,N_4174,N_6148);
or U6714 (N_6714,N_5626,N_2091);
or U6715 (N_6715,N_1805,N_6167);
xor U6716 (N_6716,N_172,N_1378);
and U6717 (N_6717,N_3684,N_2119);
nor U6718 (N_6718,N_564,N_4933);
and U6719 (N_6719,N_2981,N_1264);
or U6720 (N_6720,N_4911,N_5093);
and U6721 (N_6721,N_3839,N_4186);
nor U6722 (N_6722,N_5017,N_6090);
or U6723 (N_6723,N_1716,N_609);
nor U6724 (N_6724,N_1191,N_5328);
or U6725 (N_6725,N_5830,N_4621);
or U6726 (N_6726,N_3246,N_6249);
xnor U6727 (N_6727,N_743,N_3999);
xnor U6728 (N_6728,N_899,N_2759);
nor U6729 (N_6729,N_2295,N_4946);
and U6730 (N_6730,N_675,N_4862);
nand U6731 (N_6731,N_660,N_115);
nor U6732 (N_6732,N_2011,N_1454);
nand U6733 (N_6733,N_5157,N_535);
nand U6734 (N_6734,N_1148,N_492);
xnor U6735 (N_6735,N_3848,N_3800);
nand U6736 (N_6736,N_2771,N_5309);
and U6737 (N_6737,N_235,N_1474);
or U6738 (N_6738,N_1453,N_1119);
xor U6739 (N_6739,N_4971,N_5264);
or U6740 (N_6740,N_2742,N_4007);
and U6741 (N_6741,N_1866,N_3864);
or U6742 (N_6742,N_881,N_4993);
nand U6743 (N_6743,N_4445,N_371);
xor U6744 (N_6744,N_5435,N_1170);
nand U6745 (N_6745,N_3550,N_4950);
nor U6746 (N_6746,N_5563,N_2542);
nand U6747 (N_6747,N_2757,N_216);
or U6748 (N_6748,N_2261,N_2350);
or U6749 (N_6749,N_1894,N_673);
and U6750 (N_6750,N_4681,N_3318);
nor U6751 (N_6751,N_5132,N_416);
and U6752 (N_6752,N_6168,N_1097);
or U6753 (N_6753,N_2381,N_1816);
and U6754 (N_6754,N_6190,N_4003);
nand U6755 (N_6755,N_2125,N_724);
and U6756 (N_6756,N_2183,N_518);
nor U6757 (N_6757,N_8,N_2689);
and U6758 (N_6758,N_2629,N_77);
nor U6759 (N_6759,N_5100,N_4040);
nand U6760 (N_6760,N_71,N_6212);
nor U6761 (N_6761,N_5416,N_4630);
and U6762 (N_6762,N_2171,N_1071);
nand U6763 (N_6763,N_3121,N_1579);
nor U6764 (N_6764,N_1189,N_552);
nor U6765 (N_6765,N_6095,N_2664);
nor U6766 (N_6766,N_6233,N_357);
and U6767 (N_6767,N_4851,N_282);
nand U6768 (N_6768,N_5104,N_3209);
xor U6769 (N_6769,N_1893,N_2226);
xor U6770 (N_6770,N_1766,N_1787);
nand U6771 (N_6771,N_2243,N_5631);
or U6772 (N_6772,N_1043,N_1884);
or U6773 (N_6773,N_5058,N_1090);
xor U6774 (N_6774,N_4634,N_804);
nand U6775 (N_6775,N_3044,N_4179);
nor U6776 (N_6776,N_3517,N_4616);
and U6777 (N_6777,N_428,N_2179);
or U6778 (N_6778,N_5110,N_5824);
and U6779 (N_6779,N_353,N_1536);
and U6780 (N_6780,N_1733,N_3407);
nand U6781 (N_6781,N_4922,N_1051);
nor U6782 (N_6782,N_3858,N_178);
nor U6783 (N_6783,N_5334,N_3881);
or U6784 (N_6784,N_5307,N_2047);
and U6785 (N_6785,N_3817,N_3870);
nand U6786 (N_6786,N_1853,N_4638);
and U6787 (N_6787,N_6032,N_5813);
nor U6788 (N_6788,N_5914,N_3393);
nor U6789 (N_6789,N_43,N_5843);
and U6790 (N_6790,N_2392,N_4618);
nor U6791 (N_6791,N_2032,N_5325);
nand U6792 (N_6792,N_5327,N_5854);
nor U6793 (N_6793,N_5277,N_1503);
nand U6794 (N_6794,N_3098,N_3381);
or U6795 (N_6795,N_6087,N_3686);
and U6796 (N_6796,N_3634,N_1464);
nand U6797 (N_6797,N_3196,N_6147);
nand U6798 (N_6798,N_439,N_1985);
and U6799 (N_6799,N_4116,N_4026);
or U6800 (N_6800,N_5720,N_1301);
nor U6801 (N_6801,N_1606,N_1686);
and U6802 (N_6802,N_297,N_3053);
nor U6803 (N_6803,N_2680,N_5046);
or U6804 (N_6804,N_1268,N_1832);
nand U6805 (N_6805,N_4612,N_146);
nand U6806 (N_6806,N_4757,N_985);
or U6807 (N_6807,N_1181,N_5662);
and U6808 (N_6808,N_4341,N_1092);
nand U6809 (N_6809,N_5691,N_3788);
and U6810 (N_6810,N_710,N_5373);
and U6811 (N_6811,N_4149,N_942);
and U6812 (N_6812,N_4599,N_289);
nor U6813 (N_6813,N_2518,N_3018);
and U6814 (N_6814,N_462,N_784);
nor U6815 (N_6815,N_5314,N_3527);
and U6816 (N_6816,N_4340,N_163);
nor U6817 (N_6817,N_885,N_4472);
xnor U6818 (N_6818,N_3905,N_3225);
or U6819 (N_6819,N_2083,N_894);
and U6820 (N_6820,N_6074,N_3955);
nor U6821 (N_6821,N_3251,N_3838);
and U6822 (N_6822,N_497,N_3827);
nand U6823 (N_6823,N_923,N_3429);
nor U6824 (N_6824,N_1836,N_5202);
nor U6825 (N_6825,N_1095,N_2118);
and U6826 (N_6826,N_933,N_5650);
nand U6827 (N_6827,N_142,N_3045);
and U6828 (N_6828,N_4951,N_5937);
and U6829 (N_6829,N_4814,N_19);
or U6830 (N_6830,N_3821,N_3181);
xor U6831 (N_6831,N_6020,N_3055);
and U6832 (N_6832,N_2691,N_171);
nand U6833 (N_6833,N_6076,N_3468);
and U6834 (N_6834,N_4103,N_4059);
nand U6835 (N_6835,N_5407,N_4777);
nor U6836 (N_6836,N_132,N_2376);
nand U6837 (N_6837,N_3330,N_4694);
and U6838 (N_6838,N_2146,N_4631);
and U6839 (N_6839,N_626,N_5859);
nor U6840 (N_6840,N_5917,N_3127);
and U6841 (N_6841,N_3090,N_3808);
nor U6842 (N_6842,N_2156,N_5705);
nand U6843 (N_6843,N_967,N_6176);
nand U6844 (N_6844,N_3764,N_4206);
nand U6845 (N_6845,N_4342,N_5479);
xor U6846 (N_6846,N_1687,N_3701);
nor U6847 (N_6847,N_5648,N_3477);
nor U6848 (N_6848,N_2377,N_73);
and U6849 (N_6849,N_1298,N_1941);
nand U6850 (N_6850,N_3382,N_5423);
nor U6851 (N_6851,N_2266,N_5041);
or U6852 (N_6852,N_2885,N_5219);
or U6853 (N_6853,N_5075,N_1869);
and U6854 (N_6854,N_4705,N_4478);
or U6855 (N_6855,N_2488,N_1839);
nand U6856 (N_6856,N_4106,N_5606);
or U6857 (N_6857,N_5534,N_4254);
nor U6858 (N_6858,N_5660,N_1142);
nor U6859 (N_6859,N_2855,N_1644);
and U6860 (N_6860,N_4788,N_4002);
nor U6861 (N_6861,N_1695,N_5636);
or U6862 (N_6862,N_658,N_3137);
nand U6863 (N_6863,N_2692,N_1761);
and U6864 (N_6864,N_4760,N_1908);
xor U6865 (N_6865,N_5467,N_5002);
and U6866 (N_6866,N_5616,N_1663);
or U6867 (N_6867,N_417,N_5791);
or U6868 (N_6868,N_5470,N_3792);
and U6869 (N_6869,N_5792,N_5822);
or U6870 (N_6870,N_2443,N_5396);
nor U6871 (N_6871,N_2405,N_1398);
and U6872 (N_6872,N_4155,N_3312);
or U6873 (N_6873,N_1386,N_2955);
and U6874 (N_6874,N_5138,N_4932);
nand U6875 (N_6875,N_5740,N_4213);
nand U6876 (N_6876,N_1455,N_256);
and U6877 (N_6877,N_4650,N_3604);
or U6878 (N_6878,N_1967,N_3279);
and U6879 (N_6879,N_739,N_3666);
or U6880 (N_6880,N_2131,N_607);
nand U6881 (N_6881,N_1391,N_2042);
nor U6882 (N_6882,N_1944,N_476);
nor U6883 (N_6883,N_4888,N_3992);
and U6884 (N_6884,N_4920,N_1287);
nand U6885 (N_6885,N_3580,N_2872);
or U6886 (N_6886,N_3245,N_1403);
and U6887 (N_6887,N_4316,N_123);
nor U6888 (N_6888,N_4219,N_4531);
or U6889 (N_6889,N_3656,N_3682);
or U6890 (N_6890,N_3614,N_2791);
nand U6891 (N_6891,N_1849,N_4728);
nor U6892 (N_6892,N_3702,N_5749);
or U6893 (N_6893,N_3560,N_1540);
and U6894 (N_6894,N_3595,N_5715);
nand U6895 (N_6895,N_3732,N_3074);
or U6896 (N_6896,N_4999,N_1848);
nand U6897 (N_6897,N_5098,N_5596);
or U6898 (N_6898,N_2231,N_2976);
xnor U6899 (N_6899,N_4239,N_4602);
and U6900 (N_6900,N_5019,N_3932);
nor U6901 (N_6901,N_464,N_962);
or U6902 (N_6902,N_494,N_2519);
nand U6903 (N_6903,N_5069,N_2429);
and U6904 (N_6904,N_15,N_3657);
or U6905 (N_6905,N_262,N_2406);
nand U6906 (N_6906,N_1310,N_2806);
or U6907 (N_6907,N_5475,N_3234);
nand U6908 (N_6908,N_2494,N_1178);
and U6909 (N_6909,N_5701,N_1077);
or U6910 (N_6910,N_1722,N_723);
and U6911 (N_6911,N_1054,N_1445);
xor U6912 (N_6912,N_2320,N_4502);
nor U6913 (N_6913,N_5544,N_4683);
nand U6914 (N_6914,N_4114,N_5301);
and U6915 (N_6915,N_5406,N_596);
nand U6916 (N_6916,N_2306,N_12);
nor U6917 (N_6917,N_1107,N_5072);
xnor U6918 (N_6918,N_3818,N_109);
and U6919 (N_6919,N_3956,N_1448);
nand U6920 (N_6920,N_3984,N_1921);
and U6921 (N_6921,N_900,N_3807);
and U6922 (N_6922,N_2624,N_292);
nand U6923 (N_6923,N_5161,N_4231);
and U6924 (N_6924,N_4092,N_6026);
nand U6925 (N_6925,N_3620,N_4459);
or U6926 (N_6926,N_1764,N_118);
and U6927 (N_6927,N_2071,N_769);
nand U6928 (N_6928,N_2498,N_762);
or U6929 (N_6929,N_4891,N_852);
nor U6930 (N_6930,N_1599,N_6154);
nand U6931 (N_6931,N_78,N_5169);
nand U6932 (N_6932,N_3431,N_1727);
and U6933 (N_6933,N_3780,N_4305);
nor U6934 (N_6934,N_6063,N_3871);
nand U6935 (N_6935,N_2839,N_2636);
or U6936 (N_6936,N_2351,N_2007);
and U6937 (N_6937,N_2592,N_2263);
xor U6938 (N_6938,N_6140,N_5055);
nand U6939 (N_6939,N_3094,N_2783);
nor U6940 (N_6940,N_593,N_4447);
nand U6941 (N_6941,N_2975,N_2169);
nor U6942 (N_6942,N_5123,N_4900);
or U6943 (N_6943,N_5259,N_6019);
or U6944 (N_6944,N_3869,N_5463);
nand U6945 (N_6945,N_5029,N_2373);
nand U6946 (N_6946,N_3166,N_340);
nand U6947 (N_6947,N_587,N_6025);
and U6948 (N_6948,N_389,N_5000);
and U6949 (N_6949,N_56,N_5176);
nor U6950 (N_6950,N_2825,N_4708);
or U6951 (N_6951,N_3064,N_4390);
nor U6952 (N_6952,N_3378,N_5707);
nor U6953 (N_6953,N_653,N_6072);
xnor U6954 (N_6954,N_3062,N_2603);
nor U6955 (N_6955,N_2627,N_5295);
and U6956 (N_6956,N_2439,N_2840);
and U6957 (N_6957,N_3048,N_2416);
nor U6958 (N_6958,N_1549,N_1086);
and U6959 (N_6959,N_5690,N_4654);
nor U6960 (N_6960,N_257,N_5861);
nand U6961 (N_6961,N_2543,N_3524);
or U6962 (N_6962,N_4493,N_1571);
nand U6963 (N_6963,N_5430,N_1339);
nand U6964 (N_6964,N_4230,N_3276);
nor U6965 (N_6965,N_1520,N_3060);
and U6966 (N_6966,N_5137,N_4464);
or U6967 (N_6967,N_2907,N_742);
or U6968 (N_6968,N_2318,N_652);
or U6969 (N_6969,N_4164,N_4859);
nand U6970 (N_6970,N_6227,N_36);
or U6971 (N_6971,N_551,N_1387);
or U6972 (N_6972,N_2313,N_1331);
nand U6973 (N_6973,N_6208,N_6173);
and U6974 (N_6974,N_4208,N_498);
nand U6975 (N_6975,N_2167,N_2591);
and U6976 (N_6976,N_2345,N_3426);
and U6977 (N_6977,N_1076,N_2782);
and U6978 (N_6978,N_3015,N_1975);
and U6979 (N_6979,N_2431,N_5623);
and U6980 (N_6980,N_751,N_1422);
and U6981 (N_6981,N_355,N_3116);
xor U6982 (N_6982,N_3016,N_5823);
and U6983 (N_6983,N_4180,N_4767);
xor U6984 (N_6984,N_3713,N_598);
nand U6985 (N_6985,N_1752,N_2041);
nor U6986 (N_6986,N_4635,N_5141);
xnor U6987 (N_6987,N_5092,N_4300);
nor U6988 (N_6988,N_6052,N_2962);
xnor U6989 (N_6989,N_4210,N_4069);
or U6990 (N_6990,N_4226,N_2748);
nor U6991 (N_6991,N_5642,N_761);
nand U6992 (N_6992,N_5862,N_4376);
nor U6993 (N_6993,N_2846,N_5050);
nor U6994 (N_6994,N_1684,N_4805);
nand U6995 (N_6995,N_4279,N_2204);
or U6996 (N_6996,N_2886,N_2151);
or U6997 (N_6997,N_1276,N_4013);
nand U6998 (N_6998,N_1049,N_4844);
nand U6999 (N_6999,N_1491,N_4150);
nand U7000 (N_7000,N_667,N_6172);
and U7001 (N_7001,N_838,N_3020);
xor U7002 (N_7002,N_4205,N_4014);
nor U7003 (N_7003,N_377,N_3088);
nand U7004 (N_7004,N_6106,N_2008);
or U7005 (N_7005,N_2153,N_6189);
or U7006 (N_7006,N_3434,N_3176);
or U7007 (N_7007,N_550,N_5469);
nand U7008 (N_7008,N_6134,N_1934);
or U7009 (N_7009,N_901,N_5820);
nor U7010 (N_7010,N_2449,N_1203);
nand U7011 (N_7011,N_4012,N_349);
and U7012 (N_7012,N_768,N_2528);
or U7013 (N_7013,N_2540,N_897);
nand U7014 (N_7014,N_668,N_666);
xnor U7015 (N_7015,N_58,N_934);
nor U7016 (N_7016,N_1184,N_165);
xnor U7017 (N_7017,N_2538,N_3736);
xor U7018 (N_7018,N_3490,N_3976);
and U7019 (N_7019,N_4361,N_25);
nor U7020 (N_7020,N_2499,N_3177);
xor U7021 (N_7021,N_3644,N_5006);
xor U7022 (N_7022,N_3975,N_2722);
xnor U7023 (N_7023,N_3141,N_861);
nand U7024 (N_7024,N_4716,N_4868);
and U7025 (N_7025,N_1532,N_4086);
nor U7026 (N_7026,N_124,N_2189);
or U7027 (N_7027,N_6113,N_5773);
nand U7028 (N_7028,N_2833,N_5593);
and U7029 (N_7029,N_774,N_5944);
and U7030 (N_7030,N_4853,N_6118);
nand U7031 (N_7031,N_3583,N_3113);
nor U7032 (N_7032,N_5746,N_1167);
or U7033 (N_7033,N_1558,N_4500);
and U7034 (N_7034,N_81,N_265);
xnor U7035 (N_7035,N_830,N_4332);
or U7036 (N_7036,N_1796,N_5064);
nor U7037 (N_7037,N_3610,N_3619);
nand U7038 (N_7038,N_3650,N_99);
or U7039 (N_7039,N_3199,N_5704);
xnor U7040 (N_7040,N_4939,N_445);
xnor U7041 (N_7041,N_3144,N_1480);
and U7042 (N_7042,N_747,N_3182);
nand U7043 (N_7043,N_780,N_2447);
nor U7044 (N_7044,N_3464,N_1605);
nand U7045 (N_7045,N_4839,N_3674);
or U7046 (N_7046,N_2678,N_3716);
nand U7047 (N_7047,N_5187,N_1656);
nand U7048 (N_7048,N_2078,N_834);
xor U7049 (N_7049,N_6123,N_2253);
nand U7050 (N_7050,N_2780,N_2671);
and U7051 (N_7051,N_5607,N_2147);
and U7052 (N_7052,N_4651,N_6094);
or U7053 (N_7053,N_179,N_418);
nor U7054 (N_7054,N_3618,N_3997);
and U7055 (N_7055,N_3001,N_4479);
nor U7056 (N_7056,N_488,N_1851);
nand U7057 (N_7057,N_2048,N_2382);
nand U7058 (N_7058,N_2185,N_5224);
xor U7059 (N_7059,N_6177,N_3758);
and U7060 (N_7060,N_1369,N_1688);
or U7061 (N_7061,N_2365,N_2865);
nor U7062 (N_7062,N_4726,N_5367);
nand U7063 (N_7063,N_316,N_619);
and U7064 (N_7064,N_1743,N_2898);
nor U7065 (N_7065,N_3988,N_2176);
nor U7066 (N_7066,N_920,N_3128);
nor U7067 (N_7067,N_6092,N_3228);
and U7068 (N_7068,N_2784,N_5975);
and U7069 (N_7069,N_2695,N_5449);
and U7070 (N_7070,N_4657,N_721);
nand U7071 (N_7071,N_3909,N_4042);
nor U7072 (N_7072,N_686,N_2642);
nor U7073 (N_7073,N_3011,N_624);
and U7074 (N_7074,N_5076,N_4553);
nor U7075 (N_7075,N_3868,N_4240);
and U7076 (N_7076,N_1526,N_2953);
xnor U7077 (N_7077,N_4698,N_1209);
nand U7078 (N_7078,N_3301,N_5995);
xor U7079 (N_7079,N_2752,N_4949);
or U7080 (N_7080,N_2109,N_3454);
or U7081 (N_7081,N_1361,N_1017);
or U7082 (N_7082,N_4399,N_5628);
nand U7083 (N_7083,N_5689,N_1547);
or U7084 (N_7084,N_1040,N_1712);
or U7085 (N_7085,N_4327,N_5223);
and U7086 (N_7086,N_4441,N_273);
and U7087 (N_7087,N_4697,N_5399);
xnor U7088 (N_7088,N_2018,N_908);
xor U7089 (N_7089,N_3273,N_4809);
xnor U7090 (N_7090,N_3283,N_6064);
or U7091 (N_7091,N_310,N_3667);
and U7092 (N_7092,N_5578,N_2736);
nor U7093 (N_7093,N_6243,N_831);
nand U7094 (N_7094,N_4386,N_662);
nand U7095 (N_7095,N_1094,N_806);
and U7096 (N_7096,N_2354,N_3275);
xnor U7097 (N_7097,N_6237,N_2870);
nand U7098 (N_7098,N_1416,N_5136);
nand U7099 (N_7099,N_1831,N_421);
nand U7100 (N_7100,N_446,N_5894);
or U7101 (N_7101,N_2604,N_5574);
nor U7102 (N_7102,N_2570,N_1397);
nand U7103 (N_7103,N_601,N_2548);
and U7104 (N_7104,N_2188,N_4196);
nand U7105 (N_7105,N_5222,N_5681);
nor U7106 (N_7106,N_3058,N_2630);
or U7107 (N_7107,N_5361,N_2110);
nor U7108 (N_7108,N_2849,N_1911);
and U7109 (N_7109,N_5809,N_1212);
nor U7110 (N_7110,N_2739,N_1450);
or U7111 (N_7111,N_2393,N_2587);
nand U7112 (N_7112,N_4886,N_6050);
and U7113 (N_7113,N_105,N_6043);
and U7114 (N_7114,N_5724,N_3961);
xnor U7115 (N_7115,N_6213,N_5942);
xnor U7116 (N_7116,N_558,N_2559);
or U7117 (N_7117,N_4298,N_4987);
or U7118 (N_7118,N_162,N_961);
or U7119 (N_7119,N_3133,N_187);
xnor U7120 (N_7120,N_569,N_2371);
nor U7121 (N_7121,N_4748,N_5697);
nand U7122 (N_7122,N_2349,N_1497);
xnor U7123 (N_7123,N_3652,N_4415);
nand U7124 (N_7124,N_2248,N_4779);
or U7125 (N_7125,N_3856,N_3982);
nor U7126 (N_7126,N_6150,N_998);
nand U7127 (N_7127,N_6215,N_2658);
and U7128 (N_7128,N_1050,N_5679);
xor U7129 (N_7129,N_1004,N_4918);
or U7130 (N_7130,N_972,N_1797);
and U7131 (N_7131,N_3480,N_1507);
xor U7132 (N_7132,N_2380,N_1476);
nor U7133 (N_7133,N_1602,N_2945);
or U7134 (N_7134,N_3872,N_1355);
or U7135 (N_7135,N_1705,N_4820);
nand U7136 (N_7136,N_6018,N_5487);
nand U7137 (N_7137,N_2436,N_4801);
xnor U7138 (N_7138,N_250,N_5774);
or U7139 (N_7139,N_2106,N_4914);
or U7140 (N_7140,N_5940,N_4590);
nand U7141 (N_7141,N_735,N_1477);
and U7142 (N_7142,N_1206,N_1063);
or U7143 (N_7143,N_5556,N_2826);
nand U7144 (N_7144,N_4191,N_3047);
nand U7145 (N_7145,N_5382,N_1151);
and U7146 (N_7146,N_461,N_2977);
nand U7147 (N_7147,N_2072,N_251);
and U7148 (N_7148,N_6198,N_4586);
nand U7149 (N_7149,N_1282,N_4833);
nand U7150 (N_7150,N_4506,N_5394);
or U7151 (N_7151,N_3648,N_1924);
or U7152 (N_7152,N_3087,N_1299);
nand U7153 (N_7153,N_1283,N_4093);
nand U7154 (N_7154,N_4784,N_348);
xor U7155 (N_7155,N_863,N_902);
xor U7156 (N_7156,N_1205,N_5725);
nand U7157 (N_7157,N_18,N_3041);
or U7158 (N_7158,N_2520,N_2560);
nor U7159 (N_7159,N_2521,N_1601);
or U7160 (N_7160,N_2326,N_429);
and U7161 (N_7161,N_4047,N_4818);
nand U7162 (N_7162,N_5852,N_6205);
nor U7163 (N_7163,N_4504,N_4780);
nand U7164 (N_7164,N_4540,N_5147);
or U7165 (N_7165,N_4509,N_4543);
or U7166 (N_7166,N_2763,N_4410);
nand U7167 (N_7167,N_5562,N_2090);
and U7168 (N_7168,N_4125,N_2004);
or U7169 (N_7169,N_3388,N_1960);
nor U7170 (N_7170,N_2228,N_4194);
and U7171 (N_7171,N_5258,N_5353);
or U7172 (N_7172,N_2286,N_4295);
nor U7173 (N_7173,N_4768,N_4255);
nand U7174 (N_7174,N_1544,N_2727);
xnor U7175 (N_7175,N_4963,N_144);
nand U7176 (N_7176,N_3602,N_42);
or U7177 (N_7177,N_7,N_5674);
and U7178 (N_7178,N_3145,N_2639);
or U7179 (N_7179,N_2230,N_3467);
or U7180 (N_7180,N_3404,N_3859);
nand U7181 (N_7181,N_1829,N_1390);
nand U7182 (N_7182,N_4140,N_1199);
xnor U7183 (N_7183,N_4380,N_1616);
and U7184 (N_7184,N_5583,N_1977);
and U7185 (N_7185,N_2205,N_5872);
nor U7186 (N_7186,N_3399,N_5865);
nand U7187 (N_7187,N_1806,N_4800);
xor U7188 (N_7188,N_2961,N_4271);
nand U7189 (N_7189,N_3599,N_6013);
nor U7190 (N_7190,N_2933,N_309);
and U7191 (N_7191,N_1084,N_3866);
nand U7192 (N_7192,N_2476,N_1306);
xnor U7193 (N_7193,N_3243,N_2383);
nor U7194 (N_7194,N_2073,N_2260);
nand U7195 (N_7195,N_3315,N_5845);
and U7196 (N_7196,N_5008,N_303);
and U7197 (N_7197,N_4057,N_3298);
nor U7198 (N_7198,N_4893,N_2740);
nand U7199 (N_7199,N_423,N_5317);
nor U7200 (N_7200,N_2491,N_2735);
nand U7201 (N_7201,N_5638,N_3704);
nor U7202 (N_7202,N_4051,N_1876);
nor U7203 (N_7203,N_606,N_1225);
and U7204 (N_7204,N_2086,N_2427);
or U7205 (N_7205,N_659,N_129);
nand U7206 (N_7206,N_5060,N_5338);
and U7207 (N_7207,N_1285,N_4569);
nand U7208 (N_7208,N_1834,N_3244);
nor U7209 (N_7209,N_3293,N_3124);
nor U7210 (N_7210,N_2888,N_3427);
or U7211 (N_7211,N_5921,N_2296);
and U7212 (N_7212,N_4487,N_5051);
xnor U7213 (N_7213,N_1294,N_1701);
or U7214 (N_7214,N_5038,N_1615);
and U7215 (N_7215,N_5629,N_2772);
nand U7216 (N_7216,N_2369,N_452);
nor U7217 (N_7217,N_2223,N_2346);
nor U7218 (N_7218,N_2807,N_4710);
and U7219 (N_7219,N_4962,N_4535);
nand U7220 (N_7220,N_4991,N_2237);
nand U7221 (N_7221,N_4591,N_258);
nand U7222 (N_7222,N_4897,N_5550);
nor U7223 (N_7223,N_1843,N_5680);
and U7224 (N_7224,N_5857,N_2208);
or U7225 (N_7225,N_2502,N_1715);
and U7226 (N_7226,N_1860,N_4729);
and U7227 (N_7227,N_102,N_300);
nor U7228 (N_7228,N_2412,N_2339);
xnor U7229 (N_7229,N_1735,N_5504);
and U7230 (N_7230,N_5403,N_4636);
nand U7231 (N_7231,N_4090,N_5840);
nor U7232 (N_7232,N_1153,N_5377);
xnor U7233 (N_7233,N_5542,N_2178);
nor U7234 (N_7234,N_5632,N_5983);
nor U7235 (N_7235,N_2168,N_3723);
xnor U7236 (N_7236,N_2732,N_4741);
and U7237 (N_7237,N_487,N_3402);
or U7238 (N_7238,N_92,N_1029);
nand U7239 (N_7239,N_4244,N_576);
nand U7240 (N_7240,N_4362,N_379);
nor U7241 (N_7241,N_5344,N_4359);
and U7242 (N_7242,N_1473,N_2453);
or U7243 (N_7243,N_4727,N_3895);
nand U7244 (N_7244,N_1135,N_4243);
and U7245 (N_7245,N_5899,N_5664);
or U7246 (N_7246,N_2112,N_1781);
or U7247 (N_7247,N_3421,N_5266);
nand U7248 (N_7248,N_4496,N_157);
nand U7249 (N_7249,N_5835,N_548);
and U7250 (N_7250,N_3885,N_650);
nand U7251 (N_7251,N_3417,N_2988);
nand U7252 (N_7252,N_5456,N_3425);
nand U7253 (N_7253,N_3946,N_5381);
xnor U7254 (N_7254,N_2417,N_799);
or U7255 (N_7255,N_5150,N_5004);
nor U7256 (N_7256,N_237,N_2659);
and U7257 (N_7257,N_1169,N_3270);
nor U7258 (N_7258,N_2555,N_3445);
nor U7259 (N_7259,N_275,N_3184);
or U7260 (N_7260,N_218,N_3926);
or U7261 (N_7261,N_4216,N_717);
and U7262 (N_7262,N_3117,N_3726);
nand U7263 (N_7263,N_5644,N_459);
nor U7264 (N_7264,N_79,N_911);
or U7265 (N_7265,N_4515,N_2407);
nand U7266 (N_7266,N_5761,N_65);
nand U7267 (N_7267,N_4259,N_2127);
xnor U7268 (N_7268,N_3617,N_2879);
nand U7269 (N_7269,N_3953,N_2984);
and U7270 (N_7270,N_5717,N_6217);
nand U7271 (N_7271,N_2375,N_1846);
nand U7272 (N_7272,N_3631,N_333);
xnor U7273 (N_7273,N_5731,N_4321);
nor U7274 (N_7274,N_2837,N_3004);
and U7275 (N_7275,N_2858,N_5832);
nand U7276 (N_7276,N_5706,N_1534);
nor U7277 (N_7277,N_5217,N_528);
nand U7278 (N_7278,N_509,N_529);
or U7279 (N_7279,N_4171,N_1415);
xor U7280 (N_7280,N_1969,N_5450);
nand U7281 (N_7281,N_434,N_456);
and U7282 (N_7282,N_753,N_2397);
nand U7283 (N_7283,N_5451,N_4627);
nor U7284 (N_7284,N_3232,N_4595);
and U7285 (N_7285,N_4161,N_4608);
and U7286 (N_7286,N_3508,N_4787);
nor U7287 (N_7287,N_3379,N_5179);
nor U7288 (N_7288,N_5512,N_119);
and U7289 (N_7289,N_5035,N_6225);
and U7290 (N_7290,N_5825,N_3498);
nor U7291 (N_7291,N_4954,N_2884);
nand U7292 (N_7292,N_6175,N_4617);
nor U7293 (N_7293,N_6079,N_3546);
and U7294 (N_7294,N_80,N_4407);
nand U7295 (N_7295,N_5521,N_1418);
nor U7296 (N_7296,N_1642,N_1850);
xnor U7297 (N_7297,N_3171,N_85);
and U7298 (N_7298,N_1749,N_2940);
nand U7299 (N_7299,N_1228,N_501);
nor U7300 (N_7300,N_5429,N_3325);
or U7301 (N_7301,N_1622,N_4066);
nand U7302 (N_7302,N_4937,N_5695);
nand U7303 (N_7303,N_5103,N_1804);
and U7304 (N_7304,N_383,N_1165);
or U7305 (N_7305,N_223,N_2463);
nor U7306 (N_7306,N_61,N_4366);
xnor U7307 (N_7307,N_801,N_1751);
or U7308 (N_7308,N_1370,N_5696);
nand U7309 (N_7309,N_1986,N_4559);
and U7310 (N_7310,N_2648,N_5365);
xor U7311 (N_7311,N_30,N_5013);
or U7312 (N_7312,N_2905,N_522);
nor U7313 (N_7313,N_3677,N_5140);
and U7314 (N_7314,N_5608,N_1466);
and U7315 (N_7315,N_4798,N_3143);
nor U7316 (N_7316,N_560,N_3624);
or U7317 (N_7317,N_120,N_919);
xor U7318 (N_7318,N_4832,N_2835);
nor U7319 (N_7319,N_472,N_5278);
or U7320 (N_7320,N_5097,N_2968);
or U7321 (N_7321,N_1527,N_4425);
nor U7322 (N_7322,N_2121,N_5973);
and U7323 (N_7323,N_4734,N_5699);
nor U7324 (N_7324,N_1706,N_3691);
nor U7325 (N_7325,N_5127,N_1430);
nand U7326 (N_7326,N_1680,N_5733);
or U7327 (N_7327,N_2651,N_5347);
and U7328 (N_7328,N_5332,N_2600);
or U7329 (N_7329,N_2913,N_707);
or U7330 (N_7330,N_2148,N_3632);
nor U7331 (N_7331,N_3319,N_5719);
xnor U7332 (N_7332,N_3170,N_1514);
and U7333 (N_7333,N_4162,N_1755);
nor U7334 (N_7334,N_4062,N_1971);
xor U7335 (N_7335,N_4609,N_1257);
and U7336 (N_7336,N_5356,N_3521);
and U7337 (N_7337,N_4348,N_3156);
and U7338 (N_7338,N_2487,N_5204);
or U7339 (N_7339,N_531,N_1565);
xnor U7340 (N_7340,N_2229,N_4510);
nor U7341 (N_7341,N_409,N_3443);
and U7342 (N_7342,N_2960,N_347);
nor U7343 (N_7343,N_1679,N_5946);
nor U7344 (N_7344,N_6245,N_5977);
xnor U7345 (N_7345,N_2372,N_4045);
or U7346 (N_7346,N_1874,N_3059);
nor U7347 (N_7347,N_5811,N_4335);
nand U7348 (N_7348,N_4320,N_3973);
nor U7349 (N_7349,N_964,N_2054);
nand U7350 (N_7350,N_4632,N_3175);
nand U7351 (N_7351,N_3908,N_5622);
xnor U7352 (N_7352,N_5015,N_279);
nand U7353 (N_7353,N_971,N_4732);
nand U7354 (N_7354,N_873,N_5387);
nand U7355 (N_7355,N_3824,N_1885);
nor U7356 (N_7356,N_2776,N_912);
or U7357 (N_7357,N_1665,N_253);
nor U7358 (N_7358,N_738,N_1809);
or U7359 (N_7359,N_321,N_5146);
nand U7360 (N_7360,N_3336,N_4315);
nand U7361 (N_7361,N_4848,N_5417);
or U7362 (N_7362,N_3802,N_2293);
and U7363 (N_7363,N_4299,N_1254);
or U7364 (N_7364,N_4000,N_1154);
nor U7365 (N_7365,N_2666,N_5911);
nand U7366 (N_7366,N_2300,N_5779);
or U7367 (N_7367,N_2477,N_5905);
nor U7368 (N_7368,N_1171,N_1052);
nand U7369 (N_7369,N_749,N_2620);
and U7370 (N_7370,N_835,N_3664);
nor U7371 (N_7371,N_4730,N_5907);
nor U7372 (N_7372,N_1958,N_726);
nor U7373 (N_7373,N_2918,N_5782);
nor U7374 (N_7374,N_3472,N_3085);
nor U7375 (N_7375,N_4704,N_5021);
nor U7376 (N_7376,N_2493,N_45);
and U7377 (N_7377,N_2503,N_3898);
and U7378 (N_7378,N_1837,N_4588);
nor U7379 (N_7379,N_2744,N_4475);
xor U7380 (N_7380,N_1334,N_5061);
and U7381 (N_7381,N_966,N_2132);
or U7382 (N_7382,N_1669,N_1047);
nand U7383 (N_7383,N_4451,N_5881);
nor U7384 (N_7384,N_6186,N_6073);
and U7385 (N_7385,N_3941,N_1446);
and U7386 (N_7386,N_1333,N_2360);
nand U7387 (N_7387,N_4592,N_4587);
xnor U7388 (N_7388,N_2819,N_988);
and U7389 (N_7389,N_2534,N_4861);
and U7390 (N_7390,N_3478,N_4753);
or U7391 (N_7391,N_502,N_5546);
nand U7392 (N_7392,N_3092,N_5185);
nor U7393 (N_7393,N_2729,N_1318);
nand U7394 (N_7394,N_207,N_3711);
nor U7395 (N_7395,N_5374,N_2433);
nor U7396 (N_7396,N_4020,N_1300);
nand U7397 (N_7397,N_4241,N_5933);
or U7398 (N_7398,N_1937,N_1319);
nand U7399 (N_7399,N_3927,N_2362);
or U7400 (N_7400,N_2822,N_5956);
or U7401 (N_7401,N_699,N_217);
nand U7402 (N_7402,N_5119,N_5418);
and U7403 (N_7403,N_4282,N_3577);
nor U7404 (N_7404,N_1402,N_4197);
nor U7405 (N_7405,N_5472,N_544);
nor U7406 (N_7406,N_3458,N_4982);
xor U7407 (N_7407,N_22,N_2881);
nand U7408 (N_7408,N_2201,N_1487);
and U7409 (N_7409,N_654,N_4700);
nand U7410 (N_7410,N_4881,N_4942);
nor U7411 (N_7411,N_3576,N_6033);
xor U7412 (N_7412,N_2157,N_3310);
and U7413 (N_7413,N_2298,N_4456);
and U7414 (N_7414,N_5239,N_4262);
and U7415 (N_7415,N_3253,N_226);
and U7416 (N_7416,N_2364,N_1551);
or U7417 (N_7417,N_4435,N_1226);
or U7418 (N_7418,N_330,N_676);
or U7419 (N_7419,N_4581,N_5288);
or U7420 (N_7420,N_6224,N_6003);
or U7421 (N_7421,N_1116,N_1925);
and U7422 (N_7422,N_5063,N_4163);
or U7423 (N_7423,N_952,N_1545);
nand U7424 (N_7424,N_3056,N_2363);
nand U7425 (N_7425,N_3733,N_2685);
and U7426 (N_7426,N_5745,N_703);
or U7427 (N_7427,N_2682,N_614);
xor U7428 (N_7428,N_2022,N_4158);
nor U7429 (N_7429,N_4707,N_3046);
and U7430 (N_7430,N_2796,N_573);
and U7431 (N_7431,N_5554,N_2866);
nand U7432 (N_7432,N_5934,N_3855);
nand U7433 (N_7433,N_5459,N_3601);
or U7434 (N_7434,N_3430,N_4492);
nand U7435 (N_7435,N_1548,N_997);
nand U7436 (N_7436,N_5465,N_750);
and U7437 (N_7437,N_2754,N_403);
nor U7438 (N_7438,N_893,N_164);
nand U7439 (N_7439,N_6057,N_2026);
or U7440 (N_7440,N_4331,N_1972);
nand U7441 (N_7441,N_5592,N_1243);
or U7442 (N_7442,N_3155,N_851);
and U7443 (N_7443,N_198,N_3709);
and U7444 (N_7444,N_970,N_4766);
xnor U7445 (N_7445,N_1594,N_856);
and U7446 (N_7446,N_4526,N_1266);
nand U7447 (N_7447,N_3860,N_4437);
and U7448 (N_7448,N_1129,N_1066);
nand U7449 (N_7449,N_3854,N_3694);
or U7450 (N_7450,N_3189,N_4860);
xnor U7451 (N_7451,N_4883,N_2272);
nor U7452 (N_7452,N_4129,N_4450);
or U7453 (N_7453,N_6053,N_1692);
xor U7454 (N_7454,N_1115,N_3787);
nand U7455 (N_7455,N_3334,N_3355);
nand U7456 (N_7456,N_850,N_3627);
or U7457 (N_7457,N_1484,N_5047);
xor U7458 (N_7458,N_2302,N_2869);
or U7459 (N_7459,N_322,N_2214);
or U7460 (N_7460,N_5173,N_5565);
xor U7461 (N_7461,N_2398,N_3533);
and U7462 (N_7462,N_3008,N_134);
nand U7463 (N_7463,N_2446,N_2747);
xor U7464 (N_7464,N_5912,N_963);
nor U7465 (N_7465,N_3851,N_5789);
xor U7466 (N_7466,N_5576,N_1368);
and U7467 (N_7467,N_5659,N_3642);
nand U7468 (N_7468,N_5604,N_1649);
and U7469 (N_7469,N_4443,N_1664);
xnor U7470 (N_7470,N_1776,N_2182);
or U7471 (N_7471,N_2553,N_2430);
and U7472 (N_7472,N_213,N_1699);
or U7473 (N_7473,N_1800,N_6021);
or U7474 (N_7474,N_232,N_4597);
and U7475 (N_7475,N_2743,N_917);
nand U7476 (N_7476,N_1414,N_5641);
or U7477 (N_7477,N_3154,N_5022);
and U7478 (N_7478,N_3400,N_3769);
nor U7479 (N_7479,N_463,N_4281);
and U7480 (N_7480,N_1337,N_3949);
nand U7481 (N_7481,N_2941,N_3891);
nor U7482 (N_7482,N_201,N_4841);
and U7483 (N_7483,N_918,N_3267);
and U7484 (N_7484,N_1635,N_4455);
nand U7485 (N_7485,N_4462,N_2746);
or U7486 (N_7486,N_4491,N_3556);
nor U7487 (N_7487,N_3606,N_5891);
and U7488 (N_7488,N_5870,N_106);
or U7489 (N_7489,N_460,N_6232);
or U7490 (N_7490,N_3488,N_82);
nand U7491 (N_7491,N_5471,N_1863);
nor U7492 (N_7492,N_2951,N_3977);
nand U7493 (N_7493,N_4998,N_2473);
and U7494 (N_7494,N_5333,N_5023);
and U7495 (N_7495,N_4759,N_3963);
and U7496 (N_7496,N_5057,N_5555);
and U7497 (N_7497,N_4031,N_3506);
or U7498 (N_7498,N_3693,N_5145);
and U7499 (N_7499,N_3671,N_2394);
nand U7500 (N_7500,N_5947,N_2341);
or U7501 (N_7501,N_3823,N_3564);
nor U7502 (N_7502,N_1900,N_2238);
nand U7503 (N_7503,N_827,N_1903);
nand U7504 (N_7504,N_1785,N_1904);
nand U7505 (N_7505,N_798,N_1489);
and U7506 (N_7506,N_6195,N_6248);
nand U7507 (N_7507,N_1835,N_2906);
or U7508 (N_7508,N_3174,N_857);
xor U7509 (N_7509,N_5427,N_5115);
or U7510 (N_7510,N_3886,N_5536);
or U7511 (N_7511,N_5829,N_4633);
nor U7512 (N_7512,N_414,N_1645);
nor U7513 (N_7513,N_2983,N_1626);
or U7514 (N_7514,N_150,N_4518);
xor U7515 (N_7515,N_3022,N_2200);
nand U7516 (N_7516,N_3759,N_6108);
and U7517 (N_7517,N_3211,N_1567);
or U7518 (N_7518,N_4669,N_1);
or U7519 (N_7519,N_1126,N_2419);
nand U7520 (N_7520,N_4943,N_1657);
nand U7521 (N_7521,N_5769,N_2808);
nor U7522 (N_7522,N_5207,N_5254);
nor U7523 (N_7523,N_4996,N_2569);
xor U7524 (N_7524,N_2424,N_844);
nor U7525 (N_7525,N_1554,N_4647);
nand U7526 (N_7526,N_4131,N_3158);
xor U7527 (N_7527,N_3596,N_4611);
nor U7528 (N_7528,N_4573,N_6169);
or U7529 (N_7529,N_3698,N_1703);
or U7530 (N_7530,N_2005,N_3406);
nor U7531 (N_7531,N_3970,N_1232);
xnor U7532 (N_7532,N_2020,N_4318);
nand U7533 (N_7533,N_984,N_3383);
or U7534 (N_7534,N_4267,N_1612);
and U7535 (N_7535,N_2812,N_268);
nor U7536 (N_7536,N_5499,N_2108);
nand U7537 (N_7537,N_2335,N_2919);
and U7538 (N_7538,N_4102,N_4392);
nor U7539 (N_7539,N_3389,N_5949);
or U7540 (N_7540,N_5932,N_4799);
or U7541 (N_7541,N_1214,N_440);
and U7542 (N_7542,N_853,N_5203);
and U7543 (N_7543,N_1611,N_615);
nor U7544 (N_7544,N_5304,N_1782);
and U7545 (N_7545,N_2745,N_4660);
and U7546 (N_7546,N_4495,N_2235);
nand U7547 (N_7547,N_6102,N_4827);
and U7548 (N_7548,N_5694,N_3289);
nand U7549 (N_7549,N_2971,N_185);
nand U7550 (N_7550,N_5032,N_2797);
nand U7551 (N_7551,N_5414,N_3079);
nand U7552 (N_7552,N_2305,N_5197);
or U7553 (N_7553,N_2618,N_1886);
nor U7554 (N_7554,N_500,N_3380);
nand U7555 (N_7555,N_2871,N_2635);
and U7556 (N_7556,N_1012,N_5094);
nand U7557 (N_7557,N_5776,N_4877);
nor U7558 (N_7558,N_3653,N_5748);
or U7559 (N_7559,N_3637,N_1348);
nor U7560 (N_7560,N_5437,N_1451);
or U7561 (N_7561,N_996,N_2677);
or U7562 (N_7562,N_839,N_6191);
nand U7563 (N_7563,N_574,N_3993);
nor U7564 (N_7564,N_4123,N_3314);
nor U7565 (N_7565,N_1564,N_833);
nand U7566 (N_7566,N_199,N_981);
nand U7567 (N_7567,N_4875,N_2088);
nor U7568 (N_7568,N_4117,N_4792);
and U7569 (N_7569,N_3345,N_4220);
or U7570 (N_7570,N_3662,N_602);
nand U7571 (N_7571,N_2701,N_97);
xnor U7572 (N_7572,N_4072,N_2720);
nand U7573 (N_7573,N_6228,N_1702);
or U7574 (N_7574,N_2911,N_1179);
or U7575 (N_7575,N_3728,N_5700);
and U7576 (N_7576,N_21,N_3235);
nand U7577 (N_7577,N_2557,N_5062);
nor U7578 (N_7578,N_5003,N_5833);
nand U7579 (N_7579,N_5540,N_3603);
nand U7580 (N_7580,N_2868,N_2734);
or U7581 (N_7581,N_5348,N_5953);
or U7582 (N_7582,N_1260,N_4417);
or U7583 (N_7583,N_5313,N_5212);
nand U7584 (N_7584,N_3411,N_475);
or U7585 (N_7585,N_2733,N_4857);
or U7586 (N_7586,N_3543,N_2308);
nand U7587 (N_7587,N_3205,N_787);
nor U7588 (N_7588,N_5987,N_4141);
nand U7589 (N_7589,N_2164,N_2706);
or U7590 (N_7590,N_3582,N_4428);
xnor U7591 (N_7591,N_2094,N_2943);
nand U7592 (N_7592,N_890,N_4055);
and U7593 (N_7593,N_5492,N_6116);
xnor U7594 (N_7594,N_381,N_3612);
nor U7595 (N_7595,N_4643,N_2114);
nor U7596 (N_7596,N_4166,N_907);
nand U7597 (N_7597,N_959,N_2122);
and U7598 (N_7598,N_4625,N_4890);
and U7599 (N_7599,N_3416,N_211);
or U7600 (N_7600,N_2160,N_229);
xnor U7601 (N_7601,N_4228,N_1064);
nor U7602 (N_7602,N_5543,N_5999);
nand U7603 (N_7603,N_4721,N_4536);
nand U7604 (N_7604,N_1517,N_4744);
or U7605 (N_7605,N_2256,N_2723);
and U7606 (N_7606,N_3793,N_5948);
or U7607 (N_7607,N_3536,N_3125);
xor U7608 (N_7608,N_5812,N_5560);
or U7609 (N_7609,N_3083,N_451);
or U7610 (N_7610,N_5408,N_4793);
nand U7611 (N_7611,N_1058,N_4771);
or U7612 (N_7612,N_1589,N_4379);
or U7613 (N_7613,N_1041,N_3945);
nor U7614 (N_7614,N_155,N_2061);
nand U7615 (N_7615,N_4498,N_3916);
or U7616 (N_7616,N_1542,N_1623);
and U7617 (N_7617,N_4275,N_539);
and U7618 (N_7618,N_6109,N_4253);
nor U7619 (N_7619,N_1393,N_4438);
and U7620 (N_7620,N_5290,N_254);
nand U7621 (N_7621,N_3313,N_6179);
or U7622 (N_7622,N_4876,N_4905);
or U7623 (N_7623,N_2395,N_3608);
nor U7624 (N_7624,N_2959,N_1340);
nand U7625 (N_7625,N_4846,N_2793);
nand U7626 (N_7626,N_3009,N_4250);
or U7627 (N_7627,N_2033,N_1202);
and U7628 (N_7628,N_3588,N_5846);
nand U7629 (N_7629,N_4068,N_3248);
or U7630 (N_7630,N_2319,N_589);
or U7631 (N_7631,N_503,N_2768);
nor U7632 (N_7632,N_234,N_5397);
and U7633 (N_7633,N_5412,N_4577);
nor U7634 (N_7634,N_930,N_3080);
and U7635 (N_7635,N_4538,N_3902);
and U7636 (N_7636,N_5573,N_5297);
nand U7637 (N_7637,N_4307,N_5324);
and U7638 (N_7638,N_995,N_2596);
xnor U7639 (N_7639,N_2000,N_5436);
nor U7640 (N_7640,N_4533,N_3593);
nor U7641 (N_7641,N_2867,N_5634);
or U7642 (N_7642,N_5763,N_5765);
nand U7643 (N_7643,N_3051,N_2694);
nand U7644 (N_7644,N_4873,N_1566);
and U7645 (N_7645,N_4242,N_3850);
nand U7646 (N_7646,N_4222,N_499);
nor U7647 (N_7647,N_3339,N_5401);
xor U7648 (N_7648,N_1269,N_5447);
and U7649 (N_7649,N_5099,N_1273);
nor U7650 (N_7650,N_563,N_1256);
and U7651 (N_7651,N_1928,N_214);
and U7652 (N_7652,N_4195,N_5756);
xor U7653 (N_7653,N_128,N_6210);
nand U7654 (N_7654,N_2751,N_2159);
or U7655 (N_7655,N_1919,N_93);
nor U7656 (N_7656,N_400,N_4845);
or U7657 (N_7657,N_2514,N_1952);
or U7658 (N_7658,N_2549,N_640);
xor U7659 (N_7659,N_5777,N_4579);
or U7660 (N_7660,N_3920,N_2264);
and U7661 (N_7661,N_5319,N_4291);
and U7662 (N_7662,N_1976,N_2085);
or U7663 (N_7663,N_6047,N_1767);
nor U7664 (N_7664,N_5879,N_5461);
nand U7665 (N_7665,N_4144,N_1177);
or U7666 (N_7666,N_1738,N_1758);
or U7667 (N_7667,N_6091,N_4081);
and U7668 (N_7668,N_6048,N_788);
and U7669 (N_7669,N_1492,N_524);
nand U7670 (N_7670,N_1145,N_1760);
nor U7671 (N_7671,N_2728,N_2355);
nand U7672 (N_7672,N_493,N_5049);
nor U7673 (N_7673,N_5941,N_1218);
and U7674 (N_7674,N_634,N_4713);
or U7675 (N_7675,N_1812,N_3288);
xnor U7676 (N_7676,N_1909,N_6037);
nor U7677 (N_7677,N_3348,N_376);
nand U7678 (N_7678,N_5198,N_3518);
nor U7679 (N_7679,N_4105,N_786);
and U7680 (N_7680,N_3392,N_1949);
or U7681 (N_7681,N_2927,N_3303);
xnor U7682 (N_7682,N_2725,N_1512);
nand U7683 (N_7683,N_2472,N_5468);
or U7684 (N_7684,N_5121,N_3504);
nor U7685 (N_7685,N_1356,N_17);
nand U7686 (N_7686,N_2730,N_814);
and U7687 (N_7687,N_3118,N_3590);
nor U7688 (N_7688,N_4071,N_1109);
and U7689 (N_7689,N_4345,N_3297);
and U7690 (N_7690,N_1910,N_3401);
or U7691 (N_7691,N_623,N_957);
xor U7692 (N_7692,N_2937,N_3510);
or U7693 (N_7693,N_4743,N_3042);
nor U7694 (N_7694,N_6126,N_5422);
or U7695 (N_7695,N_4234,N_1578);
nor U7696 (N_7696,N_5354,N_4539);
nand U7697 (N_7697,N_2841,N_3123);
or U7698 (N_7698,N_2481,N_1629);
nor U7699 (N_7699,N_4044,N_5237);
and U7700 (N_7700,N_2344,N_3647);
or U7701 (N_7701,N_657,N_5775);
nor U7702 (N_7702,N_3331,N_228);
nor U7703 (N_7703,N_4807,N_3441);
nand U7704 (N_7704,N_1121,N_95);
or U7705 (N_7705,N_3761,N_5635);
nor U7706 (N_7706,N_4060,N_1309);
and U7707 (N_7707,N_621,N_2021);
nand U7708 (N_7708,N_143,N_1898);
nor U7709 (N_7709,N_2590,N_4078);
nand U7710 (N_7710,N_149,N_611);
and U7711 (N_7711,N_491,N_4442);
nor U7712 (N_7712,N_2634,N_1120);
and U7713 (N_7713,N_2883,N_915);
xnor U7714 (N_7714,N_4076,N_5339);
nor U7715 (N_7715,N_3980,N_14);
or U7716 (N_7716,N_3394,N_4);
or U7717 (N_7717,N_505,N_2152);
or U7718 (N_7718,N_4646,N_196);
or U7719 (N_7719,N_4986,N_444);
and U7720 (N_7720,N_4288,N_4689);
nand U7721 (N_7721,N_4325,N_5369);
nor U7722 (N_7722,N_5821,N_580);
and U7723 (N_7723,N_2471,N_2389);
nor U7724 (N_7724,N_3565,N_2278);
and U7725 (N_7725,N_1332,N_308);
xor U7726 (N_7726,N_1231,N_2532);
and U7727 (N_7727,N_1845,N_3791);
or U7728 (N_7728,N_1524,N_1286);
and U7729 (N_7729,N_4769,N_848);
and U7730 (N_7730,N_4187,N_3173);
and U7731 (N_7731,N_5957,N_3986);
or U7732 (N_7732,N_929,N_2457);
xor U7733 (N_7733,N_1326,N_3019);
nor U7734 (N_7734,N_3828,N_313);
or U7735 (N_7735,N_5245,N_2605);
or U7736 (N_7736,N_2480,N_1591);
xor U7737 (N_7737,N_4227,N_826);
nor U7738 (N_7738,N_135,N_90);
or U7739 (N_7739,N_3924,N_4605);
or U7740 (N_7740,N_5148,N_507);
nor U7741 (N_7741,N_692,N_1465);
nand U7742 (N_7742,N_4261,N_193);
or U7743 (N_7743,N_870,N_5081);
and U7744 (N_7744,N_2633,N_4218);
and U7745 (N_7745,N_5525,N_2513);
or U7746 (N_7746,N_670,N_2359);
nor U7747 (N_7747,N_5991,N_4711);
nor U7748 (N_7748,N_3503,N_1131);
nand U7749 (N_7749,N_3164,N_828);
nor U7750 (N_7750,N_600,N_5326);
and U7751 (N_7751,N_4831,N_5651);
or U7752 (N_7752,N_3349,N_1617);
and U7753 (N_7753,N_1349,N_1926);
nand U7754 (N_7754,N_4764,N_3921);
xor U7755 (N_7755,N_4326,N_398);
nand U7756 (N_7756,N_4296,N_4387);
or U7757 (N_7757,N_1963,N_4725);
nor U7758 (N_7758,N_183,N_4181);
xnor U7759 (N_7759,N_4659,N_796);
nand U7760 (N_7760,N_3277,N_1472);
nand U7761 (N_7761,N_5249,N_173);
nand U7762 (N_7762,N_1122,N_3549);
xor U7763 (N_7763,N_306,N_4746);
and U7764 (N_7764,N_4620,N_865);
and U7765 (N_7765,N_4879,N_2769);
nor U7766 (N_7766,N_4036,N_231);
and U7767 (N_7767,N_1509,N_6174);
and U7768 (N_7768,N_4589,N_4339);
nor U7769 (N_7769,N_4989,N_5411);
xor U7770 (N_7770,N_4701,N_4774);
nand U7771 (N_7771,N_771,N_5302);
and U7772 (N_7772,N_5280,N_121);
and U7773 (N_7773,N_5533,N_2921);
and U7774 (N_7774,N_1363,N_2165);
nand U7775 (N_7775,N_3901,N_2577);
nand U7776 (N_7776,N_2111,N_3223);
xor U7777 (N_7777,N_431,N_1127);
and U7778 (N_7778,N_3081,N_1421);
or U7779 (N_7779,N_442,N_4555);
nand U7780 (N_7780,N_2930,N_4662);
or U7781 (N_7781,N_4508,N_2824);
or U7782 (N_7782,N_671,N_4046);
xnor U7783 (N_7783,N_3720,N_3972);
or U7784 (N_7784,N_948,N_5404);
and U7785 (N_7785,N_2774,N_663);
nor U7786 (N_7786,N_5481,N_2087);
xor U7787 (N_7787,N_4367,N_3537);
nor U7788 (N_7788,N_6129,N_701);
or U7789 (N_7789,N_3917,N_4265);
and U7790 (N_7790,N_326,N_4752);
or U7791 (N_7791,N_3385,N_4394);
or U7792 (N_7792,N_3724,N_690);
and U7793 (N_7793,N_3714,N_2804);
nand U7794 (N_7794,N_3929,N_1817);
nor U7795 (N_7795,N_3741,N_323);
nor U7796 (N_7796,N_557,N_3131);
nand U7797 (N_7797,N_5101,N_111);
and U7798 (N_7798,N_5744,N_4077);
and U7799 (N_7799,N_396,N_1981);
nand U7800 (N_7800,N_1672,N_5548);
nand U7801 (N_7801,N_5124,N_4285);
and U7802 (N_7802,N_1953,N_4623);
and U7803 (N_7803,N_5960,N_4041);
nor U7804 (N_7804,N_2902,N_4446);
or U7805 (N_7805,N_1693,N_311);
nand U7806 (N_7806,N_1516,N_1500);
nor U7807 (N_7807,N_709,N_892);
nand U7808 (N_7808,N_3540,N_6068);
or U7809 (N_7809,N_3160,N_3915);
or U7810 (N_7810,N_4169,N_4402);
nand U7811 (N_7811,N_3122,N_5318);
nand U7812 (N_7812,N_2332,N_4693);
xor U7813 (N_7813,N_5980,N_1573);
nor U7814 (N_7814,N_399,N_656);
or U7815 (N_7815,N_2001,N_677);
nand U7816 (N_7816,N_2531,N_2334);
or U7817 (N_7817,N_5652,N_221);
nand U7818 (N_7818,N_757,N_6098);
or U7819 (N_7819,N_1720,N_4583);
and U7820 (N_7820,N_5073,N_714);
nor U7821 (N_7821,N_1411,N_5453);
nand U7822 (N_7822,N_1917,N_5391);
nand U7823 (N_7823,N_4022,N_3651);
and U7824 (N_7824,N_1890,N_2474);
nor U7825 (N_7825,N_2104,N_489);
nand U7826 (N_7826,N_3967,N_5350);
nand U7827 (N_7827,N_3106,N_5205);
nor U7828 (N_7828,N_4913,N_815);
or U7829 (N_7829,N_4615,N_4652);
xnor U7830 (N_7830,N_3770,N_3959);
nor U7831 (N_7831,N_4224,N_3743);
nor U7832 (N_7832,N_664,N_2556);
nor U7833 (N_7833,N_4639,N_521);
and U7834 (N_7834,N_4789,N_1089);
and U7835 (N_7835,N_4147,N_3237);
nor U7836 (N_7836,N_1014,N_4488);
or U7837 (N_7837,N_1372,N_3214);
or U7838 (N_7838,N_1730,N_5888);
or U7839 (N_7839,N_4797,N_3373);
or U7840 (N_7840,N_1608,N_5661);
and U7841 (N_7841,N_3183,N_6016);
or U7842 (N_7842,N_4409,N_1347);
or U7843 (N_7843,N_3272,N_5084);
xor U7844 (N_7844,N_3317,N_4675);
nor U7845 (N_7845,N_5702,N_3753);
and U7846 (N_7846,N_5189,N_1561);
and U7847 (N_7847,N_3740,N_1208);
nor U7848 (N_7848,N_3773,N_3197);
or U7849 (N_7849,N_2710,N_363);
nand U7850 (N_7850,N_1026,N_3484);
and U7851 (N_7851,N_1297,N_778);
or U7852 (N_7852,N_3635,N_5928);
and U7853 (N_7853,N_3474,N_4373);
or U7854 (N_7854,N_1419,N_5462);
nor U7855 (N_7855,N_1895,N_4494);
nand U7856 (N_7856,N_62,N_3140);
xor U7857 (N_7857,N_845,N_4596);
or U7858 (N_7858,N_4018,N_3559);
nand U7859 (N_7859,N_3332,N_1104);
or U7860 (N_7860,N_4690,N_5502);
nand U7861 (N_7861,N_1652,N_2079);
nor U7862 (N_7862,N_2062,N_898);
and U7863 (N_7863,N_3892,N_1943);
xor U7864 (N_7864,N_6203,N_16);
nand U7865 (N_7865,N_4984,N_1217);
and U7866 (N_7866,N_2342,N_4027);
or U7867 (N_7867,N_2705,N_3689);
xor U7868 (N_7868,N_2545,N_1556);
or U7869 (N_7869,N_2116,N_5508);
and U7870 (N_7870,N_5572,N_4958);
nor U7871 (N_7871,N_1295,N_373);
and U7872 (N_7872,N_1814,N_4554);
nand U7873 (N_7873,N_4347,N_1948);
nand U7874 (N_7874,N_3572,N_4619);
and U7875 (N_7875,N_437,N_4952);
nor U7876 (N_7876,N_4524,N_3622);
nor U7877 (N_7877,N_1322,N_2191);
xnor U7878 (N_7878,N_2737,N_2741);
nand U7879 (N_7879,N_1016,N_395);
nor U7880 (N_7880,N_3514,N_2274);
nor U7881 (N_7881,N_5088,N_2546);
nor U7882 (N_7882,N_4418,N_4201);
or U7883 (N_7883,N_879,N_3286);
nor U7884 (N_7884,N_1878,N_6103);
nand U7885 (N_7885,N_3295,N_496);
and U7886 (N_7886,N_69,N_307);
or U7887 (N_7887,N_324,N_4747);
and U7888 (N_7888,N_2414,N_4733);
and U7889 (N_7889,N_4547,N_3912);
nand U7890 (N_7890,N_5037,N_781);
and U7891 (N_7891,N_4855,N_2173);
nand U7892 (N_7892,N_2645,N_67);
nand U7893 (N_7893,N_6236,N_4997);
xor U7894 (N_7894,N_5269,N_684);
nand U7895 (N_7895,N_5723,N_2379);
nand U7896 (N_7896,N_1647,N_1947);
nand U7897 (N_7897,N_4751,N_785);
xor U7898 (N_7898,N_441,N_4233);
or U7899 (N_7899,N_410,N_5643);
nand U7900 (N_7900,N_5125,N_84);
or U7901 (N_7901,N_2246,N_2190);
or U7902 (N_7902,N_3372,N_4576);
xor U7903 (N_7903,N_5666,N_6100);
or U7904 (N_7904,N_2794,N_3326);
or U7905 (N_7905,N_1128,N_1303);
and U7906 (N_7906,N_2139,N_510);
nor U7907 (N_7907,N_2947,N_3784);
and U7908 (N_7908,N_542,N_5358);
or U7909 (N_7909,N_1858,N_3148);
nand U7910 (N_7910,N_5134,N_5675);
and U7911 (N_7911,N_2647,N_4465);
and U7912 (N_7912,N_3562,N_404);
or U7913 (N_7913,N_1223,N_5291);
and U7914 (N_7914,N_1057,N_1486);
xor U7915 (N_7915,N_4006,N_3853);
nand U7916 (N_7916,N_4967,N_478);
and U7917 (N_7917,N_1462,N_5741);
nor U7918 (N_7918,N_3960,N_3555);
xor U7919 (N_7919,N_5260,N_219);
and U7920 (N_7920,N_2500,N_1923);
nand U7921 (N_7921,N_4460,N_1330);
or U7922 (N_7922,N_3607,N_3449);
and U7923 (N_7923,N_3794,N_5996);
nand U7924 (N_7924,N_1220,N_260);
nand U7925 (N_7925,N_5787,N_3096);
nand U7926 (N_7926,N_374,N_4976);
and U7927 (N_7927,N_3418,N_1112);
nand U7928 (N_7928,N_3661,N_3934);
nor U7929 (N_7929,N_527,N_6036);
nor U7930 (N_7930,N_1428,N_269);
and U7931 (N_7931,N_5283,N_3346);
and U7932 (N_7932,N_2324,N_1019);
nand U7933 (N_7933,N_2973,N_242);
nand U7934 (N_7934,N_729,N_298);
nand U7935 (N_7935,N_2995,N_369);
nand U7936 (N_7936,N_1671,N_2512);
and U7937 (N_7937,N_4808,N_1436);
nand U7938 (N_7938,N_4336,N_1899);
nor U7939 (N_7939,N_2338,N_6070);
and U7940 (N_7940,N_2485,N_941);
xor U7941 (N_7941,N_591,N_443);
nand U7942 (N_7942,N_4926,N_6086);
nand U7943 (N_7943,N_5711,N_2896);
nor U7944 (N_7944,N_1531,N_2211);
or U7945 (N_7945,N_4120,N_5225);
nor U7946 (N_7946,N_1074,N_4916);
xor U7947 (N_7947,N_2410,N_2641);
or U7948 (N_7948,N_2174,N_4398);
nor U7949 (N_7949,N_2458,N_3172);
nand U7950 (N_7950,N_3231,N_1105);
and U7951 (N_7951,N_1676,N_519);
and U7952 (N_7952,N_1238,N_1392);
nand U7953 (N_7953,N_4405,N_4936);
xnor U7954 (N_7954,N_4849,N_4653);
xor U7955 (N_7955,N_3861,N_1396);
nor U7956 (N_7956,N_3361,N_1449);
nor U7957 (N_7957,N_5218,N_4461);
nor U7958 (N_7958,N_3007,N_360);
nand U7959 (N_7959,N_5345,N_1315);
nor U7960 (N_7960,N_5488,N_5089);
or U7961 (N_7961,N_4109,N_4190);
nand U7962 (N_7962,N_2625,N_925);
nor U7963 (N_7963,N_903,N_1609);
nand U7964 (N_7964,N_1892,N_4139);
nor U7965 (N_7965,N_3455,N_4578);
and U7966 (N_7966,N_4001,N_3673);
or U7967 (N_7967,N_2829,N_60);
and U7968 (N_7968,N_3863,N_698);
and U7969 (N_7969,N_2492,N_3918);
and U7970 (N_7970,N_1102,N_4249);
nand U7971 (N_7971,N_884,N_1255);
xnor U7972 (N_7972,N_5184,N_1481);
nand U7973 (N_7973,N_5808,N_6209);
nor U7974 (N_7974,N_2039,N_4925);
nor U7975 (N_7975,N_4738,N_5270);
and U7976 (N_7976,N_516,N_5806);
nand U7977 (N_7977,N_2276,N_4829);
nand U7978 (N_7978,N_5507,N_5402);
or U7979 (N_7979,N_772,N_2269);
and U7980 (N_7980,N_581,N_5096);
nand U7981 (N_7981,N_3910,N_1732);
nand U7982 (N_7982,N_1736,N_3163);
or U7983 (N_7983,N_4263,N_167);
or U7984 (N_7984,N_6014,N_4714);
nor U7985 (N_7985,N_5457,N_5770);
nor U7986 (N_7986,N_1175,N_5855);
or U7987 (N_7987,N_5285,N_4838);
and U7988 (N_7988,N_3075,N_1087);
nand U7989 (N_7989,N_5601,N_6222);
nand U7990 (N_7990,N_1995,N_2813);
or U7991 (N_7991,N_586,N_1235);
nand U7992 (N_7992,N_4672,N_5216);
or U7993 (N_7993,N_4593,N_4434);
and U7994 (N_7994,N_365,N_4715);
and U7995 (N_7995,N_2040,N_2916);
nor U7996 (N_7996,N_305,N_5610);
or U7997 (N_7997,N_272,N_5454);
nor U7998 (N_7998,N_3107,N_4622);
and U7999 (N_7999,N_5816,N_854);
nand U8000 (N_8000,N_3570,N_3729);
and U8001 (N_8001,N_2880,N_992);
or U8002 (N_8002,N_3847,N_4152);
nor U8003 (N_8003,N_385,N_449);
and U8004 (N_8004,N_3491,N_2490);
nand U8005 (N_8005,N_4193,N_1553);
xnor U8006 (N_8006,N_3487,N_3035);
nand U8007 (N_8007,N_3616,N_4268);
xor U8008 (N_8008,N_4346,N_1690);
nor U8009 (N_8009,N_4030,N_5982);
nor U8010 (N_8010,N_3718,N_1721);
or U8011 (N_8011,N_3535,N_33);
or U8012 (N_8012,N_4742,N_1992);
and U8013 (N_8013,N_3768,N_5693);
or U8014 (N_8014,N_2281,N_1515);
and U8015 (N_8015,N_3433,N_858);
or U8016 (N_8016,N_4551,N_32);
nand U8017 (N_8017,N_2117,N_5630);
nand U8018 (N_8018,N_4514,N_1859);
nand U8019 (N_8019,N_2496,N_2456);
nand U8020 (N_8020,N_2724,N_3940);
nor U8021 (N_8021,N_314,N_1508);
and U8022 (N_8022,N_2626,N_4919);
nor U8023 (N_8023,N_5262,N_2418);
or U8024 (N_8024,N_2015,N_3390);
xnor U8025 (N_8025,N_5352,N_4354);
nand U8026 (N_8026,N_642,N_5455);
or U8027 (N_8027,N_2029,N_5790);
nand U8028 (N_8028,N_2348,N_3819);
nor U8029 (N_8029,N_3456,N_6234);
nor U8030 (N_8030,N_909,N_2217);
nand U8031 (N_8031,N_2053,N_4928);
or U8032 (N_8032,N_1801,N_359);
xnor U8033 (N_8033,N_6170,N_1379);
and U8034 (N_8034,N_2299,N_1046);
and U8035 (N_8035,N_3738,N_4312);
nand U8036 (N_8036,N_5768,N_6028);
nand U8037 (N_8037,N_3509,N_1783);
nor U8038 (N_8038,N_6046,N_2654);
nor U8039 (N_8039,N_5915,N_3797);
nor U8040 (N_8040,N_4128,N_2030);
xnor U8041 (N_8041,N_4039,N_6223);
nor U8042 (N_8042,N_3842,N_4264);
or U8043 (N_8043,N_4289,N_1130);
and U8044 (N_8044,N_2455,N_3151);
or U8045 (N_8045,N_2031,N_2712);
or U8046 (N_8046,N_274,N_3798);
and U8047 (N_8047,N_905,N_116);
or U8048 (N_8048,N_3663,N_1631);
and U8049 (N_8049,N_3391,N_3091);
nor U8050 (N_8050,N_3358,N_1621);
nor U8051 (N_8051,N_4284,N_2882);
or U8052 (N_8052,N_2527,N_3208);
nand U8053 (N_8053,N_3966,N_3120);
nor U8054 (N_8054,N_514,N_1103);
or U8055 (N_8055,N_4626,N_4505);
and U8056 (N_8056,N_4482,N_5918);
or U8057 (N_8057,N_1889,N_4270);
nand U8058 (N_8058,N_1784,N_3447);
or U8059 (N_8059,N_2547,N_5577);
or U8060 (N_8060,N_5617,N_284);
and U8061 (N_8061,N_1068,N_4938);
xor U8062 (N_8062,N_1984,N_5703);
nand U8063 (N_8063,N_954,N_1098);
nor U8064 (N_8064,N_697,N_5421);
or U8065 (N_8065,N_776,N_1253);
and U8066 (N_8066,N_4035,N_6096);
nand U8067 (N_8067,N_2181,N_3669);
or U8068 (N_8068,N_4674,N_5897);
and U8069 (N_8069,N_755,N_1219);
or U8070 (N_8070,N_1155,N_1974);
nand U8071 (N_8071,N_2199,N_1117);
or U8072 (N_8072,N_1991,N_5486);
and U8073 (N_8073,N_4830,N_4082);
or U8074 (N_8074,N_603,N_4005);
nor U8075 (N_8075,N_4204,N_4004);
and U8076 (N_8076,N_1354,N_3259);
or U8077 (N_8077,N_2609,N_4172);
or U8078 (N_8078,N_1955,N_6142);
or U8079 (N_8079,N_4433,N_2614);
and U8080 (N_8080,N_4930,N_2708);
or U8081 (N_8081,N_4811,N_1182);
nand U8082 (N_8082,N_2096,N_5726);
or U8083 (N_8083,N_2450,N_406);
nor U8084 (N_8084,N_3485,N_4699);
nand U8085 (N_8085,N_3257,N_2386);
nand U8086 (N_8086,N_1935,N_4258);
nor U8087 (N_8087,N_3880,N_4872);
and U8088 (N_8088,N_5432,N_3302);
nor U8089 (N_8089,N_5042,N_5564);
nand U8090 (N_8090,N_1932,N_6034);
or U8091 (N_8091,N_2170,N_3799);
nand U8092 (N_8092,N_3466,N_5284);
nand U8093 (N_8093,N_4217,N_24);
nand U8094 (N_8094,N_4884,N_130);
nand U8095 (N_8095,N_1284,N_3037);
and U8096 (N_8096,N_4310,N_2010);
and U8097 (N_8097,N_3463,N_4048);
nand U8098 (N_8098,N_5386,N_2756);
or U8099 (N_8099,N_647,N_2051);
nand U8100 (N_8100,N_4924,N_3294);
and U8101 (N_8101,N_4297,N_5919);
nor U8102 (N_8102,N_869,N_4696);
nor U8103 (N_8103,N_2265,N_6038);
or U8104 (N_8104,N_1042,N_2631);
or U8105 (N_8105,N_2343,N_6002);
xnor U8106 (N_8106,N_1604,N_1978);
or U8107 (N_8107,N_693,N_3028);
and U8108 (N_8108,N_3507,N_877);
nor U8109 (N_8109,N_2234,N_1034);
and U8110 (N_8110,N_1597,N_3681);
or U8111 (N_8111,N_5767,N_3623);
xnor U8112 (N_8112,N_4931,N_4073);
or U8113 (N_8113,N_2755,N_3774);
nor U8114 (N_8114,N_1920,N_5863);
and U8115 (N_8115,N_2764,N_2388);
nand U8116 (N_8116,N_1485,N_702);
and U8117 (N_8117,N_4396,N_3825);
or U8118 (N_8118,N_5938,N_700);
and U8119 (N_8119,N_5337,N_5188);
nor U8120 (N_8120,N_2461,N_4061);
nor U8121 (N_8121,N_5882,N_255);
and U8122 (N_8122,N_5836,N_5678);
xnor U8123 (N_8123,N_4601,N_4923);
and U8124 (N_8124,N_1864,N_3937);
and U8125 (N_8125,N_1552,N_977);
and U8126 (N_8126,N_3581,N_1513);
nand U8127 (N_8127,N_3744,N_5794);
xnor U8128 (N_8128,N_5444,N_5117);
nor U8129 (N_8129,N_2938,N_1640);
nand U8130 (N_8130,N_1539,N_1827);
nor U8131 (N_8131,N_2250,N_2128);
nand U8132 (N_8132,N_5698,N_3031);
xor U8133 (N_8133,N_1133,N_3129);
nand U8134 (N_8134,N_5005,N_4251);
and U8135 (N_8135,N_2177,N_2579);
xor U8136 (N_8136,N_362,N_5810);
or U8137 (N_8137,N_2766,N_458);
nand U8138 (N_8138,N_1768,N_825);
nor U8139 (N_8139,N_2873,N_5965);
or U8140 (N_8140,N_4558,N_195);
nand U8141 (N_8141,N_3033,N_3423);
nand U8142 (N_8142,N_3571,N_5034);
or U8143 (N_8143,N_2738,N_6145);
nand U8144 (N_8144,N_5154,N_2632);
or U8145 (N_8145,N_4561,N_629);
or U8146 (N_8146,N_4175,N_425);
nand U8147 (N_8147,N_3359,N_4474);
nor U8148 (N_8148,N_252,N_4896);
or U8149 (N_8149,N_2252,N_1021);
or U8150 (N_8150,N_3224,N_4534);
and U8151 (N_8151,N_5166,N_3227);
or U8152 (N_8152,N_5106,N_4247);
or U8153 (N_8153,N_2934,N_1311);
nand U8154 (N_8154,N_3057,N_2852);
nor U8155 (N_8155,N_2561,N_1015);
and U8156 (N_8156,N_4670,N_3919);
or U8157 (N_8157,N_2301,N_1173);
and U8158 (N_8158,N_5378,N_5967);
xnor U8159 (N_8159,N_1773,N_5569);
or U8160 (N_8160,N_114,N_789);
nand U8161 (N_8161,N_4575,N_748);
xnor U8162 (N_8162,N_4334,N_5803);
xnor U8163 (N_8163,N_3403,N_2857);
and U8164 (N_8164,N_3152,N_5801);
nand U8165 (N_8165,N_2284,N_6080);
nand U8166 (N_8166,N_2584,N_2920);
nand U8167 (N_8167,N_2336,N_1059);
xnor U8168 (N_8168,N_3801,N_40);
nor U8169 (N_8169,N_921,N_4256);
nand U8170 (N_8170,N_54,N_4091);
and U8171 (N_8171,N_1769,N_1653);
xnor U8172 (N_8172,N_904,N_6196);
nand U8173 (N_8173,N_4416,N_6240);
and U8174 (N_8174,N_1650,N_2533);
or U8175 (N_8175,N_5618,N_4821);
nor U8176 (N_8176,N_4641,N_5802);
or U8177 (N_8177,N_5438,N_4212);
nand U8178 (N_8178,N_582,N_2244);
and U8179 (N_8179,N_4957,N_2134);
xor U8180 (N_8180,N_1265,N_4075);
nand U8181 (N_8181,N_2827,N_1431);
nor U8182 (N_8182,N_3783,N_1577);
and U8183 (N_8183,N_4499,N_26);
or U8184 (N_8184,N_5175,N_5474);
nor U8185 (N_8185,N_5366,N_1343);
nand U8186 (N_8186,N_1819,N_5466);
nand U8187 (N_8187,N_471,N_1980);
nand U8188 (N_8188,N_1036,N_4706);
xor U8189 (N_8189,N_5955,N_5360);
and U8190 (N_8190,N_719,N_1793);
nor U8191 (N_8191,N_4666,N_525);
nor U8192 (N_8192,N_947,N_5095);
xor U8193 (N_8193,N_191,N_1433);
nor U8194 (N_8194,N_3071,N_3413);
nand U8195 (N_8195,N_1994,N_3925);
or U8196 (N_8196,N_4823,N_3857);
and U8197 (N_8197,N_3460,N_5177);
xor U8198 (N_8198,N_3100,N_2082);
nor U8199 (N_8199,N_1954,N_3012);
or U8200 (N_8200,N_5294,N_608);
and U8201 (N_8201,N_2788,N_5043);
xor U8202 (N_8202,N_874,N_401);
and U8203 (N_8203,N_4421,N_350);
or U8204 (N_8204,N_1501,N_3989);
nor U8205 (N_8205,N_2731,N_4529);
nand U8206 (N_8206,N_5683,N_4968);
nand U8207 (N_8207,N_5501,N_1417);
nor U8208 (N_8208,N_3874,N_4722);
or U8209 (N_8209,N_5243,N_2459);
and U8210 (N_8210,N_6141,N_2792);
nor U8211 (N_8211,N_1619,N_5529);
nor U8212 (N_8212,N_3180,N_4761);
nand U8213 (N_8213,N_2811,N_555);
nor U8214 (N_8214,N_2541,N_3968);
nor U8215 (N_8215,N_5273,N_6151);
and U8216 (N_8216,N_1070,N_1717);
and U8217 (N_8217,N_4850,N_4525);
nand U8218 (N_8218,N_2197,N_276);
or U8219 (N_8219,N_5566,N_10);
nor U8220 (N_8220,N_3522,N_3675);
and U8221 (N_8221,N_990,N_5312);
and U8222 (N_8222,N_1901,N_4712);
nor U8223 (N_8223,N_4490,N_1404);
nor U8224 (N_8224,N_5954,N_577);
or U8225 (N_8225,N_5736,N_4556);
nand U8226 (N_8226,N_3024,N_1737);
nand U8227 (N_8227,N_4165,N_936);
nand U8228 (N_8228,N_1143,N_6119);
and U8229 (N_8229,N_2931,N_156);
nand U8230 (N_8230,N_5764,N_1201);
nand U8231 (N_8231,N_267,N_113);
and U8232 (N_8232,N_6200,N_1144);
nor U8233 (N_8233,N_136,N_5738);
and U8234 (N_8234,N_5384,N_4858);
nand U8235 (N_8235,N_4973,N_5215);
and U8236 (N_8236,N_3311,N_628);
nor U8237 (N_8237,N_752,N_922);
or U8238 (N_8238,N_2206,N_1082);
nand U8239 (N_8239,N_2854,N_2660);
nor U8240 (N_8240,N_6181,N_1459);
or U8241 (N_8241,N_5561,N_1198);
and U8242 (N_8242,N_4878,N_4687);
or U8243 (N_8243,N_3777,N_3457);
nand U8244 (N_8244,N_1270,N_3903);
nor U8245 (N_8245,N_4132,N_775);
and U8246 (N_8246,N_224,N_2696);
nor U8247 (N_8247,N_5246,N_3254);
xor U8248 (N_8248,N_3448,N_1613);
or U8249 (N_8249,N_688,N_5750);
nand U8250 (N_8250,N_2650,N_153);
nand U8251 (N_8251,N_2667,N_1957);
and U8252 (N_8252,N_110,N_1308);
nand U8253 (N_8253,N_4313,N_2468);
nand U8254 (N_8254,N_1125,N_1643);
and U8255 (N_8255,N_5036,N_1697);
or U8256 (N_8256,N_5068,N_4758);
and U8257 (N_8257,N_3261,N_1176);
and U8258 (N_8258,N_6075,N_5306);
nor U8259 (N_8259,N_1811,N_5510);
nand U8260 (N_8260,N_2673,N_4885);
xnor U8261 (N_8261,N_1763,N_5311);
nor U8262 (N_8262,N_4391,N_3812);
or U8263 (N_8263,N_2384,N_829);
and U8264 (N_8264,N_5557,N_4178);
nor U8265 (N_8265,N_4143,N_1584);
nor U8266 (N_8266,N_2510,N_1563);
xor U8267 (N_8267,N_212,N_3410);
nor U8268 (N_8268,N_3103,N_3432);
or U8269 (N_8269,N_4360,N_1595);
and U8270 (N_8270,N_3964,N_820);
and U8271 (N_8271,N_4146,N_793);
and U8272 (N_8272,N_3998,N_4640);
or U8273 (N_8273,N_2644,N_1038);
nor U8274 (N_8274,N_955,N_4564);
xor U8275 (N_8275,N_1028,N_5242);
nor U8276 (N_8276,N_2126,N_2914);
nor U8277 (N_8277,N_1620,N_189);
nand U8278 (N_8278,N_4308,N_3126);
and U8279 (N_8279,N_1759,N_5155);
nand U8280 (N_8280,N_2084,N_5458);
nand U8281 (N_8281,N_1365,N_3247);
nand U8282 (N_8282,N_3708,N_620);
and U8283 (N_8283,N_35,N_1639);
nor U8284 (N_8284,N_2522,N_1802);
xnor U8285 (N_8285,N_1823,N_4019);
or U8286 (N_8286,N_1078,N_5020);
nand U8287 (N_8287,N_4686,N_140);
nand U8288 (N_8288,N_5028,N_5551);
and U8289 (N_8289,N_1710,N_3615);
nand U8290 (N_8290,N_4423,N_447);
nand U8291 (N_8291,N_0,N_880);
and U8292 (N_8292,N_339,N_4852);
and U8293 (N_8293,N_2216,N_3679);
nor U8294 (N_8294,N_2221,N_3747);
nand U8295 (N_8295,N_3609,N_4215);
and U8296 (N_8296,N_951,N_540);
and U8297 (N_8297,N_2674,N_3695);
and U8298 (N_8298,N_1204,N_5231);
and U8299 (N_8299,N_5489,N_843);
nor U8300 (N_8300,N_6067,N_6015);
nand U8301 (N_8301,N_1005,N_5730);
and U8302 (N_8302,N_3374,N_3981);
nand U8303 (N_8303,N_588,N_6219);
and U8304 (N_8304,N_4378,N_2207);
nand U8305 (N_8305,N_5591,N_1772);
nor U8306 (N_8306,N_928,N_1775);
and U8307 (N_8307,N_4964,N_3551);
or U8308 (N_8308,N_3735,N_1215);
nor U8309 (N_8309,N_4834,N_5922);
or U8310 (N_8310,N_3084,N_3692);
or U8311 (N_8311,N_2785,N_2801);
or U8312 (N_8312,N_5931,N_3078);
and U8313 (N_8313,N_594,N_3159);
nor U8314 (N_8314,N_6041,N_4803);
nor U8315 (N_8315,N_5152,N_5415);
and U8316 (N_8316,N_3362,N_2024);
and U8317 (N_8317,N_2643,N_47);
and U8318 (N_8318,N_1426,N_5102);
xnor U8319 (N_8319,N_5970,N_583);
nor U8320 (N_8320,N_635,N_1562);
nor U8321 (N_8321,N_1824,N_672);
or U8322 (N_8322,N_5077,N_5158);
nand U8323 (N_8323,N_2800,N_4667);
and U8324 (N_8324,N_3574,N_1913);
and U8325 (N_8325,N_1818,N_4837);
nand U8326 (N_8326,N_3397,N_2130);
nor U8327 (N_8327,N_5923,N_4466);
nor U8328 (N_8328,N_651,N_3629);
nor U8329 (N_8329,N_1723,N_3545);
nor U8330 (N_8330,N_5668,N_2120);
and U8331 (N_8331,N_4865,N_3760);
nand U8332 (N_8332,N_4903,N_1166);
xor U8333 (N_8333,N_5310,N_809);
or U8334 (N_8334,N_5951,N_533);
nand U8335 (N_8335,N_1961,N_5059);
or U8336 (N_8336,N_131,N_5878);
nand U8337 (N_8337,N_182,N_5162);
and U8338 (N_8338,N_4527,N_2606);
nand U8339 (N_8339,N_3526,N_3888);
or U8340 (N_8340,N_3746,N_5392);
or U8341 (N_8341,N_5070,N_3203);
nand U8342 (N_8342,N_5716,N_4469);
nand U8343 (N_8343,N_2610,N_679);
and U8344 (N_8344,N_2270,N_3727);
nand U8345 (N_8345,N_1830,N_3497);
or U8346 (N_8346,N_3328,N_2580);
nand U8347 (N_8347,N_618,N_5001);
xor U8348 (N_8348,N_4192,N_1013);
or U8349 (N_8349,N_2193,N_5308);
and U8350 (N_8350,N_4511,N_3206);
nor U8351 (N_8351,N_5871,N_4658);
xor U8352 (N_8352,N_2611,N_1469);
xor U8353 (N_8353,N_504,N_2675);
and U8354 (N_8354,N_4882,N_1080);
nor U8355 (N_8355,N_578,N_5252);
nand U8356 (N_8356,N_6089,N_1405);
nor U8357 (N_8357,N_1249,N_6069);
or U8358 (N_8358,N_3296,N_3890);
or U8359 (N_8359,N_1389,N_2750);
xnor U8360 (N_8360,N_2440,N_2267);
nand U8361 (N_8361,N_4507,N_1338);
and U8362 (N_8362,N_6130,N_1241);
or U8363 (N_8363,N_4965,N_5490);
nand U8364 (N_8364,N_243,N_800);
or U8365 (N_8365,N_2465,N_939);
nand U8366 (N_8366,N_325,N_3153);
nand U8367 (N_8367,N_1423,N_2594);
nand U8368 (N_8368,N_6054,N_2102);
nor U8369 (N_8369,N_484,N_5129);
or U8370 (N_8370,N_5538,N_5524);
nor U8371 (N_8371,N_713,N_2539);
or U8372 (N_8372,N_2507,N_3061);
nand U8373 (N_8373,N_200,N_3258);
and U8374 (N_8374,N_910,N_2209);
xor U8375 (N_8375,N_3076,N_5637);
and U8376 (N_8376,N_384,N_5785);
or U8377 (N_8377,N_3598,N_2285);
or U8378 (N_8378,N_760,N_960);
or U8379 (N_8379,N_821,N_5226);
and U8380 (N_8380,N_2617,N_3420);
nand U8381 (N_8381,N_2437,N_4548);
or U8382 (N_8382,N_1118,N_3710);
or U8383 (N_8383,N_2203,N_5615);
or U8384 (N_8384,N_3367,N_991);
and U8385 (N_8385,N_4580,N_44);
or U8386 (N_8386,N_3364,N_1670);
nand U8387 (N_8387,N_1482,N_5056);
or U8388 (N_8388,N_3268,N_1460);
nor U8389 (N_8389,N_3569,N_2013);
nor U8390 (N_8390,N_732,N_5992);
nor U8391 (N_8391,N_4912,N_4736);
or U8392 (N_8392,N_2333,N_2247);
xnor U8393 (N_8393,N_5372,N_1067);
or U8394 (N_8394,N_3843,N_4813);
nand U8395 (N_8395,N_2452,N_4017);
nor U8396 (N_8396,N_4343,N_4628);
or U8397 (N_8397,N_2115,N_474);
or U8398 (N_8398,N_2982,N_2551);
nand U8399 (N_8399,N_5316,N_3292);
nor U8400 (N_8400,N_5371,N_2980);
nand U8401 (N_8401,N_5649,N_4745);
or U8402 (N_8402,N_1139,N_896);
or U8403 (N_8403,N_68,N_2291);
and U8404 (N_8404,N_5526,N_2222);
or U8405 (N_8405,N_1519,N_2262);
nand U8406 (N_8406,N_1007,N_791);
xor U8407 (N_8407,N_3032,N_1185);
nor U8408 (N_8408,N_2501,N_5165);
or U8409 (N_8409,N_5685,N_5452);
and U8410 (N_8410,N_2847,N_5182);
and U8411 (N_8411,N_808,N_1808);
nor U8412 (N_8412,N_1888,N_4024);
and U8413 (N_8413,N_706,N_1799);
and U8414 (N_8414,N_4420,N_6117);
nand U8415 (N_8415,N_520,N_822);
nor U8416 (N_8416,N_1400,N_6115);
or U8417 (N_8417,N_3375,N_4357);
and U8418 (N_8418,N_3324,N_3338);
or U8419 (N_8419,N_1862,N_3226);
nor U8420 (N_8420,N_2413,N_2544);
or U8421 (N_8421,N_3688,N_645);
nor U8422 (N_8422,N_4229,N_1504);
or U8423 (N_8423,N_5271,N_1140);
xnor U8424 (N_8424,N_3412,N_1718);
or U8425 (N_8425,N_5752,N_4272);
and U8426 (N_8426,N_4232,N_1382);
nor U8427 (N_8427,N_52,N_4613);
nor U8428 (N_8428,N_888,N_3322);
nor U8429 (N_8429,N_2434,N_1136);
and U8430 (N_8430,N_277,N_1114);
nor U8431 (N_8431,N_4584,N_4772);
xnor U8432 (N_8432,N_4892,N_3363);
and U8433 (N_8433,N_5434,N_2140);
nand U8434 (N_8434,N_849,N_1946);
and U8435 (N_8435,N_6060,N_637);
or U8436 (N_8436,N_3542,N_6107);
nor U8437 (N_8437,N_868,N_1970);
nand U8438 (N_8438,N_3586,N_5619);
and U8439 (N_8439,N_3552,N_515);
and U8440 (N_8440,N_1659,N_5440);
and U8441 (N_8441,N_2669,N_202);
nand U8442 (N_8442,N_5834,N_480);
xnor U8443 (N_8443,N_1290,N_5107);
nor U8444 (N_8444,N_5362,N_649);
xor U8445 (N_8445,N_2249,N_4058);
or U8446 (N_8446,N_3050,N_3395);
and U8447 (N_8447,N_5943,N_2081);
nor U8448 (N_8448,N_4098,N_3396);
or U8449 (N_8449,N_3849,N_2681);
nor U8450 (N_8450,N_2686,N_4424);
and U8451 (N_8451,N_4252,N_867);
nor U8452 (N_8452,N_341,N_559);
nor U8453 (N_8453,N_1998,N_2663);
and U8454 (N_8454,N_3260,N_4095);
and U8455 (N_8455,N_5426,N_2749);
xor U8456 (N_8456,N_1207,N_386);
or U8457 (N_8457,N_3745,N_1655);
xor U8458 (N_8458,N_4371,N_1725);
or U8459 (N_8459,N_3215,N_2999);
or U8460 (N_8460,N_5712,N_3405);
or U8461 (N_8461,N_5903,N_3765);
nor U8462 (N_8462,N_6192,N_4382);
nor U8463 (N_8463,N_4673,N_4921);
or U8464 (N_8464,N_4322,N_1916);
or U8465 (N_8465,N_1407,N_3877);
and U8466 (N_8466,N_5473,N_83);
nor U8467 (N_8467,N_1600,N_2391);
xnor U8468 (N_8468,N_511,N_3806);
and U8469 (N_8469,N_2150,N_3613);
xor U8470 (N_8470,N_1441,N_3789);
nand U8471 (N_8471,N_2454,N_3978);
xnor U8472 (N_8472,N_485,N_5663);
and U8473 (N_8473,N_3442,N_372);
and U8474 (N_8474,N_6231,N_694);
nand U8475 (N_8475,N_2760,N_2965);
or U8476 (N_8476,N_1658,N_3063);
or U8477 (N_8477,N_4947,N_3285);
nor U8478 (N_8478,N_4603,N_1654);
or U8479 (N_8479,N_3541,N_2936);
nor U8480 (N_8480,N_3089,N_2595);
or U8481 (N_8481,N_1881,N_2155);
and U8482 (N_8482,N_2311,N_1637);
nand U8483 (N_8483,N_506,N_1897);
or U8484 (N_8484,N_3039,N_1792);
or U8485 (N_8485,N_1789,N_1630);
or U8486 (N_8486,N_2699,N_4135);
nor U8487 (N_8487,N_427,N_75);
or U8488 (N_8488,N_725,N_2092);
nor U8489 (N_8489,N_5796,N_4765);
nor U8490 (N_8490,N_3878,N_2060);
nand U8491 (N_8491,N_1009,N_6220);
nor U8492 (N_8492,N_4400,N_2036);
xnor U8493 (N_8493,N_3233,N_2310);
and U8494 (N_8494,N_34,N_1186);
and U8495 (N_8495,N_5330,N_2987);
or U8496 (N_8496,N_3833,N_3725);
or U8497 (N_8497,N_6023,N_4412);
and U8498 (N_8498,N_2442,N_4236);
or U8499 (N_8499,N_3771,N_2969);
or U8500 (N_8500,N_2242,N_4350);
or U8501 (N_8501,N_4452,N_3638);
or U8502 (N_8502,N_1458,N_2831);
nor U8503 (N_8503,N_4513,N_1828);
nand U8504 (N_8504,N_4009,N_3195);
nor U8505 (N_8505,N_4863,N_1371);
nand U8506 (N_8506,N_3043,N_2861);
and U8507 (N_8507,N_2017,N_914);
nand U8508 (N_8508,N_3299,N_3703);
nor U8509 (N_8509,N_4324,N_5549);
nor U8510 (N_8510,N_2525,N_5133);
and U8511 (N_8511,N_5031,N_4043);
and U8512 (N_8512,N_2707,N_3660);
nand U8513 (N_8513,N_2862,N_2003);
and U8514 (N_8514,N_159,N_916);
nor U8515 (N_8515,N_5011,N_1624);
and U8516 (N_8516,N_2059,N_2568);
nand U8517 (N_8517,N_3264,N_5389);
or U8518 (N_8518,N_3646,N_4056);
nor U8519 (N_8519,N_5398,N_101);
nor U8520 (N_8520,N_2979,N_1791);
and U8521 (N_8521,N_5927,N_3557);
or U8522 (N_8522,N_5710,N_4436);
nand U8523 (N_8523,N_4972,N_6218);
or U8524 (N_8524,N_4571,N_3641);
xor U8525 (N_8525,N_5240,N_5478);
nand U8526 (N_8526,N_5600,N_4786);
or U8527 (N_8527,N_5085,N_57);
nand U8528 (N_8528,N_6165,N_3639);
nand U8529 (N_8529,N_3290,N_1810);
or U8530 (N_8530,N_3086,N_1740);
nand U8531 (N_8531,N_479,N_1252);
and U8532 (N_8532,N_1000,N_5727);
or U8533 (N_8533,N_4979,N_1020);
and U8534 (N_8534,N_1242,N_5880);
or U8535 (N_8535,N_3779,N_2714);
nor U8536 (N_8536,N_2954,N_2711);
nand U8537 (N_8537,N_6166,N_4773);
nand U8538 (N_8538,N_5889,N_2924);
nor U8539 (N_8539,N_3995,N_5988);
nor U8540 (N_8540,N_5322,N_685);
xor U8541 (N_8541,N_4624,N_1479);
or U8542 (N_8542,N_2240,N_4235);
nand U8543 (N_8543,N_126,N_432);
and U8544 (N_8544,N_1666,N_3343);
or U8545 (N_8545,N_3110,N_5869);
nor U8546 (N_8546,N_5066,N_270);
nand U8547 (N_8547,N_3287,N_6127);
and U8548 (N_8548,N_4188,N_4016);
nor U8549 (N_8549,N_5045,N_1263);
or U8550 (N_8550,N_3804,N_6008);
and U8551 (N_8551,N_3500,N_4074);
nor U8552 (N_8552,N_408,N_3150);
nand U8553 (N_8553,N_3316,N_263);
nor U8554 (N_8554,N_6226,N_1222);
nand U8555 (N_8555,N_1100,N_1197);
xor U8556 (N_8556,N_1728,N_2195);
or U8557 (N_8557,N_4550,N_4099);
nor U8558 (N_8558,N_197,N_5976);
and U8559 (N_8559,N_5053,N_5509);
nand U8560 (N_8560,N_6164,N_3398);
or U8561 (N_8561,N_4594,N_3772);
or U8562 (N_8562,N_2415,N_4198);
and U8563 (N_8563,N_1490,N_546);
and U8564 (N_8564,N_4221,N_3707);
xnor U8565 (N_8565,N_2529,N_5300);
nand U8566 (N_8566,N_2761,N_1607);
nor U8567 (N_8567,N_3589,N_2451);
nor U8568 (N_8568,N_1239,N_5961);
nor U8569 (N_8569,N_5819,N_5236);
and U8570 (N_8570,N_483,N_3826);
or U8571 (N_8571,N_3475,N_5160);
or U8572 (N_8572,N_720,N_4756);
nand U8573 (N_8573,N_943,N_632);
nand U8574 (N_8574,N_2818,N_1395);
and U8575 (N_8575,N_3350,N_4432);
and U8576 (N_8576,N_1940,N_2023);
and U8577 (N_8577,N_466,N_28);
nor U8578 (N_8578,N_5232,N_4010);
or U8579 (N_8579,N_1324,N_5413);
nand U8580 (N_8580,N_5814,N_5567);
nand U8581 (N_8581,N_2612,N_117);
nand U8582 (N_8582,N_4238,N_1312);
xor U8583 (N_8583,N_169,N_3065);
and U8584 (N_8584,N_4770,N_782);
or U8585 (N_8585,N_402,N_599);
xnor U8586 (N_8586,N_3157,N_2105);
nor U8587 (N_8587,N_1891,N_5926);
or U8588 (N_8588,N_6045,N_3730);
nand U8589 (N_8589,N_4909,N_261);
nor U8590 (N_8590,N_5747,N_4485);
or U8591 (N_8591,N_2268,N_6162);
nor U8592 (N_8592,N_3530,N_3428);
and U8593 (N_8593,N_6024,N_612);
xnor U8594 (N_8594,N_1321,N_5024);
and U8595 (N_8595,N_2065,N_1168);
xor U8596 (N_8596,N_1907,N_5611);
nand U8597 (N_8597,N_2504,N_1432);
xor U8598 (N_8598,N_5886,N_1157);
and U8599 (N_8599,N_4439,N_2136);
nor U8600 (N_8600,N_5864,N_5142);
or U8601 (N_8601,N_2277,N_5506);
nor U8602 (N_8602,N_1096,N_6121);
and U8603 (N_8603,N_4537,N_1842);
nand U8604 (N_8604,N_968,N_5523);
nand U8605 (N_8605,N_5877,N_3353);
nor U8606 (N_8606,N_1141,N_5247);
and U8607 (N_8607,N_2704,N_4702);
nor U8608 (N_8608,N_407,N_1750);
nand U8609 (N_8609,N_3274,N_4453);
xnor U8610 (N_8610,N_3119,N_6007);
nand U8611 (N_8611,N_4038,N_3938);
or U8612 (N_8612,N_1590,N_1847);
nand U8613 (N_8613,N_148,N_2009);
nor U8614 (N_8614,N_3067,N_5482);
or U8615 (N_8615,N_3958,N_4029);
nand U8616 (N_8616,N_2562,N_3697);
nand U8617 (N_8617,N_2314,N_1855);
or U8618 (N_8618,N_4790,N_5261);
or U8619 (N_8619,N_5568,N_5993);
or U8620 (N_8620,N_4101,N_886);
xnor U8621 (N_8621,N_5331,N_2325);
and U8622 (N_8622,N_2387,N_2049);
xor U8623 (N_8623,N_1079,N_6006);
nor U8624 (N_8624,N_2045,N_2554);
or U8625 (N_8625,N_5713,N_329);
nand U8626 (N_8626,N_413,N_4782);
xnor U8627 (N_8627,N_4894,N_4945);
or U8628 (N_8628,N_4867,N_315);
xnor U8629 (N_8629,N_5998,N_5496);
nand U8630 (N_8630,N_5908,N_271);
nand U8631 (N_8631,N_2721,N_5178);
and U8632 (N_8632,N_2956,N_5771);
nor U8633 (N_8633,N_1062,N_220);
nand U8634 (N_8634,N_2923,N_1826);
or U8635 (N_8635,N_5234,N_4812);
xor U8636 (N_8636,N_2613,N_5448);
and U8637 (N_8637,N_5584,N_1528);
or U8638 (N_8638,N_5598,N_938);
and U8639 (N_8639,N_5692,N_610);
nor U8640 (N_8640,N_3520,N_1467);
nand U8641 (N_8641,N_192,N_3548);
xnor U8642 (N_8642,N_1316,N_5090);
xnor U8643 (N_8643,N_2149,N_5420);
nand U8644 (N_8644,N_3049,N_3705);
or U8645 (N_8645,N_876,N_2683);
nor U8646 (N_8646,N_2628,N_3269);
and U8647 (N_8647,N_3778,N_5647);
nor U8648 (N_8648,N_2900,N_1409);
nor U8649 (N_8649,N_718,N_107);
and U8650 (N_8650,N_3785,N_5376);
nor U8651 (N_8651,N_1677,N_4679);
nand U8652 (N_8652,N_4274,N_1872);
nand U8653 (N_8653,N_5760,N_3930);
and U8654 (N_8654,N_5672,N_4089);
or U8655 (N_8655,N_210,N_266);
or U8656 (N_8656,N_5230,N_1188);
nand U8657 (N_8657,N_1582,N_2767);
nand U8658 (N_8658,N_5419,N_5818);
nand U8659 (N_8659,N_1852,N_3030);
nor U8660 (N_8660,N_2803,N_5856);
or U8661 (N_8661,N_532,N_4426);
or U8662 (N_8662,N_3347,N_1329);
nand U8663 (N_8663,N_2404,N_5120);
or U8664 (N_8664,N_5156,N_5939);
nand U8665 (N_8665,N_1236,N_2832);
and U8666 (N_8666,N_3755,N_5817);
or U8667 (N_8667,N_4688,N_3304);
nand U8668 (N_8668,N_2251,N_3386);
nand U8669 (N_8669,N_5633,N_1598);
nor U8670 (N_8670,N_1437,N_2239);
nand U8671 (N_8671,N_1902,N_4413);
nand U8672 (N_8672,N_5445,N_3829);
or U8673 (N_8673,N_5007,N_5613);
nor U8674 (N_8674,N_2564,N_2143);
nand U8675 (N_8675,N_5671,N_3207);
nor U8676 (N_8676,N_958,N_6246);
and U8677 (N_8677,N_1569,N_1673);
or U8678 (N_8678,N_2904,N_4107);
nand U8679 (N_8679,N_5441,N_4648);
and U8680 (N_8680,N_4440,N_3135);
nand U8681 (N_8681,N_5978,N_3544);
nand U8682 (N_8682,N_6005,N_4898);
nor U8683 (N_8683,N_2698,N_4908);
xnor U8684 (N_8684,N_1968,N_5083);
nor U8685 (N_8685,N_1779,N_4363);
and U8686 (N_8686,N_1374,N_767);
nor U8687 (N_8687,N_139,N_2438);
nand U8688 (N_8688,N_2192,N_2836);
or U8689 (N_8689,N_1870,N_2154);
nor U8690 (N_8690,N_1838,N_1420);
nand U8691 (N_8691,N_4541,N_5393);
and U8692 (N_8692,N_575,N_5558);
or U8693 (N_8693,N_1291,N_1293);
nor U8694 (N_8694,N_5974,N_3066);
and U8695 (N_8695,N_3600,N_4750);
nand U8696 (N_8696,N_1691,N_2929);
and U8697 (N_8697,N_5181,N_4457);
nor U8698 (N_8698,N_4565,N_883);
nand U8699 (N_8699,N_3453,N_112);
nand U8700 (N_8700,N_2903,N_2043);
and U8701 (N_8701,N_5904,N_5033);
or U8702 (N_8702,N_3194,N_1873);
and U8703 (N_8703,N_3138,N_3900);
and U8704 (N_8704,N_5655,N_3320);
nand U8705 (N_8705,N_4977,N_4995);
xnor U8706 (N_8706,N_4319,N_2802);
nor U8707 (N_8707,N_238,N_6114);
nand U8708 (N_8708,N_2374,N_3013);
nand U8709 (N_8709,N_3377,N_5762);
or U8710 (N_8710,N_422,N_4381);
xor U8711 (N_8711,N_859,N_3587);
or U8712 (N_8712,N_2,N_5645);
and U8713 (N_8713,N_380,N_1216);
xnor U8714 (N_8714,N_5646,N_2399);
nor U8715 (N_8715,N_1798,N_1039);
nand U8716 (N_8716,N_3168,N_5797);
nand U8717 (N_8717,N_4344,N_3307);
and U8718 (N_8718,N_1327,N_1636);
nand U8719 (N_8719,N_5599,N_96);
nor U8720 (N_8720,N_5511,N_2944);
xnor U8721 (N_8721,N_3676,N_4025);
nand U8722 (N_8722,N_2352,N_6135);
nor U8723 (N_8723,N_6083,N_727);
and U8724 (N_8724,N_2997,N_734);
nand U8725 (N_8725,N_3752,N_3882);
xor U8726 (N_8726,N_4023,N_2601);
or U8727 (N_8727,N_1233,N_470);
nand U8728 (N_8728,N_1581,N_1726);
nand U8729 (N_8729,N_3146,N_2810);
nand U8730 (N_8730,N_2524,N_4684);
nand U8731 (N_8731,N_5200,N_5850);
or U8732 (N_8732,N_3337,N_759);
xnor U8733 (N_8733,N_1192,N_2361);
nand U8734 (N_8734,N_4557,N_5876);
or U8735 (N_8735,N_4458,N_5804);
nor U8736 (N_8736,N_3341,N_1861);
and U8737 (N_8737,N_3899,N_2915);
nor U8738 (N_8738,N_327,N_3452);
nor U8739 (N_8739,N_1875,N_2370);
xnor U8740 (N_8740,N_5900,N_2497);
and U8741 (N_8741,N_1575,N_3451);
nand U8742 (N_8742,N_1694,N_1572);
or U8743 (N_8743,N_2257,N_4795);
nor U8744 (N_8744,N_862,N_4522);
and U8745 (N_8745,N_3479,N_1221);
nor U8746 (N_8746,N_2366,N_1929);
or U8747 (N_8747,N_6159,N_1790);
or U8748 (N_8748,N_3985,N_3284);
nor U8749 (N_8749,N_5602,N_4104);
or U8750 (N_8750,N_2616,N_5849);
and U8751 (N_8751,N_4644,N_2817);
or U8752 (N_8752,N_1048,N_3840);
nand U8753 (N_8753,N_5153,N_5446);
nand U8754 (N_8754,N_6012,N_1352);
and U8755 (N_8755,N_1681,N_4370);
nor U8756 (N_8756,N_2403,N_2444);
nand U8757 (N_8757,N_6202,N_3939);
nand U8758 (N_8758,N_3835,N_3554);
nor U8759 (N_8759,N_1008,N_3077);
or U8760 (N_8760,N_4368,N_5409);
xor U8761 (N_8761,N_926,N_5275);
nand U8762 (N_8762,N_2329,N_204);
nor U8763 (N_8763,N_412,N_6112);
nand U8764 (N_8764,N_3027,N_5966);
nand U8765 (N_8765,N_2445,N_495);
and U8766 (N_8766,N_5113,N_989);
or U8767 (N_8767,N_3097,N_3837);
and U8768 (N_8768,N_2089,N_1696);
or U8769 (N_8769,N_5670,N_5460);
nand U8770 (N_8770,N_4385,N_5962);
or U8771 (N_8771,N_944,N_3002);
or U8772 (N_8772,N_840,N_3069);
or U8773 (N_8773,N_4970,N_5575);
and U8774 (N_8774,N_2713,N_842);
or U8775 (N_8775,N_4330,N_931);
or U8776 (N_8776,N_48,N_3991);
or U8777 (N_8777,N_3654,N_5276);
and U8778 (N_8778,N_2101,N_4454);
xor U8779 (N_8779,N_4183,N_5780);
nand U8780 (N_8780,N_280,N_5627);
and U8781 (N_8781,N_2464,N_2479);
nor U8782 (N_8782,N_4283,N_2550);
and U8783 (N_8783,N_1475,N_2378);
and U8784 (N_8784,N_2077,N_1150);
xnor U8785 (N_8785,N_554,N_4422);
nor U8786 (N_8786,N_4304,N_2331);
nor U8787 (N_8787,N_1033,N_4119);
or U8788 (N_8788,N_3897,N_3904);
and U8789 (N_8789,N_2621,N_4856);
or U8790 (N_8790,N_4408,N_6197);
xor U8791 (N_8791,N_4824,N_1959);
or U8792 (N_8792,N_2863,N_2280);
nor U8793 (N_8793,N_2186,N_4692);
nor U8794 (N_8794,N_4985,N_5684);
xor U8795 (N_8795,N_1146,N_3832);
or U8796 (N_8796,N_1132,N_438);
or U8797 (N_8797,N_5323,N_1032);
and U8798 (N_8798,N_5091,N_1438);
and U8799 (N_8799,N_932,N_481);
xnor U8800 (N_8800,N_4052,N_3204);
nand U8801 (N_8801,N_2368,N_2422);
or U8802 (N_8802,N_4755,N_4323);
nor U8803 (N_8803,N_4572,N_1502);
nor U8804 (N_8804,N_758,N_4521);
and U8805 (N_8805,N_168,N_4776);
or U8806 (N_8806,N_1302,N_2227);
or U8807 (N_8807,N_5541,N_2254);
nand U8808 (N_8808,N_5433,N_5355);
nand U8809 (N_8809,N_2290,N_3250);
nand U8810 (N_8810,N_1224,N_3161);
or U8811 (N_8811,N_5196,N_5786);
or U8812 (N_8812,N_2958,N_1452);
nor U8813 (N_8813,N_1366,N_1022);
and U8814 (N_8814,N_2770,N_5858);
nand U8815 (N_8815,N_1592,N_1194);
or U8816 (N_8816,N_5012,N_5320);
nand U8817 (N_8817,N_813,N_534);
xor U8818 (N_8818,N_1840,N_1200);
nor U8819 (N_8819,N_1083,N_450);
nor U8820 (N_8820,N_1463,N_728);
nor U8821 (N_8821,N_1277,N_3335);
and U8822 (N_8822,N_206,N_4203);
xnor U8823 (N_8823,N_1262,N_4544);
nor U8824 (N_8824,N_3305,N_945);
and U8825 (N_8825,N_5516,N_5896);
nor U8826 (N_8826,N_74,N_1183);
and U8827 (N_8827,N_1113,N_4377);
or U8828 (N_8828,N_3496,N_20);
nor U8829 (N_8829,N_2411,N_5027);
and U8830 (N_8830,N_59,N_4384);
or U8831 (N_8831,N_453,N_1576);
or U8832 (N_8832,N_336,N_5990);
and U8833 (N_8833,N_5751,N_240);
nand U8834 (N_8834,N_3149,N_3611);
and U8835 (N_8835,N_2123,N_3763);
or U8836 (N_8836,N_4369,N_2283);
and U8837 (N_8837,N_4389,N_1342);
xnor U8838 (N_8838,N_1754,N_1180);
and U8839 (N_8839,N_1160,N_247);
nand U8840 (N_8840,N_783,N_2421);
xor U8841 (N_8841,N_2786,N_5612);
or U8842 (N_8842,N_3566,N_1719);
nor U8843 (N_8843,N_3625,N_5267);
and U8844 (N_8844,N_6149,N_1304);
and U8845 (N_8845,N_2175,N_1996);
nand U8846 (N_8846,N_2821,N_3327);
nor U8847 (N_8847,N_5424,N_6128);
nor U8848 (N_8848,N_5044,N_2890);
nand U8849 (N_8849,N_467,N_2874);
nor U8850 (N_8850,N_3340,N_630);
nand U8851 (N_8851,N_3376,N_882);
or U8852 (N_8852,N_1525,N_5979);
nand U8853 (N_8853,N_6049,N_716);
or U8854 (N_8854,N_1159,N_864);
nor U8855 (N_8855,N_3236,N_765);
and U8856 (N_8856,N_490,N_1137);
and U8857 (N_8857,N_6111,N_2327);
nand U8858 (N_8858,N_1027,N_3884);
nand U8859 (N_8859,N_4781,N_5778);
or U8860 (N_8860,N_4067,N_1529);
nand U8861 (N_8861,N_5800,N_4202);
nand U8862 (N_8862,N_4176,N_4955);
and U8863 (N_8863,N_2218,N_161);
nor U8864 (N_8864,N_1108,N_2845);
and U8865 (N_8865,N_4301,N_3813);
nand U8866 (N_8866,N_2753,N_4566);
and U8867 (N_8867,N_5357,N_5180);
nand U8868 (N_8868,N_1336,N_4901);
and U8869 (N_8869,N_4137,N_5930);
and U8870 (N_8870,N_976,N_5893);
xor U8871 (N_8871,N_715,N_468);
nor U8872 (N_8872,N_5299,N_6193);
or U8873 (N_8873,N_2700,N_2583);
nor U8874 (N_8874,N_4142,N_4444);
or U8875 (N_8875,N_3040,N_5676);
nor U8876 (N_8876,N_3655,N_2236);
nand U8877 (N_8877,N_3935,N_9);
and U8878 (N_8878,N_5884,N_4512);
nor U8879 (N_8879,N_3742,N_4185);
or U8880 (N_8880,N_2758,N_841);
and U8881 (N_8881,N_3147,N_3415);
or U8882 (N_8882,N_1259,N_465);
nand U8883 (N_8883,N_4372,N_2775);
or U8884 (N_8884,N_2702,N_1533);
xnor U8885 (N_8885,N_1061,N_46);
nor U8886 (N_8886,N_5315,N_5130);
nor U8887 (N_8887,N_4245,N_3165);
or U8888 (N_8888,N_1457,N_430);
and U8889 (N_8889,N_4656,N_3592);
xnor U8890 (N_8890,N_696,N_3594);
nor U8891 (N_8891,N_4980,N_1989);
or U8892 (N_8892,N_3365,N_364);
nand U8893 (N_8893,N_4337,N_5535);
xnor U8894 (N_8894,N_3831,N_3523);
or U8895 (N_8895,N_4414,N_5191);
or U8896 (N_8896,N_5183,N_2834);
nand U8897 (N_8897,N_627,N_794);
xor U8898 (N_8898,N_5233,N_2145);
nand U8899 (N_8899,N_4015,N_682);
xnor U8900 (N_8900,N_1323,N_1711);
xnor U8901 (N_8901,N_2530,N_361);
or U8902 (N_8902,N_3186,N_244);
and U8903 (N_8903,N_4468,N_5368);
nor U8904 (N_8904,N_1305,N_2076);
nor U8905 (N_8905,N_3816,N_141);
nor U8906 (N_8906,N_2828,N_6035);
or U8907 (N_8907,N_1962,N_2133);
and U8908 (N_8908,N_4731,N_5522);
and U8909 (N_8909,N_1023,N_3221);
and U8910 (N_8910,N_5168,N_4302);
and U8911 (N_8911,N_4794,N_3408);
and U8912 (N_8912,N_5959,N_4070);
xnor U8913 (N_8913,N_2058,N_5186);
or U8914 (N_8914,N_5851,N_2163);
and U8915 (N_8915,N_1412,N_6088);
nor U8916 (N_8916,N_3167,N_152);
nand U8917 (N_8917,N_4663,N_5143);
xnor U8918 (N_8918,N_5827,N_3948);
or U8919 (N_8919,N_1461,N_2599);
or U8920 (N_8920,N_1774,N_5282);
nand U8921 (N_8921,N_5614,N_4720);
and U8922 (N_8922,N_98,N_2423);
nand U8923 (N_8923,N_4546,N_285);
and U8924 (N_8924,N_127,N_1152);
xnor U8925 (N_8925,N_3942,N_878);
nand U8926 (N_8926,N_3519,N_2462);
and U8927 (N_8927,N_1499,N_4645);
nor U8928 (N_8928,N_3217,N_6184);
xor U8929 (N_8929,N_2585,N_1187);
nand U8930 (N_8930,N_4388,N_2787);
xnor U8931 (N_8931,N_2684,N_1741);
and U8932 (N_8932,N_38,N_4649);
or U8933 (N_8933,N_2340,N_4740);
nor U8934 (N_8934,N_2099,N_2064);
or U8935 (N_8935,N_3220,N_2602);
and U8936 (N_8936,N_1488,N_4709);
or U8937 (N_8937,N_6022,N_4574);
and U8938 (N_8938,N_5625,N_5349);
nor U8939 (N_8939,N_3424,N_6040);
xor U8940 (N_8940,N_949,N_2516);
nand U8941 (N_8941,N_455,N_5753);
or U8942 (N_8942,N_4582,N_3329);
and U8943 (N_8943,N_2037,N_3700);
nand U8944 (N_8944,N_2552,N_5734);
nand U8945 (N_8945,N_4411,N_3249);
nand U8946 (N_8946,N_1560,N_2535);
xor U8947 (N_8947,N_5342,N_2574);
and U8948 (N_8948,N_2034,N_1495);
and U8949 (N_8949,N_3082,N_2312);
nor U8950 (N_8950,N_337,N_5520);
xor U8951 (N_8951,N_6144,N_1044);
and U8952 (N_8952,N_6133,N_1841);
nand U8953 (N_8953,N_5139,N_5505);
nor U8954 (N_8954,N_1060,N_5682);
nor U8955 (N_8955,N_875,N_6188);
or U8956 (N_8956,N_4484,N_2805);
or U8957 (N_8957,N_4563,N_687);
and U8958 (N_8958,N_1683,N_5532);
and U8959 (N_8959,N_6183,N_5721);
nand U8960 (N_8960,N_5286,N_4154);
and U8961 (N_8961,N_3790,N_2315);
nor U8962 (N_8962,N_6081,N_5263);
and U8963 (N_8963,N_6132,N_2275);
and U8964 (N_8964,N_5375,N_1272);
nand U8965 (N_8965,N_3893,N_2321);
nand U8966 (N_8966,N_6051,N_3482);
nor U8967 (N_8967,N_3006,N_5131);
nand U8968 (N_8968,N_1072,N_2489);
and U8969 (N_8969,N_1240,N_5913);
or U8970 (N_8970,N_4549,N_2765);
and U8971 (N_8971,N_4685,N_6187);
nor U8972 (N_8972,N_6124,N_5135);
nand U8973 (N_8973,N_6030,N_3852);
nor U8974 (N_8974,N_4349,N_1056);
or U8975 (N_8975,N_91,N_1174);
and U8976 (N_8976,N_3444,N_2652);
nor U8977 (N_8977,N_3134,N_1689);
nand U8978 (N_8978,N_346,N_2623);
nor U8979 (N_8979,N_1325,N_512);
and U8980 (N_8980,N_4754,N_3515);
and U8981 (N_8981,N_4403,N_1313);
nand U8982 (N_8982,N_5211,N_5170);
and U8983 (N_8983,N_3575,N_5195);
nor U8984 (N_8984,N_708,N_328);
or U8985 (N_8985,N_4448,N_1149);
or U8986 (N_8986,N_3198,N_5757);
nor U8987 (N_8987,N_5500,N_1771);
and U8988 (N_8988,N_5590,N_2002);
nand U8989 (N_8989,N_5335,N_393);
nor U8990 (N_8990,N_5603,N_1211);
xnor U8991 (N_8991,N_2573,N_1250);
xor U8992 (N_8992,N_5194,N_4333);
nand U8993 (N_8993,N_4170,N_705);
or U8994 (N_8994,N_1912,N_2795);
nor U8995 (N_8995,N_473,N_5025);
nand U8996 (N_8996,N_486,N_4034);
xor U8997 (N_8997,N_3026,N_1383);
or U8998 (N_8998,N_2715,N_2789);
and U8999 (N_8999,N_1746,N_2070);
and U9000 (N_9000,N_4293,N_2637);
and U9001 (N_9001,N_1541,N_433);
or U9002 (N_9002,N_1377,N_2860);
and U9003 (N_9003,N_5739,N_2224);
and U9004 (N_9004,N_4096,N_3775);
and U9005 (N_9005,N_999,N_245);
or U9006 (N_9006,N_390,N_1880);
nor U9007 (N_9007,N_1493,N_2035);
or U9008 (N_9008,N_4083,N_367);
or U9009 (N_9009,N_215,N_186);
or U9010 (N_9010,N_1537,N_5722);
nand U9011 (N_9011,N_4470,N_2993);
or U9012 (N_9012,N_1045,N_2823);
and U9013 (N_9013,N_5363,N_4473);
and U9014 (N_9014,N_2162,N_5159);
nor U9015 (N_9015,N_937,N_5209);
and U9016 (N_9016,N_1156,N_4974);
xnor U9017 (N_9017,N_2172,N_1210);
and U9018 (N_9018,N_3212,N_1413);
nand U9019 (N_9019,N_2141,N_3169);
nor U9020 (N_9020,N_1341,N_4053);
nor U9021 (N_9021,N_2814,N_2893);
nor U9022 (N_9022,N_174,N_6163);
and U9023 (N_9023,N_1288,N_4309);
nand U9024 (N_9024,N_227,N_2998);
and U9025 (N_9025,N_5221,N_816);
and U9026 (N_9026,N_2475,N_2622);
or U9027 (N_9027,N_6065,N_1747);
nand U9028 (N_9028,N_2897,N_2428);
and U9029 (N_9029,N_5620,N_1124);
nor U9030 (N_9030,N_6078,N_2337);
and U9031 (N_9031,N_553,N_3584);
or U9032 (N_9032,N_2050,N_2198);
and U9033 (N_9033,N_6077,N_4351);
nand U9034 (N_9034,N_2019,N_3342);
or U9035 (N_9035,N_2448,N_2676);
xor U9036 (N_9036,N_1546,N_2506);
and U9037 (N_9037,N_4130,N_2910);
nand U9038 (N_9038,N_764,N_3690);
nor U9039 (N_9039,N_2985,N_3354);
nor U9040 (N_9040,N_5518,N_358);
xor U9041 (N_9041,N_2932,N_5380);
and U9042 (N_9042,N_4011,N_317);
or U9043 (N_9043,N_4248,N_5788);
nor U9044 (N_9044,N_2401,N_3070);
nor U9045 (N_9045,N_530,N_3643);
or U9046 (N_9046,N_1085,N_4118);
or U9047 (N_9047,N_1002,N_4084);
or U9048 (N_9048,N_3865,N_2996);
and U9049 (N_9049,N_5298,N_4822);
or U9050 (N_9050,N_122,N_288);
and U9051 (N_9051,N_138,N_241);
or U9052 (N_9052,N_6229,N_4121);
or U9053 (N_9053,N_1982,N_2566);
nand U9054 (N_9054,N_1373,N_4286);
and U9055 (N_9055,N_3933,N_2142);
nand U9056 (N_9056,N_3534,N_4278);
or U9057 (N_9057,N_2856,N_1883);
or U9058 (N_9058,N_27,N_5826);
nor U9059 (N_9059,N_3822,N_4661);
nand U9060 (N_9060,N_1380,N_543);
or U9061 (N_9061,N_2917,N_1945);
or U9062 (N_9062,N_2656,N_5766);
nand U9063 (N_9063,N_5514,N_4668);
or U9064 (N_9064,N_5383,N_2901);
nor U9065 (N_9065,N_1965,N_6084);
xnor U9066 (N_9066,N_2279,N_737);
nand U9067 (N_9067,N_665,N_4157);
and U9068 (N_9068,N_2581,N_1344);
and U9069 (N_9069,N_6104,N_4819);
and U9070 (N_9070,N_170,N_426);
and U9071 (N_9071,N_3439,N_6139);
nand U9072 (N_9072,N_4520,N_3419);
nor U9073 (N_9073,N_1328,N_1439);
nor U9074 (N_9074,N_5842,N_5289);
or U9075 (N_9075,N_836,N_5503);
nand U9076 (N_9076,N_5281,N_5528);
and U9077 (N_9077,N_4542,N_3906);
or U9078 (N_9078,N_777,N_2187);
or U9079 (N_9079,N_1906,N_2075);
and U9080 (N_9080,N_4783,N_3023);
nand U9081 (N_9081,N_5828,N_4941);
or U9082 (N_9082,N_5906,N_5935);
and U9083 (N_9083,N_6201,N_4110);
or U9084 (N_9084,N_1709,N_5172);
or U9085 (N_9085,N_1794,N_394);
nand U9086 (N_9086,N_2571,N_2067);
and U9087 (N_9087,N_6156,N_5838);
xor U9088 (N_9088,N_1557,N_2180);
nor U9089 (N_9089,N_6194,N_2607);
nor U9090 (N_9090,N_1010,N_2640);
xnor U9091 (N_9091,N_2670,N_4763);
xor U9092 (N_9092,N_5910,N_5087);
or U9093 (N_9093,N_5639,N_2820);
nor U9094 (N_9094,N_233,N_4835);
nand U9095 (N_9095,N_1053,N_5105);
and U9096 (N_9096,N_4097,N_3750);
nand U9097 (N_9097,N_125,N_2467);
nor U9098 (N_9098,N_2851,N_5873);
and U9099 (N_9099,N_1522,N_1770);
nand U9100 (N_9100,N_4735,N_3630);
or U9101 (N_9101,N_3731,N_1510);
or U9102 (N_9102,N_2144,N_3672);
or U9103 (N_9103,N_3979,N_5784);
and U9104 (N_9104,N_5883,N_76);
and U9105 (N_9105,N_3115,N_1367);
or U9106 (N_9106,N_3561,N_4610);
and U9107 (N_9107,N_4960,N_209);
and U9108 (N_9108,N_6042,N_4836);
and U9109 (N_9109,N_4303,N_3585);
and U9110 (N_9110,N_4486,N_3969);
xnor U9111 (N_9111,N_5885,N_175);
or U9112 (N_9112,N_2572,N_4151);
nor U9113 (N_9113,N_39,N_2255);
or U9114 (N_9114,N_5305,N_1518);
or U9115 (N_9115,N_3309,N_1261);
nand U9116 (N_9116,N_5984,N_3102);
or U9117 (N_9117,N_1147,N_644);
or U9118 (N_9118,N_2889,N_1538);
nand U9119 (N_9119,N_1918,N_4184);
nand U9120 (N_9120,N_2271,N_6105);
or U9121 (N_9121,N_2688,N_3495);
or U9122 (N_9122,N_1585,N_3990);
nor U9123 (N_9123,N_1523,N_351);
nand U9124 (N_9124,N_2838,N_3645);
nand U9125 (N_9125,N_5235,N_4953);
xnor U9126 (N_9126,N_661,N_5171);
nor U9127 (N_9127,N_3213,N_5026);
or U9128 (N_9128,N_5537,N_13);
or U9129 (N_9129,N_683,N_4080);
or U9130 (N_9130,N_2478,N_3621);
and U9131 (N_9131,N_1279,N_2025);
and U9132 (N_9132,N_4021,N_3962);
nor U9133 (N_9133,N_1246,N_3265);
nand U9134 (N_9134,N_1307,N_366);
xor U9135 (N_9135,N_1641,N_622);
nor U9136 (N_9136,N_278,N_6066);
nand U9137 (N_9137,N_4719,N_3873);
nor U9138 (N_9138,N_3280,N_1997);
and U9139 (N_9139,N_6011,N_1588);
nor U9140 (N_9140,N_973,N_1821);
and U9141 (N_9141,N_6009,N_6099);
nand U9142 (N_9142,N_5016,N_795);
nand U9143 (N_9143,N_3190,N_4489);
nor U9144 (N_9144,N_5126,N_1675);
nor U9145 (N_9145,N_5379,N_4266);
xnor U9146 (N_9146,N_5545,N_6214);
or U9147 (N_9147,N_1275,N_2672);
nand U9148 (N_9148,N_2288,N_1025);
nor U9149 (N_9149,N_3238,N_4523);
and U9150 (N_9150,N_3538,N_5772);
or U9151 (N_9151,N_3922,N_4940);
or U9152 (N_9152,N_295,N_605);
nand U9153 (N_9153,N_1384,N_722);
nor U9154 (N_9154,N_4199,N_3384);
and U9155 (N_9155,N_5040,N_2655);
xor U9156 (N_9156,N_1882,N_3291);
nor U9157 (N_9157,N_1753,N_3278);
nand U9158 (N_9158,N_5729,N_1625);
and U9159 (N_9159,N_3911,N_811);
or U9160 (N_9160,N_1867,N_87);
or U9161 (N_9161,N_2303,N_2582);
nor U9162 (N_9162,N_5274,N_5895);
nor U9163 (N_9163,N_817,N_2957);
xor U9164 (N_9164,N_1700,N_302);
xor U9165 (N_9165,N_154,N_3139);
nand U9166 (N_9166,N_3192,N_5677);
and U9167 (N_9167,N_807,N_344);
and U9168 (N_9168,N_5210,N_579);
nand U9169 (N_9169,N_1651,N_3529);
nand U9170 (N_9170,N_5082,N_66);
nand U9171 (N_9171,N_5343,N_5831);
xor U9172 (N_9172,N_5847,N_3010);
nor U9173 (N_9173,N_1714,N_5014);
nand U9174 (N_9174,N_1966,N_2790);
and U9175 (N_9175,N_6122,N_2426);
nand U9176 (N_9176,N_6230,N_744);
or U9177 (N_9177,N_4552,N_4724);
xor U9178 (N_9178,N_3351,N_5108);
xor U9179 (N_9179,N_5405,N_3844);
nand U9180 (N_9180,N_1267,N_2567);
nor U9181 (N_9181,N_435,N_3511);
and U9182 (N_9182,N_2990,N_3109);
nand U9183 (N_9183,N_3841,N_2435);
nor U9184 (N_9184,N_1375,N_4983);
and U9185 (N_9185,N_3957,N_2328);
nor U9186 (N_9186,N_3699,N_4871);
and U9187 (N_9187,N_6242,N_4637);
and U9188 (N_9188,N_3142,N_2006);
nor U9189 (N_9189,N_4079,N_805);
or U9190 (N_9190,N_72,N_1559);
nor U9191 (N_9191,N_2441,N_5206);
nor U9192 (N_9192,N_3216,N_3739);
xnor U9193 (N_9193,N_41,N_1424);
or U9194 (N_9194,N_5519,N_2323);
and U9195 (N_9195,N_51,N_5667);
nor U9196 (N_9196,N_2124,N_3054);
or U9197 (N_9197,N_2991,N_4501);
nor U9198 (N_9198,N_2066,N_741);
nand U9199 (N_9199,N_3862,N_5192);
nor U9200 (N_9200,N_2912,N_5388);
nand U9201 (N_9201,N_6055,N_5898);
and U9202 (N_9202,N_887,N_5425);
or U9203 (N_9203,N_5485,N_4870);
nand U9204 (N_9204,N_940,N_689);
or U9205 (N_9205,N_5963,N_1698);
nand U9206 (N_9206,N_1065,N_3105);
or U9207 (N_9207,N_2830,N_2864);
nand U9208 (N_9208,N_745,N_2844);
and U9209 (N_9209,N_1987,N_2322);
and U9210 (N_9210,N_1915,N_1505);
or U9211 (N_9211,N_5981,N_3876);
nor U9212 (N_9212,N_1922,N_5208);
and U9213 (N_9213,N_1756,N_1586);
nand U9214 (N_9214,N_3803,N_2777);
or U9215 (N_9215,N_3814,N_4358);
nand U9216 (N_9216,N_5128,N_5527);
and U9217 (N_9217,N_5336,N_296);
nor U9218 (N_9218,N_264,N_1646);
nor U9219 (N_9219,N_1877,N_2347);
xor U9220 (N_9220,N_5798,N_3502);
nand U9221 (N_9221,N_5359,N_3252);
or U9222 (N_9222,N_5476,N_4404);
or U9223 (N_9223,N_513,N_4929);
or U9224 (N_9224,N_318,N_4678);
and U9225 (N_9225,N_3722,N_3762);
or U9226 (N_9226,N_4739,N_5657);
nand U9227 (N_9227,N_3262,N_1435);
or U9228 (N_9228,N_1550,N_1444);
or U9229 (N_9229,N_1674,N_6093);
or U9230 (N_9230,N_1704,N_5969);
and U9231 (N_9231,N_3811,N_4054);
nand U9232 (N_9232,N_4944,N_4138);
and U9233 (N_9233,N_2495,N_3820);
and U9234 (N_9234,N_855,N_3567);
xor U9235 (N_9235,N_994,N_4677);
and U9236 (N_9236,N_3715,N_3951);
nor U9237 (N_9237,N_3952,N_2219);
nand U9238 (N_9238,N_570,N_342);
or U9239 (N_9239,N_4214,N_1478);
nand U9240 (N_9240,N_2726,N_482);
or U9241 (N_9241,N_3896,N_669);
and U9242 (N_9242,N_1158,N_5597);
nor U9243 (N_9243,N_2038,N_4338);
or U9244 (N_9244,N_537,N_2307);
nand U9245 (N_9245,N_6000,N_1627);
nor U9246 (N_9246,N_290,N_4159);
and U9247 (N_9247,N_5010,N_638);
nand U9248 (N_9248,N_4430,N_5111);
nand U9249 (N_9249,N_1138,N_5588);
nand U9250 (N_9250,N_1055,N_5039);
and U9251 (N_9251,N_5553,N_3974);
and U9252 (N_9252,N_5080,N_2661);
nand U9253 (N_9253,N_3987,N_5279);
and U9254 (N_9254,N_2703,N_5495);
xnor U9255 (N_9255,N_2259,N_1018);
and U9256 (N_9256,N_1006,N_5190);
nand U9257 (N_9257,N_1833,N_49);
nand U9258 (N_9258,N_177,N_3578);
and U9259 (N_9259,N_3101,N_3685);
nor U9260 (N_9260,N_103,N_3914);
nor U9261 (N_9261,N_4237,N_352);
or U9262 (N_9262,N_3649,N_4988);
and U9263 (N_9263,N_104,N_3605);
nor U9264 (N_9264,N_5916,N_2408);
nor U9265 (N_9265,N_5609,N_3786);
and U9266 (N_9266,N_2093,N_293);
xor U9267 (N_9267,N_2887,N_2526);
or U9268 (N_9268,N_4177,N_3971);
or U9269 (N_9269,N_2212,N_1440);
or U9270 (N_9270,N_4887,N_3493);
nand U9271 (N_9271,N_6152,N_4817);
nor U9272 (N_9272,N_3202,N_1359);
and U9273 (N_9273,N_4134,N_160);
nand U9274 (N_9274,N_4049,N_590);
and U9275 (N_9275,N_889,N_1278);
and U9276 (N_9276,N_1734,N_2972);
xnor U9277 (N_9277,N_158,N_5364);
nor U9278 (N_9278,N_3187,N_2052);
and U9279 (N_9279,N_3450,N_319);
nand U9280 (N_9280,N_5972,N_4033);
and U9281 (N_9281,N_860,N_2598);
and U9282 (N_9282,N_4294,N_1856);
nand U9283 (N_9283,N_304,N_4050);
xor U9284 (N_9284,N_248,N_3034);
and U9285 (N_9285,N_88,N_286);
or U9286 (N_9286,N_5144,N_2966);
nand U9287 (N_9287,N_3323,N_3670);
nor U9288 (N_9288,N_3093,N_1001);
nand U9289 (N_9289,N_1073,N_847);
nand U9290 (N_9290,N_3683,N_3636);
or U9291 (N_9291,N_3409,N_1213);
xor U9292 (N_9292,N_1668,N_1999);
nand U9293 (N_9293,N_1511,N_4854);
or U9294 (N_9294,N_1973,N_378);
and U9295 (N_9295,N_1786,N_3255);
or U9296 (N_9296,N_3512,N_2588);
and U9297 (N_9297,N_4419,N_345);
and U9298 (N_9298,N_2385,N_5570);
or U9299 (N_9299,N_779,N_375);
nor U9300 (N_9300,N_249,N_1164);
or U9301 (N_9301,N_4189,N_2892);
nor U9302 (N_9302,N_2597,N_4122);
xor U9303 (N_9303,N_2894,N_5321);
and U9304 (N_9304,N_1364,N_3242);
or U9305 (N_9305,N_6031,N_392);
nor U9306 (N_9306,N_639,N_4111);
nor U9307 (N_9307,N_2233,N_2294);
or U9308 (N_9308,N_145,N_3505);
or U9309 (N_9309,N_4329,N_4124);
and U9310 (N_9310,N_1618,N_4317);
or U9311 (N_9311,N_5079,N_6082);
nand U9312 (N_9312,N_1494,N_754);
nor U9313 (N_9313,N_5163,N_4828);
xor U9314 (N_9314,N_891,N_3633);
and U9315 (N_9315,N_6029,N_5656);
and U9316 (N_9316,N_6206,N_53);
nor U9317 (N_9317,N_1724,N_1101);
nor U9318 (N_9318,N_477,N_636);
and U9319 (N_9319,N_405,N_1345);
xnor U9320 (N_9320,N_5122,N_5901);
nor U9321 (N_9321,N_1385,N_3553);
xnor U9322 (N_9322,N_4825,N_2432);
nand U9323 (N_9323,N_2425,N_294);
and U9324 (N_9324,N_2717,N_4280);
nor U9325 (N_9325,N_3489,N_6171);
or U9326 (N_9326,N_3719,N_4691);
or U9327 (N_9327,N_4869,N_4791);
nor U9328 (N_9328,N_5781,N_567);
nand U9329 (N_9329,N_597,N_2638);
nor U9330 (N_9330,N_5989,N_523);
and U9331 (N_9331,N_766,N_1707);
nand U9332 (N_9332,N_4802,N_4127);
or U9333 (N_9333,N_3029,N_1745);
or U9334 (N_9334,N_4517,N_3547);
and U9335 (N_9335,N_5220,N_2353);
nor U9336 (N_9336,N_2356,N_1633);
xnor U9337 (N_9337,N_3072,N_1075);
xnor U9338 (N_9338,N_6216,N_2028);
nor U9339 (N_9339,N_4113,N_4431);
or U9340 (N_9340,N_2484,N_740);
nand U9341 (N_9341,N_924,N_3191);
or U9342 (N_9342,N_4276,N_2196);
nor U9343 (N_9343,N_1230,N_5868);
and U9344 (N_9344,N_4629,N_4994);
or U9345 (N_9345,N_792,N_2850);
or U9346 (N_9346,N_733,N_1914);
and U9347 (N_9347,N_147,N_4427);
and U9348 (N_9348,N_176,N_993);
nor U9349 (N_9349,N_3539,N_1931);
xor U9350 (N_9350,N_5030,N_3356);
nor U9351 (N_9351,N_3369,N_3591);
and U9352 (N_9352,N_2877,N_3640);
or U9353 (N_9353,N_6101,N_3469);
and U9354 (N_9354,N_5255,N_913);
nand U9355 (N_9355,N_184,N_6061);
or U9356 (N_9356,N_946,N_6235);
nand U9357 (N_9357,N_1648,N_4866);
nor U9358 (N_9358,N_3387,N_3095);
or U9359 (N_9359,N_6221,N_5395);
nor U9360 (N_9360,N_6110,N_133);
and U9361 (N_9361,N_457,N_5517);
and U9362 (N_9362,N_4064,N_4975);
and U9363 (N_9363,N_2161,N_4966);
and U9364 (N_9364,N_1807,N_2646);
nor U9365 (N_9365,N_4133,N_6131);
or U9366 (N_9366,N_5742,N_3836);
or U9367 (N_9367,N_1401,N_3795);
and U9368 (N_9368,N_1258,N_3188);
or U9369 (N_9369,N_31,N_2558);
or U9370 (N_9370,N_2925,N_2809);
xnor U9371 (N_9371,N_50,N_5986);
or U9372 (N_9372,N_2069,N_3907);
and U9373 (N_9373,N_4365,N_222);
nand U9374 (N_9374,N_4843,N_4156);
or U9375 (N_9375,N_2058,N_1077);
and U9376 (N_9376,N_3518,N_4540);
nand U9377 (N_9377,N_5768,N_2812);
and U9378 (N_9378,N_1394,N_5111);
nand U9379 (N_9379,N_4719,N_873);
and U9380 (N_9380,N_3302,N_1656);
or U9381 (N_9381,N_5705,N_2081);
nand U9382 (N_9382,N_1293,N_5276);
or U9383 (N_9383,N_5023,N_5352);
nor U9384 (N_9384,N_1837,N_3634);
or U9385 (N_9385,N_3288,N_3531);
or U9386 (N_9386,N_3036,N_3177);
or U9387 (N_9387,N_3137,N_1272);
and U9388 (N_9388,N_3814,N_3636);
and U9389 (N_9389,N_3715,N_4673);
and U9390 (N_9390,N_2270,N_5162);
nor U9391 (N_9391,N_5504,N_4446);
nand U9392 (N_9392,N_2926,N_72);
or U9393 (N_9393,N_3541,N_720);
nand U9394 (N_9394,N_4561,N_673);
nand U9395 (N_9395,N_4567,N_2596);
or U9396 (N_9396,N_3235,N_2448);
or U9397 (N_9397,N_5555,N_3909);
or U9398 (N_9398,N_4846,N_48);
nor U9399 (N_9399,N_2118,N_2498);
or U9400 (N_9400,N_1930,N_2546);
nor U9401 (N_9401,N_2952,N_4749);
nand U9402 (N_9402,N_1226,N_2567);
nor U9403 (N_9403,N_2694,N_5883);
nor U9404 (N_9404,N_2764,N_396);
nand U9405 (N_9405,N_4897,N_3051);
nand U9406 (N_9406,N_5343,N_4916);
and U9407 (N_9407,N_3057,N_3626);
and U9408 (N_9408,N_1717,N_5281);
and U9409 (N_9409,N_1515,N_2382);
and U9410 (N_9410,N_4760,N_2031);
nor U9411 (N_9411,N_1868,N_550);
and U9412 (N_9412,N_4062,N_4671);
nor U9413 (N_9413,N_1111,N_1262);
or U9414 (N_9414,N_2102,N_4509);
nand U9415 (N_9415,N_3104,N_3082);
nand U9416 (N_9416,N_1068,N_2024);
nand U9417 (N_9417,N_1727,N_3454);
or U9418 (N_9418,N_601,N_5283);
and U9419 (N_9419,N_5657,N_1117);
and U9420 (N_9420,N_5537,N_5339);
nand U9421 (N_9421,N_1970,N_5808);
nand U9422 (N_9422,N_4694,N_3448);
or U9423 (N_9423,N_1351,N_2681);
nor U9424 (N_9424,N_4731,N_2018);
or U9425 (N_9425,N_1085,N_5881);
or U9426 (N_9426,N_3131,N_696);
nand U9427 (N_9427,N_2253,N_1297);
nor U9428 (N_9428,N_3946,N_6064);
or U9429 (N_9429,N_644,N_2737);
or U9430 (N_9430,N_3033,N_260);
nand U9431 (N_9431,N_5542,N_1926);
or U9432 (N_9432,N_5955,N_1477);
nand U9433 (N_9433,N_4357,N_3329);
nor U9434 (N_9434,N_1215,N_2668);
and U9435 (N_9435,N_5328,N_2684);
xnor U9436 (N_9436,N_116,N_214);
or U9437 (N_9437,N_4346,N_3117);
nand U9438 (N_9438,N_3922,N_3880);
xnor U9439 (N_9439,N_3970,N_1071);
and U9440 (N_9440,N_1820,N_2925);
or U9441 (N_9441,N_3825,N_3560);
xor U9442 (N_9442,N_1615,N_1553);
and U9443 (N_9443,N_1330,N_3951);
nand U9444 (N_9444,N_2140,N_5366);
and U9445 (N_9445,N_2273,N_3553);
nor U9446 (N_9446,N_1099,N_2183);
nor U9447 (N_9447,N_5494,N_4897);
xor U9448 (N_9448,N_4982,N_1495);
nor U9449 (N_9449,N_1667,N_3161);
nand U9450 (N_9450,N_3403,N_6125);
nand U9451 (N_9451,N_5487,N_2237);
nand U9452 (N_9452,N_5242,N_4946);
nor U9453 (N_9453,N_4007,N_4694);
or U9454 (N_9454,N_3594,N_425);
or U9455 (N_9455,N_1470,N_1987);
or U9456 (N_9456,N_1327,N_6110);
and U9457 (N_9457,N_378,N_3578);
nor U9458 (N_9458,N_5043,N_5787);
xnor U9459 (N_9459,N_2707,N_4827);
or U9460 (N_9460,N_4469,N_4079);
nand U9461 (N_9461,N_5344,N_2373);
and U9462 (N_9462,N_2273,N_3941);
and U9463 (N_9463,N_4865,N_3033);
and U9464 (N_9464,N_5501,N_4663);
and U9465 (N_9465,N_4402,N_3178);
nand U9466 (N_9466,N_1446,N_4549);
nand U9467 (N_9467,N_4834,N_655);
nor U9468 (N_9468,N_5003,N_2534);
and U9469 (N_9469,N_3468,N_87);
or U9470 (N_9470,N_2916,N_1160);
and U9471 (N_9471,N_5891,N_95);
nand U9472 (N_9472,N_2999,N_5784);
or U9473 (N_9473,N_3423,N_849);
or U9474 (N_9474,N_4708,N_4807);
xor U9475 (N_9475,N_6055,N_4605);
and U9476 (N_9476,N_1658,N_2906);
or U9477 (N_9477,N_6203,N_239);
nand U9478 (N_9478,N_2040,N_1598);
nand U9479 (N_9479,N_2374,N_5345);
nand U9480 (N_9480,N_2545,N_1483);
or U9481 (N_9481,N_3522,N_1136);
xnor U9482 (N_9482,N_6036,N_3620);
and U9483 (N_9483,N_2922,N_4650);
xnor U9484 (N_9484,N_5222,N_5406);
xor U9485 (N_9485,N_2982,N_5310);
nor U9486 (N_9486,N_3594,N_2984);
nor U9487 (N_9487,N_259,N_1146);
and U9488 (N_9488,N_2955,N_5094);
nor U9489 (N_9489,N_4802,N_591);
nor U9490 (N_9490,N_6104,N_1066);
nor U9491 (N_9491,N_4165,N_3478);
or U9492 (N_9492,N_3709,N_6146);
nor U9493 (N_9493,N_3463,N_951);
or U9494 (N_9494,N_5778,N_2591);
nor U9495 (N_9495,N_5715,N_4295);
nand U9496 (N_9496,N_2702,N_4216);
and U9497 (N_9497,N_4918,N_1164);
and U9498 (N_9498,N_3548,N_412);
or U9499 (N_9499,N_6045,N_4020);
or U9500 (N_9500,N_4517,N_3370);
or U9501 (N_9501,N_1404,N_4780);
xor U9502 (N_9502,N_3359,N_1543);
xnor U9503 (N_9503,N_1736,N_3450);
nand U9504 (N_9504,N_3661,N_1688);
and U9505 (N_9505,N_932,N_2264);
nor U9506 (N_9506,N_5259,N_1134);
nor U9507 (N_9507,N_1556,N_2768);
or U9508 (N_9508,N_958,N_3265);
xnor U9509 (N_9509,N_4437,N_3065);
or U9510 (N_9510,N_1679,N_4172);
nor U9511 (N_9511,N_779,N_762);
and U9512 (N_9512,N_456,N_2689);
or U9513 (N_9513,N_1930,N_1612);
and U9514 (N_9514,N_2891,N_3647);
and U9515 (N_9515,N_2052,N_3386);
nor U9516 (N_9516,N_724,N_2655);
nand U9517 (N_9517,N_6086,N_3398);
nor U9518 (N_9518,N_1782,N_2409);
nand U9519 (N_9519,N_6184,N_2316);
xor U9520 (N_9520,N_1245,N_2609);
nand U9521 (N_9521,N_884,N_267);
or U9522 (N_9522,N_6114,N_3721);
and U9523 (N_9523,N_2038,N_1372);
and U9524 (N_9524,N_4154,N_3563);
and U9525 (N_9525,N_784,N_2295);
nand U9526 (N_9526,N_2259,N_1386);
xnor U9527 (N_9527,N_5573,N_2911);
nand U9528 (N_9528,N_1614,N_5111);
and U9529 (N_9529,N_1894,N_1515);
nor U9530 (N_9530,N_1339,N_4136);
and U9531 (N_9531,N_3943,N_5232);
xnor U9532 (N_9532,N_3789,N_4118);
or U9533 (N_9533,N_2489,N_5721);
nand U9534 (N_9534,N_3536,N_2439);
nand U9535 (N_9535,N_3696,N_4501);
nand U9536 (N_9536,N_412,N_4563);
and U9537 (N_9537,N_4954,N_558);
or U9538 (N_9538,N_4559,N_4801);
xnor U9539 (N_9539,N_3896,N_4275);
or U9540 (N_9540,N_5813,N_5807);
nor U9541 (N_9541,N_425,N_6111);
and U9542 (N_9542,N_1118,N_4650);
nand U9543 (N_9543,N_2382,N_4240);
nor U9544 (N_9544,N_3471,N_3662);
nor U9545 (N_9545,N_4364,N_5284);
nand U9546 (N_9546,N_1277,N_2132);
or U9547 (N_9547,N_505,N_449);
nand U9548 (N_9548,N_3653,N_3143);
and U9549 (N_9549,N_5186,N_5683);
or U9550 (N_9550,N_4078,N_5524);
or U9551 (N_9551,N_4725,N_1787);
nand U9552 (N_9552,N_5017,N_4064);
or U9553 (N_9553,N_1165,N_2493);
xnor U9554 (N_9554,N_5812,N_5247);
nand U9555 (N_9555,N_146,N_2970);
nor U9556 (N_9556,N_3779,N_3441);
nor U9557 (N_9557,N_2154,N_2671);
nand U9558 (N_9558,N_5722,N_3148);
nor U9559 (N_9559,N_922,N_3403);
and U9560 (N_9560,N_2093,N_5366);
and U9561 (N_9561,N_1499,N_1032);
and U9562 (N_9562,N_3632,N_3394);
nor U9563 (N_9563,N_5921,N_5908);
xnor U9564 (N_9564,N_4858,N_2855);
nor U9565 (N_9565,N_3984,N_1829);
or U9566 (N_9566,N_4047,N_2272);
xnor U9567 (N_9567,N_1905,N_517);
nor U9568 (N_9568,N_1044,N_4967);
and U9569 (N_9569,N_891,N_294);
nand U9570 (N_9570,N_5000,N_4998);
nor U9571 (N_9571,N_4584,N_4603);
xnor U9572 (N_9572,N_698,N_2259);
and U9573 (N_9573,N_5948,N_194);
nor U9574 (N_9574,N_1330,N_1015);
or U9575 (N_9575,N_3673,N_5631);
nand U9576 (N_9576,N_6135,N_6221);
and U9577 (N_9577,N_1751,N_293);
and U9578 (N_9578,N_918,N_3330);
and U9579 (N_9579,N_1839,N_3831);
nand U9580 (N_9580,N_1820,N_833);
nor U9581 (N_9581,N_2788,N_4811);
nand U9582 (N_9582,N_4844,N_5179);
and U9583 (N_9583,N_4030,N_5910);
nand U9584 (N_9584,N_5338,N_849);
nor U9585 (N_9585,N_3745,N_3350);
and U9586 (N_9586,N_941,N_1998);
xnor U9587 (N_9587,N_2065,N_4338);
nor U9588 (N_9588,N_3187,N_3565);
nor U9589 (N_9589,N_5268,N_2309);
and U9590 (N_9590,N_2880,N_773);
or U9591 (N_9591,N_3114,N_1429);
nand U9592 (N_9592,N_1839,N_2938);
or U9593 (N_9593,N_4775,N_3170);
or U9594 (N_9594,N_5548,N_900);
xor U9595 (N_9595,N_2420,N_1862);
nor U9596 (N_9596,N_5207,N_2130);
nand U9597 (N_9597,N_3557,N_2606);
and U9598 (N_9598,N_4717,N_2101);
and U9599 (N_9599,N_5865,N_3592);
xnor U9600 (N_9600,N_3332,N_6234);
nor U9601 (N_9601,N_3429,N_78);
and U9602 (N_9602,N_5086,N_1933);
or U9603 (N_9603,N_1086,N_4938);
or U9604 (N_9604,N_4605,N_4391);
or U9605 (N_9605,N_2383,N_5034);
or U9606 (N_9606,N_3703,N_1106);
nand U9607 (N_9607,N_2300,N_1217);
or U9608 (N_9608,N_4245,N_6011);
and U9609 (N_9609,N_733,N_310);
nand U9610 (N_9610,N_5180,N_2389);
nor U9611 (N_9611,N_1453,N_1619);
and U9612 (N_9612,N_3158,N_4176);
nand U9613 (N_9613,N_5594,N_5686);
xor U9614 (N_9614,N_372,N_368);
or U9615 (N_9615,N_5387,N_3429);
xor U9616 (N_9616,N_2595,N_315);
nor U9617 (N_9617,N_4814,N_2354);
xor U9618 (N_9618,N_3916,N_3104);
nor U9619 (N_9619,N_2012,N_3998);
xor U9620 (N_9620,N_5417,N_2437);
or U9621 (N_9621,N_6221,N_1087);
and U9622 (N_9622,N_2178,N_5393);
and U9623 (N_9623,N_5186,N_3822);
and U9624 (N_9624,N_3109,N_4711);
nand U9625 (N_9625,N_1461,N_2792);
or U9626 (N_9626,N_5354,N_4213);
and U9627 (N_9627,N_3841,N_554);
or U9628 (N_9628,N_981,N_3582);
or U9629 (N_9629,N_4486,N_4858);
and U9630 (N_9630,N_610,N_1405);
or U9631 (N_9631,N_1673,N_4950);
or U9632 (N_9632,N_5279,N_2566);
nor U9633 (N_9633,N_5527,N_2987);
nor U9634 (N_9634,N_1548,N_2391);
and U9635 (N_9635,N_361,N_1629);
and U9636 (N_9636,N_2125,N_5144);
nand U9637 (N_9637,N_5688,N_4796);
or U9638 (N_9638,N_5040,N_1516);
nand U9639 (N_9639,N_3353,N_2487);
nor U9640 (N_9640,N_2114,N_4336);
and U9641 (N_9641,N_5255,N_3520);
xor U9642 (N_9642,N_1995,N_1926);
or U9643 (N_9643,N_5401,N_1706);
and U9644 (N_9644,N_5107,N_835);
nand U9645 (N_9645,N_6100,N_2037);
or U9646 (N_9646,N_2305,N_3404);
nor U9647 (N_9647,N_6137,N_4364);
or U9648 (N_9648,N_2028,N_3730);
nand U9649 (N_9649,N_5825,N_5863);
nand U9650 (N_9650,N_5320,N_2682);
nand U9651 (N_9651,N_4209,N_4256);
nand U9652 (N_9652,N_3756,N_4773);
or U9653 (N_9653,N_6202,N_3109);
and U9654 (N_9654,N_3035,N_4796);
or U9655 (N_9655,N_3451,N_250);
nand U9656 (N_9656,N_5094,N_2379);
and U9657 (N_9657,N_6070,N_5658);
and U9658 (N_9658,N_5372,N_558);
xor U9659 (N_9659,N_6011,N_5508);
xnor U9660 (N_9660,N_1935,N_5422);
or U9661 (N_9661,N_4673,N_1486);
xor U9662 (N_9662,N_5351,N_3905);
nand U9663 (N_9663,N_5670,N_3240);
or U9664 (N_9664,N_1951,N_665);
and U9665 (N_9665,N_4642,N_3617);
or U9666 (N_9666,N_5556,N_1068);
and U9667 (N_9667,N_3275,N_3368);
xor U9668 (N_9668,N_2534,N_1402);
nand U9669 (N_9669,N_3614,N_46);
or U9670 (N_9670,N_6170,N_107);
or U9671 (N_9671,N_4164,N_2515);
xor U9672 (N_9672,N_4817,N_2001);
and U9673 (N_9673,N_3809,N_1882);
nand U9674 (N_9674,N_5378,N_4061);
or U9675 (N_9675,N_2146,N_5207);
xor U9676 (N_9676,N_5545,N_1922);
nor U9677 (N_9677,N_3253,N_2967);
nor U9678 (N_9678,N_2095,N_1798);
nand U9679 (N_9679,N_1200,N_1649);
nand U9680 (N_9680,N_2287,N_5511);
and U9681 (N_9681,N_2385,N_4893);
nor U9682 (N_9682,N_538,N_4163);
or U9683 (N_9683,N_791,N_210);
or U9684 (N_9684,N_4919,N_3007);
nand U9685 (N_9685,N_3414,N_1419);
nor U9686 (N_9686,N_3894,N_13);
or U9687 (N_9687,N_6099,N_4504);
nor U9688 (N_9688,N_3634,N_5724);
nand U9689 (N_9689,N_6131,N_5621);
nand U9690 (N_9690,N_4894,N_3114);
or U9691 (N_9691,N_6010,N_1896);
nor U9692 (N_9692,N_2600,N_589);
xnor U9693 (N_9693,N_578,N_1139);
xor U9694 (N_9694,N_4133,N_1163);
nor U9695 (N_9695,N_5033,N_825);
or U9696 (N_9696,N_5231,N_81);
nor U9697 (N_9697,N_5159,N_1540);
or U9698 (N_9698,N_4888,N_2954);
nand U9699 (N_9699,N_84,N_4468);
and U9700 (N_9700,N_2798,N_963);
nand U9701 (N_9701,N_46,N_33);
xor U9702 (N_9702,N_1221,N_1505);
and U9703 (N_9703,N_5497,N_1766);
nor U9704 (N_9704,N_4529,N_5558);
and U9705 (N_9705,N_3999,N_4215);
nor U9706 (N_9706,N_818,N_3684);
or U9707 (N_9707,N_3475,N_4068);
and U9708 (N_9708,N_5230,N_291);
and U9709 (N_9709,N_5868,N_5736);
and U9710 (N_9710,N_3946,N_3313);
nor U9711 (N_9711,N_5127,N_5847);
nor U9712 (N_9712,N_3722,N_2935);
nor U9713 (N_9713,N_5637,N_4482);
nand U9714 (N_9714,N_3313,N_2322);
or U9715 (N_9715,N_3129,N_4598);
nand U9716 (N_9716,N_3715,N_685);
and U9717 (N_9717,N_5493,N_6222);
and U9718 (N_9718,N_1904,N_5055);
and U9719 (N_9719,N_101,N_3440);
or U9720 (N_9720,N_3057,N_2468);
and U9721 (N_9721,N_5858,N_2422);
or U9722 (N_9722,N_3978,N_6152);
and U9723 (N_9723,N_990,N_2403);
and U9724 (N_9724,N_5750,N_1218);
nand U9725 (N_9725,N_2131,N_5558);
and U9726 (N_9726,N_205,N_1791);
or U9727 (N_9727,N_1679,N_1055);
nand U9728 (N_9728,N_2133,N_1838);
xor U9729 (N_9729,N_3211,N_6096);
nand U9730 (N_9730,N_5335,N_3569);
or U9731 (N_9731,N_3804,N_5647);
and U9732 (N_9732,N_5014,N_3448);
nor U9733 (N_9733,N_1127,N_2637);
or U9734 (N_9734,N_4093,N_5135);
or U9735 (N_9735,N_5336,N_5595);
and U9736 (N_9736,N_2167,N_2445);
or U9737 (N_9737,N_4153,N_1033);
nand U9738 (N_9738,N_3760,N_488);
or U9739 (N_9739,N_2024,N_487);
or U9740 (N_9740,N_2152,N_3562);
xor U9741 (N_9741,N_405,N_4216);
nand U9742 (N_9742,N_2177,N_1654);
nand U9743 (N_9743,N_4360,N_70);
nor U9744 (N_9744,N_423,N_1148);
or U9745 (N_9745,N_6023,N_2148);
nor U9746 (N_9746,N_2362,N_131);
and U9747 (N_9747,N_148,N_3739);
or U9748 (N_9748,N_2301,N_4494);
xnor U9749 (N_9749,N_3103,N_1492);
or U9750 (N_9750,N_3237,N_4616);
nor U9751 (N_9751,N_5902,N_1012);
and U9752 (N_9752,N_1262,N_3773);
nand U9753 (N_9753,N_1852,N_1038);
or U9754 (N_9754,N_187,N_4412);
and U9755 (N_9755,N_2508,N_1038);
nand U9756 (N_9756,N_4636,N_3244);
and U9757 (N_9757,N_4164,N_2236);
xnor U9758 (N_9758,N_841,N_4555);
nand U9759 (N_9759,N_5413,N_2721);
and U9760 (N_9760,N_4740,N_5159);
nand U9761 (N_9761,N_186,N_6223);
or U9762 (N_9762,N_2845,N_2957);
nor U9763 (N_9763,N_2642,N_5177);
and U9764 (N_9764,N_1515,N_5736);
xor U9765 (N_9765,N_3896,N_1348);
xnor U9766 (N_9766,N_4601,N_599);
or U9767 (N_9767,N_243,N_2555);
or U9768 (N_9768,N_4090,N_4021);
and U9769 (N_9769,N_6053,N_3515);
or U9770 (N_9770,N_871,N_3247);
nand U9771 (N_9771,N_5851,N_5119);
or U9772 (N_9772,N_6054,N_5799);
nand U9773 (N_9773,N_4296,N_2170);
xor U9774 (N_9774,N_1157,N_1117);
and U9775 (N_9775,N_1657,N_484);
nor U9776 (N_9776,N_6150,N_5582);
or U9777 (N_9777,N_1311,N_5379);
and U9778 (N_9778,N_5465,N_1892);
nand U9779 (N_9779,N_5576,N_3468);
and U9780 (N_9780,N_4210,N_3924);
xnor U9781 (N_9781,N_1178,N_2052);
xor U9782 (N_9782,N_4158,N_5337);
nor U9783 (N_9783,N_1931,N_1724);
or U9784 (N_9784,N_53,N_4910);
nor U9785 (N_9785,N_872,N_4224);
xor U9786 (N_9786,N_1951,N_5034);
and U9787 (N_9787,N_4121,N_1462);
and U9788 (N_9788,N_3680,N_333);
nor U9789 (N_9789,N_4891,N_2839);
and U9790 (N_9790,N_4485,N_5287);
or U9791 (N_9791,N_1827,N_959);
or U9792 (N_9792,N_1645,N_3550);
nor U9793 (N_9793,N_2544,N_1518);
and U9794 (N_9794,N_3840,N_774);
and U9795 (N_9795,N_2388,N_2574);
nand U9796 (N_9796,N_5352,N_4951);
or U9797 (N_9797,N_2097,N_1861);
nor U9798 (N_9798,N_2617,N_741);
or U9799 (N_9799,N_1586,N_5261);
nor U9800 (N_9800,N_1454,N_5927);
nand U9801 (N_9801,N_2345,N_71);
and U9802 (N_9802,N_4876,N_240);
nand U9803 (N_9803,N_184,N_3620);
and U9804 (N_9804,N_4958,N_3337);
nand U9805 (N_9805,N_345,N_3152);
and U9806 (N_9806,N_1184,N_4721);
xor U9807 (N_9807,N_2874,N_3288);
nor U9808 (N_9808,N_4725,N_542);
nor U9809 (N_9809,N_2164,N_255);
and U9810 (N_9810,N_5537,N_5250);
nand U9811 (N_9811,N_2116,N_442);
nor U9812 (N_9812,N_4388,N_4822);
xor U9813 (N_9813,N_1519,N_2028);
and U9814 (N_9814,N_1906,N_5445);
or U9815 (N_9815,N_5153,N_67);
and U9816 (N_9816,N_2949,N_415);
or U9817 (N_9817,N_5225,N_6038);
or U9818 (N_9818,N_3718,N_6182);
xnor U9819 (N_9819,N_4092,N_5695);
nor U9820 (N_9820,N_5290,N_5317);
nor U9821 (N_9821,N_2958,N_2957);
or U9822 (N_9822,N_1996,N_3428);
and U9823 (N_9823,N_5303,N_1349);
and U9824 (N_9824,N_1682,N_1512);
xnor U9825 (N_9825,N_5229,N_5787);
xnor U9826 (N_9826,N_174,N_3565);
nor U9827 (N_9827,N_5557,N_5235);
or U9828 (N_9828,N_2460,N_5562);
nor U9829 (N_9829,N_2139,N_461);
or U9830 (N_9830,N_1071,N_4397);
and U9831 (N_9831,N_1486,N_5190);
nor U9832 (N_9832,N_66,N_2038);
and U9833 (N_9833,N_3966,N_1065);
or U9834 (N_9834,N_3415,N_4205);
nor U9835 (N_9835,N_2862,N_828);
xnor U9836 (N_9836,N_2511,N_5734);
xor U9837 (N_9837,N_2112,N_1428);
nand U9838 (N_9838,N_1429,N_3827);
nand U9839 (N_9839,N_4699,N_1653);
or U9840 (N_9840,N_4060,N_1442);
nand U9841 (N_9841,N_1348,N_3599);
or U9842 (N_9842,N_5236,N_2668);
xor U9843 (N_9843,N_1593,N_5061);
nand U9844 (N_9844,N_5256,N_4627);
nand U9845 (N_9845,N_758,N_5626);
nand U9846 (N_9846,N_5770,N_2406);
nand U9847 (N_9847,N_2217,N_4385);
nand U9848 (N_9848,N_5313,N_3017);
or U9849 (N_9849,N_1562,N_3199);
xnor U9850 (N_9850,N_5881,N_5044);
nor U9851 (N_9851,N_2225,N_3735);
nor U9852 (N_9852,N_2961,N_4865);
and U9853 (N_9853,N_2808,N_160);
nand U9854 (N_9854,N_6219,N_5513);
nor U9855 (N_9855,N_3848,N_6022);
nand U9856 (N_9856,N_1796,N_2848);
nor U9857 (N_9857,N_2116,N_3250);
nor U9858 (N_9858,N_1071,N_6041);
xor U9859 (N_9859,N_5874,N_5523);
or U9860 (N_9860,N_1134,N_3375);
and U9861 (N_9861,N_2484,N_2512);
and U9862 (N_9862,N_1481,N_3350);
or U9863 (N_9863,N_1084,N_579);
nor U9864 (N_9864,N_2101,N_230);
nand U9865 (N_9865,N_3092,N_4887);
xor U9866 (N_9866,N_1506,N_4927);
or U9867 (N_9867,N_6052,N_5946);
and U9868 (N_9868,N_4091,N_6234);
nor U9869 (N_9869,N_3971,N_254);
and U9870 (N_9870,N_4562,N_3524);
and U9871 (N_9871,N_2448,N_744);
or U9872 (N_9872,N_1593,N_2645);
or U9873 (N_9873,N_4848,N_454);
and U9874 (N_9874,N_5102,N_1459);
and U9875 (N_9875,N_2085,N_5658);
or U9876 (N_9876,N_3325,N_579);
nor U9877 (N_9877,N_1469,N_2968);
nand U9878 (N_9878,N_467,N_2615);
nor U9879 (N_9879,N_2769,N_4061);
nor U9880 (N_9880,N_4589,N_3591);
or U9881 (N_9881,N_684,N_3740);
and U9882 (N_9882,N_5486,N_3265);
xor U9883 (N_9883,N_1151,N_918);
nor U9884 (N_9884,N_1590,N_3781);
nor U9885 (N_9885,N_4199,N_122);
xnor U9886 (N_9886,N_2774,N_1024);
or U9887 (N_9887,N_83,N_5736);
and U9888 (N_9888,N_3502,N_1552);
nor U9889 (N_9889,N_1035,N_4452);
nand U9890 (N_9890,N_655,N_6149);
nand U9891 (N_9891,N_2639,N_3334);
or U9892 (N_9892,N_2795,N_1280);
nand U9893 (N_9893,N_4519,N_2453);
nand U9894 (N_9894,N_3334,N_36);
xor U9895 (N_9895,N_1215,N_1322);
or U9896 (N_9896,N_3980,N_1792);
nor U9897 (N_9897,N_279,N_5640);
and U9898 (N_9898,N_1486,N_3059);
xnor U9899 (N_9899,N_1666,N_2810);
xnor U9900 (N_9900,N_3909,N_619);
and U9901 (N_9901,N_4846,N_396);
or U9902 (N_9902,N_2435,N_5953);
xor U9903 (N_9903,N_3000,N_5200);
or U9904 (N_9904,N_2583,N_306);
nand U9905 (N_9905,N_3041,N_893);
xnor U9906 (N_9906,N_2534,N_645);
and U9907 (N_9907,N_2348,N_3839);
nand U9908 (N_9908,N_3286,N_5439);
xor U9909 (N_9909,N_5870,N_5919);
and U9910 (N_9910,N_4701,N_1560);
and U9911 (N_9911,N_5136,N_1329);
and U9912 (N_9912,N_2582,N_482);
xnor U9913 (N_9913,N_4719,N_398);
or U9914 (N_9914,N_4758,N_2048);
nor U9915 (N_9915,N_2051,N_4809);
xnor U9916 (N_9916,N_1204,N_2622);
nand U9917 (N_9917,N_2094,N_4043);
nand U9918 (N_9918,N_4328,N_402);
nand U9919 (N_9919,N_5870,N_6045);
and U9920 (N_9920,N_5123,N_609);
nand U9921 (N_9921,N_3033,N_3162);
nand U9922 (N_9922,N_694,N_2049);
or U9923 (N_9923,N_3702,N_3606);
xnor U9924 (N_9924,N_996,N_1103);
or U9925 (N_9925,N_1072,N_317);
and U9926 (N_9926,N_4272,N_2340);
or U9927 (N_9927,N_1736,N_1545);
and U9928 (N_9928,N_4131,N_842);
and U9929 (N_9929,N_6198,N_1030);
or U9930 (N_9930,N_963,N_3285);
or U9931 (N_9931,N_4880,N_5759);
or U9932 (N_9932,N_860,N_973);
and U9933 (N_9933,N_993,N_5610);
nand U9934 (N_9934,N_4914,N_887);
or U9935 (N_9935,N_3405,N_2404);
nor U9936 (N_9936,N_1449,N_1986);
nor U9937 (N_9937,N_1979,N_3247);
xor U9938 (N_9938,N_5935,N_3770);
nand U9939 (N_9939,N_4193,N_3766);
nand U9940 (N_9940,N_4761,N_4001);
nor U9941 (N_9941,N_2668,N_6163);
or U9942 (N_9942,N_3663,N_5863);
and U9943 (N_9943,N_2342,N_4944);
and U9944 (N_9944,N_3889,N_3004);
nor U9945 (N_9945,N_5612,N_2984);
or U9946 (N_9946,N_1372,N_4463);
and U9947 (N_9947,N_929,N_3354);
nor U9948 (N_9948,N_1492,N_5341);
nand U9949 (N_9949,N_329,N_1858);
nand U9950 (N_9950,N_6166,N_1558);
nor U9951 (N_9951,N_4202,N_3984);
nand U9952 (N_9952,N_4146,N_5833);
nand U9953 (N_9953,N_5150,N_361);
and U9954 (N_9954,N_2682,N_903);
or U9955 (N_9955,N_2812,N_2103);
nor U9956 (N_9956,N_464,N_2877);
and U9957 (N_9957,N_786,N_6173);
or U9958 (N_9958,N_2511,N_954);
and U9959 (N_9959,N_5676,N_5927);
nor U9960 (N_9960,N_6125,N_4980);
nor U9961 (N_9961,N_1185,N_1666);
xor U9962 (N_9962,N_1413,N_634);
nor U9963 (N_9963,N_5226,N_1236);
nand U9964 (N_9964,N_4157,N_2436);
or U9965 (N_9965,N_2099,N_5665);
or U9966 (N_9966,N_5210,N_5615);
and U9967 (N_9967,N_1963,N_681);
or U9968 (N_9968,N_5287,N_4177);
xnor U9969 (N_9969,N_5788,N_6132);
and U9970 (N_9970,N_337,N_5317);
and U9971 (N_9971,N_3209,N_6080);
nor U9972 (N_9972,N_5465,N_3774);
nor U9973 (N_9973,N_1964,N_3529);
xnor U9974 (N_9974,N_2152,N_410);
or U9975 (N_9975,N_3719,N_708);
nand U9976 (N_9976,N_252,N_3325);
or U9977 (N_9977,N_2240,N_1356);
nand U9978 (N_9978,N_5764,N_5516);
and U9979 (N_9979,N_346,N_2122);
nor U9980 (N_9980,N_1302,N_3986);
and U9981 (N_9981,N_4792,N_2023);
and U9982 (N_9982,N_4089,N_5762);
or U9983 (N_9983,N_1032,N_131);
and U9984 (N_9984,N_1638,N_2642);
nor U9985 (N_9985,N_1223,N_3281);
and U9986 (N_9986,N_2170,N_1176);
nor U9987 (N_9987,N_4256,N_2635);
nand U9988 (N_9988,N_1465,N_978);
xor U9989 (N_9989,N_5624,N_6123);
nor U9990 (N_9990,N_2695,N_1680);
nor U9991 (N_9991,N_2113,N_1251);
nor U9992 (N_9992,N_447,N_5275);
and U9993 (N_9993,N_1883,N_1524);
or U9994 (N_9994,N_845,N_3680);
or U9995 (N_9995,N_2306,N_3193);
nand U9996 (N_9996,N_1031,N_4633);
or U9997 (N_9997,N_4302,N_6030);
or U9998 (N_9998,N_1735,N_2334);
and U9999 (N_9999,N_5848,N_1808);
or U10000 (N_10000,N_4321,N_3070);
and U10001 (N_10001,N_5587,N_1939);
or U10002 (N_10002,N_3424,N_1942);
nand U10003 (N_10003,N_120,N_5586);
xnor U10004 (N_10004,N_5517,N_2808);
or U10005 (N_10005,N_5608,N_1533);
xor U10006 (N_10006,N_4292,N_3556);
or U10007 (N_10007,N_4036,N_3712);
or U10008 (N_10008,N_178,N_4316);
or U10009 (N_10009,N_4144,N_753);
nor U10010 (N_10010,N_1235,N_5563);
nand U10011 (N_10011,N_3079,N_5308);
and U10012 (N_10012,N_1591,N_4358);
or U10013 (N_10013,N_5892,N_5639);
nor U10014 (N_10014,N_4280,N_4709);
nor U10015 (N_10015,N_1398,N_1980);
and U10016 (N_10016,N_5900,N_2109);
or U10017 (N_10017,N_559,N_1002);
and U10018 (N_10018,N_3684,N_4958);
or U10019 (N_10019,N_1085,N_5386);
nor U10020 (N_10020,N_2302,N_3550);
nand U10021 (N_10021,N_568,N_3338);
and U10022 (N_10022,N_1050,N_1202);
nand U10023 (N_10023,N_3943,N_2476);
or U10024 (N_10024,N_1512,N_1123);
and U10025 (N_10025,N_1438,N_2400);
xnor U10026 (N_10026,N_123,N_2024);
or U10027 (N_10027,N_1711,N_3874);
and U10028 (N_10028,N_2294,N_3316);
and U10029 (N_10029,N_4387,N_748);
nand U10030 (N_10030,N_763,N_1002);
and U10031 (N_10031,N_4948,N_3499);
nor U10032 (N_10032,N_602,N_4128);
nand U10033 (N_10033,N_4973,N_428);
or U10034 (N_10034,N_4024,N_1184);
nor U10035 (N_10035,N_296,N_4078);
nor U10036 (N_10036,N_3622,N_2790);
or U10037 (N_10037,N_4174,N_3542);
xor U10038 (N_10038,N_4231,N_3817);
nand U10039 (N_10039,N_3033,N_698);
and U10040 (N_10040,N_5499,N_517);
or U10041 (N_10041,N_1369,N_206);
nor U10042 (N_10042,N_5296,N_4117);
and U10043 (N_10043,N_3348,N_3319);
and U10044 (N_10044,N_3230,N_5953);
and U10045 (N_10045,N_425,N_5006);
xnor U10046 (N_10046,N_6103,N_2524);
and U10047 (N_10047,N_4914,N_2804);
nand U10048 (N_10048,N_2194,N_568);
or U10049 (N_10049,N_2490,N_67);
or U10050 (N_10050,N_357,N_4257);
nand U10051 (N_10051,N_6209,N_4102);
nand U10052 (N_10052,N_4436,N_481);
xnor U10053 (N_10053,N_261,N_4134);
nor U10054 (N_10054,N_5203,N_4837);
or U10055 (N_10055,N_5911,N_252);
nor U10056 (N_10056,N_2361,N_1520);
nand U10057 (N_10057,N_1244,N_1235);
nor U10058 (N_10058,N_5185,N_4229);
and U10059 (N_10059,N_4868,N_2500);
and U10060 (N_10060,N_5630,N_5576);
nor U10061 (N_10061,N_6175,N_3192);
or U10062 (N_10062,N_2947,N_4811);
nand U10063 (N_10063,N_504,N_5581);
and U10064 (N_10064,N_1024,N_2060);
nor U10065 (N_10065,N_3,N_2055);
nor U10066 (N_10066,N_550,N_5219);
or U10067 (N_10067,N_5585,N_5619);
and U10068 (N_10068,N_6054,N_5424);
and U10069 (N_10069,N_3625,N_4623);
nand U10070 (N_10070,N_270,N_518);
nand U10071 (N_10071,N_5517,N_1062);
nor U10072 (N_10072,N_5344,N_3115);
nor U10073 (N_10073,N_1195,N_1312);
and U10074 (N_10074,N_5197,N_138);
and U10075 (N_10075,N_4995,N_1086);
or U10076 (N_10076,N_5324,N_3080);
and U10077 (N_10077,N_5286,N_473);
nand U10078 (N_10078,N_3456,N_2592);
nand U10079 (N_10079,N_2443,N_5719);
nand U10080 (N_10080,N_4454,N_1907);
xor U10081 (N_10081,N_5783,N_2706);
nand U10082 (N_10082,N_461,N_3563);
nor U10083 (N_10083,N_3662,N_78);
or U10084 (N_10084,N_2453,N_978);
xor U10085 (N_10085,N_250,N_2820);
xor U10086 (N_10086,N_3197,N_2995);
and U10087 (N_10087,N_5191,N_2339);
nor U10088 (N_10088,N_6225,N_5559);
nand U10089 (N_10089,N_4562,N_2278);
or U10090 (N_10090,N_6158,N_4551);
nand U10091 (N_10091,N_280,N_5897);
nand U10092 (N_10092,N_1821,N_859);
or U10093 (N_10093,N_4502,N_1814);
and U10094 (N_10094,N_4595,N_4856);
nor U10095 (N_10095,N_3,N_1897);
or U10096 (N_10096,N_4701,N_1999);
nor U10097 (N_10097,N_4232,N_5435);
nand U10098 (N_10098,N_2058,N_1355);
nor U10099 (N_10099,N_3227,N_5172);
xnor U10100 (N_10100,N_312,N_1805);
nand U10101 (N_10101,N_5260,N_1430);
and U10102 (N_10102,N_4847,N_5172);
nand U10103 (N_10103,N_896,N_2019);
or U10104 (N_10104,N_2797,N_3355);
xnor U10105 (N_10105,N_3642,N_5752);
or U10106 (N_10106,N_4322,N_1614);
xnor U10107 (N_10107,N_1610,N_2842);
or U10108 (N_10108,N_5914,N_4573);
or U10109 (N_10109,N_3666,N_3300);
or U10110 (N_10110,N_384,N_2436);
xnor U10111 (N_10111,N_3949,N_1602);
and U10112 (N_10112,N_1165,N_5687);
nand U10113 (N_10113,N_4243,N_5716);
xor U10114 (N_10114,N_4756,N_4396);
nor U10115 (N_10115,N_6236,N_3677);
nor U10116 (N_10116,N_3937,N_2581);
or U10117 (N_10117,N_5423,N_5237);
nor U10118 (N_10118,N_1134,N_806);
or U10119 (N_10119,N_645,N_1578);
nand U10120 (N_10120,N_2913,N_3948);
nand U10121 (N_10121,N_4262,N_3931);
or U10122 (N_10122,N_1543,N_2585);
nand U10123 (N_10123,N_5597,N_698);
nand U10124 (N_10124,N_1887,N_522);
or U10125 (N_10125,N_3254,N_1152);
or U10126 (N_10126,N_2496,N_3501);
nand U10127 (N_10127,N_860,N_3324);
nand U10128 (N_10128,N_437,N_2987);
nand U10129 (N_10129,N_1444,N_4753);
xor U10130 (N_10130,N_3747,N_302);
nor U10131 (N_10131,N_2008,N_1651);
and U10132 (N_10132,N_3792,N_5744);
and U10133 (N_10133,N_6212,N_5063);
nand U10134 (N_10134,N_4840,N_380);
xnor U10135 (N_10135,N_125,N_2028);
xnor U10136 (N_10136,N_5200,N_6005);
nand U10137 (N_10137,N_4525,N_3696);
and U10138 (N_10138,N_1339,N_900);
nand U10139 (N_10139,N_1099,N_2225);
nor U10140 (N_10140,N_3544,N_6047);
xnor U10141 (N_10141,N_4032,N_726);
or U10142 (N_10142,N_6246,N_3758);
nor U10143 (N_10143,N_5629,N_3102);
and U10144 (N_10144,N_633,N_5898);
and U10145 (N_10145,N_3033,N_1509);
and U10146 (N_10146,N_5729,N_5069);
or U10147 (N_10147,N_6164,N_5924);
nor U10148 (N_10148,N_3028,N_1241);
and U10149 (N_10149,N_4303,N_2808);
xor U10150 (N_10150,N_2966,N_3761);
nand U10151 (N_10151,N_3110,N_3984);
nor U10152 (N_10152,N_3219,N_5931);
and U10153 (N_10153,N_180,N_2724);
nand U10154 (N_10154,N_2699,N_6182);
nor U10155 (N_10155,N_2287,N_2013);
nor U10156 (N_10156,N_2506,N_5441);
nor U10157 (N_10157,N_6045,N_5195);
and U10158 (N_10158,N_2599,N_4773);
nand U10159 (N_10159,N_1010,N_4818);
and U10160 (N_10160,N_570,N_5145);
nor U10161 (N_10161,N_4240,N_5233);
nor U10162 (N_10162,N_2342,N_3967);
nand U10163 (N_10163,N_5255,N_4989);
nor U10164 (N_10164,N_2075,N_3031);
or U10165 (N_10165,N_2249,N_5997);
nor U10166 (N_10166,N_5787,N_2823);
nor U10167 (N_10167,N_4150,N_1481);
and U10168 (N_10168,N_814,N_5731);
xor U10169 (N_10169,N_310,N_2103);
and U10170 (N_10170,N_2420,N_1209);
nor U10171 (N_10171,N_4912,N_6047);
nand U10172 (N_10172,N_2036,N_2561);
or U10173 (N_10173,N_6155,N_1056);
nand U10174 (N_10174,N_1460,N_1139);
or U10175 (N_10175,N_5688,N_1381);
nor U10176 (N_10176,N_807,N_3714);
and U10177 (N_10177,N_4452,N_2116);
or U10178 (N_10178,N_770,N_5250);
or U10179 (N_10179,N_5398,N_3201);
nor U10180 (N_10180,N_681,N_5501);
nand U10181 (N_10181,N_1656,N_4609);
nor U10182 (N_10182,N_5006,N_1123);
nand U10183 (N_10183,N_3649,N_2331);
or U10184 (N_10184,N_734,N_5928);
nand U10185 (N_10185,N_4714,N_3908);
and U10186 (N_10186,N_5626,N_2770);
and U10187 (N_10187,N_2576,N_2196);
nor U10188 (N_10188,N_1780,N_1441);
and U10189 (N_10189,N_3732,N_334);
nand U10190 (N_10190,N_5669,N_857);
nand U10191 (N_10191,N_2311,N_6067);
xnor U10192 (N_10192,N_5099,N_3089);
or U10193 (N_10193,N_2949,N_4739);
or U10194 (N_10194,N_5433,N_765);
xor U10195 (N_10195,N_3227,N_1334);
nor U10196 (N_10196,N_4457,N_4232);
and U10197 (N_10197,N_5346,N_4931);
xor U10198 (N_10198,N_5851,N_6134);
nand U10199 (N_10199,N_2500,N_4849);
or U10200 (N_10200,N_333,N_3137);
nand U10201 (N_10201,N_4452,N_5930);
nand U10202 (N_10202,N_4530,N_4777);
nor U10203 (N_10203,N_2010,N_3107);
nand U10204 (N_10204,N_1940,N_622);
and U10205 (N_10205,N_4636,N_4650);
nor U10206 (N_10206,N_2098,N_1520);
or U10207 (N_10207,N_374,N_1082);
or U10208 (N_10208,N_1565,N_640);
and U10209 (N_10209,N_4504,N_2034);
xor U10210 (N_10210,N_4035,N_514);
nor U10211 (N_10211,N_2838,N_2095);
and U10212 (N_10212,N_5790,N_203);
or U10213 (N_10213,N_330,N_556);
and U10214 (N_10214,N_1658,N_5337);
or U10215 (N_10215,N_4406,N_2947);
or U10216 (N_10216,N_79,N_740);
or U10217 (N_10217,N_5140,N_2211);
nor U10218 (N_10218,N_5483,N_1666);
nand U10219 (N_10219,N_5148,N_3314);
nand U10220 (N_10220,N_3076,N_3623);
nor U10221 (N_10221,N_2966,N_4572);
xnor U10222 (N_10222,N_3585,N_4431);
nand U10223 (N_10223,N_1097,N_3825);
and U10224 (N_10224,N_774,N_833);
and U10225 (N_10225,N_4730,N_1024);
or U10226 (N_10226,N_4820,N_2844);
and U10227 (N_10227,N_4835,N_5506);
nand U10228 (N_10228,N_3668,N_3784);
or U10229 (N_10229,N_4709,N_2188);
nor U10230 (N_10230,N_963,N_2333);
or U10231 (N_10231,N_1981,N_5881);
nand U10232 (N_10232,N_5860,N_1837);
or U10233 (N_10233,N_4999,N_1333);
and U10234 (N_10234,N_4324,N_3840);
nor U10235 (N_10235,N_5231,N_4381);
or U10236 (N_10236,N_2682,N_3003);
nand U10237 (N_10237,N_4189,N_3172);
or U10238 (N_10238,N_4408,N_6153);
and U10239 (N_10239,N_5505,N_5530);
and U10240 (N_10240,N_2369,N_4768);
nand U10241 (N_10241,N_2289,N_5995);
nor U10242 (N_10242,N_72,N_2035);
nor U10243 (N_10243,N_912,N_3006);
or U10244 (N_10244,N_5257,N_2847);
and U10245 (N_10245,N_694,N_34);
nor U10246 (N_10246,N_1581,N_775);
nand U10247 (N_10247,N_2493,N_5019);
and U10248 (N_10248,N_1219,N_1083);
nand U10249 (N_10249,N_6085,N_4188);
nor U10250 (N_10250,N_394,N_4305);
nor U10251 (N_10251,N_3799,N_3383);
or U10252 (N_10252,N_3469,N_4482);
nand U10253 (N_10253,N_2623,N_4078);
nor U10254 (N_10254,N_1264,N_1749);
nor U10255 (N_10255,N_4025,N_3108);
and U10256 (N_10256,N_2756,N_481);
xnor U10257 (N_10257,N_3120,N_2732);
or U10258 (N_10258,N_3254,N_5376);
and U10259 (N_10259,N_4705,N_2231);
or U10260 (N_10260,N_5013,N_2900);
and U10261 (N_10261,N_550,N_6042);
nand U10262 (N_10262,N_1523,N_1318);
nor U10263 (N_10263,N_5827,N_5255);
or U10264 (N_10264,N_1982,N_5308);
or U10265 (N_10265,N_5806,N_1782);
nand U10266 (N_10266,N_1645,N_5837);
nor U10267 (N_10267,N_2752,N_4051);
and U10268 (N_10268,N_3637,N_1413);
or U10269 (N_10269,N_3521,N_1339);
nand U10270 (N_10270,N_2180,N_1756);
nor U10271 (N_10271,N_1,N_753);
nand U10272 (N_10272,N_2114,N_4606);
xnor U10273 (N_10273,N_3905,N_2885);
nor U10274 (N_10274,N_5148,N_5873);
or U10275 (N_10275,N_1666,N_425);
nand U10276 (N_10276,N_5744,N_957);
or U10277 (N_10277,N_2762,N_4018);
or U10278 (N_10278,N_3786,N_2172);
nand U10279 (N_10279,N_6021,N_258);
and U10280 (N_10280,N_2086,N_6174);
nor U10281 (N_10281,N_2508,N_2650);
and U10282 (N_10282,N_875,N_4440);
nor U10283 (N_10283,N_1675,N_37);
and U10284 (N_10284,N_3794,N_5180);
and U10285 (N_10285,N_4291,N_259);
nand U10286 (N_10286,N_715,N_4228);
nand U10287 (N_10287,N_2325,N_2962);
or U10288 (N_10288,N_2139,N_495);
nor U10289 (N_10289,N_4146,N_1144);
and U10290 (N_10290,N_2441,N_1955);
and U10291 (N_10291,N_3895,N_2618);
and U10292 (N_10292,N_202,N_4107);
nor U10293 (N_10293,N_2853,N_2253);
and U10294 (N_10294,N_4398,N_1106);
nand U10295 (N_10295,N_3726,N_4779);
or U10296 (N_10296,N_600,N_4540);
and U10297 (N_10297,N_5758,N_6085);
nor U10298 (N_10298,N_3961,N_1863);
or U10299 (N_10299,N_5972,N_2821);
nand U10300 (N_10300,N_4902,N_2911);
nor U10301 (N_10301,N_1865,N_1625);
nand U10302 (N_10302,N_4696,N_5167);
nor U10303 (N_10303,N_3017,N_169);
and U10304 (N_10304,N_5690,N_6144);
nand U10305 (N_10305,N_1434,N_4599);
and U10306 (N_10306,N_4259,N_1027);
nor U10307 (N_10307,N_4541,N_4366);
nand U10308 (N_10308,N_5444,N_4799);
or U10309 (N_10309,N_5958,N_1888);
nand U10310 (N_10310,N_5184,N_1575);
and U10311 (N_10311,N_352,N_5824);
nand U10312 (N_10312,N_2861,N_2105);
and U10313 (N_10313,N_4935,N_2920);
and U10314 (N_10314,N_1198,N_4054);
nand U10315 (N_10315,N_5895,N_1908);
nand U10316 (N_10316,N_4478,N_5387);
nor U10317 (N_10317,N_6013,N_5990);
or U10318 (N_10318,N_5373,N_848);
and U10319 (N_10319,N_700,N_356);
and U10320 (N_10320,N_5412,N_3080);
nand U10321 (N_10321,N_2652,N_2269);
nand U10322 (N_10322,N_5482,N_4886);
or U10323 (N_10323,N_1275,N_3373);
nor U10324 (N_10324,N_1086,N_3846);
xor U10325 (N_10325,N_5310,N_2850);
and U10326 (N_10326,N_4047,N_1434);
and U10327 (N_10327,N_4014,N_4155);
nor U10328 (N_10328,N_3300,N_2088);
and U10329 (N_10329,N_2082,N_3222);
nor U10330 (N_10330,N_4277,N_2198);
nor U10331 (N_10331,N_2514,N_2529);
nor U10332 (N_10332,N_2691,N_3945);
or U10333 (N_10333,N_5363,N_6163);
xor U10334 (N_10334,N_1626,N_1409);
and U10335 (N_10335,N_2232,N_3184);
and U10336 (N_10336,N_4263,N_1048);
nand U10337 (N_10337,N_5666,N_2714);
nand U10338 (N_10338,N_3705,N_3925);
nor U10339 (N_10339,N_6209,N_1221);
nand U10340 (N_10340,N_3571,N_734);
and U10341 (N_10341,N_2138,N_5834);
or U10342 (N_10342,N_4088,N_1375);
and U10343 (N_10343,N_5726,N_4766);
nand U10344 (N_10344,N_4877,N_4354);
xnor U10345 (N_10345,N_1417,N_4170);
nor U10346 (N_10346,N_1663,N_5965);
or U10347 (N_10347,N_2462,N_3207);
or U10348 (N_10348,N_4085,N_4971);
or U10349 (N_10349,N_3513,N_5838);
nor U10350 (N_10350,N_5660,N_1053);
nand U10351 (N_10351,N_5765,N_5485);
and U10352 (N_10352,N_3320,N_1024);
xnor U10353 (N_10353,N_2019,N_5164);
nand U10354 (N_10354,N_5354,N_5104);
nand U10355 (N_10355,N_2623,N_3861);
or U10356 (N_10356,N_3281,N_3382);
and U10357 (N_10357,N_4961,N_3993);
nand U10358 (N_10358,N_4815,N_774);
and U10359 (N_10359,N_577,N_1723);
nor U10360 (N_10360,N_790,N_2246);
and U10361 (N_10361,N_1422,N_1362);
nand U10362 (N_10362,N_4815,N_1613);
or U10363 (N_10363,N_4236,N_1655);
or U10364 (N_10364,N_1134,N_4962);
or U10365 (N_10365,N_1655,N_6066);
or U10366 (N_10366,N_4406,N_4636);
or U10367 (N_10367,N_1804,N_5024);
or U10368 (N_10368,N_5238,N_2477);
xnor U10369 (N_10369,N_4962,N_2971);
and U10370 (N_10370,N_2150,N_3367);
and U10371 (N_10371,N_2101,N_4618);
nor U10372 (N_10372,N_4688,N_5518);
nor U10373 (N_10373,N_4530,N_2980);
nand U10374 (N_10374,N_5214,N_3930);
nor U10375 (N_10375,N_3104,N_1289);
and U10376 (N_10376,N_2170,N_2785);
xnor U10377 (N_10377,N_4904,N_2899);
or U10378 (N_10378,N_4223,N_265);
nand U10379 (N_10379,N_1573,N_3299);
or U10380 (N_10380,N_6201,N_199);
nor U10381 (N_10381,N_69,N_74);
nand U10382 (N_10382,N_812,N_5382);
and U10383 (N_10383,N_141,N_2120);
nand U10384 (N_10384,N_1587,N_5646);
nor U10385 (N_10385,N_5708,N_2845);
nand U10386 (N_10386,N_1533,N_3346);
and U10387 (N_10387,N_1396,N_1678);
nor U10388 (N_10388,N_2255,N_795);
nor U10389 (N_10389,N_2114,N_1663);
nor U10390 (N_10390,N_4995,N_2173);
and U10391 (N_10391,N_312,N_714);
nand U10392 (N_10392,N_366,N_1862);
nand U10393 (N_10393,N_1467,N_5995);
and U10394 (N_10394,N_4115,N_6011);
nand U10395 (N_10395,N_2925,N_3681);
or U10396 (N_10396,N_2600,N_4272);
or U10397 (N_10397,N_1864,N_1198);
and U10398 (N_10398,N_2215,N_1530);
or U10399 (N_10399,N_6033,N_5235);
and U10400 (N_10400,N_3138,N_6159);
nand U10401 (N_10401,N_5198,N_1330);
nor U10402 (N_10402,N_4439,N_4208);
nand U10403 (N_10403,N_827,N_1655);
nand U10404 (N_10404,N_4833,N_2895);
nor U10405 (N_10405,N_1704,N_4461);
and U10406 (N_10406,N_2383,N_5533);
and U10407 (N_10407,N_2565,N_3461);
or U10408 (N_10408,N_3974,N_2118);
nor U10409 (N_10409,N_617,N_964);
nand U10410 (N_10410,N_2184,N_3118);
nor U10411 (N_10411,N_2596,N_2090);
nor U10412 (N_10412,N_5357,N_5992);
nand U10413 (N_10413,N_2615,N_1679);
and U10414 (N_10414,N_3231,N_601);
nand U10415 (N_10415,N_3718,N_6055);
nand U10416 (N_10416,N_3193,N_214);
nor U10417 (N_10417,N_3676,N_988);
nand U10418 (N_10418,N_4215,N_5888);
xor U10419 (N_10419,N_4380,N_4146);
nand U10420 (N_10420,N_4158,N_2201);
nor U10421 (N_10421,N_3944,N_4171);
or U10422 (N_10422,N_211,N_892);
and U10423 (N_10423,N_3639,N_3602);
nand U10424 (N_10424,N_4298,N_4625);
or U10425 (N_10425,N_969,N_5085);
nand U10426 (N_10426,N_4618,N_64);
and U10427 (N_10427,N_3453,N_3757);
or U10428 (N_10428,N_3842,N_5127);
xor U10429 (N_10429,N_3207,N_2445);
or U10430 (N_10430,N_5271,N_5957);
xor U10431 (N_10431,N_5905,N_3031);
xor U10432 (N_10432,N_4542,N_3155);
or U10433 (N_10433,N_2382,N_3232);
nor U10434 (N_10434,N_850,N_844);
and U10435 (N_10435,N_2917,N_634);
nand U10436 (N_10436,N_2547,N_929);
nand U10437 (N_10437,N_3854,N_5436);
xnor U10438 (N_10438,N_1182,N_2554);
and U10439 (N_10439,N_3960,N_3996);
or U10440 (N_10440,N_5883,N_2369);
nand U10441 (N_10441,N_3525,N_2762);
xnor U10442 (N_10442,N_3016,N_4379);
or U10443 (N_10443,N_386,N_5200);
and U10444 (N_10444,N_5716,N_5631);
or U10445 (N_10445,N_5581,N_3271);
nand U10446 (N_10446,N_127,N_4947);
nor U10447 (N_10447,N_4141,N_5630);
and U10448 (N_10448,N_3856,N_2162);
nand U10449 (N_10449,N_1169,N_2169);
nand U10450 (N_10450,N_5762,N_3426);
nor U10451 (N_10451,N_5798,N_3344);
nor U10452 (N_10452,N_52,N_629);
or U10453 (N_10453,N_3850,N_6235);
nor U10454 (N_10454,N_5189,N_4563);
nand U10455 (N_10455,N_2455,N_3974);
and U10456 (N_10456,N_3064,N_3208);
nand U10457 (N_10457,N_51,N_1314);
and U10458 (N_10458,N_567,N_5545);
or U10459 (N_10459,N_4107,N_3953);
or U10460 (N_10460,N_4856,N_2894);
or U10461 (N_10461,N_2928,N_1461);
and U10462 (N_10462,N_924,N_1526);
nor U10463 (N_10463,N_1802,N_5463);
nor U10464 (N_10464,N_2601,N_2014);
and U10465 (N_10465,N_942,N_1247);
nand U10466 (N_10466,N_728,N_6151);
xor U10467 (N_10467,N_4256,N_3671);
and U10468 (N_10468,N_1582,N_6165);
or U10469 (N_10469,N_2513,N_2025);
nand U10470 (N_10470,N_3552,N_1531);
and U10471 (N_10471,N_5550,N_2691);
or U10472 (N_10472,N_6188,N_5078);
or U10473 (N_10473,N_2926,N_3009);
nand U10474 (N_10474,N_3372,N_693);
nand U10475 (N_10475,N_5285,N_5860);
and U10476 (N_10476,N_2700,N_5649);
nand U10477 (N_10477,N_638,N_5850);
or U10478 (N_10478,N_4782,N_2816);
and U10479 (N_10479,N_1427,N_3361);
or U10480 (N_10480,N_4574,N_3123);
nand U10481 (N_10481,N_5595,N_6135);
nand U10482 (N_10482,N_1165,N_960);
nor U10483 (N_10483,N_3333,N_3366);
and U10484 (N_10484,N_3913,N_1079);
xnor U10485 (N_10485,N_2087,N_2825);
xor U10486 (N_10486,N_50,N_3617);
or U10487 (N_10487,N_4826,N_5824);
or U10488 (N_10488,N_3206,N_5543);
or U10489 (N_10489,N_3470,N_2204);
and U10490 (N_10490,N_6091,N_1320);
nor U10491 (N_10491,N_5024,N_2053);
or U10492 (N_10492,N_5637,N_4618);
nor U10493 (N_10493,N_5125,N_6110);
nor U10494 (N_10494,N_5111,N_281);
nand U10495 (N_10495,N_2202,N_3259);
nand U10496 (N_10496,N_3073,N_802);
nor U10497 (N_10497,N_2847,N_4879);
or U10498 (N_10498,N_3550,N_2814);
nor U10499 (N_10499,N_3716,N_3187);
or U10500 (N_10500,N_1313,N_184);
nor U10501 (N_10501,N_4390,N_404);
nor U10502 (N_10502,N_4764,N_4685);
nor U10503 (N_10503,N_3300,N_4663);
nor U10504 (N_10504,N_1157,N_2673);
nand U10505 (N_10505,N_2410,N_1722);
and U10506 (N_10506,N_3952,N_1872);
nand U10507 (N_10507,N_3124,N_4456);
xnor U10508 (N_10508,N_889,N_4526);
nor U10509 (N_10509,N_5177,N_3038);
nor U10510 (N_10510,N_3304,N_52);
nor U10511 (N_10511,N_1389,N_5461);
and U10512 (N_10512,N_5862,N_3717);
nor U10513 (N_10513,N_2903,N_1432);
nand U10514 (N_10514,N_1440,N_2382);
nand U10515 (N_10515,N_295,N_1803);
xnor U10516 (N_10516,N_2029,N_1822);
or U10517 (N_10517,N_599,N_6211);
and U10518 (N_10518,N_3248,N_2649);
or U10519 (N_10519,N_2417,N_5268);
nand U10520 (N_10520,N_3033,N_1105);
or U10521 (N_10521,N_4842,N_5236);
nor U10522 (N_10522,N_5186,N_6203);
nand U10523 (N_10523,N_2623,N_4596);
nor U10524 (N_10524,N_6193,N_310);
nor U10525 (N_10525,N_4198,N_2543);
nor U10526 (N_10526,N_1876,N_364);
nand U10527 (N_10527,N_1806,N_3075);
nand U10528 (N_10528,N_3402,N_1944);
and U10529 (N_10529,N_677,N_1704);
xnor U10530 (N_10530,N_66,N_5214);
nor U10531 (N_10531,N_4894,N_2841);
and U10532 (N_10532,N_3180,N_4505);
xnor U10533 (N_10533,N_6144,N_1704);
or U10534 (N_10534,N_473,N_5272);
xor U10535 (N_10535,N_1359,N_4526);
and U10536 (N_10536,N_5513,N_487);
nor U10537 (N_10537,N_4196,N_1366);
nor U10538 (N_10538,N_1717,N_363);
or U10539 (N_10539,N_6061,N_1887);
nor U10540 (N_10540,N_378,N_903);
and U10541 (N_10541,N_4151,N_5331);
and U10542 (N_10542,N_116,N_5012);
xnor U10543 (N_10543,N_687,N_4636);
nand U10544 (N_10544,N_2817,N_4480);
nor U10545 (N_10545,N_3457,N_1010);
nand U10546 (N_10546,N_1654,N_1072);
or U10547 (N_10547,N_3492,N_4874);
and U10548 (N_10548,N_2259,N_232);
and U10549 (N_10549,N_3217,N_2167);
nor U10550 (N_10550,N_1269,N_3862);
nand U10551 (N_10551,N_6133,N_380);
or U10552 (N_10552,N_4405,N_219);
or U10553 (N_10553,N_4928,N_6039);
nor U10554 (N_10554,N_3535,N_3787);
or U10555 (N_10555,N_1174,N_2519);
xor U10556 (N_10556,N_5789,N_685);
and U10557 (N_10557,N_3185,N_4427);
nor U10558 (N_10558,N_503,N_2085);
nor U10559 (N_10559,N_4038,N_1852);
or U10560 (N_10560,N_534,N_495);
or U10561 (N_10561,N_1907,N_1827);
and U10562 (N_10562,N_3359,N_5033);
or U10563 (N_10563,N_431,N_1800);
or U10564 (N_10564,N_4986,N_5681);
and U10565 (N_10565,N_5290,N_3815);
xor U10566 (N_10566,N_853,N_2548);
or U10567 (N_10567,N_556,N_2793);
nor U10568 (N_10568,N_829,N_5943);
nand U10569 (N_10569,N_4074,N_6196);
xor U10570 (N_10570,N_1882,N_3060);
and U10571 (N_10571,N_5744,N_895);
nand U10572 (N_10572,N_5716,N_5070);
or U10573 (N_10573,N_3077,N_5366);
and U10574 (N_10574,N_4666,N_2754);
nor U10575 (N_10575,N_3353,N_3493);
nor U10576 (N_10576,N_4824,N_1444);
nor U10577 (N_10577,N_4932,N_4818);
or U10578 (N_10578,N_1028,N_5166);
or U10579 (N_10579,N_5198,N_5961);
xnor U10580 (N_10580,N_2092,N_416);
nand U10581 (N_10581,N_4424,N_3431);
nand U10582 (N_10582,N_1782,N_4332);
nand U10583 (N_10583,N_1991,N_3354);
xnor U10584 (N_10584,N_5978,N_693);
nor U10585 (N_10585,N_6217,N_1379);
nor U10586 (N_10586,N_3685,N_4592);
nand U10587 (N_10587,N_1198,N_3529);
and U10588 (N_10588,N_1236,N_4340);
nand U10589 (N_10589,N_275,N_4374);
nor U10590 (N_10590,N_5400,N_4807);
and U10591 (N_10591,N_3697,N_2872);
or U10592 (N_10592,N_1568,N_1283);
or U10593 (N_10593,N_5164,N_5297);
and U10594 (N_10594,N_2542,N_3797);
and U10595 (N_10595,N_3164,N_1279);
nor U10596 (N_10596,N_5962,N_1984);
or U10597 (N_10597,N_4508,N_2340);
nand U10598 (N_10598,N_3329,N_467);
xor U10599 (N_10599,N_3420,N_1807);
and U10600 (N_10600,N_4891,N_6076);
nand U10601 (N_10601,N_4111,N_4928);
nand U10602 (N_10602,N_5386,N_5471);
and U10603 (N_10603,N_1681,N_4690);
or U10604 (N_10604,N_1781,N_5542);
or U10605 (N_10605,N_2177,N_1416);
or U10606 (N_10606,N_1313,N_4593);
nand U10607 (N_10607,N_4254,N_2904);
or U10608 (N_10608,N_662,N_4039);
or U10609 (N_10609,N_2557,N_1870);
or U10610 (N_10610,N_924,N_736);
xnor U10611 (N_10611,N_4684,N_4807);
nand U10612 (N_10612,N_3698,N_2953);
and U10613 (N_10613,N_3969,N_2464);
nand U10614 (N_10614,N_2575,N_1860);
nand U10615 (N_10615,N_6153,N_2877);
and U10616 (N_10616,N_1118,N_107);
nor U10617 (N_10617,N_824,N_141);
nand U10618 (N_10618,N_1872,N_3898);
nor U10619 (N_10619,N_1375,N_3659);
nor U10620 (N_10620,N_2848,N_3127);
nand U10621 (N_10621,N_4757,N_5121);
and U10622 (N_10622,N_4048,N_3176);
or U10623 (N_10623,N_3576,N_1336);
nor U10624 (N_10624,N_1137,N_2218);
nor U10625 (N_10625,N_5792,N_5873);
nor U10626 (N_10626,N_5264,N_1422);
nand U10627 (N_10627,N_5365,N_587);
or U10628 (N_10628,N_1745,N_3320);
or U10629 (N_10629,N_4059,N_3586);
nor U10630 (N_10630,N_870,N_323);
or U10631 (N_10631,N_2137,N_2740);
or U10632 (N_10632,N_5010,N_5898);
nand U10633 (N_10633,N_3008,N_5677);
nand U10634 (N_10634,N_4317,N_6105);
nand U10635 (N_10635,N_3351,N_1462);
xnor U10636 (N_10636,N_4601,N_3347);
nor U10637 (N_10637,N_4691,N_54);
nand U10638 (N_10638,N_2925,N_4294);
nand U10639 (N_10639,N_4934,N_174);
xor U10640 (N_10640,N_5719,N_3415);
nor U10641 (N_10641,N_1037,N_1087);
nand U10642 (N_10642,N_5123,N_1039);
or U10643 (N_10643,N_3948,N_1863);
nand U10644 (N_10644,N_1627,N_3799);
nand U10645 (N_10645,N_5415,N_1376);
nor U10646 (N_10646,N_4334,N_763);
xnor U10647 (N_10647,N_4856,N_3234);
nand U10648 (N_10648,N_1615,N_6047);
and U10649 (N_10649,N_2082,N_829);
nor U10650 (N_10650,N_4534,N_4204);
or U10651 (N_10651,N_6034,N_2513);
and U10652 (N_10652,N_1647,N_355);
or U10653 (N_10653,N_4064,N_4067);
xor U10654 (N_10654,N_989,N_303);
nor U10655 (N_10655,N_3598,N_2642);
and U10656 (N_10656,N_5002,N_4706);
nand U10657 (N_10657,N_5441,N_688);
nor U10658 (N_10658,N_706,N_945);
nand U10659 (N_10659,N_4830,N_3770);
or U10660 (N_10660,N_6228,N_914);
nand U10661 (N_10661,N_5657,N_3119);
nor U10662 (N_10662,N_6105,N_5928);
xor U10663 (N_10663,N_3559,N_3878);
and U10664 (N_10664,N_4514,N_4080);
nand U10665 (N_10665,N_5342,N_1945);
or U10666 (N_10666,N_5984,N_2984);
or U10667 (N_10667,N_734,N_2058);
or U10668 (N_10668,N_6107,N_5958);
xnor U10669 (N_10669,N_2140,N_3584);
xor U10670 (N_10670,N_3961,N_4371);
nand U10671 (N_10671,N_3864,N_611);
and U10672 (N_10672,N_406,N_6141);
and U10673 (N_10673,N_3882,N_5231);
or U10674 (N_10674,N_5314,N_5988);
or U10675 (N_10675,N_181,N_5396);
nand U10676 (N_10676,N_5793,N_3066);
and U10677 (N_10677,N_2817,N_2515);
and U10678 (N_10678,N_4882,N_5918);
nand U10679 (N_10679,N_3957,N_448);
and U10680 (N_10680,N_171,N_113);
or U10681 (N_10681,N_5504,N_1370);
xor U10682 (N_10682,N_746,N_2138);
and U10683 (N_10683,N_4730,N_4607);
and U10684 (N_10684,N_3027,N_743);
nand U10685 (N_10685,N_1505,N_1401);
or U10686 (N_10686,N_3519,N_2532);
nand U10687 (N_10687,N_4443,N_930);
or U10688 (N_10688,N_2228,N_1033);
nor U10689 (N_10689,N_509,N_500);
nor U10690 (N_10690,N_3879,N_561);
or U10691 (N_10691,N_6149,N_5348);
and U10692 (N_10692,N_3985,N_5706);
nor U10693 (N_10693,N_3704,N_2590);
nor U10694 (N_10694,N_2242,N_3033);
nand U10695 (N_10695,N_3409,N_1671);
nand U10696 (N_10696,N_4964,N_5103);
and U10697 (N_10697,N_5991,N_2865);
or U10698 (N_10698,N_1850,N_76);
xor U10699 (N_10699,N_2257,N_3926);
nand U10700 (N_10700,N_4698,N_1708);
or U10701 (N_10701,N_4203,N_3819);
and U10702 (N_10702,N_1951,N_4491);
nor U10703 (N_10703,N_5231,N_4565);
or U10704 (N_10704,N_3626,N_1785);
nor U10705 (N_10705,N_5919,N_4587);
nand U10706 (N_10706,N_3404,N_3933);
or U10707 (N_10707,N_1394,N_3164);
nand U10708 (N_10708,N_5125,N_3394);
and U10709 (N_10709,N_1964,N_5015);
or U10710 (N_10710,N_4481,N_1492);
or U10711 (N_10711,N_3060,N_75);
nor U10712 (N_10712,N_2243,N_4496);
nand U10713 (N_10713,N_3635,N_2392);
nand U10714 (N_10714,N_3532,N_3607);
xnor U10715 (N_10715,N_1975,N_2889);
and U10716 (N_10716,N_5200,N_2196);
and U10717 (N_10717,N_3973,N_2117);
xor U10718 (N_10718,N_4263,N_3444);
xor U10719 (N_10719,N_5477,N_5916);
and U10720 (N_10720,N_4772,N_402);
nand U10721 (N_10721,N_3429,N_5278);
nor U10722 (N_10722,N_3952,N_3408);
xor U10723 (N_10723,N_4280,N_1080);
nor U10724 (N_10724,N_5671,N_5032);
nor U10725 (N_10725,N_765,N_3582);
nand U10726 (N_10726,N_2411,N_2052);
nand U10727 (N_10727,N_2849,N_5451);
xor U10728 (N_10728,N_2802,N_889);
and U10729 (N_10729,N_2014,N_6013);
and U10730 (N_10730,N_2200,N_2899);
or U10731 (N_10731,N_6067,N_4936);
nand U10732 (N_10732,N_5778,N_1944);
and U10733 (N_10733,N_6062,N_4828);
nor U10734 (N_10734,N_1397,N_529);
nor U10735 (N_10735,N_3204,N_2281);
or U10736 (N_10736,N_1082,N_5197);
or U10737 (N_10737,N_2420,N_5729);
or U10738 (N_10738,N_1071,N_1259);
nor U10739 (N_10739,N_2871,N_572);
or U10740 (N_10740,N_2586,N_3397);
nand U10741 (N_10741,N_4861,N_5248);
and U10742 (N_10742,N_4319,N_4356);
xnor U10743 (N_10743,N_4695,N_3694);
and U10744 (N_10744,N_4499,N_993);
and U10745 (N_10745,N_4322,N_1948);
or U10746 (N_10746,N_605,N_3120);
or U10747 (N_10747,N_2361,N_2650);
nand U10748 (N_10748,N_948,N_1287);
and U10749 (N_10749,N_1846,N_5147);
and U10750 (N_10750,N_3024,N_4617);
or U10751 (N_10751,N_2653,N_876);
nand U10752 (N_10752,N_2128,N_2815);
nand U10753 (N_10753,N_1548,N_1515);
or U10754 (N_10754,N_3835,N_3508);
nand U10755 (N_10755,N_4166,N_5727);
nor U10756 (N_10756,N_1456,N_2768);
and U10757 (N_10757,N_5333,N_3955);
or U10758 (N_10758,N_788,N_3953);
nand U10759 (N_10759,N_5633,N_1243);
and U10760 (N_10760,N_3694,N_1301);
nor U10761 (N_10761,N_5113,N_720);
nand U10762 (N_10762,N_4485,N_5111);
or U10763 (N_10763,N_3993,N_97);
xor U10764 (N_10764,N_910,N_4779);
nand U10765 (N_10765,N_4465,N_5445);
nor U10766 (N_10766,N_5607,N_1388);
nand U10767 (N_10767,N_3152,N_4086);
nand U10768 (N_10768,N_2006,N_1182);
and U10769 (N_10769,N_4566,N_3373);
or U10770 (N_10770,N_3243,N_3228);
nand U10771 (N_10771,N_5159,N_3657);
and U10772 (N_10772,N_781,N_283);
nor U10773 (N_10773,N_3820,N_1796);
and U10774 (N_10774,N_3290,N_4045);
nand U10775 (N_10775,N_3849,N_5554);
and U10776 (N_10776,N_217,N_5910);
and U10777 (N_10777,N_4608,N_5166);
or U10778 (N_10778,N_3703,N_4711);
nor U10779 (N_10779,N_5277,N_3055);
nor U10780 (N_10780,N_3214,N_850);
nor U10781 (N_10781,N_98,N_1304);
or U10782 (N_10782,N_3017,N_1973);
nor U10783 (N_10783,N_1475,N_1570);
and U10784 (N_10784,N_4369,N_2082);
or U10785 (N_10785,N_5140,N_528);
nand U10786 (N_10786,N_5126,N_29);
or U10787 (N_10787,N_1102,N_376);
xnor U10788 (N_10788,N_454,N_5957);
nor U10789 (N_10789,N_6243,N_2235);
xnor U10790 (N_10790,N_1884,N_3355);
or U10791 (N_10791,N_3595,N_3801);
nand U10792 (N_10792,N_2867,N_3845);
nand U10793 (N_10793,N_346,N_1955);
nand U10794 (N_10794,N_3772,N_1729);
xor U10795 (N_10795,N_4329,N_2144);
xor U10796 (N_10796,N_4210,N_4795);
nand U10797 (N_10797,N_1029,N_921);
or U10798 (N_10798,N_2039,N_2575);
nor U10799 (N_10799,N_378,N_1537);
nand U10800 (N_10800,N_2496,N_594);
nand U10801 (N_10801,N_1686,N_941);
or U10802 (N_10802,N_5907,N_1293);
and U10803 (N_10803,N_190,N_2550);
nand U10804 (N_10804,N_2823,N_4010);
nand U10805 (N_10805,N_2513,N_2793);
nand U10806 (N_10806,N_4213,N_1178);
nor U10807 (N_10807,N_3974,N_1062);
nand U10808 (N_10808,N_1147,N_5416);
and U10809 (N_10809,N_4507,N_1746);
and U10810 (N_10810,N_2637,N_1921);
xnor U10811 (N_10811,N_2682,N_6018);
and U10812 (N_10812,N_2641,N_4896);
nor U10813 (N_10813,N_4105,N_3488);
nor U10814 (N_10814,N_597,N_278);
nand U10815 (N_10815,N_3988,N_6201);
nor U10816 (N_10816,N_2439,N_3258);
xor U10817 (N_10817,N_1962,N_3065);
or U10818 (N_10818,N_2270,N_1482);
and U10819 (N_10819,N_5369,N_3585);
nor U10820 (N_10820,N_5041,N_4093);
xor U10821 (N_10821,N_4307,N_1291);
or U10822 (N_10822,N_1834,N_5333);
xnor U10823 (N_10823,N_3993,N_5418);
or U10824 (N_10824,N_3128,N_5);
and U10825 (N_10825,N_849,N_3066);
nand U10826 (N_10826,N_3088,N_1599);
nor U10827 (N_10827,N_59,N_2397);
or U10828 (N_10828,N_5068,N_5833);
nand U10829 (N_10829,N_4376,N_3648);
nand U10830 (N_10830,N_5784,N_4938);
or U10831 (N_10831,N_4790,N_973);
nor U10832 (N_10832,N_160,N_6083);
or U10833 (N_10833,N_111,N_3333);
and U10834 (N_10834,N_4019,N_5623);
nor U10835 (N_10835,N_1163,N_1048);
nand U10836 (N_10836,N_3198,N_3433);
nor U10837 (N_10837,N_215,N_4364);
nor U10838 (N_10838,N_3673,N_200);
nor U10839 (N_10839,N_2514,N_4813);
or U10840 (N_10840,N_6047,N_2062);
xnor U10841 (N_10841,N_5083,N_4038);
and U10842 (N_10842,N_4115,N_3177);
and U10843 (N_10843,N_4213,N_2970);
nand U10844 (N_10844,N_301,N_6066);
and U10845 (N_10845,N_6106,N_5183);
and U10846 (N_10846,N_2922,N_2488);
or U10847 (N_10847,N_3012,N_451);
and U10848 (N_10848,N_4995,N_4181);
xor U10849 (N_10849,N_4590,N_1872);
nand U10850 (N_10850,N_583,N_4081);
or U10851 (N_10851,N_5069,N_4172);
and U10852 (N_10852,N_2263,N_2715);
nor U10853 (N_10853,N_5443,N_1596);
and U10854 (N_10854,N_1705,N_5046);
and U10855 (N_10855,N_4315,N_5586);
nand U10856 (N_10856,N_5074,N_4920);
or U10857 (N_10857,N_140,N_5266);
nor U10858 (N_10858,N_30,N_4952);
nor U10859 (N_10859,N_4695,N_2354);
and U10860 (N_10860,N_1201,N_551);
nand U10861 (N_10861,N_667,N_2094);
and U10862 (N_10862,N_3003,N_43);
or U10863 (N_10863,N_4110,N_1131);
or U10864 (N_10864,N_745,N_4782);
or U10865 (N_10865,N_2535,N_6018);
or U10866 (N_10866,N_4903,N_2030);
nand U10867 (N_10867,N_3076,N_2182);
or U10868 (N_10868,N_679,N_3486);
nor U10869 (N_10869,N_1856,N_5387);
and U10870 (N_10870,N_1500,N_2102);
nand U10871 (N_10871,N_3889,N_1655);
or U10872 (N_10872,N_434,N_496);
nor U10873 (N_10873,N_979,N_3409);
or U10874 (N_10874,N_475,N_4385);
and U10875 (N_10875,N_5882,N_1732);
nor U10876 (N_10876,N_5615,N_2701);
nand U10877 (N_10877,N_1965,N_1968);
or U10878 (N_10878,N_4682,N_1485);
nand U10879 (N_10879,N_1734,N_1634);
or U10880 (N_10880,N_6245,N_1583);
xor U10881 (N_10881,N_2207,N_2181);
and U10882 (N_10882,N_791,N_3312);
and U10883 (N_10883,N_5487,N_1417);
or U10884 (N_10884,N_2970,N_964);
nand U10885 (N_10885,N_1614,N_4754);
nor U10886 (N_10886,N_3387,N_3377);
and U10887 (N_10887,N_628,N_5784);
nand U10888 (N_10888,N_4096,N_176);
nor U10889 (N_10889,N_4052,N_861);
nand U10890 (N_10890,N_6146,N_3673);
nand U10891 (N_10891,N_848,N_608);
nor U10892 (N_10892,N_4609,N_4176);
nor U10893 (N_10893,N_5085,N_4715);
xor U10894 (N_10894,N_1122,N_5318);
nand U10895 (N_10895,N_5044,N_2772);
or U10896 (N_10896,N_238,N_735);
nand U10897 (N_10897,N_928,N_4086);
or U10898 (N_10898,N_1779,N_1922);
and U10899 (N_10899,N_65,N_5249);
nand U10900 (N_10900,N_3420,N_3188);
nor U10901 (N_10901,N_16,N_805);
or U10902 (N_10902,N_946,N_4688);
and U10903 (N_10903,N_3558,N_4978);
or U10904 (N_10904,N_374,N_2202);
or U10905 (N_10905,N_4168,N_1669);
or U10906 (N_10906,N_5288,N_3516);
or U10907 (N_10907,N_1194,N_3970);
or U10908 (N_10908,N_2945,N_1255);
nand U10909 (N_10909,N_1263,N_6095);
nand U10910 (N_10910,N_4536,N_721);
nor U10911 (N_10911,N_1482,N_5763);
or U10912 (N_10912,N_2353,N_3012);
xor U10913 (N_10913,N_437,N_5546);
nor U10914 (N_10914,N_2960,N_5862);
nand U10915 (N_10915,N_5216,N_761);
nand U10916 (N_10916,N_1085,N_3668);
or U10917 (N_10917,N_5047,N_3228);
and U10918 (N_10918,N_5722,N_1463);
nor U10919 (N_10919,N_5677,N_4891);
nand U10920 (N_10920,N_4517,N_4172);
nand U10921 (N_10921,N_2870,N_5320);
nand U10922 (N_10922,N_4816,N_655);
or U10923 (N_10923,N_2516,N_1489);
nand U10924 (N_10924,N_6208,N_4388);
xnor U10925 (N_10925,N_293,N_5832);
or U10926 (N_10926,N_3037,N_495);
xnor U10927 (N_10927,N_4828,N_2948);
nand U10928 (N_10928,N_3095,N_165);
nand U10929 (N_10929,N_3979,N_119);
nand U10930 (N_10930,N_3542,N_26);
and U10931 (N_10931,N_1861,N_3985);
and U10932 (N_10932,N_3137,N_3074);
xnor U10933 (N_10933,N_38,N_3311);
xor U10934 (N_10934,N_734,N_1498);
or U10935 (N_10935,N_5514,N_2439);
or U10936 (N_10936,N_4022,N_3268);
xor U10937 (N_10937,N_4775,N_377);
nand U10938 (N_10938,N_4671,N_3331);
nand U10939 (N_10939,N_4797,N_1768);
or U10940 (N_10940,N_4973,N_3257);
and U10941 (N_10941,N_4134,N_5008);
nand U10942 (N_10942,N_5874,N_5742);
nand U10943 (N_10943,N_4214,N_1656);
or U10944 (N_10944,N_6173,N_147);
nand U10945 (N_10945,N_2853,N_3656);
or U10946 (N_10946,N_4486,N_2871);
nor U10947 (N_10947,N_4011,N_2928);
or U10948 (N_10948,N_5338,N_4308);
or U10949 (N_10949,N_2856,N_3969);
nor U10950 (N_10950,N_1492,N_2300);
nand U10951 (N_10951,N_2750,N_2989);
nor U10952 (N_10952,N_5136,N_5292);
nand U10953 (N_10953,N_3691,N_4892);
nor U10954 (N_10954,N_3128,N_2974);
nor U10955 (N_10955,N_267,N_4033);
and U10956 (N_10956,N_4389,N_4501);
and U10957 (N_10957,N_1226,N_211);
xnor U10958 (N_10958,N_4043,N_2613);
and U10959 (N_10959,N_4840,N_2182);
nand U10960 (N_10960,N_3209,N_372);
nand U10961 (N_10961,N_861,N_3409);
nand U10962 (N_10962,N_3610,N_5452);
xnor U10963 (N_10963,N_3729,N_2020);
xor U10964 (N_10964,N_4408,N_4673);
or U10965 (N_10965,N_5262,N_4126);
nor U10966 (N_10966,N_331,N_5183);
and U10967 (N_10967,N_5819,N_5011);
nor U10968 (N_10968,N_5108,N_5621);
nor U10969 (N_10969,N_868,N_5425);
nand U10970 (N_10970,N_1037,N_104);
nand U10971 (N_10971,N_2195,N_4304);
xor U10972 (N_10972,N_2914,N_6019);
and U10973 (N_10973,N_3210,N_1815);
and U10974 (N_10974,N_4501,N_5816);
and U10975 (N_10975,N_1149,N_3115);
xnor U10976 (N_10976,N_4363,N_396);
nand U10977 (N_10977,N_2360,N_391);
or U10978 (N_10978,N_5514,N_6113);
or U10979 (N_10979,N_876,N_5227);
nand U10980 (N_10980,N_18,N_4672);
or U10981 (N_10981,N_3127,N_6058);
or U10982 (N_10982,N_4852,N_4646);
and U10983 (N_10983,N_1564,N_3423);
or U10984 (N_10984,N_3115,N_2900);
or U10985 (N_10985,N_670,N_134);
and U10986 (N_10986,N_4837,N_1884);
and U10987 (N_10987,N_2813,N_2894);
nor U10988 (N_10988,N_4096,N_562);
nor U10989 (N_10989,N_2763,N_2808);
nor U10990 (N_10990,N_2032,N_3079);
xnor U10991 (N_10991,N_5593,N_462);
and U10992 (N_10992,N_1406,N_3685);
or U10993 (N_10993,N_5169,N_2531);
or U10994 (N_10994,N_4926,N_2689);
nand U10995 (N_10995,N_6199,N_375);
nand U10996 (N_10996,N_464,N_3882);
nand U10997 (N_10997,N_312,N_5829);
nor U10998 (N_10998,N_4239,N_5078);
and U10999 (N_10999,N_5222,N_1314);
and U11000 (N_11000,N_4412,N_2672);
and U11001 (N_11001,N_3444,N_4112);
nor U11002 (N_11002,N_5245,N_1582);
nand U11003 (N_11003,N_4516,N_5031);
or U11004 (N_11004,N_5007,N_25);
nor U11005 (N_11005,N_1057,N_413);
nor U11006 (N_11006,N_1592,N_6244);
nand U11007 (N_11007,N_968,N_4712);
nor U11008 (N_11008,N_5023,N_1749);
or U11009 (N_11009,N_5404,N_2578);
or U11010 (N_11010,N_1567,N_2556);
and U11011 (N_11011,N_2088,N_1408);
nand U11012 (N_11012,N_2581,N_5457);
or U11013 (N_11013,N_1345,N_837);
nor U11014 (N_11014,N_5781,N_4459);
nor U11015 (N_11015,N_1494,N_6065);
and U11016 (N_11016,N_3669,N_4699);
xor U11017 (N_11017,N_4700,N_819);
and U11018 (N_11018,N_1013,N_3393);
nor U11019 (N_11019,N_4849,N_565);
nand U11020 (N_11020,N_4330,N_3124);
nor U11021 (N_11021,N_5923,N_1952);
or U11022 (N_11022,N_45,N_1362);
nor U11023 (N_11023,N_5302,N_3038);
or U11024 (N_11024,N_3250,N_4767);
nor U11025 (N_11025,N_3858,N_2562);
nand U11026 (N_11026,N_2429,N_819);
nand U11027 (N_11027,N_1958,N_5798);
and U11028 (N_11028,N_1687,N_2020);
nor U11029 (N_11029,N_2851,N_3464);
and U11030 (N_11030,N_1575,N_1337);
or U11031 (N_11031,N_1552,N_4381);
or U11032 (N_11032,N_5185,N_5671);
xnor U11033 (N_11033,N_4361,N_5468);
xnor U11034 (N_11034,N_5955,N_4936);
or U11035 (N_11035,N_2336,N_3064);
xnor U11036 (N_11036,N_1127,N_788);
nor U11037 (N_11037,N_402,N_4616);
or U11038 (N_11038,N_3834,N_928);
xnor U11039 (N_11039,N_4881,N_5290);
nor U11040 (N_11040,N_2383,N_1815);
and U11041 (N_11041,N_4297,N_5876);
nor U11042 (N_11042,N_3819,N_1405);
and U11043 (N_11043,N_2758,N_4534);
nor U11044 (N_11044,N_196,N_404);
nor U11045 (N_11045,N_301,N_2249);
or U11046 (N_11046,N_3793,N_878);
and U11047 (N_11047,N_5263,N_3453);
nand U11048 (N_11048,N_3672,N_5073);
nand U11049 (N_11049,N_1837,N_2494);
and U11050 (N_11050,N_1721,N_4008);
or U11051 (N_11051,N_1458,N_3962);
nor U11052 (N_11052,N_2870,N_2513);
nor U11053 (N_11053,N_708,N_1200);
or U11054 (N_11054,N_6011,N_2607);
or U11055 (N_11055,N_5129,N_5097);
nand U11056 (N_11056,N_4878,N_270);
nand U11057 (N_11057,N_4326,N_6018);
nor U11058 (N_11058,N_4121,N_4354);
and U11059 (N_11059,N_577,N_5560);
nor U11060 (N_11060,N_1551,N_77);
xor U11061 (N_11061,N_5052,N_3096);
xor U11062 (N_11062,N_4382,N_3335);
and U11063 (N_11063,N_3127,N_3720);
and U11064 (N_11064,N_6187,N_4833);
and U11065 (N_11065,N_5647,N_2690);
and U11066 (N_11066,N_4653,N_4898);
nand U11067 (N_11067,N_3354,N_5468);
and U11068 (N_11068,N_1319,N_3058);
nor U11069 (N_11069,N_1499,N_5879);
and U11070 (N_11070,N_6149,N_231);
nor U11071 (N_11071,N_2478,N_6218);
nand U11072 (N_11072,N_5566,N_1742);
nor U11073 (N_11073,N_392,N_3564);
or U11074 (N_11074,N_2473,N_4212);
nor U11075 (N_11075,N_4103,N_2002);
xor U11076 (N_11076,N_4558,N_3988);
and U11077 (N_11077,N_1992,N_964);
and U11078 (N_11078,N_676,N_25);
and U11079 (N_11079,N_4266,N_1784);
and U11080 (N_11080,N_148,N_2423);
nand U11081 (N_11081,N_3598,N_3733);
or U11082 (N_11082,N_1550,N_993);
and U11083 (N_11083,N_246,N_2930);
or U11084 (N_11084,N_1649,N_3430);
nand U11085 (N_11085,N_912,N_2640);
nor U11086 (N_11086,N_3319,N_4090);
nor U11087 (N_11087,N_1043,N_795);
or U11088 (N_11088,N_793,N_1229);
and U11089 (N_11089,N_5904,N_3786);
and U11090 (N_11090,N_3730,N_4565);
nor U11091 (N_11091,N_1385,N_5085);
nor U11092 (N_11092,N_4493,N_5970);
or U11093 (N_11093,N_4890,N_4674);
nand U11094 (N_11094,N_2059,N_1342);
nor U11095 (N_11095,N_832,N_5323);
nand U11096 (N_11096,N_88,N_1666);
xor U11097 (N_11097,N_5462,N_1244);
nand U11098 (N_11098,N_5059,N_6169);
and U11099 (N_11099,N_2806,N_1176);
or U11100 (N_11100,N_2015,N_4081);
nand U11101 (N_11101,N_522,N_107);
xnor U11102 (N_11102,N_5306,N_1956);
or U11103 (N_11103,N_4727,N_6079);
xnor U11104 (N_11104,N_1768,N_4407);
xor U11105 (N_11105,N_3101,N_3366);
nor U11106 (N_11106,N_5357,N_4556);
or U11107 (N_11107,N_2931,N_1054);
nand U11108 (N_11108,N_1936,N_2699);
or U11109 (N_11109,N_1921,N_2748);
and U11110 (N_11110,N_3834,N_5812);
nor U11111 (N_11111,N_2339,N_1028);
nand U11112 (N_11112,N_4158,N_3610);
and U11113 (N_11113,N_2752,N_3866);
and U11114 (N_11114,N_2883,N_4241);
nor U11115 (N_11115,N_5916,N_1859);
nor U11116 (N_11116,N_244,N_3624);
nor U11117 (N_11117,N_4120,N_2936);
nor U11118 (N_11118,N_964,N_800);
nand U11119 (N_11119,N_1031,N_5553);
xnor U11120 (N_11120,N_5911,N_2265);
or U11121 (N_11121,N_2959,N_1207);
nand U11122 (N_11122,N_6010,N_108);
or U11123 (N_11123,N_4459,N_5432);
nor U11124 (N_11124,N_408,N_945);
nand U11125 (N_11125,N_4511,N_3538);
nand U11126 (N_11126,N_4330,N_914);
and U11127 (N_11127,N_1400,N_1940);
nor U11128 (N_11128,N_5894,N_985);
or U11129 (N_11129,N_5176,N_436);
or U11130 (N_11130,N_485,N_3309);
nand U11131 (N_11131,N_1670,N_2058);
nand U11132 (N_11132,N_2694,N_3125);
or U11133 (N_11133,N_955,N_3507);
nand U11134 (N_11134,N_2248,N_5054);
or U11135 (N_11135,N_2073,N_3489);
and U11136 (N_11136,N_6155,N_100);
nor U11137 (N_11137,N_2172,N_3227);
nand U11138 (N_11138,N_1219,N_5116);
or U11139 (N_11139,N_2092,N_4937);
nand U11140 (N_11140,N_607,N_4512);
nor U11141 (N_11141,N_466,N_1465);
nand U11142 (N_11142,N_2199,N_2269);
or U11143 (N_11143,N_5602,N_3362);
or U11144 (N_11144,N_2201,N_1138);
nand U11145 (N_11145,N_3008,N_3646);
or U11146 (N_11146,N_2404,N_4341);
nor U11147 (N_11147,N_5360,N_978);
nand U11148 (N_11148,N_1848,N_3460);
and U11149 (N_11149,N_3927,N_1872);
xnor U11150 (N_11150,N_5749,N_2357);
nand U11151 (N_11151,N_1808,N_5489);
or U11152 (N_11152,N_5089,N_4214);
and U11153 (N_11153,N_5837,N_280);
nand U11154 (N_11154,N_688,N_2093);
or U11155 (N_11155,N_5244,N_2427);
nand U11156 (N_11156,N_0,N_3749);
and U11157 (N_11157,N_139,N_3280);
nand U11158 (N_11158,N_3149,N_4131);
or U11159 (N_11159,N_4271,N_6080);
nor U11160 (N_11160,N_3065,N_3564);
and U11161 (N_11161,N_2292,N_5663);
nor U11162 (N_11162,N_1072,N_983);
nor U11163 (N_11163,N_3182,N_2844);
nand U11164 (N_11164,N_3973,N_1269);
or U11165 (N_11165,N_1349,N_1679);
xnor U11166 (N_11166,N_369,N_5943);
nor U11167 (N_11167,N_1106,N_5199);
nor U11168 (N_11168,N_1686,N_2560);
and U11169 (N_11169,N_5422,N_4805);
xnor U11170 (N_11170,N_3591,N_3004);
nor U11171 (N_11171,N_5659,N_336);
or U11172 (N_11172,N_4070,N_1714);
nor U11173 (N_11173,N_4137,N_2850);
and U11174 (N_11174,N_4953,N_3675);
nor U11175 (N_11175,N_3829,N_5953);
and U11176 (N_11176,N_405,N_2677);
nor U11177 (N_11177,N_6217,N_5355);
nor U11178 (N_11178,N_761,N_6055);
nor U11179 (N_11179,N_3964,N_746);
nand U11180 (N_11180,N_42,N_3466);
nand U11181 (N_11181,N_2870,N_116);
nor U11182 (N_11182,N_4455,N_361);
and U11183 (N_11183,N_42,N_920);
or U11184 (N_11184,N_1315,N_3538);
or U11185 (N_11185,N_2514,N_922);
nor U11186 (N_11186,N_2890,N_1940);
and U11187 (N_11187,N_5659,N_3582);
nor U11188 (N_11188,N_1290,N_2438);
and U11189 (N_11189,N_3056,N_4336);
and U11190 (N_11190,N_74,N_558);
nand U11191 (N_11191,N_2928,N_4138);
xnor U11192 (N_11192,N_3783,N_4691);
nand U11193 (N_11193,N_428,N_1224);
nor U11194 (N_11194,N_5156,N_235);
nor U11195 (N_11195,N_1943,N_2315);
or U11196 (N_11196,N_5801,N_3549);
or U11197 (N_11197,N_4845,N_1722);
nand U11198 (N_11198,N_2003,N_4888);
and U11199 (N_11199,N_4424,N_252);
nor U11200 (N_11200,N_823,N_6196);
or U11201 (N_11201,N_360,N_2847);
and U11202 (N_11202,N_5111,N_4137);
xnor U11203 (N_11203,N_5433,N_3966);
or U11204 (N_11204,N_4905,N_545);
or U11205 (N_11205,N_3177,N_4106);
nand U11206 (N_11206,N_4012,N_3559);
and U11207 (N_11207,N_4431,N_2106);
nor U11208 (N_11208,N_2070,N_947);
nand U11209 (N_11209,N_5141,N_2093);
and U11210 (N_11210,N_2189,N_2934);
nor U11211 (N_11211,N_3970,N_2903);
or U11212 (N_11212,N_158,N_3475);
nor U11213 (N_11213,N_1082,N_10);
nor U11214 (N_11214,N_2426,N_640);
or U11215 (N_11215,N_513,N_1151);
and U11216 (N_11216,N_5578,N_4799);
nor U11217 (N_11217,N_1589,N_2983);
xnor U11218 (N_11218,N_44,N_997);
and U11219 (N_11219,N_273,N_6059);
or U11220 (N_11220,N_6226,N_6146);
nor U11221 (N_11221,N_2666,N_3859);
nand U11222 (N_11222,N_176,N_2252);
nand U11223 (N_11223,N_1794,N_1490);
and U11224 (N_11224,N_4291,N_1407);
and U11225 (N_11225,N_4139,N_1820);
and U11226 (N_11226,N_449,N_4988);
nand U11227 (N_11227,N_3141,N_140);
or U11228 (N_11228,N_3580,N_4446);
nor U11229 (N_11229,N_252,N_886);
nor U11230 (N_11230,N_6169,N_3496);
nor U11231 (N_11231,N_833,N_1182);
nor U11232 (N_11232,N_2972,N_275);
nor U11233 (N_11233,N_1767,N_5402);
and U11234 (N_11234,N_5778,N_4221);
nor U11235 (N_11235,N_2712,N_3337);
or U11236 (N_11236,N_1889,N_4768);
and U11237 (N_11237,N_4254,N_497);
nand U11238 (N_11238,N_2036,N_1391);
xor U11239 (N_11239,N_1880,N_1254);
nand U11240 (N_11240,N_188,N_5216);
xnor U11241 (N_11241,N_2184,N_5418);
and U11242 (N_11242,N_472,N_813);
or U11243 (N_11243,N_2532,N_1052);
nand U11244 (N_11244,N_247,N_3108);
nor U11245 (N_11245,N_1397,N_2635);
or U11246 (N_11246,N_4629,N_3460);
or U11247 (N_11247,N_4645,N_5584);
and U11248 (N_11248,N_3530,N_4291);
xor U11249 (N_11249,N_2371,N_115);
nor U11250 (N_11250,N_2652,N_5318);
and U11251 (N_11251,N_2729,N_3868);
xor U11252 (N_11252,N_1565,N_4640);
and U11253 (N_11253,N_5030,N_676);
and U11254 (N_11254,N_615,N_2802);
xor U11255 (N_11255,N_345,N_4154);
nand U11256 (N_11256,N_4767,N_4068);
and U11257 (N_11257,N_4148,N_2753);
or U11258 (N_11258,N_3137,N_1591);
and U11259 (N_11259,N_1587,N_6172);
nor U11260 (N_11260,N_5991,N_2348);
nor U11261 (N_11261,N_5009,N_3406);
nand U11262 (N_11262,N_6123,N_1788);
and U11263 (N_11263,N_2178,N_3896);
or U11264 (N_11264,N_4746,N_5021);
or U11265 (N_11265,N_3392,N_36);
xnor U11266 (N_11266,N_5477,N_1726);
nand U11267 (N_11267,N_4797,N_770);
and U11268 (N_11268,N_3723,N_4062);
or U11269 (N_11269,N_3768,N_3250);
xor U11270 (N_11270,N_5025,N_2922);
or U11271 (N_11271,N_3008,N_450);
xnor U11272 (N_11272,N_403,N_1966);
and U11273 (N_11273,N_4721,N_801);
nand U11274 (N_11274,N_1360,N_4186);
and U11275 (N_11275,N_866,N_3517);
nand U11276 (N_11276,N_5580,N_3541);
nor U11277 (N_11277,N_3495,N_934);
nand U11278 (N_11278,N_6234,N_1454);
nand U11279 (N_11279,N_341,N_4774);
xnor U11280 (N_11280,N_1362,N_2288);
or U11281 (N_11281,N_4845,N_4938);
nand U11282 (N_11282,N_477,N_5667);
and U11283 (N_11283,N_5827,N_4237);
and U11284 (N_11284,N_5276,N_3828);
nand U11285 (N_11285,N_6108,N_4891);
nand U11286 (N_11286,N_3414,N_3517);
nor U11287 (N_11287,N_434,N_4589);
nor U11288 (N_11288,N_1246,N_2361);
nand U11289 (N_11289,N_6204,N_741);
nor U11290 (N_11290,N_2714,N_2293);
xor U11291 (N_11291,N_3712,N_5509);
and U11292 (N_11292,N_1743,N_2826);
nand U11293 (N_11293,N_483,N_1573);
and U11294 (N_11294,N_3701,N_647);
nand U11295 (N_11295,N_5466,N_3817);
nand U11296 (N_11296,N_5663,N_4285);
nor U11297 (N_11297,N_569,N_4681);
and U11298 (N_11298,N_2901,N_1860);
and U11299 (N_11299,N_5957,N_859);
or U11300 (N_11300,N_3225,N_5581);
or U11301 (N_11301,N_2384,N_4158);
nor U11302 (N_11302,N_1874,N_3549);
nand U11303 (N_11303,N_1728,N_636);
nor U11304 (N_11304,N_3880,N_3515);
nand U11305 (N_11305,N_207,N_398);
and U11306 (N_11306,N_227,N_74);
nor U11307 (N_11307,N_2688,N_817);
and U11308 (N_11308,N_909,N_1262);
or U11309 (N_11309,N_6112,N_1062);
nor U11310 (N_11310,N_4282,N_402);
and U11311 (N_11311,N_5633,N_4521);
nand U11312 (N_11312,N_191,N_1967);
nand U11313 (N_11313,N_637,N_2964);
or U11314 (N_11314,N_5428,N_4766);
and U11315 (N_11315,N_4881,N_5764);
and U11316 (N_11316,N_2012,N_6080);
nor U11317 (N_11317,N_2621,N_2678);
and U11318 (N_11318,N_3721,N_5130);
nor U11319 (N_11319,N_818,N_6144);
nand U11320 (N_11320,N_2239,N_79);
or U11321 (N_11321,N_4664,N_1423);
and U11322 (N_11322,N_2078,N_4113);
and U11323 (N_11323,N_961,N_2948);
xor U11324 (N_11324,N_1380,N_2011);
nand U11325 (N_11325,N_4215,N_3629);
nor U11326 (N_11326,N_5694,N_2756);
nand U11327 (N_11327,N_1277,N_5566);
nor U11328 (N_11328,N_1213,N_2701);
nand U11329 (N_11329,N_3630,N_748);
nor U11330 (N_11330,N_3045,N_3358);
and U11331 (N_11331,N_2342,N_4628);
nand U11332 (N_11332,N_3831,N_4444);
nor U11333 (N_11333,N_1723,N_3788);
xor U11334 (N_11334,N_3154,N_2911);
xnor U11335 (N_11335,N_1949,N_336);
nand U11336 (N_11336,N_732,N_1489);
xor U11337 (N_11337,N_1154,N_3488);
nor U11338 (N_11338,N_2568,N_1844);
nand U11339 (N_11339,N_3475,N_164);
nand U11340 (N_11340,N_3838,N_2339);
nor U11341 (N_11341,N_2464,N_1505);
nor U11342 (N_11342,N_5614,N_521);
nor U11343 (N_11343,N_5547,N_6093);
xnor U11344 (N_11344,N_5294,N_2345);
nor U11345 (N_11345,N_5104,N_645);
and U11346 (N_11346,N_4022,N_4955);
nand U11347 (N_11347,N_3689,N_540);
nor U11348 (N_11348,N_1085,N_3599);
and U11349 (N_11349,N_4859,N_672);
and U11350 (N_11350,N_5291,N_5142);
nor U11351 (N_11351,N_1896,N_2990);
and U11352 (N_11352,N_2852,N_1191);
nand U11353 (N_11353,N_4529,N_5752);
xnor U11354 (N_11354,N_1455,N_5083);
and U11355 (N_11355,N_1467,N_2615);
nor U11356 (N_11356,N_3915,N_1738);
and U11357 (N_11357,N_709,N_2332);
nand U11358 (N_11358,N_5286,N_1252);
nand U11359 (N_11359,N_5090,N_305);
and U11360 (N_11360,N_5242,N_1434);
nor U11361 (N_11361,N_5371,N_2561);
or U11362 (N_11362,N_2820,N_3971);
nor U11363 (N_11363,N_3193,N_2881);
nor U11364 (N_11364,N_5813,N_3304);
or U11365 (N_11365,N_5660,N_3976);
nor U11366 (N_11366,N_3154,N_948);
nor U11367 (N_11367,N_5964,N_1772);
and U11368 (N_11368,N_4465,N_5403);
nor U11369 (N_11369,N_5449,N_4870);
and U11370 (N_11370,N_5260,N_2134);
and U11371 (N_11371,N_1056,N_4490);
or U11372 (N_11372,N_2196,N_5468);
nand U11373 (N_11373,N_6114,N_5202);
nand U11374 (N_11374,N_11,N_322);
or U11375 (N_11375,N_773,N_5523);
and U11376 (N_11376,N_6065,N_4578);
or U11377 (N_11377,N_1320,N_6153);
and U11378 (N_11378,N_483,N_1121);
nand U11379 (N_11379,N_4190,N_2721);
or U11380 (N_11380,N_1924,N_4439);
xor U11381 (N_11381,N_2665,N_2356);
xnor U11382 (N_11382,N_2584,N_1231);
nand U11383 (N_11383,N_3373,N_4495);
and U11384 (N_11384,N_3781,N_519);
nor U11385 (N_11385,N_5751,N_1979);
or U11386 (N_11386,N_6004,N_3313);
and U11387 (N_11387,N_2957,N_4467);
nor U11388 (N_11388,N_779,N_1749);
nand U11389 (N_11389,N_2610,N_1827);
or U11390 (N_11390,N_121,N_2194);
nor U11391 (N_11391,N_2666,N_5535);
nor U11392 (N_11392,N_1411,N_6044);
nor U11393 (N_11393,N_3243,N_1146);
and U11394 (N_11394,N_679,N_1272);
and U11395 (N_11395,N_713,N_1116);
or U11396 (N_11396,N_4236,N_814);
nand U11397 (N_11397,N_5081,N_2127);
or U11398 (N_11398,N_1700,N_5713);
nand U11399 (N_11399,N_4654,N_1564);
nor U11400 (N_11400,N_5849,N_5053);
nand U11401 (N_11401,N_1909,N_9);
or U11402 (N_11402,N_2644,N_3567);
xnor U11403 (N_11403,N_3869,N_1230);
or U11404 (N_11404,N_2250,N_5608);
and U11405 (N_11405,N_2892,N_4313);
nor U11406 (N_11406,N_3073,N_4250);
and U11407 (N_11407,N_30,N_3874);
nor U11408 (N_11408,N_4886,N_561);
or U11409 (N_11409,N_5152,N_872);
nor U11410 (N_11410,N_559,N_43);
nor U11411 (N_11411,N_2284,N_4757);
xnor U11412 (N_11412,N_3772,N_6151);
and U11413 (N_11413,N_5322,N_3766);
xnor U11414 (N_11414,N_2281,N_1361);
and U11415 (N_11415,N_17,N_5925);
nor U11416 (N_11416,N_4538,N_54);
nor U11417 (N_11417,N_4831,N_4951);
or U11418 (N_11418,N_6233,N_4634);
and U11419 (N_11419,N_141,N_1824);
nor U11420 (N_11420,N_1733,N_652);
nor U11421 (N_11421,N_6224,N_4195);
or U11422 (N_11422,N_3795,N_3153);
xnor U11423 (N_11423,N_4463,N_854);
and U11424 (N_11424,N_304,N_245);
nand U11425 (N_11425,N_2937,N_222);
or U11426 (N_11426,N_3722,N_1431);
and U11427 (N_11427,N_5346,N_5530);
and U11428 (N_11428,N_5663,N_3856);
or U11429 (N_11429,N_6025,N_5595);
nand U11430 (N_11430,N_3429,N_2646);
nand U11431 (N_11431,N_804,N_4884);
or U11432 (N_11432,N_3965,N_2545);
nand U11433 (N_11433,N_5942,N_3510);
nand U11434 (N_11434,N_3623,N_2958);
or U11435 (N_11435,N_2390,N_790);
nor U11436 (N_11436,N_5507,N_2479);
xnor U11437 (N_11437,N_587,N_5373);
nor U11438 (N_11438,N_2831,N_4383);
or U11439 (N_11439,N_4119,N_5613);
or U11440 (N_11440,N_4009,N_1325);
nand U11441 (N_11441,N_3979,N_3643);
nand U11442 (N_11442,N_3073,N_4974);
or U11443 (N_11443,N_1696,N_903);
nor U11444 (N_11444,N_3074,N_5475);
and U11445 (N_11445,N_3848,N_83);
or U11446 (N_11446,N_2882,N_1855);
or U11447 (N_11447,N_2169,N_3678);
nor U11448 (N_11448,N_3540,N_4663);
nor U11449 (N_11449,N_1002,N_1729);
or U11450 (N_11450,N_4254,N_4085);
nor U11451 (N_11451,N_5814,N_4423);
and U11452 (N_11452,N_3970,N_101);
nor U11453 (N_11453,N_2051,N_5197);
xnor U11454 (N_11454,N_5173,N_641);
nand U11455 (N_11455,N_5789,N_736);
nand U11456 (N_11456,N_1986,N_4921);
and U11457 (N_11457,N_6049,N_871);
and U11458 (N_11458,N_4946,N_373);
or U11459 (N_11459,N_4529,N_3989);
or U11460 (N_11460,N_4475,N_4923);
and U11461 (N_11461,N_5797,N_4279);
nor U11462 (N_11462,N_4587,N_4396);
nand U11463 (N_11463,N_2547,N_4408);
nand U11464 (N_11464,N_4535,N_2000);
and U11465 (N_11465,N_5029,N_614);
nor U11466 (N_11466,N_1762,N_5756);
nand U11467 (N_11467,N_3606,N_4651);
nand U11468 (N_11468,N_3870,N_2439);
or U11469 (N_11469,N_1204,N_2087);
and U11470 (N_11470,N_3438,N_6171);
nor U11471 (N_11471,N_5028,N_224);
or U11472 (N_11472,N_3322,N_2249);
or U11473 (N_11473,N_4032,N_2058);
or U11474 (N_11474,N_2405,N_5516);
and U11475 (N_11475,N_3764,N_5341);
or U11476 (N_11476,N_1332,N_1628);
or U11477 (N_11477,N_5297,N_995);
nand U11478 (N_11478,N_3013,N_4622);
nand U11479 (N_11479,N_731,N_3323);
and U11480 (N_11480,N_3902,N_2082);
nand U11481 (N_11481,N_4214,N_6145);
nor U11482 (N_11482,N_4832,N_1219);
and U11483 (N_11483,N_118,N_3801);
nor U11484 (N_11484,N_2916,N_1336);
nand U11485 (N_11485,N_5502,N_5604);
or U11486 (N_11486,N_2626,N_14);
or U11487 (N_11487,N_137,N_3191);
and U11488 (N_11488,N_2025,N_1443);
xnor U11489 (N_11489,N_4555,N_2987);
xnor U11490 (N_11490,N_4167,N_5816);
and U11491 (N_11491,N_438,N_5170);
nand U11492 (N_11492,N_501,N_5497);
xor U11493 (N_11493,N_4748,N_5316);
nand U11494 (N_11494,N_175,N_2096);
and U11495 (N_11495,N_1081,N_2231);
and U11496 (N_11496,N_5460,N_4192);
and U11497 (N_11497,N_4253,N_2169);
and U11498 (N_11498,N_3121,N_3821);
or U11499 (N_11499,N_268,N_2931);
xor U11500 (N_11500,N_2411,N_5748);
nand U11501 (N_11501,N_591,N_2734);
or U11502 (N_11502,N_1771,N_13);
and U11503 (N_11503,N_1169,N_3671);
and U11504 (N_11504,N_4311,N_1028);
nor U11505 (N_11505,N_5531,N_5796);
and U11506 (N_11506,N_3211,N_3439);
nor U11507 (N_11507,N_2949,N_1310);
nor U11508 (N_11508,N_987,N_586);
nor U11509 (N_11509,N_2916,N_3790);
and U11510 (N_11510,N_4361,N_817);
or U11511 (N_11511,N_3765,N_2630);
and U11512 (N_11512,N_3552,N_2559);
and U11513 (N_11513,N_1716,N_1727);
or U11514 (N_11514,N_1466,N_583);
nand U11515 (N_11515,N_4987,N_1618);
or U11516 (N_11516,N_5396,N_2855);
nand U11517 (N_11517,N_2186,N_3440);
nand U11518 (N_11518,N_1984,N_4075);
and U11519 (N_11519,N_3103,N_2092);
or U11520 (N_11520,N_2502,N_3185);
nor U11521 (N_11521,N_4940,N_372);
or U11522 (N_11522,N_5019,N_3290);
nor U11523 (N_11523,N_2097,N_3297);
or U11524 (N_11524,N_29,N_3405);
or U11525 (N_11525,N_3195,N_3578);
and U11526 (N_11526,N_5652,N_6080);
or U11527 (N_11527,N_4607,N_2516);
nor U11528 (N_11528,N_5337,N_2323);
and U11529 (N_11529,N_6069,N_5958);
or U11530 (N_11530,N_2700,N_4419);
nand U11531 (N_11531,N_3711,N_2355);
nand U11532 (N_11532,N_4690,N_3729);
nand U11533 (N_11533,N_3915,N_5600);
or U11534 (N_11534,N_381,N_1126);
nand U11535 (N_11535,N_2252,N_1413);
nand U11536 (N_11536,N_3508,N_4459);
nand U11537 (N_11537,N_5869,N_2140);
nand U11538 (N_11538,N_192,N_737);
nor U11539 (N_11539,N_2756,N_2479);
or U11540 (N_11540,N_6155,N_4401);
and U11541 (N_11541,N_3232,N_3925);
and U11542 (N_11542,N_2048,N_2144);
or U11543 (N_11543,N_2170,N_4778);
and U11544 (N_11544,N_4677,N_5298);
and U11545 (N_11545,N_5868,N_2110);
nand U11546 (N_11546,N_2686,N_22);
and U11547 (N_11547,N_4214,N_272);
and U11548 (N_11548,N_147,N_2933);
or U11549 (N_11549,N_4426,N_4078);
or U11550 (N_11550,N_4763,N_3891);
and U11551 (N_11551,N_1469,N_1066);
and U11552 (N_11552,N_2195,N_705);
and U11553 (N_11553,N_4070,N_5867);
and U11554 (N_11554,N_3577,N_1041);
or U11555 (N_11555,N_5034,N_5548);
and U11556 (N_11556,N_1771,N_2513);
or U11557 (N_11557,N_1556,N_3070);
nor U11558 (N_11558,N_960,N_2242);
and U11559 (N_11559,N_2675,N_6230);
and U11560 (N_11560,N_1661,N_4311);
or U11561 (N_11561,N_985,N_571);
nand U11562 (N_11562,N_4308,N_1917);
xor U11563 (N_11563,N_1648,N_3316);
or U11564 (N_11564,N_4107,N_5330);
nand U11565 (N_11565,N_1255,N_3235);
nand U11566 (N_11566,N_2519,N_1740);
or U11567 (N_11567,N_1581,N_5800);
and U11568 (N_11568,N_5784,N_4429);
nor U11569 (N_11569,N_1436,N_1790);
nor U11570 (N_11570,N_3029,N_587);
or U11571 (N_11571,N_390,N_2073);
or U11572 (N_11572,N_5631,N_5774);
and U11573 (N_11573,N_2367,N_4469);
xnor U11574 (N_11574,N_417,N_4085);
nand U11575 (N_11575,N_3454,N_2673);
nand U11576 (N_11576,N_5251,N_2787);
nand U11577 (N_11577,N_1663,N_2279);
or U11578 (N_11578,N_3237,N_2139);
and U11579 (N_11579,N_4416,N_1597);
xnor U11580 (N_11580,N_3860,N_3545);
nor U11581 (N_11581,N_4538,N_5813);
nand U11582 (N_11582,N_3426,N_3915);
or U11583 (N_11583,N_3864,N_5167);
nand U11584 (N_11584,N_866,N_1493);
xor U11585 (N_11585,N_1059,N_4033);
and U11586 (N_11586,N_4727,N_4491);
and U11587 (N_11587,N_5999,N_1578);
nor U11588 (N_11588,N_1646,N_3460);
or U11589 (N_11589,N_5182,N_1543);
and U11590 (N_11590,N_2483,N_5885);
and U11591 (N_11591,N_2792,N_5908);
nor U11592 (N_11592,N_3972,N_6102);
and U11593 (N_11593,N_592,N_3122);
nand U11594 (N_11594,N_5798,N_915);
nand U11595 (N_11595,N_3944,N_1697);
and U11596 (N_11596,N_2737,N_3277);
nand U11597 (N_11597,N_991,N_3638);
nand U11598 (N_11598,N_1791,N_3685);
nor U11599 (N_11599,N_3269,N_3455);
and U11600 (N_11600,N_3440,N_4885);
and U11601 (N_11601,N_2103,N_6221);
nand U11602 (N_11602,N_5870,N_5290);
or U11603 (N_11603,N_572,N_1465);
xor U11604 (N_11604,N_3132,N_3696);
nand U11605 (N_11605,N_3158,N_2708);
and U11606 (N_11606,N_2640,N_5927);
nand U11607 (N_11607,N_1862,N_5101);
and U11608 (N_11608,N_5937,N_2819);
and U11609 (N_11609,N_1525,N_2188);
nand U11610 (N_11610,N_257,N_3004);
and U11611 (N_11611,N_6243,N_2533);
and U11612 (N_11612,N_5961,N_1881);
nand U11613 (N_11613,N_1709,N_4873);
nor U11614 (N_11614,N_5959,N_4103);
nor U11615 (N_11615,N_1391,N_5050);
nor U11616 (N_11616,N_835,N_2850);
or U11617 (N_11617,N_2728,N_4656);
or U11618 (N_11618,N_5681,N_4829);
nand U11619 (N_11619,N_3581,N_4375);
or U11620 (N_11620,N_768,N_5293);
and U11621 (N_11621,N_1654,N_5116);
nand U11622 (N_11622,N_1553,N_5633);
and U11623 (N_11623,N_4327,N_3955);
nand U11624 (N_11624,N_729,N_3183);
and U11625 (N_11625,N_5248,N_375);
or U11626 (N_11626,N_5320,N_4298);
or U11627 (N_11627,N_3530,N_6234);
and U11628 (N_11628,N_3524,N_3609);
and U11629 (N_11629,N_991,N_5200);
or U11630 (N_11630,N_4262,N_3570);
xnor U11631 (N_11631,N_2331,N_1115);
or U11632 (N_11632,N_1709,N_2985);
nor U11633 (N_11633,N_3411,N_1721);
and U11634 (N_11634,N_5597,N_1567);
and U11635 (N_11635,N_2785,N_6187);
nor U11636 (N_11636,N_361,N_2655);
nand U11637 (N_11637,N_4321,N_753);
nor U11638 (N_11638,N_3533,N_4839);
and U11639 (N_11639,N_4348,N_2494);
and U11640 (N_11640,N_814,N_3040);
and U11641 (N_11641,N_1438,N_1282);
nand U11642 (N_11642,N_461,N_3823);
nor U11643 (N_11643,N_3806,N_5827);
nor U11644 (N_11644,N_5183,N_1354);
nor U11645 (N_11645,N_1746,N_1239);
nand U11646 (N_11646,N_315,N_2681);
xor U11647 (N_11647,N_3482,N_2157);
xor U11648 (N_11648,N_3695,N_2242);
nand U11649 (N_11649,N_6026,N_3947);
nor U11650 (N_11650,N_4034,N_4509);
and U11651 (N_11651,N_3601,N_1452);
xor U11652 (N_11652,N_222,N_4442);
or U11653 (N_11653,N_2780,N_4438);
and U11654 (N_11654,N_5877,N_4681);
nor U11655 (N_11655,N_1735,N_2672);
nand U11656 (N_11656,N_3800,N_2650);
nand U11657 (N_11657,N_2122,N_1437);
and U11658 (N_11658,N_5663,N_1619);
and U11659 (N_11659,N_2240,N_1071);
and U11660 (N_11660,N_1488,N_5099);
or U11661 (N_11661,N_70,N_3483);
nor U11662 (N_11662,N_200,N_2345);
nand U11663 (N_11663,N_5899,N_1430);
nor U11664 (N_11664,N_6133,N_5202);
nand U11665 (N_11665,N_337,N_1920);
nand U11666 (N_11666,N_316,N_4591);
nor U11667 (N_11667,N_78,N_5397);
nand U11668 (N_11668,N_3112,N_3457);
and U11669 (N_11669,N_1333,N_5705);
or U11670 (N_11670,N_2670,N_988);
xor U11671 (N_11671,N_3232,N_1968);
or U11672 (N_11672,N_1687,N_1829);
and U11673 (N_11673,N_5974,N_4422);
and U11674 (N_11674,N_5475,N_822);
and U11675 (N_11675,N_2721,N_1731);
or U11676 (N_11676,N_856,N_2214);
nand U11677 (N_11677,N_1341,N_4657);
nand U11678 (N_11678,N_6078,N_3629);
or U11679 (N_11679,N_5180,N_6190);
xnor U11680 (N_11680,N_3632,N_2962);
nand U11681 (N_11681,N_1082,N_1213);
nor U11682 (N_11682,N_3011,N_4205);
xnor U11683 (N_11683,N_5806,N_2597);
and U11684 (N_11684,N_757,N_584);
or U11685 (N_11685,N_2145,N_1162);
nand U11686 (N_11686,N_258,N_4020);
nand U11687 (N_11687,N_1136,N_1754);
and U11688 (N_11688,N_1879,N_1736);
and U11689 (N_11689,N_2489,N_1506);
and U11690 (N_11690,N_3523,N_2091);
and U11691 (N_11691,N_627,N_2263);
and U11692 (N_11692,N_131,N_5692);
and U11693 (N_11693,N_1537,N_2788);
nor U11694 (N_11694,N_5767,N_2167);
or U11695 (N_11695,N_5170,N_3434);
nor U11696 (N_11696,N_5673,N_2347);
nand U11697 (N_11697,N_4518,N_587);
nand U11698 (N_11698,N_5670,N_3413);
and U11699 (N_11699,N_6232,N_3127);
nor U11700 (N_11700,N_5193,N_4101);
nand U11701 (N_11701,N_5259,N_521);
or U11702 (N_11702,N_3826,N_5510);
xor U11703 (N_11703,N_248,N_3682);
nor U11704 (N_11704,N_1909,N_5525);
nor U11705 (N_11705,N_411,N_914);
or U11706 (N_11706,N_2052,N_5924);
xnor U11707 (N_11707,N_1655,N_4052);
nor U11708 (N_11708,N_6064,N_1156);
and U11709 (N_11709,N_4516,N_5587);
nor U11710 (N_11710,N_1157,N_4313);
and U11711 (N_11711,N_4455,N_2606);
nand U11712 (N_11712,N_2140,N_3634);
nor U11713 (N_11713,N_5365,N_5395);
xor U11714 (N_11714,N_6091,N_728);
nand U11715 (N_11715,N_207,N_162);
or U11716 (N_11716,N_514,N_3944);
or U11717 (N_11717,N_5288,N_2418);
or U11718 (N_11718,N_3494,N_902);
and U11719 (N_11719,N_4949,N_1186);
and U11720 (N_11720,N_5638,N_5356);
and U11721 (N_11721,N_2604,N_4056);
nand U11722 (N_11722,N_5794,N_1664);
nor U11723 (N_11723,N_3120,N_3619);
or U11724 (N_11724,N_746,N_2900);
nor U11725 (N_11725,N_3037,N_3572);
nor U11726 (N_11726,N_3964,N_1892);
xor U11727 (N_11727,N_1150,N_770);
xnor U11728 (N_11728,N_3041,N_3142);
nor U11729 (N_11729,N_104,N_2864);
nand U11730 (N_11730,N_5990,N_1602);
nand U11731 (N_11731,N_3771,N_3769);
and U11732 (N_11732,N_1235,N_5001);
nor U11733 (N_11733,N_1472,N_2095);
or U11734 (N_11734,N_1994,N_5261);
nand U11735 (N_11735,N_1232,N_1345);
nand U11736 (N_11736,N_5361,N_5529);
nor U11737 (N_11737,N_4118,N_1343);
xnor U11738 (N_11738,N_1826,N_5297);
nor U11739 (N_11739,N_874,N_4477);
or U11740 (N_11740,N_2288,N_4273);
nand U11741 (N_11741,N_3009,N_1521);
nor U11742 (N_11742,N_1478,N_1582);
nand U11743 (N_11743,N_4097,N_1160);
and U11744 (N_11744,N_2776,N_935);
nor U11745 (N_11745,N_2125,N_5602);
nor U11746 (N_11746,N_4191,N_4556);
or U11747 (N_11747,N_3616,N_3478);
or U11748 (N_11748,N_3285,N_3583);
or U11749 (N_11749,N_5097,N_3175);
nand U11750 (N_11750,N_1143,N_4242);
or U11751 (N_11751,N_5940,N_2512);
or U11752 (N_11752,N_490,N_1156);
nand U11753 (N_11753,N_5712,N_3133);
or U11754 (N_11754,N_343,N_4949);
or U11755 (N_11755,N_4202,N_1530);
and U11756 (N_11756,N_5684,N_2687);
nand U11757 (N_11757,N_633,N_201);
and U11758 (N_11758,N_3058,N_4210);
nor U11759 (N_11759,N_709,N_909);
or U11760 (N_11760,N_2759,N_2030);
and U11761 (N_11761,N_709,N_228);
nand U11762 (N_11762,N_1580,N_4680);
nor U11763 (N_11763,N_5915,N_609);
nor U11764 (N_11764,N_3632,N_6006);
nand U11765 (N_11765,N_1653,N_5262);
and U11766 (N_11766,N_1498,N_2802);
and U11767 (N_11767,N_92,N_3608);
nand U11768 (N_11768,N_2936,N_4064);
nand U11769 (N_11769,N_5954,N_703);
nand U11770 (N_11770,N_2973,N_4277);
and U11771 (N_11771,N_2621,N_3323);
and U11772 (N_11772,N_3725,N_427);
nor U11773 (N_11773,N_2630,N_2595);
nor U11774 (N_11774,N_1083,N_3634);
nand U11775 (N_11775,N_4041,N_839);
or U11776 (N_11776,N_4326,N_2986);
or U11777 (N_11777,N_5162,N_4798);
or U11778 (N_11778,N_1930,N_1673);
and U11779 (N_11779,N_3180,N_5968);
nand U11780 (N_11780,N_4249,N_2939);
and U11781 (N_11781,N_1458,N_3954);
nor U11782 (N_11782,N_2137,N_102);
nand U11783 (N_11783,N_3261,N_1661);
nor U11784 (N_11784,N_3887,N_1828);
and U11785 (N_11785,N_3299,N_2613);
or U11786 (N_11786,N_5540,N_1359);
or U11787 (N_11787,N_511,N_3125);
nand U11788 (N_11788,N_4864,N_4956);
nor U11789 (N_11789,N_2020,N_5139);
or U11790 (N_11790,N_1345,N_2920);
nand U11791 (N_11791,N_4777,N_3855);
nand U11792 (N_11792,N_6086,N_4149);
nand U11793 (N_11793,N_2212,N_3614);
or U11794 (N_11794,N_1937,N_2901);
nor U11795 (N_11795,N_3956,N_3582);
and U11796 (N_11796,N_1594,N_2483);
nand U11797 (N_11797,N_3402,N_548);
and U11798 (N_11798,N_888,N_3726);
nor U11799 (N_11799,N_3152,N_5241);
or U11800 (N_11800,N_5017,N_4131);
nor U11801 (N_11801,N_3963,N_2227);
or U11802 (N_11802,N_832,N_2377);
nand U11803 (N_11803,N_382,N_5561);
and U11804 (N_11804,N_651,N_3991);
and U11805 (N_11805,N_5690,N_1365);
and U11806 (N_11806,N_3276,N_4034);
nand U11807 (N_11807,N_5297,N_2167);
nand U11808 (N_11808,N_4591,N_5012);
or U11809 (N_11809,N_2994,N_1190);
and U11810 (N_11810,N_5384,N_6245);
nor U11811 (N_11811,N_2314,N_563);
nor U11812 (N_11812,N_1436,N_6119);
or U11813 (N_11813,N_2550,N_79);
and U11814 (N_11814,N_896,N_5451);
xnor U11815 (N_11815,N_3686,N_5268);
xnor U11816 (N_11816,N_2104,N_421);
and U11817 (N_11817,N_3777,N_5061);
nor U11818 (N_11818,N_4504,N_5757);
nor U11819 (N_11819,N_1769,N_3985);
nand U11820 (N_11820,N_3259,N_3606);
xor U11821 (N_11821,N_2154,N_2187);
nand U11822 (N_11822,N_3686,N_3222);
nand U11823 (N_11823,N_4131,N_6118);
or U11824 (N_11824,N_6084,N_59);
nand U11825 (N_11825,N_5771,N_833);
nand U11826 (N_11826,N_2189,N_536);
nand U11827 (N_11827,N_3067,N_1186);
xor U11828 (N_11828,N_5962,N_2228);
or U11829 (N_11829,N_1615,N_2883);
and U11830 (N_11830,N_410,N_6231);
or U11831 (N_11831,N_1682,N_4901);
nand U11832 (N_11832,N_5937,N_37);
and U11833 (N_11833,N_3190,N_5153);
nor U11834 (N_11834,N_4732,N_3741);
or U11835 (N_11835,N_6087,N_5291);
and U11836 (N_11836,N_2679,N_2697);
nand U11837 (N_11837,N_547,N_6138);
nor U11838 (N_11838,N_3883,N_5563);
nor U11839 (N_11839,N_5702,N_2630);
nand U11840 (N_11840,N_2812,N_1599);
nor U11841 (N_11841,N_2233,N_4944);
or U11842 (N_11842,N_4361,N_2521);
nand U11843 (N_11843,N_1599,N_2600);
xnor U11844 (N_11844,N_2002,N_598);
nand U11845 (N_11845,N_4355,N_3806);
or U11846 (N_11846,N_3944,N_5251);
or U11847 (N_11847,N_1485,N_5691);
and U11848 (N_11848,N_4424,N_5742);
and U11849 (N_11849,N_3425,N_2104);
and U11850 (N_11850,N_1526,N_510);
xnor U11851 (N_11851,N_4126,N_3346);
or U11852 (N_11852,N_3292,N_4783);
and U11853 (N_11853,N_1023,N_5076);
xor U11854 (N_11854,N_1541,N_983);
or U11855 (N_11855,N_4465,N_2697);
and U11856 (N_11856,N_2441,N_4300);
and U11857 (N_11857,N_5328,N_4297);
or U11858 (N_11858,N_1076,N_4147);
or U11859 (N_11859,N_5561,N_1934);
nand U11860 (N_11860,N_6081,N_5995);
xnor U11861 (N_11861,N_4754,N_3707);
nand U11862 (N_11862,N_1552,N_3491);
or U11863 (N_11863,N_5884,N_5592);
and U11864 (N_11864,N_4254,N_4566);
and U11865 (N_11865,N_2335,N_1262);
xor U11866 (N_11866,N_5293,N_2321);
nor U11867 (N_11867,N_728,N_5727);
xor U11868 (N_11868,N_2240,N_2211);
and U11869 (N_11869,N_3127,N_4910);
nand U11870 (N_11870,N_2185,N_2053);
and U11871 (N_11871,N_4118,N_4142);
nor U11872 (N_11872,N_4901,N_2085);
nor U11873 (N_11873,N_4909,N_4996);
or U11874 (N_11874,N_5705,N_1434);
or U11875 (N_11875,N_3214,N_4373);
or U11876 (N_11876,N_1984,N_2923);
nand U11877 (N_11877,N_4524,N_4258);
nand U11878 (N_11878,N_3677,N_1892);
nor U11879 (N_11879,N_957,N_2239);
and U11880 (N_11880,N_6220,N_1753);
and U11881 (N_11881,N_4740,N_243);
and U11882 (N_11882,N_884,N_5929);
and U11883 (N_11883,N_5988,N_2233);
nor U11884 (N_11884,N_3628,N_543);
nor U11885 (N_11885,N_1838,N_1452);
nor U11886 (N_11886,N_3536,N_5661);
or U11887 (N_11887,N_5112,N_546);
nand U11888 (N_11888,N_5238,N_3469);
or U11889 (N_11889,N_3079,N_1807);
and U11890 (N_11890,N_3266,N_4406);
xor U11891 (N_11891,N_5610,N_1143);
nor U11892 (N_11892,N_1315,N_2801);
and U11893 (N_11893,N_3759,N_2839);
xor U11894 (N_11894,N_956,N_2086);
nand U11895 (N_11895,N_5511,N_2982);
nor U11896 (N_11896,N_3044,N_4468);
nor U11897 (N_11897,N_1126,N_6157);
and U11898 (N_11898,N_4065,N_2090);
xor U11899 (N_11899,N_2262,N_3894);
nor U11900 (N_11900,N_3490,N_3175);
nor U11901 (N_11901,N_275,N_2358);
and U11902 (N_11902,N_3743,N_95);
or U11903 (N_11903,N_2821,N_3842);
and U11904 (N_11904,N_2090,N_3012);
or U11905 (N_11905,N_5652,N_698);
and U11906 (N_11906,N_3606,N_3769);
or U11907 (N_11907,N_4386,N_176);
nor U11908 (N_11908,N_4643,N_3179);
nand U11909 (N_11909,N_296,N_1505);
nor U11910 (N_11910,N_1583,N_3932);
xnor U11911 (N_11911,N_6134,N_2536);
nand U11912 (N_11912,N_5889,N_1745);
or U11913 (N_11913,N_5947,N_1479);
and U11914 (N_11914,N_2024,N_1979);
nor U11915 (N_11915,N_5371,N_2812);
and U11916 (N_11916,N_1426,N_6098);
and U11917 (N_11917,N_3114,N_4953);
nor U11918 (N_11918,N_5965,N_1119);
nor U11919 (N_11919,N_1453,N_3244);
and U11920 (N_11920,N_3910,N_947);
and U11921 (N_11921,N_4857,N_426);
nor U11922 (N_11922,N_5161,N_2550);
and U11923 (N_11923,N_5140,N_3964);
or U11924 (N_11924,N_2870,N_3126);
nor U11925 (N_11925,N_402,N_5660);
nand U11926 (N_11926,N_4979,N_360);
nor U11927 (N_11927,N_2425,N_3359);
nor U11928 (N_11928,N_2765,N_5385);
nor U11929 (N_11929,N_2751,N_1208);
xnor U11930 (N_11930,N_1519,N_1426);
nand U11931 (N_11931,N_3972,N_4991);
nand U11932 (N_11932,N_5003,N_3644);
and U11933 (N_11933,N_34,N_2052);
nor U11934 (N_11934,N_2172,N_2703);
or U11935 (N_11935,N_4632,N_3356);
nor U11936 (N_11936,N_4557,N_4474);
and U11937 (N_11937,N_3993,N_6021);
nor U11938 (N_11938,N_878,N_4842);
and U11939 (N_11939,N_2437,N_1868);
nand U11940 (N_11940,N_651,N_5906);
and U11941 (N_11941,N_2447,N_1843);
nor U11942 (N_11942,N_438,N_4710);
or U11943 (N_11943,N_5452,N_331);
nor U11944 (N_11944,N_5189,N_6225);
and U11945 (N_11945,N_2152,N_146);
or U11946 (N_11946,N_367,N_2571);
and U11947 (N_11947,N_2915,N_5910);
or U11948 (N_11948,N_1790,N_5630);
xnor U11949 (N_11949,N_4680,N_695);
xor U11950 (N_11950,N_5622,N_1209);
and U11951 (N_11951,N_660,N_2131);
xnor U11952 (N_11952,N_1554,N_30);
and U11953 (N_11953,N_5131,N_4369);
and U11954 (N_11954,N_1734,N_128);
and U11955 (N_11955,N_5781,N_2899);
nand U11956 (N_11956,N_3471,N_4762);
and U11957 (N_11957,N_2656,N_6187);
nand U11958 (N_11958,N_3462,N_5258);
xnor U11959 (N_11959,N_1782,N_2781);
or U11960 (N_11960,N_2552,N_3891);
nand U11961 (N_11961,N_2321,N_1882);
and U11962 (N_11962,N_5347,N_6235);
or U11963 (N_11963,N_6172,N_2889);
nor U11964 (N_11964,N_1069,N_2927);
nor U11965 (N_11965,N_3876,N_4988);
and U11966 (N_11966,N_3064,N_1432);
nand U11967 (N_11967,N_216,N_1019);
or U11968 (N_11968,N_1552,N_5013);
nor U11969 (N_11969,N_2207,N_3180);
or U11970 (N_11970,N_3562,N_2888);
xnor U11971 (N_11971,N_2572,N_2155);
or U11972 (N_11972,N_5644,N_2418);
or U11973 (N_11973,N_3989,N_22);
and U11974 (N_11974,N_4570,N_1334);
nor U11975 (N_11975,N_55,N_5504);
and U11976 (N_11976,N_4618,N_1170);
and U11977 (N_11977,N_4686,N_5696);
nand U11978 (N_11978,N_4094,N_6195);
nand U11979 (N_11979,N_6079,N_2126);
or U11980 (N_11980,N_2515,N_1486);
xor U11981 (N_11981,N_1069,N_5068);
nor U11982 (N_11982,N_3966,N_512);
nor U11983 (N_11983,N_6140,N_303);
nor U11984 (N_11984,N_3720,N_892);
or U11985 (N_11985,N_6178,N_2097);
nand U11986 (N_11986,N_786,N_5980);
nand U11987 (N_11987,N_2969,N_4986);
nor U11988 (N_11988,N_1825,N_3831);
and U11989 (N_11989,N_1917,N_6207);
nand U11990 (N_11990,N_2722,N_403);
nor U11991 (N_11991,N_1978,N_5118);
and U11992 (N_11992,N_2881,N_4235);
nor U11993 (N_11993,N_4039,N_2971);
nor U11994 (N_11994,N_876,N_1029);
xnor U11995 (N_11995,N_2455,N_805);
or U11996 (N_11996,N_239,N_4358);
nor U11997 (N_11997,N_2062,N_1600);
or U11998 (N_11998,N_49,N_5419);
and U11999 (N_11999,N_2630,N_732);
and U12000 (N_12000,N_5778,N_561);
nand U12001 (N_12001,N_1542,N_4618);
nor U12002 (N_12002,N_167,N_3869);
xor U12003 (N_12003,N_5298,N_4913);
nor U12004 (N_12004,N_5625,N_3176);
nand U12005 (N_12005,N_4003,N_6097);
nor U12006 (N_12006,N_4088,N_2291);
and U12007 (N_12007,N_3706,N_3479);
nor U12008 (N_12008,N_3570,N_421);
and U12009 (N_12009,N_2341,N_647);
and U12010 (N_12010,N_1839,N_3123);
nand U12011 (N_12011,N_4177,N_5431);
nand U12012 (N_12012,N_4368,N_4778);
xor U12013 (N_12013,N_3938,N_6088);
nand U12014 (N_12014,N_5556,N_3431);
nor U12015 (N_12015,N_5907,N_2741);
and U12016 (N_12016,N_1035,N_5495);
nor U12017 (N_12017,N_5087,N_566);
xnor U12018 (N_12018,N_3872,N_3651);
or U12019 (N_12019,N_1456,N_2743);
nand U12020 (N_12020,N_2822,N_6088);
and U12021 (N_12021,N_470,N_1796);
xnor U12022 (N_12022,N_640,N_5755);
nand U12023 (N_12023,N_3675,N_4968);
or U12024 (N_12024,N_503,N_74);
and U12025 (N_12025,N_5340,N_132);
and U12026 (N_12026,N_2728,N_446);
and U12027 (N_12027,N_5764,N_5567);
nor U12028 (N_12028,N_4371,N_769);
nor U12029 (N_12029,N_4099,N_5402);
and U12030 (N_12030,N_866,N_1734);
nor U12031 (N_12031,N_870,N_5047);
xnor U12032 (N_12032,N_1350,N_4674);
or U12033 (N_12033,N_3831,N_3364);
nor U12034 (N_12034,N_4327,N_3318);
nand U12035 (N_12035,N_41,N_2146);
nand U12036 (N_12036,N_4488,N_4058);
nand U12037 (N_12037,N_2454,N_1446);
and U12038 (N_12038,N_4184,N_2679);
and U12039 (N_12039,N_3086,N_4118);
nor U12040 (N_12040,N_733,N_3843);
and U12041 (N_12041,N_3771,N_4947);
nand U12042 (N_12042,N_529,N_5101);
or U12043 (N_12043,N_883,N_5129);
nand U12044 (N_12044,N_2866,N_193);
or U12045 (N_12045,N_1591,N_5425);
nand U12046 (N_12046,N_4013,N_4504);
nor U12047 (N_12047,N_730,N_4200);
and U12048 (N_12048,N_4496,N_111);
nor U12049 (N_12049,N_4797,N_823);
nand U12050 (N_12050,N_219,N_5499);
nor U12051 (N_12051,N_4362,N_1222);
and U12052 (N_12052,N_5437,N_122);
nand U12053 (N_12053,N_5909,N_5409);
xor U12054 (N_12054,N_1983,N_1608);
nor U12055 (N_12055,N_1124,N_4487);
nor U12056 (N_12056,N_1890,N_4201);
nand U12057 (N_12057,N_4644,N_6223);
nor U12058 (N_12058,N_4323,N_572);
or U12059 (N_12059,N_6240,N_779);
nor U12060 (N_12060,N_4567,N_4946);
nand U12061 (N_12061,N_1520,N_118);
and U12062 (N_12062,N_5591,N_5651);
nor U12063 (N_12063,N_4378,N_323);
and U12064 (N_12064,N_362,N_1136);
or U12065 (N_12065,N_146,N_3034);
and U12066 (N_12066,N_5884,N_532);
or U12067 (N_12067,N_2573,N_3610);
nand U12068 (N_12068,N_4426,N_2178);
and U12069 (N_12069,N_1674,N_5625);
and U12070 (N_12070,N_4091,N_2000);
nor U12071 (N_12071,N_4731,N_5485);
or U12072 (N_12072,N_2172,N_736);
and U12073 (N_12073,N_5558,N_417);
nor U12074 (N_12074,N_255,N_4983);
nand U12075 (N_12075,N_2302,N_6106);
nor U12076 (N_12076,N_5561,N_2915);
nor U12077 (N_12077,N_2981,N_5790);
nor U12078 (N_12078,N_6062,N_1190);
nand U12079 (N_12079,N_2833,N_2388);
or U12080 (N_12080,N_4839,N_5599);
nor U12081 (N_12081,N_4780,N_2675);
nor U12082 (N_12082,N_4880,N_2085);
and U12083 (N_12083,N_592,N_3341);
nand U12084 (N_12084,N_180,N_5517);
or U12085 (N_12085,N_834,N_363);
xor U12086 (N_12086,N_2966,N_4905);
nor U12087 (N_12087,N_5978,N_2091);
nand U12088 (N_12088,N_2520,N_3373);
nand U12089 (N_12089,N_2642,N_4755);
and U12090 (N_12090,N_5035,N_6248);
xnor U12091 (N_12091,N_1891,N_2297);
nor U12092 (N_12092,N_900,N_2296);
nand U12093 (N_12093,N_6074,N_453);
and U12094 (N_12094,N_5557,N_1395);
xor U12095 (N_12095,N_3083,N_4310);
nor U12096 (N_12096,N_4538,N_43);
or U12097 (N_12097,N_2210,N_1701);
and U12098 (N_12098,N_949,N_3283);
nand U12099 (N_12099,N_681,N_3028);
xor U12100 (N_12100,N_3012,N_3768);
nor U12101 (N_12101,N_965,N_4520);
and U12102 (N_12102,N_4781,N_485);
nor U12103 (N_12103,N_3706,N_4543);
or U12104 (N_12104,N_5948,N_415);
or U12105 (N_12105,N_4904,N_5763);
nor U12106 (N_12106,N_341,N_1284);
or U12107 (N_12107,N_1506,N_3504);
nor U12108 (N_12108,N_2894,N_4261);
or U12109 (N_12109,N_3205,N_1844);
or U12110 (N_12110,N_2155,N_3453);
and U12111 (N_12111,N_188,N_3465);
xnor U12112 (N_12112,N_2558,N_6128);
nand U12113 (N_12113,N_2550,N_4930);
nor U12114 (N_12114,N_366,N_4817);
or U12115 (N_12115,N_1031,N_4928);
or U12116 (N_12116,N_2782,N_2071);
nand U12117 (N_12117,N_2632,N_5489);
and U12118 (N_12118,N_5602,N_4325);
nor U12119 (N_12119,N_3371,N_2210);
nand U12120 (N_12120,N_6057,N_3952);
or U12121 (N_12121,N_3092,N_199);
nand U12122 (N_12122,N_2809,N_2760);
nor U12123 (N_12123,N_413,N_2177);
nand U12124 (N_12124,N_2651,N_2800);
and U12125 (N_12125,N_2346,N_2691);
or U12126 (N_12126,N_1546,N_805);
nor U12127 (N_12127,N_1961,N_5076);
and U12128 (N_12128,N_6148,N_1997);
or U12129 (N_12129,N_4275,N_3103);
nor U12130 (N_12130,N_3087,N_3138);
and U12131 (N_12131,N_3693,N_4738);
xnor U12132 (N_12132,N_3213,N_4368);
and U12133 (N_12133,N_3155,N_1502);
and U12134 (N_12134,N_226,N_3994);
nand U12135 (N_12135,N_2112,N_293);
nor U12136 (N_12136,N_3347,N_6083);
nand U12137 (N_12137,N_5384,N_1429);
and U12138 (N_12138,N_4011,N_201);
xor U12139 (N_12139,N_1503,N_4647);
and U12140 (N_12140,N_1877,N_1350);
or U12141 (N_12141,N_6063,N_5643);
or U12142 (N_12142,N_801,N_5648);
or U12143 (N_12143,N_1796,N_1793);
or U12144 (N_12144,N_492,N_5899);
nor U12145 (N_12145,N_4751,N_2272);
nor U12146 (N_12146,N_4918,N_3717);
nand U12147 (N_12147,N_1437,N_3840);
nand U12148 (N_12148,N_2954,N_4470);
nor U12149 (N_12149,N_3942,N_3714);
or U12150 (N_12150,N_2577,N_4013);
nand U12151 (N_12151,N_3989,N_5756);
nor U12152 (N_12152,N_5959,N_2708);
or U12153 (N_12153,N_2118,N_2761);
nand U12154 (N_12154,N_1122,N_4075);
or U12155 (N_12155,N_1032,N_2927);
nand U12156 (N_12156,N_4624,N_4502);
or U12157 (N_12157,N_5097,N_5862);
nor U12158 (N_12158,N_5845,N_1492);
and U12159 (N_12159,N_2175,N_4016);
nor U12160 (N_12160,N_4023,N_2405);
and U12161 (N_12161,N_3594,N_1749);
or U12162 (N_12162,N_5922,N_2101);
and U12163 (N_12163,N_4011,N_5769);
and U12164 (N_12164,N_3123,N_4935);
nand U12165 (N_12165,N_724,N_3608);
or U12166 (N_12166,N_2043,N_2576);
or U12167 (N_12167,N_1751,N_4394);
nand U12168 (N_12168,N_4711,N_1987);
nand U12169 (N_12169,N_4660,N_2839);
nand U12170 (N_12170,N_5347,N_104);
nand U12171 (N_12171,N_156,N_1055);
nor U12172 (N_12172,N_4137,N_1950);
nand U12173 (N_12173,N_6103,N_6027);
nor U12174 (N_12174,N_1594,N_5780);
or U12175 (N_12175,N_3441,N_1931);
nor U12176 (N_12176,N_3149,N_4863);
nor U12177 (N_12177,N_4045,N_4681);
nand U12178 (N_12178,N_1697,N_5414);
or U12179 (N_12179,N_2621,N_1572);
and U12180 (N_12180,N_2382,N_2790);
or U12181 (N_12181,N_5133,N_1338);
xor U12182 (N_12182,N_1868,N_3590);
and U12183 (N_12183,N_2386,N_5572);
nand U12184 (N_12184,N_1363,N_5347);
or U12185 (N_12185,N_2055,N_42);
nand U12186 (N_12186,N_2644,N_2309);
or U12187 (N_12187,N_5010,N_3981);
xor U12188 (N_12188,N_2653,N_3269);
nor U12189 (N_12189,N_1872,N_1724);
and U12190 (N_12190,N_3877,N_4527);
or U12191 (N_12191,N_4735,N_5551);
nor U12192 (N_12192,N_5933,N_4532);
nor U12193 (N_12193,N_1178,N_3117);
nor U12194 (N_12194,N_6007,N_4138);
or U12195 (N_12195,N_1867,N_3949);
nor U12196 (N_12196,N_2625,N_1435);
xnor U12197 (N_12197,N_2831,N_2479);
and U12198 (N_12198,N_2496,N_5377);
nand U12199 (N_12199,N_1377,N_2456);
xnor U12200 (N_12200,N_3738,N_4612);
nand U12201 (N_12201,N_4997,N_5213);
and U12202 (N_12202,N_1088,N_560);
nand U12203 (N_12203,N_3800,N_668);
xnor U12204 (N_12204,N_3467,N_2649);
and U12205 (N_12205,N_6065,N_1053);
and U12206 (N_12206,N_4502,N_5594);
nor U12207 (N_12207,N_2324,N_3390);
nor U12208 (N_12208,N_1031,N_5446);
or U12209 (N_12209,N_1973,N_687);
nand U12210 (N_12210,N_4598,N_4033);
nor U12211 (N_12211,N_3074,N_709);
xor U12212 (N_12212,N_5742,N_1813);
nand U12213 (N_12213,N_5166,N_3736);
nand U12214 (N_12214,N_1137,N_1534);
and U12215 (N_12215,N_910,N_5061);
and U12216 (N_12216,N_440,N_3956);
nor U12217 (N_12217,N_1817,N_2903);
or U12218 (N_12218,N_4659,N_900);
nand U12219 (N_12219,N_3232,N_5502);
nor U12220 (N_12220,N_3929,N_2417);
nand U12221 (N_12221,N_915,N_2288);
and U12222 (N_12222,N_2887,N_5045);
nand U12223 (N_12223,N_5419,N_249);
or U12224 (N_12224,N_2630,N_5713);
and U12225 (N_12225,N_2233,N_6088);
and U12226 (N_12226,N_421,N_2144);
nor U12227 (N_12227,N_5104,N_3206);
and U12228 (N_12228,N_3789,N_4727);
nand U12229 (N_12229,N_2170,N_4450);
or U12230 (N_12230,N_4020,N_3034);
or U12231 (N_12231,N_5003,N_132);
and U12232 (N_12232,N_3565,N_4671);
nor U12233 (N_12233,N_4616,N_5388);
nand U12234 (N_12234,N_2358,N_2476);
nor U12235 (N_12235,N_5886,N_4705);
and U12236 (N_12236,N_5778,N_401);
xor U12237 (N_12237,N_1780,N_103);
or U12238 (N_12238,N_1938,N_1953);
nand U12239 (N_12239,N_4711,N_5026);
xor U12240 (N_12240,N_5594,N_5176);
nor U12241 (N_12241,N_285,N_839);
and U12242 (N_12242,N_5637,N_5294);
nor U12243 (N_12243,N_344,N_3577);
xor U12244 (N_12244,N_4228,N_3643);
xor U12245 (N_12245,N_141,N_44);
xnor U12246 (N_12246,N_1687,N_6169);
nor U12247 (N_12247,N_264,N_5028);
xor U12248 (N_12248,N_4210,N_650);
and U12249 (N_12249,N_4630,N_2151);
and U12250 (N_12250,N_3379,N_1604);
or U12251 (N_12251,N_2159,N_4534);
nand U12252 (N_12252,N_1228,N_4737);
or U12253 (N_12253,N_492,N_5384);
or U12254 (N_12254,N_603,N_2371);
or U12255 (N_12255,N_5904,N_5002);
nor U12256 (N_12256,N_4227,N_2318);
and U12257 (N_12257,N_6094,N_4383);
nand U12258 (N_12258,N_3661,N_4401);
or U12259 (N_12259,N_677,N_4491);
nor U12260 (N_12260,N_4549,N_4090);
and U12261 (N_12261,N_4703,N_5054);
and U12262 (N_12262,N_4599,N_25);
and U12263 (N_12263,N_1386,N_6162);
or U12264 (N_12264,N_720,N_49);
xor U12265 (N_12265,N_4654,N_4083);
nor U12266 (N_12266,N_3912,N_3977);
or U12267 (N_12267,N_1182,N_2919);
nand U12268 (N_12268,N_1998,N_5808);
or U12269 (N_12269,N_1197,N_1050);
xor U12270 (N_12270,N_1240,N_1982);
or U12271 (N_12271,N_2520,N_3861);
and U12272 (N_12272,N_1410,N_2151);
nor U12273 (N_12273,N_2271,N_2135);
or U12274 (N_12274,N_1681,N_1668);
nor U12275 (N_12275,N_6074,N_3550);
or U12276 (N_12276,N_2354,N_5611);
nand U12277 (N_12277,N_805,N_4342);
nand U12278 (N_12278,N_56,N_3062);
and U12279 (N_12279,N_5197,N_5156);
and U12280 (N_12280,N_163,N_1920);
xor U12281 (N_12281,N_697,N_5520);
nor U12282 (N_12282,N_1658,N_3549);
and U12283 (N_12283,N_5746,N_5437);
or U12284 (N_12284,N_5130,N_2976);
nor U12285 (N_12285,N_2939,N_2583);
and U12286 (N_12286,N_2057,N_3615);
and U12287 (N_12287,N_385,N_2649);
and U12288 (N_12288,N_3312,N_4387);
nand U12289 (N_12289,N_4713,N_3178);
nand U12290 (N_12290,N_3509,N_1260);
or U12291 (N_12291,N_3048,N_678);
nand U12292 (N_12292,N_1945,N_227);
or U12293 (N_12293,N_1449,N_3396);
and U12294 (N_12294,N_5095,N_5656);
and U12295 (N_12295,N_4131,N_1172);
nand U12296 (N_12296,N_1998,N_2000);
nor U12297 (N_12297,N_3325,N_4724);
nor U12298 (N_12298,N_3212,N_3934);
or U12299 (N_12299,N_508,N_1649);
or U12300 (N_12300,N_3655,N_1804);
and U12301 (N_12301,N_675,N_2036);
or U12302 (N_12302,N_5397,N_3348);
and U12303 (N_12303,N_2326,N_2640);
nand U12304 (N_12304,N_3538,N_3493);
nand U12305 (N_12305,N_1586,N_5110);
nor U12306 (N_12306,N_550,N_692);
nand U12307 (N_12307,N_5977,N_4156);
or U12308 (N_12308,N_4490,N_5558);
or U12309 (N_12309,N_1273,N_3934);
nand U12310 (N_12310,N_2847,N_5044);
and U12311 (N_12311,N_2586,N_3245);
nor U12312 (N_12312,N_2638,N_1031);
nand U12313 (N_12313,N_1422,N_1667);
and U12314 (N_12314,N_4037,N_5908);
or U12315 (N_12315,N_937,N_760);
nor U12316 (N_12316,N_7,N_5179);
and U12317 (N_12317,N_2079,N_411);
and U12318 (N_12318,N_4895,N_5111);
nor U12319 (N_12319,N_582,N_1389);
nand U12320 (N_12320,N_974,N_4483);
or U12321 (N_12321,N_3937,N_6107);
nor U12322 (N_12322,N_5942,N_2115);
nor U12323 (N_12323,N_2804,N_4693);
or U12324 (N_12324,N_3958,N_938);
nor U12325 (N_12325,N_3855,N_1668);
and U12326 (N_12326,N_4516,N_1921);
and U12327 (N_12327,N_3103,N_5551);
and U12328 (N_12328,N_6185,N_4903);
nor U12329 (N_12329,N_4767,N_5017);
or U12330 (N_12330,N_4434,N_3249);
or U12331 (N_12331,N_1251,N_5185);
or U12332 (N_12332,N_3002,N_5317);
nor U12333 (N_12333,N_2778,N_158);
nor U12334 (N_12334,N_4380,N_604);
nand U12335 (N_12335,N_1631,N_5730);
and U12336 (N_12336,N_875,N_1897);
nor U12337 (N_12337,N_3718,N_2053);
nand U12338 (N_12338,N_5121,N_3326);
nor U12339 (N_12339,N_3468,N_3459);
nand U12340 (N_12340,N_6247,N_3167);
xor U12341 (N_12341,N_4405,N_3606);
and U12342 (N_12342,N_4616,N_2145);
nand U12343 (N_12343,N_5686,N_2406);
or U12344 (N_12344,N_3818,N_53);
nor U12345 (N_12345,N_1664,N_3515);
nor U12346 (N_12346,N_2808,N_5277);
or U12347 (N_12347,N_354,N_2823);
nand U12348 (N_12348,N_1696,N_5102);
or U12349 (N_12349,N_5189,N_2325);
nor U12350 (N_12350,N_3340,N_3330);
or U12351 (N_12351,N_1613,N_4390);
nor U12352 (N_12352,N_4951,N_2776);
nand U12353 (N_12353,N_5223,N_772);
or U12354 (N_12354,N_4406,N_657);
and U12355 (N_12355,N_2594,N_5769);
nor U12356 (N_12356,N_365,N_2898);
or U12357 (N_12357,N_5123,N_3938);
or U12358 (N_12358,N_4533,N_5832);
or U12359 (N_12359,N_3276,N_365);
and U12360 (N_12360,N_3711,N_4513);
nor U12361 (N_12361,N_4221,N_3964);
nand U12362 (N_12362,N_5966,N_3018);
nor U12363 (N_12363,N_3557,N_5969);
xnor U12364 (N_12364,N_3523,N_2691);
nor U12365 (N_12365,N_3435,N_208);
nor U12366 (N_12366,N_3187,N_794);
xor U12367 (N_12367,N_889,N_4009);
nand U12368 (N_12368,N_3270,N_3982);
and U12369 (N_12369,N_5889,N_3453);
or U12370 (N_12370,N_4207,N_2654);
and U12371 (N_12371,N_717,N_4871);
or U12372 (N_12372,N_3262,N_5775);
nor U12373 (N_12373,N_3308,N_5531);
xor U12374 (N_12374,N_4449,N_2022);
xor U12375 (N_12375,N_773,N_881);
or U12376 (N_12376,N_5584,N_4741);
xor U12377 (N_12377,N_5309,N_5567);
nor U12378 (N_12378,N_5889,N_3371);
nand U12379 (N_12379,N_5472,N_6130);
or U12380 (N_12380,N_1722,N_1118);
nor U12381 (N_12381,N_1900,N_4561);
nor U12382 (N_12382,N_1332,N_58);
nor U12383 (N_12383,N_1861,N_2020);
or U12384 (N_12384,N_5665,N_5352);
and U12385 (N_12385,N_4003,N_4760);
nor U12386 (N_12386,N_430,N_5426);
xnor U12387 (N_12387,N_3250,N_2175);
nor U12388 (N_12388,N_6246,N_1713);
nand U12389 (N_12389,N_3165,N_5276);
and U12390 (N_12390,N_3156,N_6234);
nand U12391 (N_12391,N_2372,N_1593);
and U12392 (N_12392,N_3709,N_551);
nor U12393 (N_12393,N_1989,N_5507);
and U12394 (N_12394,N_4344,N_3665);
nand U12395 (N_12395,N_3737,N_1388);
or U12396 (N_12396,N_1662,N_373);
or U12397 (N_12397,N_1216,N_29);
or U12398 (N_12398,N_2025,N_2349);
nor U12399 (N_12399,N_4683,N_5320);
xor U12400 (N_12400,N_1231,N_3650);
nand U12401 (N_12401,N_2489,N_5225);
nor U12402 (N_12402,N_1937,N_55);
and U12403 (N_12403,N_3802,N_5531);
xor U12404 (N_12404,N_4238,N_2953);
xnor U12405 (N_12405,N_5453,N_950);
or U12406 (N_12406,N_4159,N_6061);
and U12407 (N_12407,N_3594,N_5732);
and U12408 (N_12408,N_1621,N_723);
and U12409 (N_12409,N_3653,N_1978);
nand U12410 (N_12410,N_4800,N_5306);
and U12411 (N_12411,N_5006,N_436);
nand U12412 (N_12412,N_5800,N_667);
or U12413 (N_12413,N_4618,N_1269);
or U12414 (N_12414,N_2322,N_972);
nor U12415 (N_12415,N_4578,N_312);
and U12416 (N_12416,N_4209,N_5771);
or U12417 (N_12417,N_3777,N_2071);
or U12418 (N_12418,N_3479,N_3564);
or U12419 (N_12419,N_3286,N_4299);
nor U12420 (N_12420,N_5045,N_20);
nand U12421 (N_12421,N_4079,N_2532);
and U12422 (N_12422,N_4337,N_452);
or U12423 (N_12423,N_4065,N_2784);
and U12424 (N_12424,N_1216,N_662);
and U12425 (N_12425,N_5047,N_4665);
nand U12426 (N_12426,N_6189,N_1413);
nand U12427 (N_12427,N_3609,N_3656);
nor U12428 (N_12428,N_4176,N_2003);
xnor U12429 (N_12429,N_110,N_757);
or U12430 (N_12430,N_5365,N_5706);
nor U12431 (N_12431,N_6144,N_5145);
or U12432 (N_12432,N_1220,N_4930);
xor U12433 (N_12433,N_3270,N_4359);
nor U12434 (N_12434,N_5075,N_5649);
or U12435 (N_12435,N_902,N_1579);
nand U12436 (N_12436,N_5457,N_5806);
and U12437 (N_12437,N_6084,N_1429);
or U12438 (N_12438,N_4665,N_5745);
nand U12439 (N_12439,N_2090,N_993);
nand U12440 (N_12440,N_2054,N_573);
and U12441 (N_12441,N_1101,N_4317);
and U12442 (N_12442,N_5540,N_5979);
or U12443 (N_12443,N_336,N_5573);
and U12444 (N_12444,N_1291,N_3291);
nand U12445 (N_12445,N_4018,N_5982);
nand U12446 (N_12446,N_4159,N_3785);
nand U12447 (N_12447,N_4227,N_1033);
nand U12448 (N_12448,N_1425,N_5924);
or U12449 (N_12449,N_641,N_1987);
and U12450 (N_12450,N_522,N_3137);
nand U12451 (N_12451,N_5433,N_5609);
xor U12452 (N_12452,N_2729,N_4668);
or U12453 (N_12453,N_4825,N_67);
and U12454 (N_12454,N_5998,N_2576);
xnor U12455 (N_12455,N_2579,N_6185);
nand U12456 (N_12456,N_4172,N_3895);
or U12457 (N_12457,N_3086,N_2061);
or U12458 (N_12458,N_1465,N_5942);
or U12459 (N_12459,N_686,N_398);
or U12460 (N_12460,N_5249,N_470);
nand U12461 (N_12461,N_5539,N_6185);
nand U12462 (N_12462,N_1217,N_5001);
nor U12463 (N_12463,N_5484,N_3907);
nand U12464 (N_12464,N_2414,N_2972);
or U12465 (N_12465,N_5969,N_493);
nand U12466 (N_12466,N_5863,N_4884);
nor U12467 (N_12467,N_1495,N_3837);
nor U12468 (N_12468,N_6006,N_4320);
or U12469 (N_12469,N_6005,N_4437);
or U12470 (N_12470,N_1909,N_1589);
and U12471 (N_12471,N_2456,N_3716);
nor U12472 (N_12472,N_2706,N_1637);
nand U12473 (N_12473,N_2371,N_5314);
nand U12474 (N_12474,N_4604,N_3940);
nor U12475 (N_12475,N_4483,N_1920);
nand U12476 (N_12476,N_1692,N_1354);
or U12477 (N_12477,N_5294,N_1081);
and U12478 (N_12478,N_4375,N_555);
nand U12479 (N_12479,N_5133,N_1550);
and U12480 (N_12480,N_6108,N_5162);
nor U12481 (N_12481,N_4370,N_4981);
nor U12482 (N_12482,N_3196,N_4307);
and U12483 (N_12483,N_582,N_2719);
or U12484 (N_12484,N_4745,N_3063);
nor U12485 (N_12485,N_4559,N_3274);
and U12486 (N_12486,N_3119,N_4161);
nor U12487 (N_12487,N_3727,N_5339);
xor U12488 (N_12488,N_1779,N_343);
nor U12489 (N_12489,N_895,N_2668);
xnor U12490 (N_12490,N_3083,N_1117);
nand U12491 (N_12491,N_4002,N_5018);
nand U12492 (N_12492,N_5460,N_1959);
and U12493 (N_12493,N_2576,N_1940);
or U12494 (N_12494,N_2207,N_3418);
and U12495 (N_12495,N_566,N_3239);
or U12496 (N_12496,N_2021,N_1956);
or U12497 (N_12497,N_3913,N_5976);
nand U12498 (N_12498,N_3884,N_2892);
and U12499 (N_12499,N_480,N_2301);
nor U12500 (N_12500,N_7439,N_9900);
or U12501 (N_12501,N_11700,N_8733);
nor U12502 (N_12502,N_12397,N_11007);
and U12503 (N_12503,N_6453,N_10816);
nor U12504 (N_12504,N_10727,N_10643);
and U12505 (N_12505,N_7717,N_9394);
nor U12506 (N_12506,N_8009,N_9163);
nand U12507 (N_12507,N_9144,N_8753);
and U12508 (N_12508,N_7932,N_9807);
or U12509 (N_12509,N_9249,N_12351);
nor U12510 (N_12510,N_10887,N_10258);
or U12511 (N_12511,N_10626,N_7804);
or U12512 (N_12512,N_11555,N_8583);
nand U12513 (N_12513,N_11520,N_8664);
or U12514 (N_12514,N_6285,N_8377);
and U12515 (N_12515,N_6553,N_9878);
nand U12516 (N_12516,N_8053,N_6624);
and U12517 (N_12517,N_11536,N_8737);
and U12518 (N_12518,N_6944,N_9182);
and U12519 (N_12519,N_7003,N_6673);
and U12520 (N_12520,N_8078,N_7939);
and U12521 (N_12521,N_6578,N_10325);
and U12522 (N_12522,N_6813,N_9419);
nand U12523 (N_12523,N_9872,N_6282);
xnor U12524 (N_12524,N_9861,N_11634);
nor U12525 (N_12525,N_11599,N_6460);
and U12526 (N_12526,N_6381,N_11571);
and U12527 (N_12527,N_8002,N_6412);
nor U12528 (N_12528,N_6716,N_9921);
nor U12529 (N_12529,N_9659,N_10430);
nand U12530 (N_12530,N_12042,N_8092);
nor U12531 (N_12531,N_11426,N_8613);
or U12532 (N_12532,N_8847,N_8765);
and U12533 (N_12533,N_8924,N_12186);
or U12534 (N_12534,N_9162,N_7445);
or U12535 (N_12535,N_10227,N_9142);
nor U12536 (N_12536,N_11296,N_8005);
nor U12537 (N_12537,N_9964,N_10685);
or U12538 (N_12538,N_6949,N_7603);
or U12539 (N_12539,N_8418,N_6939);
nand U12540 (N_12540,N_6845,N_7409);
and U12541 (N_12541,N_7336,N_10590);
nor U12542 (N_12542,N_9539,N_10424);
and U12543 (N_12543,N_8342,N_12079);
xor U12544 (N_12544,N_7375,N_11318);
nand U12545 (N_12545,N_8080,N_11613);
and U12546 (N_12546,N_10295,N_11250);
and U12547 (N_12547,N_8543,N_10157);
or U12548 (N_12548,N_8244,N_10622);
nor U12549 (N_12549,N_6514,N_9828);
nand U12550 (N_12550,N_7056,N_7590);
or U12551 (N_12551,N_8191,N_7339);
nor U12552 (N_12552,N_8360,N_11858);
or U12553 (N_12553,N_10608,N_10870);
nor U12554 (N_12554,N_8718,N_9343);
and U12555 (N_12555,N_7167,N_12404);
and U12556 (N_12556,N_8778,N_11937);
or U12557 (N_12557,N_10237,N_7547);
or U12558 (N_12558,N_9688,N_8468);
and U12559 (N_12559,N_7184,N_11800);
nor U12560 (N_12560,N_8103,N_9228);
nor U12561 (N_12561,N_10079,N_9545);
nor U12562 (N_12562,N_6958,N_9436);
and U12563 (N_12563,N_6953,N_11444);
or U12564 (N_12564,N_9440,N_11224);
nor U12565 (N_12565,N_11397,N_11080);
and U12566 (N_12566,N_6929,N_10603);
nand U12567 (N_12567,N_9957,N_6942);
nor U12568 (N_12568,N_8795,N_6456);
nand U12569 (N_12569,N_6569,N_7933);
or U12570 (N_12570,N_12483,N_6422);
nand U12571 (N_12571,N_7483,N_7566);
nand U12572 (N_12572,N_11311,N_12032);
or U12573 (N_12573,N_8365,N_11704);
nor U12574 (N_12574,N_9227,N_9225);
nor U12575 (N_12575,N_11871,N_7032);
nand U12576 (N_12576,N_7641,N_7394);
or U12577 (N_12577,N_10060,N_8238);
and U12578 (N_12578,N_12211,N_9752);
nand U12579 (N_12579,N_10264,N_10156);
xor U12580 (N_12580,N_6516,N_7903);
nor U12581 (N_12581,N_6725,N_9986);
or U12582 (N_12582,N_11717,N_11506);
or U12583 (N_12583,N_9180,N_11764);
xor U12584 (N_12584,N_6973,N_9973);
and U12585 (N_12585,N_10007,N_6336);
and U12586 (N_12586,N_11331,N_9628);
nor U12587 (N_12587,N_6964,N_7661);
nand U12588 (N_12588,N_9818,N_9393);
and U12589 (N_12589,N_12461,N_10881);
and U12590 (N_12590,N_10330,N_7260);
and U12591 (N_12591,N_12136,N_11026);
or U12592 (N_12592,N_12279,N_10143);
nand U12593 (N_12593,N_9617,N_7769);
or U12594 (N_12594,N_8735,N_7606);
or U12595 (N_12595,N_9885,N_11779);
and U12596 (N_12596,N_9522,N_7503);
nand U12597 (N_12597,N_8391,N_11676);
nand U12598 (N_12598,N_8046,N_7005);
and U12599 (N_12599,N_10843,N_8650);
and U12600 (N_12600,N_10538,N_7656);
nor U12601 (N_12601,N_11649,N_11344);
xor U12602 (N_12602,N_11616,N_6656);
xnor U12603 (N_12603,N_11057,N_11452);
or U12604 (N_12604,N_6357,N_7529);
nor U12605 (N_12605,N_9363,N_9198);
and U12606 (N_12606,N_7887,N_9199);
xnor U12607 (N_12607,N_11125,N_12329);
nor U12608 (N_12608,N_8827,N_7436);
xnor U12609 (N_12609,N_9210,N_6909);
nor U12610 (N_12610,N_9262,N_10819);
and U12611 (N_12611,N_6831,N_8123);
nor U12612 (N_12612,N_9757,N_7826);
or U12613 (N_12613,N_6626,N_10838);
nand U12614 (N_12614,N_10188,N_7113);
and U12615 (N_12615,N_9884,N_12242);
nand U12616 (N_12616,N_7139,N_8281);
or U12617 (N_12617,N_9481,N_9640);
xor U12618 (N_12618,N_10630,N_10797);
or U12619 (N_12619,N_8370,N_12400);
or U12620 (N_12620,N_6521,N_11580);
xor U12621 (N_12621,N_7466,N_9226);
nand U12622 (N_12622,N_11809,N_6284);
nand U12623 (N_12623,N_8974,N_11041);
nor U12624 (N_12624,N_7240,N_11622);
nand U12625 (N_12625,N_9068,N_8136);
and U12626 (N_12626,N_8663,N_8399);
and U12627 (N_12627,N_9511,N_10020);
xor U12628 (N_12628,N_6264,N_10768);
nor U12629 (N_12629,N_10491,N_10922);
nor U12630 (N_12630,N_8781,N_8866);
nor U12631 (N_12631,N_9204,N_11639);
nor U12632 (N_12632,N_11354,N_8705);
nor U12633 (N_12633,N_12266,N_7512);
nor U12634 (N_12634,N_12278,N_11647);
nor U12635 (N_12635,N_9887,N_6443);
or U12636 (N_12636,N_10397,N_8100);
or U12637 (N_12637,N_7971,N_12235);
nand U12638 (N_12638,N_6853,N_10914);
nor U12639 (N_12639,N_11200,N_10339);
nand U12640 (N_12640,N_7385,N_11998);
nand U12641 (N_12641,N_7674,N_12244);
nand U12642 (N_12642,N_9954,N_7435);
nor U12643 (N_12643,N_11699,N_7233);
xnor U12644 (N_12644,N_7210,N_12363);
and U12645 (N_12645,N_7276,N_6948);
nor U12646 (N_12646,N_9220,N_11440);
nor U12647 (N_12647,N_8511,N_9050);
nor U12648 (N_12648,N_7713,N_10578);
and U12649 (N_12649,N_12233,N_6997);
nand U12650 (N_12650,N_7083,N_10971);
nand U12651 (N_12651,N_10288,N_7346);
and U12652 (N_12652,N_9085,N_8873);
nand U12653 (N_12653,N_11011,N_11606);
and U12654 (N_12654,N_7657,N_8722);
nand U12655 (N_12655,N_8751,N_10271);
nand U12656 (N_12656,N_8324,N_11417);
and U12657 (N_12657,N_10220,N_7076);
or U12658 (N_12658,N_11798,N_10885);
nand U12659 (N_12659,N_6532,N_6549);
and U12660 (N_12660,N_11890,N_11640);
or U12661 (N_12661,N_11027,N_6685);
nor U12662 (N_12662,N_10111,N_10400);
or U12663 (N_12663,N_7371,N_6846);
nor U12664 (N_12664,N_9264,N_10828);
nand U12665 (N_12665,N_10531,N_11975);
or U12666 (N_12666,N_10080,N_11177);
nand U12667 (N_12667,N_8604,N_12046);
xnor U12668 (N_12668,N_10522,N_8265);
nor U12669 (N_12669,N_7685,N_10806);
nand U12670 (N_12670,N_8150,N_10070);
nor U12671 (N_12671,N_11138,N_7935);
or U12672 (N_12672,N_11892,N_11349);
nand U12673 (N_12673,N_9505,N_6375);
and U12674 (N_12674,N_7373,N_9924);
nand U12675 (N_12675,N_8079,N_8177);
xor U12676 (N_12676,N_11005,N_6747);
nand U12677 (N_12677,N_8233,N_7227);
nand U12678 (N_12678,N_11235,N_11448);
and U12679 (N_12679,N_9766,N_6826);
nor U12680 (N_12680,N_10517,N_7490);
or U12681 (N_12681,N_7464,N_10337);
and U12682 (N_12682,N_8285,N_8372);
or U12683 (N_12683,N_9896,N_7636);
and U12684 (N_12684,N_9983,N_9045);
nor U12685 (N_12685,N_10557,N_11399);
nor U12686 (N_12686,N_9477,N_9214);
and U12687 (N_12687,N_6695,N_9493);
nor U12688 (N_12688,N_11329,N_9217);
nand U12689 (N_12689,N_6650,N_10159);
and U12690 (N_12690,N_12255,N_8585);
and U12691 (N_12691,N_7515,N_6991);
nand U12692 (N_12692,N_10285,N_12298);
and U12693 (N_12693,N_9408,N_11566);
nand U12694 (N_12694,N_7881,N_12445);
and U12695 (N_12695,N_10406,N_7427);
nor U12696 (N_12696,N_10435,N_9356);
xor U12697 (N_12697,N_8498,N_9132);
or U12698 (N_12698,N_7992,N_7431);
nand U12699 (N_12699,N_10734,N_6303);
nand U12700 (N_12700,N_10647,N_12470);
xor U12701 (N_12701,N_9403,N_7649);
or U12702 (N_12702,N_12037,N_11462);
and U12703 (N_12703,N_9750,N_10026);
and U12704 (N_12704,N_7397,N_10107);
or U12705 (N_12705,N_11186,N_12360);
nand U12706 (N_12706,N_7170,N_9920);
xor U12707 (N_12707,N_6374,N_8895);
nand U12708 (N_12708,N_11960,N_7715);
nand U12709 (N_12709,N_11554,N_12127);
nor U12710 (N_12710,N_6993,N_9473);
nand U12711 (N_12711,N_7390,N_12081);
and U12712 (N_12712,N_11419,N_9251);
nand U12713 (N_12713,N_6817,N_12054);
or U12714 (N_12714,N_10165,N_10327);
or U12715 (N_12715,N_10729,N_7075);
nand U12716 (N_12716,N_10864,N_6433);
or U12717 (N_12717,N_8772,N_7671);
and U12718 (N_12718,N_8215,N_8368);
and U12719 (N_12719,N_11865,N_7964);
nor U12720 (N_12720,N_8149,N_7403);
or U12721 (N_12721,N_7865,N_8470);
nand U12722 (N_12722,N_9839,N_10112);
or U12723 (N_12723,N_8556,N_8193);
and U12724 (N_12724,N_7960,N_7745);
xnor U12725 (N_12725,N_7965,N_9443);
or U12726 (N_12726,N_10284,N_6508);
nor U12727 (N_12727,N_10292,N_9178);
nor U12728 (N_12728,N_9177,N_10758);
nand U12729 (N_12729,N_12172,N_6529);
xnor U12730 (N_12730,N_6862,N_9348);
or U12731 (N_12731,N_10945,N_6880);
nand U12732 (N_12732,N_7013,N_7355);
and U12733 (N_12733,N_8589,N_11753);
nor U12734 (N_12734,N_6296,N_8862);
and U12735 (N_12735,N_9232,N_9529);
or U12736 (N_12736,N_11909,N_9751);
nor U12737 (N_12737,N_6739,N_9292);
and U12738 (N_12738,N_7369,N_12464);
or U12739 (N_12739,N_10166,N_6393);
nand U12740 (N_12740,N_11662,N_8623);
xnor U12741 (N_12741,N_10584,N_7559);
and U12742 (N_12742,N_11423,N_9923);
and U12743 (N_12743,N_10038,N_10323);
nand U12744 (N_12744,N_11014,N_7222);
and U12745 (N_12745,N_6490,N_8967);
xor U12746 (N_12746,N_8709,N_7738);
nand U12747 (N_12747,N_7300,N_7796);
and U12748 (N_12748,N_8657,N_10674);
and U12749 (N_12749,N_11076,N_7533);
and U12750 (N_12750,N_11651,N_10209);
nor U12751 (N_12751,N_8118,N_11724);
or U12752 (N_12752,N_9653,N_11213);
or U12753 (N_12753,N_10103,N_8447);
xor U12754 (N_12754,N_10167,N_9349);
nand U12755 (N_12755,N_6506,N_9479);
and U12756 (N_12756,N_7918,N_12080);
nand U12757 (N_12757,N_9095,N_6451);
or U12758 (N_12758,N_8959,N_11525);
nor U12759 (N_12759,N_9320,N_9535);
and U12760 (N_12760,N_9655,N_11316);
nand U12761 (N_12761,N_7228,N_10089);
and U12762 (N_12762,N_7395,N_11194);
nand U12763 (N_12763,N_8581,N_11490);
or U12764 (N_12764,N_7502,N_9078);
xnor U12765 (N_12765,N_8813,N_7760);
or U12766 (N_12766,N_9105,N_11010);
or U12767 (N_12767,N_9079,N_7597);
xor U12768 (N_12768,N_8534,N_8647);
nand U12769 (N_12769,N_9362,N_9851);
xnor U12770 (N_12770,N_11075,N_10207);
and U12771 (N_12771,N_6629,N_8653);
and U12772 (N_12772,N_12379,N_7066);
nand U12773 (N_12773,N_8550,N_11114);
nor U12774 (N_12774,N_9347,N_6671);
or U12775 (N_12775,N_8205,N_11726);
nor U12776 (N_12776,N_6388,N_7521);
xor U12777 (N_12777,N_6930,N_7873);
nor U12778 (N_12778,N_11617,N_10123);
or U12779 (N_12779,N_11196,N_8077);
nor U12780 (N_12780,N_10027,N_11680);
or U12781 (N_12781,N_7697,N_10996);
or U12782 (N_12782,N_10579,N_11404);
nand U12783 (N_12783,N_11152,N_7430);
nor U12784 (N_12784,N_6888,N_10074);
and U12785 (N_12785,N_8806,N_10558);
and U12786 (N_12786,N_11987,N_9502);
nor U12787 (N_12787,N_11124,N_8274);
nor U12788 (N_12788,N_6358,N_9006);
and U12789 (N_12789,N_8108,N_9294);
and U12790 (N_12790,N_9538,N_8738);
and U12791 (N_12791,N_9612,N_6734);
or U12792 (N_12792,N_6628,N_7095);
xor U12793 (N_12793,N_8247,N_11363);
nand U12794 (N_12794,N_10704,N_7362);
and U12795 (N_12795,N_9181,N_7572);
nand U12796 (N_12796,N_8923,N_6705);
and U12797 (N_12797,N_10360,N_11908);
nand U12798 (N_12798,N_11790,N_11782);
xnor U12799 (N_12799,N_12467,N_9597);
nor U12800 (N_12800,N_6766,N_10487);
nor U12801 (N_12801,N_7710,N_9483);
and U12802 (N_12802,N_7561,N_8702);
and U12803 (N_12803,N_9243,N_8054);
or U12804 (N_12804,N_7585,N_7911);
or U12805 (N_12805,N_12371,N_10463);
nor U12806 (N_12806,N_12016,N_6584);
nand U12807 (N_12807,N_10662,N_10917);
and U12808 (N_12808,N_6694,N_11916);
and U12809 (N_12809,N_9241,N_8460);
nand U12810 (N_12810,N_12044,N_7347);
or U12811 (N_12811,N_9763,N_6919);
xor U12812 (N_12812,N_7312,N_7744);
nor U12813 (N_12813,N_10155,N_8344);
xnor U12814 (N_12814,N_8970,N_7983);
nand U12815 (N_12815,N_10983,N_9387);
nand U12816 (N_12816,N_7716,N_11643);
nor U12817 (N_12817,N_8485,N_11070);
nand U12818 (N_12818,N_11523,N_7562);
nand U12819 (N_12819,N_12189,N_12203);
nor U12820 (N_12820,N_7757,N_8367);
and U12821 (N_12821,N_8710,N_6679);
nor U12822 (N_12822,N_11336,N_11965);
xor U12823 (N_12823,N_8278,N_11961);
and U12824 (N_12824,N_11888,N_11876);
and U12825 (N_12825,N_10287,N_8266);
nand U12826 (N_12826,N_10222,N_8075);
nand U12827 (N_12827,N_8170,N_10342);
and U12828 (N_12828,N_9916,N_9350);
nor U12829 (N_12829,N_9879,N_7705);
and U12830 (N_12830,N_6833,N_11775);
and U12831 (N_12831,N_6408,N_10733);
nor U12832 (N_12832,N_6921,N_8541);
xnor U12833 (N_12833,N_9675,N_6339);
nand U12834 (N_12834,N_6652,N_9175);
nand U12835 (N_12835,N_12344,N_6789);
nand U12836 (N_12836,N_7631,N_7322);
and U12837 (N_12837,N_11646,N_10378);
and U12838 (N_12838,N_10450,N_8384);
nand U12839 (N_12839,N_7247,N_8106);
or U12840 (N_12840,N_9461,N_10989);
nor U12841 (N_12841,N_9600,N_12246);
nand U12842 (N_12842,N_11577,N_10362);
and U12843 (N_12843,N_8938,N_6327);
nor U12844 (N_12844,N_9867,N_10582);
nand U12845 (N_12845,N_8320,N_8198);
or U12846 (N_12846,N_6421,N_10318);
nand U12847 (N_12847,N_7213,N_10289);
and U12848 (N_12848,N_7135,N_8909);
xor U12849 (N_12849,N_8067,N_7831);
nor U12850 (N_12850,N_7401,N_11439);
and U12851 (N_12851,N_7297,N_7955);
or U12852 (N_12852,N_8893,N_11656);
or U12853 (N_12853,N_6276,N_11247);
nor U12854 (N_12854,N_10030,N_7237);
and U12855 (N_12855,N_8831,N_8685);
and U12856 (N_12856,N_7140,N_11414);
xnor U12857 (N_12857,N_12366,N_12380);
and U12858 (N_12858,N_12144,N_10499);
xnor U12859 (N_12859,N_8417,N_11037);
and U12860 (N_12860,N_6602,N_6825);
or U12861 (N_12861,N_9938,N_12070);
xor U12862 (N_12862,N_11697,N_10306);
nand U12863 (N_12863,N_10479,N_8502);
or U12864 (N_12864,N_8039,N_6479);
or U12865 (N_12865,N_12124,N_9007);
and U12866 (N_12866,N_9882,N_7316);
or U12867 (N_12867,N_7341,N_10416);
nand U12868 (N_12868,N_11610,N_11441);
xor U12869 (N_12869,N_10871,N_7772);
nand U12870 (N_12870,N_9455,N_8514);
nand U12871 (N_12871,N_6420,N_6261);
xor U12872 (N_12872,N_12125,N_6379);
nor U12873 (N_12873,N_7894,N_8984);
and U12874 (N_12874,N_6588,N_11474);
nand U12875 (N_12875,N_9824,N_11304);
nor U12876 (N_12876,N_9713,N_7141);
xnor U12877 (N_12877,N_8848,N_7456);
or U12878 (N_12878,N_9367,N_7406);
nor U12879 (N_12879,N_12139,N_8995);
or U12880 (N_12880,N_7354,N_8121);
and U12881 (N_12881,N_8293,N_7775);
or U12882 (N_12882,N_7532,N_6523);
nand U12883 (N_12883,N_8254,N_8257);
nor U12884 (N_12884,N_10006,N_11216);
or U12885 (N_12885,N_7156,N_8260);
nor U12886 (N_12886,N_6938,N_10540);
nand U12887 (N_12887,N_12448,N_11003);
xnor U12888 (N_12888,N_11768,N_12430);
and U12889 (N_12889,N_6927,N_9153);
and U12890 (N_12890,N_10617,N_7499);
nor U12891 (N_12891,N_11154,N_11645);
and U12892 (N_12892,N_6649,N_8981);
nand U12893 (N_12893,N_12480,N_12085);
and U12894 (N_12894,N_10057,N_7432);
xnor U12895 (N_12895,N_11083,N_8522);
nand U12896 (N_12896,N_7012,N_7851);
xor U12897 (N_12897,N_8476,N_11334);
nor U12898 (N_12898,N_11155,N_8048);
and U12899 (N_12899,N_9891,N_7845);
nor U12900 (N_12900,N_8698,N_8815);
or U12901 (N_12901,N_8646,N_12334);
and U12902 (N_12902,N_12185,N_9598);
and U12903 (N_12903,N_12253,N_7351);
nor U12904 (N_12904,N_6328,N_7175);
nor U12905 (N_12905,N_10134,N_7880);
nor U12906 (N_12906,N_7179,N_7506);
xnor U12907 (N_12907,N_8206,N_11945);
nand U12908 (N_12908,N_12208,N_8746);
and U12909 (N_12909,N_6400,N_12022);
or U12910 (N_12910,N_7197,N_9696);
nand U12911 (N_12911,N_8307,N_8779);
or U12912 (N_12912,N_12270,N_9985);
or U12913 (N_12913,N_9042,N_9100);
nor U12914 (N_12914,N_9892,N_8347);
nor U12915 (N_12915,N_9936,N_9028);
or U12916 (N_12916,N_6860,N_6287);
nor U12917 (N_12917,N_10997,N_7137);
nand U12918 (N_12918,N_10908,N_11741);
nor U12919 (N_12919,N_12038,N_6267);
nor U12920 (N_12920,N_6802,N_9491);
and U12921 (N_12921,N_7206,N_11882);
or U12922 (N_12922,N_9772,N_6768);
and U12923 (N_12923,N_9097,N_11207);
or U12924 (N_12924,N_11302,N_9253);
nor U12925 (N_12925,N_9681,N_10095);
nor U12926 (N_12926,N_7062,N_7613);
nand U12927 (N_12927,N_10699,N_12090);
nor U12928 (N_12928,N_9883,N_12014);
xnor U12929 (N_12929,N_10328,N_8013);
nand U12930 (N_12930,N_8015,N_11923);
or U12931 (N_12931,N_11491,N_12294);
and U12932 (N_12932,N_6913,N_10176);
nor U12933 (N_12933,N_6666,N_8394);
or U12934 (N_12934,N_9301,N_10099);
xnor U12935 (N_12935,N_8436,N_11552);
or U12936 (N_12936,N_10200,N_7163);
and U12937 (N_12937,N_9312,N_10692);
nand U12938 (N_12938,N_8505,N_8532);
or U12939 (N_12939,N_7734,N_10605);
nand U12940 (N_12940,N_7361,N_8072);
or U12941 (N_12941,N_8579,N_6410);
or U12942 (N_12942,N_8849,N_10902);
and U12943 (N_12943,N_10927,N_9278);
or U12944 (N_12944,N_8699,N_10709);
nand U12945 (N_12945,N_10154,N_8410);
xor U12946 (N_12946,N_11055,N_11305);
nand U12947 (N_12947,N_8922,N_8566);
nor U12948 (N_12948,N_7474,N_11201);
nand U12949 (N_12949,N_7189,N_10407);
xor U12950 (N_12950,N_11060,N_7616);
or U12951 (N_12951,N_6906,N_9293);
and U12952 (N_12952,N_10869,N_8161);
nand U12953 (N_12953,N_6442,N_11557);
or U12954 (N_12954,N_11339,N_7096);
nand U12955 (N_12955,N_9252,N_11562);
nand U12956 (N_12956,N_10347,N_7150);
nor U12957 (N_12957,N_8886,N_10610);
xnor U12958 (N_12958,N_11377,N_9478);
xor U12959 (N_12959,N_9183,N_6533);
or U12960 (N_12960,N_9322,N_8572);
nor U12961 (N_12961,N_6554,N_8830);
and U12962 (N_12962,N_12147,N_8715);
and U12963 (N_12963,N_11256,N_6801);
nand U12964 (N_12964,N_10461,N_10068);
or U12965 (N_12965,N_7011,N_8567);
xnor U12966 (N_12966,N_7450,N_8478);
nand U12967 (N_12967,N_6297,N_10206);
nor U12968 (N_12968,N_6617,N_7584);
nor U12969 (N_12969,N_8258,N_11832);
nor U12970 (N_12970,N_7626,N_7223);
or U12971 (N_12971,N_7821,N_9092);
and U12972 (N_12972,N_9521,N_7281);
xor U12973 (N_12973,N_12015,N_7967);
nor U12974 (N_12974,N_10369,N_6990);
or U12975 (N_12975,N_12062,N_8226);
nor U12976 (N_12976,N_11298,N_8091);
and U12977 (N_12977,N_10304,N_7234);
or U12978 (N_12978,N_8162,N_7882);
or U12979 (N_12979,N_10067,N_11150);
nand U12980 (N_12980,N_8620,N_11980);
nand U12981 (N_12981,N_10262,N_8188);
or U12982 (N_12982,N_7670,N_6722);
nand U12983 (N_12983,N_7017,N_6823);
and U12984 (N_12984,N_7089,N_8289);
nor U12985 (N_12985,N_9158,N_7743);
nand U12986 (N_12986,N_11460,N_10760);
nor U12987 (N_12987,N_11817,N_7266);
nor U12988 (N_12988,N_8340,N_11178);
nor U12989 (N_12989,N_7041,N_11099);
nor U12990 (N_12990,N_6968,N_9282);
nor U12991 (N_12991,N_9031,N_9447);
or U12992 (N_12992,N_9325,N_11219);
nand U12993 (N_12993,N_8277,N_12035);
and U12994 (N_12994,N_10319,N_12076);
and U12995 (N_12995,N_9632,N_6385);
nand U12996 (N_12996,N_6555,N_10373);
or U12997 (N_12997,N_7500,N_7752);
nand U12998 (N_12998,N_9704,N_8661);
xnor U12999 (N_12999,N_9578,N_10351);
and U13000 (N_13000,N_11572,N_8402);
and U13001 (N_13001,N_10629,N_7165);
nand U13002 (N_13002,N_10822,N_7687);
or U13003 (N_13003,N_6797,N_9984);
nand U13004 (N_13004,N_11725,N_7632);
and U13005 (N_13005,N_11664,N_10075);
nor U13006 (N_13006,N_9421,N_10833);
or U13007 (N_13007,N_9471,N_12063);
or U13008 (N_13008,N_10942,N_7271);
nor U13009 (N_13009,N_8382,N_10554);
nor U13010 (N_13010,N_8444,N_7193);
nand U13011 (N_13011,N_11660,N_11245);
or U13012 (N_13012,N_12342,N_7437);
xnor U13013 (N_13013,N_8056,N_9074);
nor U13014 (N_13014,N_10210,N_12365);
xor U13015 (N_13015,N_9556,N_8428);
or U13016 (N_13016,N_6609,N_12433);
and U13017 (N_13017,N_9561,N_11333);
and U13018 (N_13018,N_10723,N_10928);
nand U13019 (N_13019,N_10649,N_6605);
nand U13020 (N_13020,N_8796,N_12327);
nor U13021 (N_13021,N_10310,N_10639);
or U13022 (N_13022,N_9852,N_11291);
xnor U13023 (N_13023,N_10710,N_7134);
and U13024 (N_13024,N_11018,N_8336);
nor U13025 (N_13025,N_9592,N_7100);
or U13026 (N_13026,N_9275,N_7869);
and U13027 (N_13027,N_6314,N_10523);
or U13028 (N_13028,N_9370,N_8179);
and U13029 (N_13029,N_8596,N_7055);
nand U13030 (N_13030,N_8898,N_11432);
or U13031 (N_13031,N_10794,N_9943);
xor U13032 (N_13032,N_8770,N_9524);
and U13033 (N_13033,N_7797,N_7920);
or U13034 (N_13034,N_7224,N_11812);
xor U13035 (N_13035,N_9229,N_9218);
nor U13036 (N_13036,N_9519,N_10722);
nand U13037 (N_13037,N_6638,N_6407);
and U13038 (N_13038,N_12094,N_11137);
and U13039 (N_13039,N_11170,N_11828);
or U13040 (N_13040,N_7493,N_11594);
and U13041 (N_13041,N_8271,N_7793);
or U13042 (N_13042,N_6418,N_7610);
or U13043 (N_13043,N_10139,N_7287);
nand U13044 (N_13044,N_8635,N_10128);
nor U13045 (N_13045,N_9570,N_7438);
and U13046 (N_13046,N_7818,N_6795);
nor U13047 (N_13047,N_11761,N_12417);
and U13048 (N_13048,N_6515,N_8619);
nor U13049 (N_13049,N_8524,N_8124);
or U13050 (N_13050,N_9672,N_9038);
and U13051 (N_13051,N_12082,N_8434);
nand U13052 (N_13052,N_9494,N_10356);
or U13053 (N_13053,N_8202,N_7808);
nand U13054 (N_13054,N_11184,N_7919);
and U13055 (N_13055,N_9553,N_10349);
nand U13056 (N_13056,N_9799,N_7091);
xor U13057 (N_13057,N_8721,N_7673);
xnor U13058 (N_13058,N_11507,N_6423);
and U13059 (N_13059,N_8098,N_11901);
or U13060 (N_13060,N_7998,N_11074);
or U13061 (N_13061,N_7644,N_10876);
nand U13062 (N_13062,N_9464,N_6960);
nand U13063 (N_13063,N_9119,N_8939);
nand U13064 (N_13064,N_9422,N_7201);
nand U13065 (N_13065,N_10151,N_6636);
and U13066 (N_13066,N_6403,N_9552);
or U13067 (N_13067,N_9992,N_9895);
nor U13068 (N_13068,N_7008,N_9206);
nand U13069 (N_13069,N_11781,N_7121);
nand U13070 (N_13070,N_8793,N_11345);
or U13071 (N_13071,N_7975,N_9490);
or U13072 (N_13072,N_12163,N_6278);
or U13073 (N_13073,N_7741,N_10995);
and U13074 (N_13074,N_8241,N_7204);
nor U13075 (N_13075,N_6733,N_11564);
and U13076 (N_13076,N_11477,N_8679);
and U13077 (N_13077,N_7261,N_7387);
nand U13078 (N_13078,N_7872,N_9555);
and U13079 (N_13079,N_8359,N_10098);
nand U13080 (N_13080,N_10213,N_7756);
nand U13081 (N_13081,N_7381,N_6644);
xnor U13082 (N_13082,N_7836,N_11636);
and U13083 (N_13083,N_10387,N_10656);
or U13084 (N_13084,N_11442,N_10478);
nor U13085 (N_13085,N_11757,N_12143);
nor U13086 (N_13086,N_9098,N_6757);
xor U13087 (N_13087,N_9678,N_8408);
nand U13088 (N_13088,N_8726,N_7258);
nand U13089 (N_13089,N_6432,N_8499);
and U13090 (N_13090,N_11472,N_7974);
nand U13091 (N_13091,N_10975,N_7739);
nand U13092 (N_13092,N_9888,N_6917);
nand U13093 (N_13093,N_11585,N_8020);
and U13094 (N_13094,N_8742,N_9968);
or U13095 (N_13095,N_6714,N_6466);
and U13096 (N_13096,N_8376,N_6512);
and U13097 (N_13097,N_10429,N_8346);
and U13098 (N_13098,N_8832,N_10031);
and U13099 (N_13099,N_12313,N_6436);
xor U13100 (N_13100,N_10314,N_8861);
xnor U13101 (N_13101,N_8010,N_8707);
nor U13102 (N_13102,N_9248,N_10528);
nor U13103 (N_13103,N_11521,N_10383);
or U13104 (N_13104,N_6773,N_11719);
and U13105 (N_13105,N_11783,N_11830);
and U13106 (N_13106,N_9037,N_7033);
and U13107 (N_13107,N_8357,N_12011);
nor U13108 (N_13108,N_8516,N_11276);
nand U13109 (N_13109,N_9259,N_8263);
xor U13110 (N_13110,N_7116,N_8315);
nand U13111 (N_13111,N_12426,N_9975);
or U13112 (N_13112,N_7429,N_9360);
xor U13113 (N_13113,N_9285,N_9140);
nor U13114 (N_13114,N_8243,N_8798);
xnor U13115 (N_13115,N_10382,N_10379);
or U13116 (N_13116,N_7061,N_10668);
nand U13117 (N_13117,N_8252,N_10270);
and U13118 (N_13118,N_10787,N_10793);
and U13119 (N_13119,N_8919,N_7482);
xor U13120 (N_13120,N_6536,N_11835);
nand U13121 (N_13121,N_11361,N_6530);
or U13122 (N_13122,N_11535,N_11601);
or U13123 (N_13123,N_7356,N_8085);
and U13124 (N_13124,N_8627,N_8767);
and U13125 (N_13125,N_8291,N_9376);
xor U13126 (N_13126,N_6724,N_9151);
nor U13127 (N_13127,N_11957,N_6292);
nor U13128 (N_13128,N_11638,N_11860);
nor U13129 (N_13129,N_8901,N_8745);
nor U13130 (N_13130,N_8932,N_10140);
and U13131 (N_13131,N_8890,N_8638);
or U13132 (N_13132,N_11197,N_12440);
and U13133 (N_13133,N_6304,N_10803);
nor U13134 (N_13134,N_7809,N_8407);
and U13135 (N_13135,N_9454,N_6824);
nand U13136 (N_13136,N_9503,N_9515);
and U13137 (N_13137,N_8771,N_8225);
and U13138 (N_13138,N_10841,N_6367);
nor U13139 (N_13139,N_7914,N_12000);
nand U13140 (N_13140,N_6346,N_10978);
or U13141 (N_13141,N_10896,N_7145);
nor U13142 (N_13142,N_6535,N_7220);
nor U13143 (N_13143,N_7658,N_11451);
or U13144 (N_13144,N_10524,N_7151);
or U13145 (N_13145,N_6946,N_8947);
nor U13146 (N_13146,N_8624,N_9149);
xor U13147 (N_13147,N_12179,N_9107);
or U13148 (N_13148,N_11427,N_7177);
and U13149 (N_13149,N_7768,N_10849);
nand U13150 (N_13150,N_9299,N_10321);
nor U13151 (N_13151,N_12191,N_10253);
nand U13152 (N_13152,N_8871,N_9734);
and U13153 (N_13153,N_8228,N_6478);
nand U13154 (N_13154,N_8692,N_7290);
or U13155 (N_13155,N_10754,N_7039);
nand U13156 (N_13156,N_9375,N_10861);
nand U13157 (N_13157,N_9993,N_7132);
nand U13158 (N_13158,N_6873,N_9550);
xnor U13159 (N_13159,N_12401,N_10968);
nand U13160 (N_13160,N_11158,N_9819);
or U13161 (N_13161,N_9838,N_10469);
or U13162 (N_13162,N_7782,N_8038);
xnor U13163 (N_13163,N_10619,N_11218);
nor U13164 (N_13164,N_7377,N_11454);
nor U13165 (N_13165,N_10316,N_11161);
or U13166 (N_13166,N_12256,N_7418);
and U13167 (N_13167,N_11642,N_7087);
and U13168 (N_13168,N_7459,N_10298);
or U13169 (N_13169,N_9815,N_9949);
and U13170 (N_13170,N_11038,N_6592);
nand U13171 (N_13171,N_9609,N_10724);
or U13172 (N_13172,N_9207,N_10418);
and U13173 (N_13173,N_12117,N_10903);
nand U13174 (N_13174,N_11933,N_6470);
nor U13175 (N_13175,N_6748,N_11984);
or U13176 (N_13176,N_9135,N_10807);
xor U13177 (N_13177,N_8561,N_10307);
nor U13178 (N_13178,N_9365,N_8301);
nor U13179 (N_13179,N_7310,N_11253);
xor U13180 (N_13180,N_6613,N_10411);
xnor U13181 (N_13181,N_10009,N_10632);
nor U13182 (N_13182,N_11878,N_10663);
nor U13183 (N_13183,N_8069,N_9903);
or U13184 (N_13184,N_8095,N_11582);
xor U13185 (N_13185,N_7683,N_8211);
xor U13186 (N_13186,N_7637,N_6956);
nor U13187 (N_13187,N_6511,N_9754);
or U13188 (N_13188,N_7396,N_10686);
nor U13189 (N_13189,N_12299,N_12116);
or U13190 (N_13190,N_11893,N_9319);
xor U13191 (N_13191,N_11072,N_7392);
nor U13192 (N_13192,N_10771,N_9065);
nor U13193 (N_13193,N_10925,N_10689);
xor U13194 (N_13194,N_8560,N_10212);
nor U13195 (N_13195,N_11458,N_9735);
nand U13196 (N_13196,N_9814,N_6627);
and U13197 (N_13197,N_6986,N_12039);
nor U13198 (N_13198,N_7832,N_12096);
nand U13199 (N_13199,N_8598,N_11587);
and U13200 (N_13200,N_9689,N_9513);
nor U13201 (N_13201,N_8262,N_9056);
nor U13202 (N_13202,N_8775,N_7953);
or U13203 (N_13203,N_9244,N_11802);
and U13204 (N_13204,N_10792,N_9517);
and U13205 (N_13205,N_9196,N_9499);
and U13206 (N_13206,N_6852,N_7930);
and U13207 (N_13207,N_12409,N_12262);
or U13208 (N_13208,N_8486,N_12154);
nand U13209 (N_13209,N_11118,N_6484);
nor U13210 (N_13210,N_12173,N_7798);
and U13211 (N_13211,N_8345,N_9804);
nand U13212 (N_13212,N_8972,N_7862);
nand U13213 (N_13213,N_10338,N_9417);
or U13214 (N_13214,N_6955,N_8144);
and U13215 (N_13215,N_11384,N_9749);
nor U13216 (N_13216,N_8892,N_6674);
or U13217 (N_13217,N_6427,N_11248);
and U13218 (N_13218,N_11824,N_7412);
xnor U13219 (N_13219,N_9361,N_6899);
or U13220 (N_13220,N_11192,N_8876);
nand U13221 (N_13221,N_11408,N_9512);
and U13222 (N_13222,N_8720,N_11721);
and U13223 (N_13223,N_11698,N_11856);
and U13224 (N_13224,N_12222,N_6641);
and U13225 (N_13225,N_10505,N_9761);
nor U13226 (N_13226,N_6752,N_8375);
or U13227 (N_13227,N_11708,N_10390);
nor U13228 (N_13228,N_7026,N_10029);
nand U13229 (N_13229,N_11227,N_7043);
xnor U13230 (N_13230,N_7317,N_9131);
nor U13231 (N_13231,N_10789,N_6816);
nor U13232 (N_13232,N_6784,N_11791);
nor U13233 (N_13233,N_8788,N_8107);
nor U13234 (N_13234,N_6577,N_7444);
nand U13235 (N_13235,N_6778,N_12310);
nand U13236 (N_13236,N_9514,N_8668);
or U13237 (N_13237,N_7122,N_8232);
or U13238 (N_13238,N_7492,N_9369);
or U13239 (N_13239,N_8641,N_7042);
nand U13240 (N_13240,N_10417,N_11723);
or U13241 (N_13241,N_6257,N_8554);
or U13242 (N_13242,N_7969,N_9638);
nor U13243 (N_13243,N_6709,N_8551);
or U13244 (N_13244,N_9240,N_6343);
nand U13245 (N_13245,N_10835,N_12451);
or U13246 (N_13246,N_8383,N_8988);
nand U13247 (N_13247,N_10402,N_6985);
nor U13248 (N_13248,N_12423,N_11926);
nand U13249 (N_13249,N_10108,N_10982);
xnor U13250 (N_13250,N_11198,N_9418);
nor U13251 (N_13251,N_7740,N_6762);
nor U13252 (N_13252,N_6348,N_7343);
nand U13253 (N_13253,N_6892,N_8614);
or U13254 (N_13254,N_10854,N_6890);
nor U13255 (N_13255,N_8264,N_8304);
nor U13256 (N_13256,N_11625,N_6546);
or U13257 (N_13257,N_7301,N_11977);
or U13258 (N_13258,N_12045,N_9221);
xnor U13259 (N_13259,N_6896,N_9165);
nor U13260 (N_13260,N_11350,N_10431);
nor U13261 (N_13261,N_6362,N_7183);
nor U13262 (N_13262,N_11996,N_10045);
and U13263 (N_13263,N_12374,N_6524);
or U13264 (N_13264,N_7313,N_7672);
nand U13265 (N_13265,N_9245,N_10249);
or U13266 (N_13266,N_7353,N_10180);
nand U13267 (N_13267,N_11825,N_10624);
nand U13268 (N_13268,N_10051,N_7800);
nor U13269 (N_13269,N_9691,N_10230);
nand U13270 (N_13270,N_10534,N_12068);
and U13271 (N_13271,N_9411,N_6793);
nand U13272 (N_13272,N_10657,N_10569);
nand U13273 (N_13273,N_11379,N_6962);
nand U13274 (N_13274,N_7563,N_10786);
and U13275 (N_13275,N_11097,N_7917);
and U13276 (N_13276,N_9205,N_8094);
xor U13277 (N_13277,N_7906,N_12072);
nor U13278 (N_13278,N_10913,N_7124);
nand U13279 (N_13279,N_10274,N_8242);
nor U13280 (N_13280,N_10530,N_9746);
nor U13281 (N_13281,N_12010,N_10974);
or U13282 (N_13282,N_9019,N_7360);
and U13283 (N_13283,N_7830,N_7045);
or U13284 (N_13284,N_7980,N_10415);
nand U13285 (N_13285,N_7038,N_7899);
xor U13286 (N_13286,N_12003,N_11259);
nand U13287 (N_13287,N_7458,N_9064);
xor U13288 (N_13288,N_12353,N_9366);
nand U13289 (N_13289,N_8902,N_8081);
and U13290 (N_13290,N_10320,N_10192);
or U13291 (N_13291,N_9917,N_8850);
xnor U13292 (N_13292,N_10050,N_8378);
xnor U13293 (N_13293,N_11230,N_10300);
nor U13294 (N_13294,N_12418,N_8025);
xnor U13295 (N_13295,N_10679,N_7380);
and U13296 (N_13296,N_10242,N_8600);
nand U13297 (N_13297,N_9886,N_12155);
and U13298 (N_13298,N_10817,N_6932);
nor U13299 (N_13299,N_11789,N_11315);
and U13300 (N_13300,N_7105,N_9508);
and U13301 (N_13301,N_11895,N_9324);
nand U13302 (N_13302,N_6730,N_9260);
nor U13303 (N_13303,N_10086,N_9309);
and U13304 (N_13304,N_10969,N_8165);
and U13305 (N_13305,N_6908,N_10421);
nor U13306 (N_13306,N_7959,N_6542);
nor U13307 (N_13307,N_11281,N_7303);
nor U13308 (N_13308,N_8363,N_9542);
or U13309 (N_13309,N_9146,N_8859);
or U13310 (N_13310,N_10780,N_6806);
nand U13311 (N_13311,N_11483,N_7689);
nor U13312 (N_13312,N_11189,N_6562);
nand U13313 (N_13313,N_11778,N_11567);
nor U13314 (N_13314,N_8634,N_10273);
xnor U13315 (N_13315,N_7733,N_11479);
and U13316 (N_13316,N_10963,N_12128);
nor U13317 (N_13317,N_11744,N_11792);
nand U13318 (N_13318,N_7634,N_6847);
xor U13319 (N_13319,N_10077,N_12131);
or U13320 (N_13320,N_6526,N_7404);
nand U13321 (N_13321,N_11972,N_9703);
xor U13322 (N_13322,N_10782,N_8356);
nor U13323 (N_13323,N_8270,N_12129);
nand U13324 (N_13324,N_8329,N_10567);
nand U13325 (N_13325,N_7591,N_8594);
or U13326 (N_13326,N_6589,N_10223);
and U13327 (N_13327,N_7185,N_10219);
nand U13328 (N_13328,N_9005,N_11844);
nor U13329 (N_13329,N_11851,N_11063);
or U13330 (N_13330,N_10994,N_12214);
nor U13331 (N_13331,N_10751,N_11543);
nand U13332 (N_13332,N_10602,N_9875);
nand U13333 (N_13333,N_9702,N_11707);
nand U13334 (N_13334,N_9156,N_10475);
nand U13335 (N_13335,N_9959,N_12415);
and U13336 (N_13336,N_10892,N_11470);
nor U13337 (N_13337,N_10818,N_11461);
or U13338 (N_13338,N_11071,N_7388);
nand U13339 (N_13339,N_7545,N_8099);
and U13340 (N_13340,N_12453,N_12484);
and U13341 (N_13341,N_7049,N_11934);
nor U13342 (N_13342,N_6496,N_8500);
or U13343 (N_13343,N_8350,N_10149);
or U13344 (N_13344,N_9290,N_11309);
or U13345 (N_13345,N_10813,N_10990);
or U13346 (N_13346,N_8204,N_8513);
nor U13347 (N_13347,N_11434,N_10615);
nand U13348 (N_13348,N_9453,N_9758);
nand U13349 (N_13349,N_7622,N_11292);
nor U13350 (N_13350,N_12050,N_8033);
xnor U13351 (N_13351,N_10081,N_10269);
nand U13352 (N_13352,N_6294,N_7662);
xnor U13353 (N_13353,N_10642,N_7536);
and U13354 (N_13354,N_7024,N_11973);
xor U13355 (N_13355,N_10637,N_8529);
and U13356 (N_13356,N_10900,N_11689);
and U13357 (N_13357,N_7647,N_10510);
xnor U13358 (N_13358,N_10846,N_10954);
nand U13359 (N_13359,N_12372,N_7025);
nor U13360 (N_13360,N_7238,N_10520);
nand U13361 (N_13361,N_9099,N_6329);
or U13362 (N_13362,N_11595,N_12487);
or U13363 (N_13363,N_6575,N_11358);
nand U13364 (N_13364,N_11720,N_11413);
and U13365 (N_13365,N_9338,N_12280);
nor U13366 (N_13366,N_8684,N_10991);
and U13367 (N_13367,N_10420,N_6324);
nand U13368 (N_13368,N_8683,N_11728);
or U13369 (N_13369,N_8894,N_12319);
nor U13370 (N_13370,N_8531,N_6634);
or U13371 (N_13371,N_8269,N_10943);
and U13372 (N_13372,N_11096,N_6591);
nor U13373 (N_13373,N_8259,N_8481);
nor U13374 (N_13374,N_8783,N_7093);
nor U13375 (N_13375,N_6788,N_10441);
or U13376 (N_13376,N_8275,N_10714);
xor U13377 (N_13377,N_10721,N_9341);
nand U13378 (N_13378,N_9745,N_10353);
or U13379 (N_13379,N_6936,N_11369);
nor U13380 (N_13380,N_8986,N_10218);
nand U13381 (N_13381,N_8729,N_10678);
xor U13382 (N_13382,N_7065,N_7190);
nand U13383 (N_13383,N_8160,N_6338);
or U13384 (N_13384,N_10129,N_7006);
or U13385 (N_13385,N_9340,N_11569);
or U13386 (N_13386,N_7885,N_8740);
nor U13387 (N_13387,N_12287,N_6580);
nor U13388 (N_13388,N_11028,N_8665);
xnor U13389 (N_13389,N_6272,N_9877);
and U13390 (N_13390,N_9790,N_9715);
or U13391 (N_13391,N_6646,N_10700);
or U13392 (N_13392,N_8472,N_10701);
or U13393 (N_13393,N_10755,N_9261);
and U13394 (N_13394,N_6377,N_10529);
nor U13395 (N_13395,N_6746,N_9414);
and U13396 (N_13396,N_6978,N_8423);
nand U13397 (N_13397,N_11574,N_6548);
nor U13398 (N_13398,N_9276,N_12254);
and U13399 (N_13399,N_7028,N_11269);
nor U13400 (N_13400,N_10498,N_11755);
and U13401 (N_13401,N_11255,N_6414);
or U13402 (N_13402,N_10966,N_12281);
nand U13403 (N_13403,N_8605,N_9559);
nand U13404 (N_13404,N_6781,N_7852);
nand U13405 (N_13405,N_9496,N_10092);
and U13406 (N_13406,N_11848,N_10747);
and U13407 (N_13407,N_11238,N_8469);
nor U13408 (N_13408,N_9035,N_9641);
nor U13409 (N_13409,N_6796,N_10085);
and U13410 (N_13410,N_7593,N_7289);
or U13411 (N_13411,N_8451,N_6309);
nor U13412 (N_13412,N_7665,N_12007);
nand U13413 (N_13413,N_10281,N_9739);
nand U13414 (N_13414,N_6434,N_6482);
and U13415 (N_13415,N_11955,N_8730);
nor U13416 (N_13416,N_7101,N_6614);
or U13417 (N_13417,N_9998,N_7550);
or U13418 (N_13418,N_8821,N_7538);
or U13419 (N_13419,N_10189,N_8992);
and U13420 (N_13420,N_9601,N_11701);
or U13421 (N_13421,N_8944,N_12271);
or U13422 (N_13422,N_8537,N_7767);
and U13423 (N_13423,N_10117,N_7440);
or U13424 (N_13424,N_11581,N_7252);
nor U13425 (N_13425,N_10741,N_8128);
nor U13426 (N_13426,N_7877,N_7178);
nor U13427 (N_13427,N_10810,N_10254);
nand U13428 (N_13428,N_6874,N_9756);
nor U13429 (N_13429,N_8130,N_7577);
and U13430 (N_13430,N_7046,N_6897);
or U13431 (N_13431,N_9811,N_9671);
and U13432 (N_13432,N_12476,N_11469);
and U13433 (N_13433,N_9665,N_10361);
xor U13434 (N_13434,N_7451,N_9652);
and U13435 (N_13435,N_11683,N_7358);
and U13436 (N_13436,N_10766,N_7274);
and U13437 (N_13437,N_11655,N_12479);
or U13438 (N_13438,N_11385,N_6799);
nand U13439 (N_13439,N_8752,N_9942);
nand U13440 (N_13440,N_7805,N_11563);
and U13441 (N_13441,N_11619,N_12364);
nor U13442 (N_13442,N_9381,N_10756);
or U13443 (N_13443,N_8414,N_12383);
nand U13444 (N_13444,N_10062,N_7084);
or U13445 (N_13445,N_12238,N_12025);
and U13446 (N_13446,N_10052,N_10033);
xor U13447 (N_13447,N_11409,N_7520);
and U13448 (N_13448,N_9645,N_7315);
and U13449 (N_13449,N_10509,N_10120);
xnor U13450 (N_13450,N_12200,N_12413);
and U13451 (N_13451,N_7706,N_7221);
and U13452 (N_13452,N_9820,N_9743);
and U13453 (N_13453,N_10322,N_10865);
xor U13454 (N_13454,N_6404,N_11559);
and U13455 (N_13455,N_10744,N_7495);
or U13456 (N_13456,N_9543,N_11593);
or U13457 (N_13457,N_11279,N_8875);
nand U13458 (N_13458,N_9929,N_9607);
nor U13459 (N_13459,N_7417,N_9339);
and U13460 (N_13460,N_8509,N_12064);
or U13461 (N_13461,N_7094,N_6499);
and U13462 (N_13462,N_12292,N_8785);
nor U13463 (N_13463,N_8145,N_10518);
or U13464 (N_13464,N_8762,N_9518);
or U13465 (N_13465,N_10153,N_6402);
or U13466 (N_13466,N_6376,N_10664);
nand U13467 (N_13467,N_8690,N_8210);
nand U13468 (N_13468,N_8777,N_8558);
nor U13469 (N_13469,N_11185,N_9018);
nor U13470 (N_13470,N_11529,N_11738);
or U13471 (N_13471,N_10711,N_7217);
nor U13472 (N_13472,N_11515,N_6571);
nand U13473 (N_13473,N_11839,N_10546);
nand U13474 (N_13474,N_12387,N_11635);
and U13475 (N_13475,N_9934,N_9802);
and U13476 (N_13476,N_10366,N_8086);
nor U13477 (N_13477,N_10293,N_7040);
nand U13478 (N_13478,N_9297,N_12486);
nand U13479 (N_13479,N_7609,N_11769);
nor U13480 (N_13480,N_11431,N_11089);
or U13481 (N_13481,N_7963,N_12378);
and U13482 (N_13482,N_11611,N_7604);
nand U13483 (N_13483,N_7791,N_11445);
nor U13484 (N_13484,N_7810,N_11914);
or U13485 (N_13485,N_12263,N_7926);
nand U13486 (N_13486,N_6468,N_11589);
or U13487 (N_13487,N_6677,N_6485);
nor U13488 (N_13488,N_11297,N_9438);
or U13489 (N_13489,N_9208,N_7425);
nor U13490 (N_13490,N_8231,N_9379);
and U13491 (N_13491,N_7664,N_8131);
nand U13492 (N_13492,N_8917,N_9008);
xor U13493 (N_13493,N_7254,N_10930);
xnor U13494 (N_13494,N_12403,N_10276);
nor U13495 (N_13495,N_11356,N_9610);
and U13496 (N_13496,N_12285,N_8380);
nand U13497 (N_13497,N_9572,N_11176);
or U13498 (N_13498,N_12103,N_8446);
and U13499 (N_13499,N_11278,N_7126);
xnor U13500 (N_13500,N_9574,N_8942);
or U13501 (N_13501,N_7895,N_6622);
and U13502 (N_13502,N_9452,N_7022);
nand U13503 (N_13503,N_9088,N_7389);
or U13504 (N_13504,N_10198,N_8227);
nand U13505 (N_13505,N_9303,N_10472);
and U13506 (N_13506,N_12111,N_7159);
nand U13507 (N_13507,N_6446,N_6750);
and U13508 (N_13508,N_6441,N_11912);
nor U13509 (N_13509,N_10344,N_8521);
nand U13510 (N_13510,N_10055,N_6764);
and U13511 (N_13511,N_8854,N_10960);
xor U13512 (N_13512,N_7838,N_6416);
nor U13513 (N_13513,N_11511,N_7448);
or U13514 (N_13514,N_9716,N_12243);
nand U13515 (N_13515,N_11869,N_10681);
nand U13516 (N_13516,N_6543,N_9306);
and U13517 (N_13517,N_7940,N_12455);
nand U13518 (N_13518,N_11633,N_6676);
nand U13519 (N_13519,N_9630,N_10847);
or U13520 (N_13520,N_11542,N_6790);
or U13521 (N_13521,N_11983,N_9822);
or U13522 (N_13522,N_8419,N_9981);
nor U13523 (N_13523,N_11237,N_7736);
and U13524 (N_13524,N_8576,N_9087);
or U13525 (N_13525,N_6349,N_8109);
nand U13526 (N_13526,N_6320,N_9122);
or U13527 (N_13527,N_9765,N_7703);
or U13528 (N_13528,N_12322,N_11352);
or U13529 (N_13529,N_11182,N_11864);
nor U13530 (N_13530,N_9271,N_10097);
xor U13531 (N_13531,N_10395,N_8178);
nor U13532 (N_13532,N_10381,N_9041);
nand U13533 (N_13533,N_6544,N_10589);
and U13534 (N_13534,N_10388,N_9796);
nor U13535 (N_13535,N_10735,N_11254);
nand U13536 (N_13536,N_8140,N_8115);
and U13537 (N_13537,N_9732,N_8542);
nor U13538 (N_13538,N_10466,N_8825);
nor U13539 (N_13539,N_7789,N_11261);
nor U13540 (N_13540,N_12106,N_11314);
nand U13541 (N_13541,N_10245,N_8681);
nand U13542 (N_13542,N_6770,N_7861);
nand U13543 (N_13543,N_11514,N_12393);
or U13544 (N_13544,N_10251,N_10599);
xnor U13545 (N_13545,N_12078,N_8713);
nand U13546 (N_13546,N_10834,N_9673);
and U13547 (N_13547,N_8997,N_11522);
nand U13548 (N_13548,N_12097,N_12074);
or U13549 (N_13549,N_11365,N_11737);
nand U13550 (N_13550,N_10611,N_6323);
nor U13551 (N_13551,N_10560,N_9901);
nand U13552 (N_13552,N_9138,N_9314);
and U13553 (N_13553,N_10916,N_10363);
nand U13554 (N_13554,N_9566,N_6539);
and U13555 (N_13555,N_6473,N_7200);
nor U13556 (N_13556,N_11986,N_6313);
or U13557 (N_13557,N_9168,N_11142);
nand U13558 (N_13558,N_6717,N_10303);
nand U13559 (N_13559,N_7776,N_6266);
nand U13560 (N_13560,N_6449,N_10951);
or U13561 (N_13561,N_12257,N_11872);
nand U13562 (N_13562,N_7944,N_9372);
nand U13563 (N_13563,N_9781,N_6859);
or U13564 (N_13564,N_6517,N_10224);
nand U13565 (N_13565,N_8495,N_7915);
and U13566 (N_13566,N_6463,N_6642);
xor U13567 (N_13567,N_6518,N_7333);
nor U13568 (N_13568,N_10317,N_9125);
nor U13569 (N_13569,N_7455,N_12320);
nor U13570 (N_13570,N_9582,N_8083);
nor U13571 (N_13571,N_11002,N_6424);
or U13572 (N_13572,N_10404,N_9785);
and U13573 (N_13573,N_9442,N_8868);
or U13574 (N_13574,N_9234,N_7516);
nand U13575 (N_13575,N_6661,N_7929);
or U13576 (N_13576,N_11064,N_7293);
and U13577 (N_13577,N_7931,N_6361);
or U13578 (N_13578,N_7368,N_6707);
nand U13579 (N_13579,N_11214,N_8487);
and U13580 (N_13580,N_6830,N_9072);
nor U13581 (N_13581,N_10453,N_8592);
nor U13582 (N_13582,N_9127,N_10146);
and U13583 (N_13583,N_7594,N_9332);
nor U13584 (N_13584,N_6281,N_11686);
nand U13585 (N_13585,N_6280,N_6625);
or U13586 (N_13586,N_7372,N_6435);
or U13587 (N_13587,N_9915,N_12170);
or U13588 (N_13588,N_7212,N_9709);
nor U13589 (N_13589,N_11578,N_8749);
or U13590 (N_13590,N_10895,N_10315);
xnor U13591 (N_13591,N_9837,N_11504);
or U13592 (N_13592,N_9893,N_8031);
nor U13593 (N_13593,N_10480,N_9109);
and U13594 (N_13594,N_6672,N_7079);
or U13595 (N_13595,N_7618,N_11406);
nand U13596 (N_13596,N_10391,N_9961);
or U13597 (N_13597,N_7166,N_8457);
nand U13598 (N_13598,N_7549,N_9971);
and U13599 (N_13599,N_6277,N_12033);
or U13600 (N_13600,N_9160,N_8617);
or U13601 (N_13601,N_11243,N_11322);
or U13602 (N_13602,N_7507,N_7086);
and U13603 (N_13603,N_7311,N_7292);
or U13604 (N_13604,N_8548,N_10329);
nand U13605 (N_13605,N_6972,N_10958);
or U13606 (N_13606,N_8218,N_6450);
or U13607 (N_13607,N_9615,N_10265);
or U13608 (N_13608,N_10114,N_10376);
or U13609 (N_13609,N_8148,N_7477);
and U13610 (N_13610,N_11874,N_7608);
nand U13611 (N_13611,N_6616,N_11777);
nand U13612 (N_13612,N_7893,N_8719);
and U13613 (N_13613,N_7378,N_7218);
nor U13614 (N_13614,N_8037,N_6270);
nor U13615 (N_13615,N_7555,N_8867);
nand U13616 (N_13616,N_6923,N_6711);
nor U13617 (N_13617,N_9933,N_12223);
and U13618 (N_13618,N_11433,N_8637);
and U13619 (N_13619,N_11272,N_7837);
or U13620 (N_13620,N_10170,N_7645);
nor U13621 (N_13621,N_6683,N_10588);
or U13622 (N_13622,N_12228,N_6561);
nor U13623 (N_13623,N_11159,N_10941);
nor U13624 (N_13624,N_12259,N_11881);
or U13625 (N_13625,N_10939,N_10805);
xor U13626 (N_13626,N_7910,N_10078);
or U13627 (N_13627,N_11576,N_7936);
xor U13628 (N_13628,N_10820,N_6680);
nor U13629 (N_13629,N_9594,N_9602);
nor U13630 (N_13630,N_12348,N_8180);
nor U13631 (N_13631,N_6386,N_6970);
nor U13632 (N_13632,N_10909,N_8978);
nand U13633 (N_13633,N_9777,N_8962);
nand U13634 (N_13634,N_7857,N_10646);
nand U13635 (N_13635,N_11772,N_8309);
xor U13636 (N_13636,N_12110,N_8286);
and U13637 (N_13637,N_10752,N_7321);
nor U13638 (N_13638,N_10194,N_11685);
and U13639 (N_13639,N_6996,N_7676);
and U13640 (N_13640,N_7195,N_10508);
and U13641 (N_13641,N_11025,N_8907);
nand U13642 (N_13642,N_9427,N_9059);
or U13643 (N_13643,N_7326,N_8017);
xnor U13644 (N_13644,N_8639,N_7709);
nand U13645 (N_13645,N_8484,N_7433);
and U13646 (N_13646,N_8064,N_7627);
nand U13647 (N_13647,N_9956,N_6810);
nor U13648 (N_13648,N_9626,N_7411);
nand U13649 (N_13649,N_11950,N_12058);
nand U13650 (N_13650,N_8750,N_10640);
nand U13651 (N_13651,N_11140,N_9584);
xnor U13652 (N_13652,N_12498,N_6269);
and U13653 (N_13653,N_7754,N_6572);
xor U13654 (N_13654,N_8110,N_8949);
nand U13655 (N_13655,N_8881,N_9480);
nand U13656 (N_13656,N_11061,N_12161);
nand U13657 (N_13657,N_11803,N_8463);
or U13658 (N_13658,N_11742,N_6256);
or U13659 (N_13659,N_9826,N_10412);
or U13660 (N_13660,N_8332,N_6415);
and U13661 (N_13661,N_9618,N_6957);
or U13662 (N_13662,N_6318,N_7788);
xor U13663 (N_13663,N_11691,N_10059);
nor U13664 (N_13664,N_9359,N_10715);
or U13665 (N_13665,N_8879,N_7272);
xor U13666 (N_13666,N_10827,N_7270);
nand U13667 (N_13667,N_10234,N_8491);
nand U13668 (N_13668,N_11362,N_8137);
nor U13669 (N_13669,N_10177,N_6618);
nand U13670 (N_13670,N_9979,N_6447);
and U13671 (N_13671,N_7023,N_10495);
nand U13672 (N_13672,N_12169,N_9385);
nand U13673 (N_13673,N_12463,N_7279);
and U13674 (N_13674,N_9462,N_6920);
nand U13675 (N_13675,N_10460,N_9291);
nor U13676 (N_13676,N_7750,N_7623);
nor U13677 (N_13677,N_6298,N_11065);
and U13678 (N_13678,N_9213,N_12207);
nor U13679 (N_13679,N_12332,N_10526);
nor U13680 (N_13680,N_7148,N_12267);
or U13681 (N_13681,N_9242,N_6459);
nor U13682 (N_13682,N_7762,N_8076);
or U13683 (N_13683,N_10147,N_7080);
or U13684 (N_13684,N_6567,N_7306);
nor U13685 (N_13685,N_7250,N_6871);
nor U13686 (N_13686,N_10386,N_11880);
nor U13687 (N_13687,N_8957,N_6856);
or U13688 (N_13688,N_7871,N_10795);
or U13689 (N_13689,N_7074,N_8147);
nor U13690 (N_13690,N_8222,N_7103);
and U13691 (N_13691,N_7067,N_6775);
nand U13692 (N_13692,N_10444,N_11180);
or U13693 (N_13693,N_11641,N_10545);
nand U13694 (N_13694,N_9378,N_6692);
nor U13695 (N_13695,N_9223,N_6534);
or U13696 (N_13696,N_7878,N_9263);
and U13697 (N_13697,N_12301,N_12152);
and U13698 (N_13698,N_7391,N_10591);
nand U13699 (N_13699,N_9426,N_12194);
nand U13700 (N_13700,N_11845,N_6537);
and U13701 (N_13701,N_9203,N_10173);
nor U13702 (N_13702,N_9279,N_7219);
nand U13703 (N_13703,N_12296,N_11940);
or U13704 (N_13704,N_7778,N_8985);
nand U13705 (N_13705,N_10215,N_6693);
nor U13706 (N_13706,N_10083,N_11268);
nor U13707 (N_13707,N_10506,N_9586);
or U13708 (N_13708,N_8442,N_8609);
or U13709 (N_13709,N_9769,N_11968);
nand U13710 (N_13710,N_9631,N_11539);
and U13711 (N_13711,N_9869,N_8640);
nand U13712 (N_13712,N_10644,N_11620);
xnor U13713 (N_13713,N_8201,N_7946);
and U13714 (N_13714,N_10326,N_6645);
and U13715 (N_13715,N_9906,N_10428);
or U13716 (N_13716,N_7162,N_6783);
or U13717 (N_13717,N_9498,N_12122);
nand U13718 (N_13718,N_8573,N_9733);
or U13719 (N_13719,N_11814,N_6941);
nand U13720 (N_13720,N_10464,N_10500);
nor U13721 (N_13721,N_10163,N_11524);
and U13722 (N_13722,N_7471,N_7073);
and U13723 (N_13723,N_11942,N_12457);
or U13724 (N_13724,N_10439,N_8915);
nand U13725 (N_13725,N_11215,N_11342);
nor U13726 (N_13726,N_9188,N_12165);
or U13727 (N_13727,N_10105,N_11449);
nor U13728 (N_13728,N_9423,N_10905);
nand U13729 (N_13729,N_10867,N_11813);
nor U13730 (N_13730,N_9111,N_11967);
nand U13731 (N_13731,N_9698,N_12362);
nor U13732 (N_13732,N_11338,N_9076);
nor U13733 (N_13733,N_7251,N_8322);
xor U13734 (N_13734,N_10467,N_6979);
nor U13735 (N_13735,N_11712,N_8007);
and U13736 (N_13736,N_10684,N_9424);
nand U13737 (N_13737,N_8885,N_10924);
nand U13738 (N_13738,N_10821,N_10614);
nand U13739 (N_13739,N_9413,N_10332);
nand U13740 (N_13740,N_8236,N_11797);
or U13741 (N_13741,N_6828,N_6299);
nand U13742 (N_13742,N_10986,N_7273);
xnor U13743 (N_13743,N_12428,N_9429);
and U13744 (N_13744,N_6341,N_12031);
nor U13745 (N_13745,N_7587,N_10043);
or U13746 (N_13746,N_8946,N_9269);
nor U13747 (N_13747,N_8088,N_12311);
or U13748 (N_13748,N_8396,N_11592);
nand U13749 (N_13749,N_7248,N_12005);
nand U13750 (N_13750,N_11732,N_11375);
nand U13751 (N_13751,N_11516,N_8282);
nor U13752 (N_13752,N_12352,N_7557);
and U13753 (N_13753,N_8104,N_8882);
nor U13754 (N_13754,N_7226,N_9355);
nor U13755 (N_13755,N_11949,N_6380);
nand U13756 (N_13756,N_9845,N_6965);
nand U13757 (N_13757,N_10888,N_11135);
nor U13758 (N_13758,N_8787,N_11471);
xor U13759 (N_13759,N_12066,N_10859);
xor U13760 (N_13760,N_7332,N_7699);
or U13761 (N_13761,N_7196,N_9976);
and U13762 (N_13762,N_9685,N_11226);
nand U13763 (N_13763,N_11767,N_12021);
xnor U13764 (N_13764,N_6513,N_9969);
nor U13765 (N_13765,N_11095,N_11713);
nand U13766 (N_13766,N_6767,N_9139);
nand U13767 (N_13767,N_12305,N_6704);
nand U13768 (N_13768,N_7749,N_11293);
nor U13769 (N_13769,N_10228,N_9030);
xnor U13770 (N_13770,N_12306,N_6334);
xor U13771 (N_13771,N_6777,N_12112);
and U13772 (N_13772,N_11282,N_11733);
nor U13773 (N_13773,N_11225,N_7323);
or U13774 (N_13774,N_9313,N_8755);
xnor U13775 (N_13775,N_10042,N_11032);
or U13776 (N_13776,N_11212,N_11335);
or U13777 (N_13777,N_11922,N_7607);
or U13778 (N_13778,N_10680,N_7379);
nand U13779 (N_13779,N_10576,N_6454);
nor U13780 (N_13780,N_10001,N_8601);
nand U13781 (N_13781,N_11257,N_11706);
nor U13782 (N_13782,N_10426,N_8811);
and U13783 (N_13783,N_9212,N_8809);
or U13784 (N_13784,N_6330,N_11715);
or U13785 (N_13785,N_9925,N_10183);
xnor U13786 (N_13786,N_8675,N_10458);
and U13787 (N_13787,N_9482,N_11280);
nand U13788 (N_13788,N_9287,N_7528);
and U13789 (N_13789,N_11951,N_7399);
or U13790 (N_13790,N_10427,N_6980);
xor U13791 (N_13791,N_11684,N_9912);
nand U13792 (N_13792,N_6437,N_11999);
nand U13793 (N_13793,N_9124,N_6895);
and U13794 (N_13794,N_7467,N_7950);
nor U13795 (N_13795,N_10489,N_10661);
nor U13796 (N_13796,N_10595,N_8716);
nand U13797 (N_13797,N_7948,N_11126);
nand U13798 (N_13798,N_7823,N_6751);
and U13799 (N_13799,N_7484,N_8659);
and U13800 (N_13800,N_7724,N_8784);
nand U13801 (N_13801,N_9446,N_7575);
nor U13802 (N_13802,N_9862,N_6827);
and U13803 (N_13803,N_10076,N_12183);
and U13804 (N_13804,N_11228,N_7841);
xor U13805 (N_13805,N_10765,N_11818);
nand U13806 (N_13806,N_11275,N_11884);
nand U13807 (N_13807,N_8908,N_10174);
nor U13808 (N_13808,N_8786,N_12040);
or U13809 (N_13809,N_9648,N_11650);
and U13810 (N_13810,N_7541,N_8799);
or U13811 (N_13811,N_9352,N_9712);
xnor U13812 (N_13812,N_11103,N_9090);
and U13813 (N_13813,N_11015,N_8817);
nor U13814 (N_13814,N_11598,N_10573);
nand U13815 (N_13815,N_11299,N_7414);
nor U13816 (N_13816,N_6794,N_10940);
nor U13817 (N_13817,N_8208,N_8493);
nor U13818 (N_13818,N_11959,N_12151);
and U13819 (N_13819,N_11001,N_7422);
nand U13820 (N_13820,N_11752,N_11475);
or U13821 (N_13821,N_7169,N_10348);
nor U13822 (N_13822,N_9627,N_8126);
nor U13823 (N_13823,N_7682,N_6872);
and U13824 (N_13824,N_12252,N_12260);
and U13825 (N_13825,N_8686,N_11793);
nor U13826 (N_13826,N_8029,N_9996);
xor U13827 (N_13827,N_8117,N_11992);
and U13828 (N_13828,N_12391,N_11560);
or U13829 (N_13829,N_11929,N_10145);
nand U13830 (N_13830,N_11924,N_6916);
nand U13831 (N_13831,N_11747,N_10127);
xnor U13832 (N_13832,N_10046,N_11659);
or U13833 (N_13833,N_11120,N_12258);
and U13834 (N_13834,N_11758,N_12308);
or U13835 (N_13835,N_9742,N_10898);
nand U13836 (N_13836,N_8187,N_8113);
nor U13837 (N_13837,N_12184,N_9701);
nand U13838 (N_13838,N_9988,N_7513);
or U13839 (N_13839,N_10762,N_10158);
or U13840 (N_13840,N_11478,N_6819);
or U13841 (N_13841,N_11164,N_6780);
or U13842 (N_13842,N_11969,N_12026);
or U13843 (N_13843,N_6718,N_12006);
nor U13844 (N_13844,N_8189,N_11586);
nor U13845 (N_13845,N_10948,N_9536);
or U13846 (N_13846,N_7690,N_11435);
or U13847 (N_13847,N_7639,N_10447);
or U13848 (N_13848,N_12102,N_7510);
nand U13849 (N_13849,N_7413,N_6785);
or U13850 (N_13850,N_12138,N_11234);
or U13851 (N_13851,N_10454,N_8976);
nor U13852 (N_13852,N_7393,N_10121);
and U13853 (N_13853,N_6702,N_8030);
nor U13854 (N_13854,N_11819,N_12358);
nor U13855 (N_13855,N_12229,N_10455);
nor U13856 (N_13856,N_6868,N_8358);
and U13857 (N_13857,N_10054,N_6505);
or U13858 (N_13858,N_9466,N_10345);
nand U13859 (N_13859,N_11932,N_11389);
nand U13860 (N_13860,N_7890,N_11455);
and U13861 (N_13861,N_10539,N_7921);
nor U13862 (N_13862,N_6703,N_7868);
nor U13863 (N_13863,N_10124,N_10208);
and U13864 (N_13864,N_6836,N_10759);
nor U13865 (N_13865,N_12176,N_10312);
nand U13866 (N_13866,N_7384,N_9722);
nand U13867 (N_13867,N_8615,N_7242);
or U13868 (N_13868,N_10459,N_9907);
or U13869 (N_13869,N_10770,N_8302);
or U13870 (N_13870,N_8734,N_11222);
xor U13871 (N_13871,N_11168,N_9908);
and U13872 (N_13872,N_9952,N_12095);
nor U13873 (N_13873,N_10587,N_7344);
nor U13874 (N_13874,N_7580,N_8688);
nor U13875 (N_13875,N_10801,N_7498);
and U13876 (N_13876,N_11353,N_10482);
or U13877 (N_13877,N_9880,N_8488);
nor U13878 (N_13878,N_10944,N_10513);
nor U13879 (N_13879,N_7815,N_9130);
or U13880 (N_13880,N_9793,N_8459);
nand U13881 (N_13881,N_9250,N_10773);
and U13882 (N_13882,N_9345,N_7398);
xnor U13883 (N_13883,N_9186,N_11868);
nor U13884 (N_13884,N_7319,N_6867);
and U13885 (N_13885,N_10434,N_8805);
or U13886 (N_13886,N_7548,N_6570);
nand U13887 (N_13887,N_6945,N_11907);
and U13888 (N_13888,N_10065,N_10788);
and U13889 (N_13889,N_12330,N_9682);
and U13890 (N_13890,N_8433,N_10002);
or U13891 (N_13891,N_6712,N_10142);
or U13892 (N_13892,N_8374,N_11705);
nand U13893 (N_13893,N_7900,N_10236);
and U13894 (N_13894,N_7556,N_7263);
nor U13895 (N_13895,N_8364,N_10625);
or U13896 (N_13896,N_12024,N_11144);
nor U13897 (N_13897,N_8660,N_8517);
or U13898 (N_13898,N_10620,N_8166);
and U13899 (N_13899,N_9530,N_6630);
nand U13900 (N_13900,N_6623,N_7376);
nor U13901 (N_13901,N_9805,N_9004);
xnor U13902 (N_13902,N_9714,N_9995);
nand U13903 (N_13903,N_9333,N_9579);
and U13904 (N_13904,N_11091,N_12316);
and U13905 (N_13905,N_7888,N_6984);
or U13906 (N_13906,N_8158,N_7090);
nand U13907 (N_13907,N_6759,N_8087);
nor U13908 (N_13908,N_9532,N_8630);
and U13909 (N_13909,N_6659,N_11545);
and U13910 (N_13910,N_9654,N_6383);
xnor U13911 (N_13911,N_7460,N_12345);
nand U13912 (N_13912,N_11600,N_7839);
nand U13913 (N_13913,N_11553,N_7472);
and U13914 (N_13914,N_10277,N_11887);
xor U13915 (N_13915,N_10660,N_6723);
nor U13916 (N_13916,N_7583,N_8042);
nor U13917 (N_13917,N_6971,N_12069);
and U13918 (N_13918,N_8035,N_10109);
or U13919 (N_13919,N_8887,N_9449);
or U13920 (N_13920,N_10064,N_11608);
or U13921 (N_13921,N_7951,N_11773);
or U13922 (N_13922,N_7158,N_9767);
or U13923 (N_13923,N_10690,N_7617);
xor U13924 (N_13924,N_10443,N_9344);
and U13925 (N_13925,N_9873,N_6901);
nand U13926 (N_13926,N_10179,N_8438);
and U13927 (N_13927,N_12073,N_8135);
or U13928 (N_13928,N_6870,N_8838);
nand U13929 (N_13929,N_7202,N_12315);
nor U13930 (N_13930,N_9928,N_9791);
and U13931 (N_13931,N_9459,N_8477);
nor U13932 (N_13932,N_9706,N_9084);
nor U13933 (N_13933,N_11332,N_11058);
nand U13934 (N_13934,N_6798,N_7307);
nor U13935 (N_13935,N_11357,N_9718);
nand U13936 (N_13936,N_7803,N_9143);
nand U13937 (N_13937,N_11799,N_7907);
nand U13938 (N_13938,N_6606,N_8164);
and U13939 (N_13939,N_9284,N_10703);
and U13940 (N_13940,N_11486,N_10831);
nand U13941 (N_13941,N_9965,N_11795);
and U13942 (N_13942,N_8327,N_7481);
or U13943 (N_13943,N_7784,N_10492);
and U13944 (N_13944,N_12326,N_10536);
nor U13945 (N_13945,N_11855,N_7712);
nor U13946 (N_13946,N_9946,N_6738);
and U13947 (N_13947,N_10574,N_6665);
and U13948 (N_13948,N_11694,N_6934);
or U13949 (N_13949,N_10931,N_12239);
nand U13950 (N_13950,N_9391,N_7730);
or U13951 (N_13951,N_9762,N_10343);
or U13952 (N_13952,N_8426,N_8878);
nand U13953 (N_13953,N_7407,N_7721);
and U13954 (N_13954,N_7517,N_8965);
and U13955 (N_13955,N_10239,N_6565);
nor U13956 (N_13956,N_11837,N_9770);
xor U13957 (N_13957,N_11088,N_9202);
or U13958 (N_13958,N_12120,N_12338);
and U13959 (N_13959,N_12056,N_8482);
xnor U13960 (N_13960,N_11928,N_12053);
and U13961 (N_13961,N_12192,N_9795);
or U13962 (N_13962,N_7304,N_6507);
nor U13963 (N_13963,N_8395,N_11736);
or U13964 (N_13964,N_7526,N_11401);
nand U13965 (N_13965,N_11665,N_12475);
and U13966 (N_13966,N_11690,N_10044);
xnor U13967 (N_13967,N_9368,N_10830);
nand U13968 (N_13968,N_8479,N_9604);
xnor U13969 (N_13969,N_10072,N_11136);
or U13970 (N_13970,N_11763,N_7728);
nor U13971 (N_13971,N_11134,N_8626);
nand U13972 (N_13972,N_6975,N_8142);
or U13973 (N_13973,N_10796,N_6924);
or U13974 (N_13974,N_7854,N_10247);
nor U13975 (N_13975,N_6731,N_10354);
nor U13976 (N_13976,N_7523,N_10053);
nor U13977 (N_13977,N_7152,N_11415);
and U13978 (N_13978,N_10113,N_11012);
or U13979 (N_13979,N_9788,N_10774);
nor U13980 (N_13980,N_11862,N_9237);
and U13981 (N_13981,N_9023,N_7684);
nor U13982 (N_13982,N_9666,N_7722);
or U13983 (N_13983,N_11749,N_9497);
nand U13984 (N_13984,N_11510,N_6654);
or U13985 (N_13985,N_6754,N_6387);
nor U13986 (N_13986,N_8385,N_6316);
nor U13987 (N_13987,N_12369,N_9451);
nor U13988 (N_13988,N_9342,N_7060);
or U13989 (N_13989,N_10845,N_11251);
nand U13990 (N_13990,N_9281,N_6710);
and U13991 (N_13991,N_8768,N_10899);
nand U13992 (N_13992,N_8297,N_7324);
nor U13993 (N_13993,N_6818,N_12098);
and U13994 (N_13994,N_11376,N_8127);
nor U13995 (N_13995,N_8475,N_8888);
nand U13996 (N_13996,N_9909,N_11989);
and U13997 (N_13997,N_10504,N_11815);
xor U13998 (N_13998,N_11836,N_11740);
nand U13999 (N_13999,N_7957,N_11081);
nor U14000 (N_14000,N_11632,N_11232);
or U14001 (N_14001,N_12291,N_8186);
nand U14002 (N_14002,N_7701,N_10753);
or U14003 (N_14003,N_7773,N_10169);
nor U14004 (N_14004,N_11271,N_11696);
nand U14005 (N_14005,N_9897,N_10749);
nand U14006 (N_14006,N_6419,N_9026);
xor U14007 (N_14007,N_11416,N_7452);
and U14008 (N_14008,N_9569,N_9606);
nand U14009 (N_14009,N_10185,N_6480);
and U14010 (N_14010,N_8864,N_6283);
and U14011 (N_14011,N_6809,N_9067);
and U14012 (N_14012,N_11463,N_10437);
and U14013 (N_14013,N_7153,N_11867);
nand U14014 (N_14014,N_10866,N_7650);
xor U14015 (N_14015,N_6837,N_12067);
nand U14016 (N_14016,N_12389,N_7211);
nand U14017 (N_14017,N_8658,N_10240);
nand U14018 (N_14018,N_8445,N_9978);
or U14019 (N_14019,N_8518,N_6982);
nor U14020 (N_14020,N_7479,N_11290);
and U14021 (N_14021,N_12126,N_9289);
or U14022 (N_14022,N_10814,N_8021);
nand U14023 (N_14023,N_9268,N_11205);
and U14024 (N_14024,N_12088,N_10705);
or U14025 (N_14025,N_7186,N_11502);
xor U14026 (N_14026,N_12331,N_6519);
or U14027 (N_14027,N_9060,N_10204);
nand U14028 (N_14028,N_11391,N_12162);
xnor U14029 (N_14029,N_8063,N_6690);
nor U14030 (N_14030,N_6504,N_6310);
and U14031 (N_14031,N_8250,N_7679);
and U14032 (N_14032,N_7172,N_10949);
nor U14033 (N_14033,N_6844,N_11807);
nor U14034 (N_14034,N_12084,N_8712);
and U14035 (N_14035,N_7719,N_6931);
nor U14036 (N_14036,N_11771,N_9801);
nor U14037 (N_14037,N_10061,N_10533);
and U14038 (N_14038,N_12087,N_11591);
xnor U14039 (N_14039,N_10718,N_6406);
and U14040 (N_14040,N_12130,N_8192);
or U14041 (N_14041,N_11565,N_8465);
and U14042 (N_14042,N_7434,N_8588);
xor U14043 (N_14043,N_11437,N_9554);
and U14044 (N_14044,N_10221,N_6776);
nand U14045 (N_14045,N_12123,N_11588);
nor U14046 (N_14046,N_6951,N_9945);
nand U14047 (N_14047,N_7295,N_10798);
nand U14048 (N_14048,N_6302,N_8853);
nand U14049 (N_14049,N_7473,N_7265);
xor U14050 (N_14050,N_9150,N_8526);
or U14051 (N_14051,N_10628,N_9782);
or U14052 (N_14052,N_12442,N_10309);
and U14053 (N_14053,N_12385,N_11424);
xor U14054 (N_14054,N_7802,N_7508);
and U14055 (N_14055,N_9719,N_7742);
nand U14056 (N_14056,N_11324,N_8824);
and U14057 (N_14057,N_10372,N_10875);
nor U14058 (N_14058,N_6452,N_8758);
and U14059 (N_14059,N_8404,N_6743);
and U14060 (N_14060,N_8559,N_10659);
or U14061 (N_14061,N_9114,N_11473);
nor U14062 (N_14062,N_6706,N_11496);
or U14063 (N_14063,N_11319,N_12324);
or U14064 (N_14064,N_12001,N_8004);
nor U14065 (N_14065,N_11666,N_7970);
nor U14066 (N_14066,N_7941,N_10241);
nand U14067 (N_14067,N_10305,N_7092);
nand U14068 (N_14068,N_7746,N_8330);
or U14069 (N_14069,N_12234,N_8335);
nor U14070 (N_14070,N_6366,N_6359);
nand U14071 (N_14071,N_12240,N_9692);
nand U14072 (N_14072,N_8133,N_9926);
nand U14073 (N_14073,N_6839,N_6401);
or U14074 (N_14074,N_9197,N_6295);
nor U14075 (N_14075,N_12145,N_8643);
or U14076 (N_14076,N_8448,N_8371);
and U14077 (N_14077,N_7104,N_9346);
xnor U14078 (N_14078,N_6321,N_9546);
nand U14079 (N_14079,N_8306,N_12167);
and U14080 (N_14080,N_7128,N_12065);
nor U14081 (N_14081,N_9725,N_9235);
nand U14082 (N_14082,N_10653,N_9812);
or U14083 (N_14083,N_6440,N_6803);
nand U14084 (N_14084,N_8756,N_6658);
xor U14085 (N_14085,N_6720,N_8759);
nor U14086 (N_14086,N_8951,N_7859);
and U14087 (N_14087,N_10932,N_8822);
and U14088 (N_14088,N_9977,N_7081);
xnor U14089 (N_14089,N_8456,N_11476);
xnor U14090 (N_14090,N_10261,N_6356);
or U14091 (N_14091,N_7133,N_6428);
and U14092 (N_14092,N_11877,N_9668);
nor U14093 (N_14093,N_9433,N_11568);
and U14094 (N_14094,N_10993,N_10278);
or U14095 (N_14095,N_10405,N_7794);
or U14096 (N_14096,N_11383,N_10606);
nand U14097 (N_14097,N_6884,N_8687);
nand U14098 (N_14098,N_9409,N_8068);
xnor U14099 (N_14099,N_9302,N_7131);
nor U14100 (N_14100,N_9775,N_11745);
or U14101 (N_14101,N_7589,N_9439);
or U14102 (N_14102,N_12264,N_11300);
nand U14103 (N_14103,N_12497,N_6345);
nand U14104 (N_14104,N_11853,N_11988);
nand U14105 (N_14105,N_6352,N_6579);
and U14106 (N_14106,N_11906,N_9152);
and U14107 (N_14107,N_11087,N_10465);
xnor U14108 (N_14108,N_9526,N_9540);
nor U14109 (N_14109,N_10401,N_6353);
nor U14110 (N_14110,N_8328,N_10135);
and U14111 (N_14111,N_7305,N_7904);
or U14112 (N_14112,N_9786,N_10280);
and U14113 (N_14113,N_11575,N_9686);
and U14114 (N_14114,N_11457,N_6576);
nand U14115 (N_14115,N_11450,N_10548);
or U14116 (N_14116,N_11146,N_11497);
nor U14117 (N_14117,N_8101,N_6761);
nor U14118 (N_14118,N_9460,N_7282);
nor U14119 (N_14119,N_11829,N_11894);
or U14120 (N_14120,N_9940,N_7402);
nor U14121 (N_14121,N_6755,N_8453);
nor U14122 (N_14122,N_12441,N_9022);
or U14123 (N_14123,N_11386,N_11347);
nand U14124 (N_14124,N_10324,N_8267);
and U14125 (N_14125,N_9910,N_8857);
nand U14126 (N_14126,N_10357,N_10162);
nor U14127 (N_14127,N_7984,N_9982);
and U14128 (N_14128,N_9469,N_7867);
or U14129 (N_14129,N_6639,N_6471);
and U14130 (N_14130,N_7828,N_11838);
xnor U14131 (N_14131,N_7720,N_10359);
and U14132 (N_14132,N_9075,N_9736);
nor U14133 (N_14133,N_11368,N_9200);
and U14134 (N_14134,N_8443,N_12290);
and U14135 (N_14135,N_11693,N_9779);
nand U14136 (N_14136,N_7981,N_8872);
nand U14137 (N_14137,N_8012,N_12075);
xor U14138 (N_14138,N_9816,N_9315);
and U14139 (N_14139,N_8230,N_7696);
or U14140 (N_14140,N_6655,N_7751);
and U14141 (N_14141,N_9395,N_11077);
nand U14142 (N_14142,N_6372,N_8096);
nand U14143 (N_14143,N_12427,N_11962);
or U14144 (N_14144,N_9062,N_9858);
nand U14145 (N_14145,N_12197,N_10457);
and U14146 (N_14146,N_6887,N_9288);
or U14147 (N_14147,N_9024,N_7164);
nand U14148 (N_14148,N_11242,N_8883);
nand U14149 (N_14149,N_9404,N_10613);
nor U14150 (N_14150,N_10049,N_12236);
or U14151 (N_14151,N_6462,N_7870);
or U14152 (N_14152,N_6727,N_7648);
nor U14153 (N_14153,N_12361,N_6667);
nor U14154 (N_14154,N_6354,N_11583);
or U14155 (N_14155,N_12273,N_8797);
nor U14156 (N_14156,N_9525,N_11127);
nand U14157 (N_14157,N_8711,N_12137);
or U14158 (N_14158,N_8424,N_7363);
xor U14159 (N_14159,N_11743,N_8856);
nand U14160 (N_14160,N_7816,N_10003);
and U14161 (N_14161,N_6559,N_7048);
and U14162 (N_14162,N_7476,N_8546);
nor U14163 (N_14163,N_9358,N_9357);
xnor U14164 (N_14164,N_6263,N_10231);
nand U14165 (N_14165,N_9846,N_7286);
or U14166 (N_14166,N_10367,N_7611);
and U14167 (N_14167,N_11985,N_6560);
and U14168 (N_14168,N_11501,N_9389);
or U14169 (N_14169,N_6332,N_10965);
and U14170 (N_14170,N_6319,N_11930);
nand U14171 (N_14171,N_12247,N_6925);
or U14172 (N_14172,N_11105,N_9305);
and U14173 (N_14173,N_8754,N_9211);
and U14174 (N_14174,N_8993,N_11609);
nand U14175 (N_14175,N_9527,N_6465);
or U14176 (N_14176,N_9932,N_11631);
nor U14177 (N_14177,N_7766,N_8791);
nand U14178 (N_14178,N_10084,N_10580);
nor U14179 (N_14179,N_12249,N_11612);
or U14180 (N_14180,N_8184,N_6863);
or U14181 (N_14181,N_6525,N_10255);
or U14182 (N_14182,N_11172,N_6664);
and U14183 (N_14183,N_11122,N_6581);
or U14184 (N_14184,N_11661,N_12304);
nor U14185 (N_14185,N_7230,N_8152);
nor U14186 (N_14186,N_10957,N_12251);
and U14187 (N_14187,N_9803,N_6331);
and U14188 (N_14188,N_7518,N_11570);
and U14189 (N_14189,N_7161,N_10512);
nand U14190 (N_14190,N_10737,N_7127);
nand U14191 (N_14191,N_7934,N_7735);
nand U14192 (N_14192,N_10616,N_7007);
and U14193 (N_14193,N_8926,N_7958);
nor U14194 (N_14194,N_10365,N_7995);
nand U14195 (N_14195,N_8835,N_6382);
nand U14196 (N_14196,N_7494,N_6774);
nor U14197 (N_14197,N_6877,N_9402);
nor U14198 (N_14198,N_11313,N_10873);
or U14199 (N_14199,N_11936,N_11069);
nand U14200 (N_14200,N_9857,N_11013);
nor U14201 (N_14201,N_10921,N_8966);
nand U14202 (N_14202,N_10551,N_11590);
nand U14203 (N_14203,N_6370,N_6697);
or U14204 (N_14204,N_11517,N_12495);
and U14205 (N_14205,N_7069,N_7786);
and U14206 (N_14206,N_10449,N_10947);
nand U14207 (N_14207,N_8381,N_12108);
xor U14208 (N_14208,N_12134,N_6907);
and U14209 (N_14209,N_10100,N_10384);
nor U14210 (N_14210,N_10106,N_9081);
nor U14211 (N_14211,N_7997,N_10313);
and U14212 (N_14212,N_10268,N_9334);
nand U14213 (N_14213,N_12443,N_9987);
or U14214 (N_14214,N_11340,N_7488);
nand U14215 (N_14215,N_10745,N_10874);
xor U14216 (N_14216,N_10889,N_8388);
and U14217 (N_14217,N_11169,N_9484);
or U14218 (N_14218,N_11209,N_10776);
nor U14219 (N_14219,N_11231,N_10152);
nor U14220 (N_14220,N_12171,N_6687);
nand U14221 (N_14221,N_9307,N_11759);
and U14222 (N_14222,N_10725,N_9405);
or U14223 (N_14223,N_12437,N_7382);
xor U14224 (N_14224,N_8023,N_8844);
xnor U14225 (N_14225,N_8648,N_7537);
xnor U14226 (N_14226,N_10884,N_10063);
or U14227 (N_14227,N_9768,N_9835);
xor U14228 (N_14228,N_6696,N_9711);
and U14229 (N_14229,N_8845,N_12346);
nor U14230 (N_14230,N_9049,N_8489);
or U14231 (N_14231,N_10370,N_8973);
xnor U14232 (N_14232,N_11082,N_10633);
xnor U14233 (N_14233,N_6842,N_6489);
nor U14234 (N_14234,N_9495,N_8975);
nor U14235 (N_14235,N_9082,N_8507);
nor U14236 (N_14236,N_8935,N_11113);
or U14237 (N_14237,N_8217,N_6337);
and U14238 (N_14238,N_9167,N_8743);
nand U14239 (N_14239,N_7198,N_12187);
or U14240 (N_14240,N_8836,N_11131);
xor U14241 (N_14241,N_8466,N_8948);
nor U14242 (N_14242,N_12013,N_8934);
xnor U14243 (N_14243,N_6851,N_10433);
nand U14244 (N_14244,N_9562,N_9937);
nand U14245 (N_14245,N_10477,N_8880);
or U14246 (N_14246,N_11108,N_11043);
and U14247 (N_14247,N_8818,N_8245);
and U14248 (N_14248,N_8387,N_6728);
and U14249 (N_14249,N_7147,N_8379);
or U14250 (N_14250,N_9070,N_6841);
or U14251 (N_14251,N_9595,N_12411);
and U14252 (N_14252,N_8288,N_7654);
and U14253 (N_14253,N_9710,N_11668);
nand U14254 (N_14254,N_7138,N_7843);
and U14255 (N_14255,N_6959,N_12274);
and U14256 (N_14256,N_6483,N_9509);
nor U14257 (N_14257,N_12420,N_9780);
or U14258 (N_14258,N_6643,N_8316);
or U14259 (N_14259,N_12283,N_10593);
xnor U14260 (N_14260,N_8051,N_6815);
and U14261 (N_14261,N_8931,N_9123);
xnor U14262 (N_14262,N_8070,N_9316);
nand U14263 (N_14263,N_6582,N_11709);
nor U14264 (N_14264,N_7640,N_8190);
nand U14265 (N_14265,N_6807,N_10110);
and U14266 (N_14266,N_11337,N_7423);
or U14267 (N_14267,N_10023,N_7688);
or U14268 (N_14268,N_7916,N_8044);
nand U14269 (N_14269,N_11954,N_9565);
and U14270 (N_14270,N_8920,N_8134);
nor U14271 (N_14271,N_10882,N_9247);
nand U14272 (N_14272,N_6522,N_7937);
nor U14273 (N_14273,N_9794,N_6557);
nand U14274 (N_14274,N_7928,N_11321);
nor U14275 (N_14275,N_7491,N_9534);
nor U14276 (N_14276,N_6804,N_6933);
nor U14277 (N_14277,N_9658,N_7774);
xor U14278 (N_14278,N_8728,N_8508);
xnor U14279 (N_14279,N_7829,N_10713);
nor U14280 (N_14280,N_9428,N_7819);
nor U14281 (N_14281,N_10823,N_12323);
nor U14282 (N_14282,N_8652,N_9747);
and U14283 (N_14283,N_8111,N_6820);
xnor U14284 (N_14284,N_8896,N_12230);
and U14285 (N_14285,N_9117,N_6351);
nor U14286 (N_14286,N_6966,N_12435);
nor U14287 (N_14287,N_6426,N_11550);
and U14288 (N_14288,N_11044,N_9720);
nand U14289 (N_14289,N_6668,N_10058);
or U14290 (N_14290,N_6600,N_11139);
nand U14291 (N_14291,N_9589,N_6255);
nand U14292 (N_14292,N_9724,N_7525);
nor U14293 (N_14293,N_9813,N_7660);
xnor U14294 (N_14294,N_7812,N_11090);
and U14295 (N_14295,N_6760,N_9435);
and U14296 (N_14296,N_10585,N_9599);
and U14297 (N_14297,N_6350,N_12210);
xor U14298 (N_14298,N_6371,N_10597);
nand U14299 (N_14299,N_6274,N_11786);
xnor U14300 (N_14300,N_8747,N_6317);
nand U14301 (N_14301,N_8504,N_8940);
and U14302 (N_14302,N_8055,N_11367);
nor U14303 (N_14303,N_10811,N_9864);
or U14304 (N_14304,N_10175,N_10848);
and U14305 (N_14305,N_11306,N_10150);
nand U14306 (N_14306,N_8082,N_10137);
or U14307 (N_14307,N_8891,N_7187);
or U14308 (N_14308,N_10398,N_10812);
nand U14309 (N_14309,N_9061,N_9966);
xnor U14310 (N_14310,N_9649,N_8610);
nand U14311 (N_14311,N_7350,N_10195);
nor U14312 (N_14312,N_7364,N_10389);
nand U14313 (N_14313,N_11049,N_11411);
and U14314 (N_14314,N_10743,N_11605);
nand U14315 (N_14315,N_8151,N_7077);
or U14316 (N_14316,N_6861,N_11174);
nor U14317 (N_14317,N_10826,N_7180);
xor U14318 (N_14318,N_6265,N_11692);
or U14319 (N_14319,N_7047,N_11722);
or U14320 (N_14320,N_9377,N_8303);
or U14321 (N_14321,N_6461,N_9806);
xor U14322 (N_14322,N_7764,N_11687);
or U14323 (N_14323,N_11735,N_11695);
and U14324 (N_14324,N_11947,N_11551);
nand U14325 (N_14325,N_8874,N_7692);
and U14326 (N_14326,N_11388,N_8943);
and U14327 (N_14327,N_7348,N_11841);
xor U14328 (N_14328,N_7942,N_11050);
or U14329 (N_14329,N_9432,N_7973);
or U14330 (N_14330,N_11163,N_8941);
or U14331 (N_14331,N_10929,N_10706);
nor U14332 (N_14332,N_9773,N_11627);
nand U14333 (N_14333,N_7863,N_10636);
or U14334 (N_14334,N_10217,N_6843);
nand U14335 (N_14335,N_7383,N_7072);
and U14336 (N_14336,N_10984,N_10432);
or U14337 (N_14337,N_7825,N_12146);
xnor U14338 (N_14338,N_10036,N_8741);
nor U14339 (N_14339,N_12190,N_8221);
and U14340 (N_14340,N_12048,N_10800);
and U14341 (N_14341,N_10012,N_12318);
nor U14342 (N_14342,N_7173,N_10471);
or U14343 (N_14343,N_11756,N_9541);
nor U14344 (N_14344,N_9195,N_8415);
nand U14345 (N_14345,N_10671,N_7335);
nand U14346 (N_14346,N_8790,N_7771);
or U14347 (N_14347,N_8764,N_10962);
and U14348 (N_14348,N_8139,N_8961);
or U14349 (N_14349,N_7996,N_11252);
nor U14350 (N_14350,N_11784,N_10645);
nand U14351 (N_14351,N_8994,N_11098);
nor U14352 (N_14352,N_8049,N_8693);
or U14353 (N_14353,N_10257,N_11482);
or U14354 (N_14354,N_7702,N_10122);
and U14355 (N_14355,N_10440,N_12288);
nor U14356 (N_14356,N_12148,N_6686);
nor U14357 (N_14357,N_8739,N_8528);
nor U14358 (N_14358,N_7883,N_10675);
xnor U14359 (N_14359,N_8084,N_9412);
and U14360 (N_14360,N_12219,N_7449);
nor U14361 (N_14361,N_12356,N_9441);
and U14362 (N_14362,N_9071,N_9955);
xnor U14363 (N_14363,N_10004,N_10815);
nor U14364 (N_14364,N_11221,N_8337);
nor U14365 (N_14365,N_7535,N_8936);
or U14366 (N_14366,N_10171,N_9564);
nor U14367 (N_14367,N_7544,N_6699);
and U14368 (N_14368,N_12388,N_11875);
and U14369 (N_14369,N_7130,N_7765);
and U14370 (N_14370,N_9809,N_11285);
and U14371 (N_14371,N_11053,N_11801);
nor U14372 (N_14372,N_10141,N_11653);
and U14373 (N_14373,N_8968,N_11716);
nand U14374 (N_14374,N_10226,N_7146);
nand U14375 (N_14375,N_11056,N_12248);
nand U14376 (N_14376,N_6903,N_8331);
nand U14377 (N_14377,N_8998,N_6952);
and U14378 (N_14378,N_11438,N_9273);
and U14379 (N_14379,N_7519,N_11500);
or U14380 (N_14380,N_7553,N_11941);
or U14381 (N_14381,N_7232,N_9015);
or U14382 (N_14382,N_10682,N_7269);
and U14383 (N_14383,N_9690,N_7424);
nand U14384 (N_14384,N_6399,N_12339);
nor U14385 (N_14385,N_9465,N_7667);
nor U14386 (N_14386,N_9283,N_7889);
or U14387 (N_14387,N_6312,N_11644);
and U14388 (N_14388,N_6429,N_8449);
and U14389 (N_14389,N_11045,N_9633);
nor U14390 (N_14390,N_11270,N_10252);
nand U14391 (N_14391,N_10350,N_10377);
xor U14392 (N_14392,N_8155,N_7540);
nor U14393 (N_14393,N_8422,N_8452);
nand U14394 (N_14394,N_7497,N_7806);
and U14395 (N_14395,N_11372,N_7898);
nor U14396 (N_14396,N_8553,N_11240);
nor U14397 (N_14397,N_7283,N_11277);
xnor U14398 (N_14398,N_8480,N_9133);
nor U14399 (N_14399,N_10808,N_8450);
and U14400 (N_14400,N_11035,N_11284);
xor U14401 (N_14401,N_10331,N_8802);
and U14402 (N_14402,N_12381,N_10371);
nand U14403 (N_14403,N_8240,N_8953);
xor U14404 (N_14404,N_9764,N_7988);
or U14405 (N_14405,N_12317,N_6786);
nor U14406 (N_14406,N_11183,N_7199);
nor U14407 (N_14407,N_8629,N_8501);
nor U14408 (N_14408,N_7554,N_7334);
and U14409 (N_14409,N_6306,N_11673);
and U14410 (N_14410,N_7119,N_8954);
xor U14411 (N_14411,N_10851,N_7108);
and U14412 (N_14412,N_8389,N_10677);
or U14413 (N_14413,N_10832,N_8525);
nand U14414 (N_14414,N_10485,N_7125);
xnor U14415 (N_14415,N_10037,N_7082);
or U14416 (N_14416,N_7592,N_8536);
nand U14417 (N_14417,N_11670,N_9089);
or U14418 (N_14418,N_7531,N_12168);
nand U14419 (N_14419,N_8952,N_8833);
and U14420 (N_14420,N_7675,N_10017);
xnor U14421 (N_14421,N_9258,N_6342);
and U14422 (N_14422,N_6378,N_12303);
nand U14423 (N_14423,N_12049,N_9102);
nor U14424 (N_14424,N_11052,N_10071);
or U14425 (N_14425,N_11173,N_9069);
nor U14426 (N_14426,N_11104,N_11148);
and U14427 (N_14427,N_8568,N_6678);
nand U14428 (N_14428,N_6891,N_10101);
nand U14429 (N_14429,N_12386,N_6904);
xnor U14430 (N_14430,N_10933,N_9500);
or U14431 (N_14431,N_9680,N_10178);
and U14432 (N_14432,N_8175,N_9185);
and U14433 (N_14433,N_11274,N_10511);
nor U14434 (N_14434,N_12019,N_9058);
nand U14435 (N_14435,N_7990,N_7194);
nor U14436 (N_14436,N_10853,N_10093);
nand U14437 (N_14437,N_9318,N_9834);
and U14438 (N_14438,N_7419,N_8182);
nor U14439 (N_14439,N_9636,N_6347);
and U14440 (N_14440,N_11487,N_8283);
nor U14441 (N_14441,N_7849,N_10654);
xnor U14442 (N_14442,N_9999,N_10842);
or U14443 (N_14443,N_10658,N_8812);
and U14444 (N_14444,N_7118,N_9406);
or U14445 (N_14445,N_12218,N_6438);
and U14446 (N_14446,N_10953,N_9296);
and U14447 (N_14447,N_8565,N_10738);
and U14448 (N_14448,N_6647,N_8744);
or U14449 (N_14449,N_11821,N_10872);
and U14450 (N_14450,N_11499,N_8587);
xnor U14451 (N_14451,N_10981,N_10676);
nand U14452 (N_14452,N_9576,N_6763);
xnor U14453 (N_14453,N_9039,N_7288);
or U14454 (N_14454,N_6821,N_8437);
nor U14455 (N_14455,N_9487,N_6476);
nand U14456 (N_14456,N_7833,N_11982);
or U14457 (N_14457,N_7416,N_10333);
and U14458 (N_14458,N_9120,N_10785);
xor U14459 (N_14459,N_12193,N_8691);
nor U14460 (N_14460,N_11378,N_7824);
and U14461 (N_14461,N_10041,N_9947);
xnor U14462 (N_14462,N_9587,N_6883);
nor U14463 (N_14463,N_7020,N_8319);
nand U14464 (N_14464,N_8800,N_6850);
nor U14465 (N_14465,N_10205,N_9789);
nor U14466 (N_14466,N_10761,N_10604);
nor U14467 (N_14467,N_9660,N_11488);
nor U14468 (N_14468,N_7264,N_12416);
and U14469 (N_14469,N_11760,N_7136);
and U14470 (N_14470,N_7850,N_11165);
or U14471 (N_14471,N_6947,N_8839);
and U14472 (N_14472,N_8386,N_10040);
nor U14473 (N_14473,N_11119,N_7694);
nor U14474 (N_14474,N_6736,N_11428);
and U14475 (N_14475,N_10346,N_11392);
and U14476 (N_14476,N_11308,N_10868);
and U14477 (N_14477,N_7098,N_7925);
nor U14478 (N_14478,N_12343,N_12297);
or U14479 (N_14479,N_7820,N_8996);
nor U14480 (N_14480,N_11489,N_8026);
and U14481 (N_14481,N_11187,N_8584);
nor U14482 (N_14482,N_6333,N_9563);
nand U14483 (N_14483,N_9184,N_7783);
or U14484 (N_14484,N_9323,N_10025);
and U14485 (N_14485,N_6305,N_7982);
or U14486 (N_14486,N_7182,N_10197);
and U14487 (N_14487,N_9771,N_8860);
nand U14488 (N_14488,N_11718,N_8490);
xnor U14489 (N_14489,N_11702,N_11746);
and U14490 (N_14490,N_11711,N_9667);
or U14491 (N_14491,N_9951,N_7262);
or U14492 (N_14492,N_11294,N_11109);
xor U14493 (N_14493,N_7913,N_6268);
and U14494 (N_14494,N_8129,N_11116);
xor U14495 (N_14495,N_8982,N_7848);
xor U14496 (N_14496,N_12196,N_7962);
and U14497 (N_14497,N_9697,N_10863);
or U14498 (N_14498,N_11886,N_11233);
or U14499 (N_14499,N_8914,N_9646);
nand U14500 (N_14500,N_11017,N_6413);
and U14501 (N_14501,N_11162,N_8918);
nand U14502 (N_14502,N_11614,N_8990);
nor U14503 (N_14503,N_11330,N_12008);
or U14504 (N_14504,N_12347,N_7718);
nand U14505 (N_14505,N_7181,N_7352);
or U14506 (N_14506,N_8656,N_10732);
and U14507 (N_14507,N_8780,N_8625);
or U14508 (N_14508,N_11537,N_9571);
nor U14509 (N_14509,N_10781,N_9468);
or U14510 (N_14510,N_10263,N_10010);
nand U14511 (N_14511,N_9962,N_9670);
and U14512 (N_14512,N_8870,N_7284);
nor U14513 (N_14513,N_10409,N_8577);
and U14514 (N_14514,N_9842,N_10556);
nor U14515 (N_14515,N_11303,N_10246);
and U14516 (N_14516,N_11307,N_11770);
and U14517 (N_14517,N_11398,N_10130);
and U14518 (N_14518,N_11467,N_8977);
and U14519 (N_14519,N_12160,N_9905);
and U14520 (N_14520,N_8510,N_8392);
nor U14521 (N_14521,N_7987,N_9267);
and U14522 (N_14522,N_6391,N_9335);
nor U14523 (N_14523,N_7598,N_7567);
nand U14524 (N_14524,N_9783,N_10201);
and U14525 (N_14525,N_7652,N_7000);
nand U14526 (N_14526,N_10486,N_7642);
nand U14527 (N_14527,N_11534,N_9159);
or U14528 (N_14528,N_6998,N_12030);
nand U14529 (N_14529,N_8731,N_8343);
nand U14530 (N_14530,N_6918,N_6905);
xor U14531 (N_14531,N_10956,N_9958);
xor U14532 (N_14532,N_9927,N_8473);
or U14533 (N_14533,N_7574,N_9017);
and U14534 (N_14534,N_11558,N_12225);
nand U14535 (N_14535,N_8694,N_11151);
nand U14536 (N_14536,N_11288,N_7070);
and U14537 (N_14537,N_10772,N_9729);
and U14538 (N_14538,N_6633,N_7956);
nand U14539 (N_14539,N_11456,N_8207);
and U14540 (N_14540,N_10087,N_10393);
or U14541 (N_14541,N_8032,N_9677);
nand U14542 (N_14542,N_8689,N_10161);
nor U14543 (N_14543,N_8841,N_8290);
or U14544 (N_14544,N_11264,N_7330);
or U14545 (N_14545,N_8398,N_9246);
nand U14546 (N_14546,N_8578,N_6501);
nor U14547 (N_14547,N_11948,N_8714);
xor U14548 (N_14548,N_9523,N_11897);
nor U14549 (N_14549,N_7801,N_9504);
nor U14550 (N_14550,N_7447,N_7879);
and U14551 (N_14551,N_8631,N_12113);
nand U14552 (N_14552,N_9583,N_8571);
or U14553 (N_14553,N_7314,N_9104);
xnor U14554 (N_14554,N_9972,N_8317);
nand U14555 (N_14555,N_11153,N_9415);
nor U14556 (N_14556,N_7588,N_11446);
nand U14557 (N_14557,N_6787,N_10094);
nor U14558 (N_14558,N_10850,N_9744);
and U14559 (N_14559,N_8431,N_9012);
or U14560 (N_14560,N_7568,N_9239);
xor U14561 (N_14561,N_9083,N_7253);
and U14562 (N_14562,N_7732,N_12009);
nor U14563 (N_14563,N_11073,N_9331);
or U14564 (N_14564,N_10799,N_10403);
or U14565 (N_14565,N_8003,N_11420);
nor U14566 (N_14566,N_7621,N_8018);
or U14567 (N_14567,N_8483,N_8708);
nor U14568 (N_14568,N_8041,N_9472);
and U14569 (N_14569,N_7847,N_7912);
or U14570 (N_14570,N_11787,N_7267);
or U14571 (N_14571,N_10474,N_9994);
or U14572 (N_14572,N_7666,N_10519);
nor U14573 (N_14573,N_8562,N_12027);
nand U14574 (N_14574,N_7102,N_11822);
nor U14575 (N_14575,N_8602,N_10641);
nor U14576 (N_14576,N_9266,N_9622);
and U14577 (N_14577,N_9116,N_9148);
nand U14578 (N_14578,N_11513,N_7338);
or U14579 (N_14579,N_7475,N_7781);
or U14580 (N_14580,N_9643,N_6475);
nand U14581 (N_14581,N_11854,N_10503);
or U14582 (N_14582,N_10862,N_8313);
nand U14583 (N_14583,N_9970,N_8606);
nand U14584 (N_14584,N_8945,N_8174);
nand U14585 (N_14585,N_10937,N_9963);
nand U14586 (N_14586,N_7678,N_8564);
xnor U14587 (N_14587,N_6271,N_11394);
xnor U14588 (N_14588,N_8937,N_7927);
and U14589 (N_14589,N_6344,N_7714);
nor U14590 (N_14590,N_9110,N_6782);
nor U14591 (N_14591,N_12394,N_12216);
nand U14592 (N_14592,N_12034,N_8636);
or U14593 (N_14593,N_8276,N_8539);
and U14594 (N_14594,N_8971,N_6749);
or U14595 (N_14595,N_9614,N_11905);
or U14596 (N_14596,N_11364,N_10750);
nand U14597 (N_14597,N_8406,N_6373);
and U14598 (N_14598,N_8199,N_10413);
and U14599 (N_14599,N_7037,N_8591);
nand U14600 (N_14600,N_10196,N_11885);
and U14601 (N_14601,N_11453,N_12473);
nand U14602 (N_14602,N_7188,N_7625);
and U14603 (N_14603,N_8826,N_8353);
nor U14604 (N_14604,N_7680,N_8732);
and U14605 (N_14605,N_12384,N_10980);
nand U14606 (N_14606,N_8458,N_7725);
nor U14607 (N_14607,N_9695,N_8090);
nand U14608 (N_14608,N_8467,N_9010);
nand U14609 (N_14609,N_7638,N_9634);
nor U14610 (N_14610,N_6832,N_11866);
and U14611 (N_14611,N_9944,N_11846);
nor U14612 (N_14612,N_10470,N_11346);
nor U14613 (N_14613,N_10267,N_7892);
nor U14614 (N_14614,N_9215,N_9844);
or U14615 (N_14615,N_9760,N_10119);
nand U14616 (N_14616,N_10572,N_6876);
nand U14617 (N_14617,N_11762,N_8284);
or U14618 (N_14618,N_8065,N_12209);
nand U14619 (N_14619,N_8906,N_6657);
or U14620 (N_14620,N_8904,N_7514);
nand U14621 (N_14621,N_6493,N_10266);
nor U14622 (N_14622,N_8305,N_12447);
nor U14623 (N_14623,N_7453,N_7357);
xnor U14624 (N_14624,N_12177,N_7770);
nor U14625 (N_14625,N_8736,N_8851);
and U14626 (N_14626,N_8538,N_10282);
or U14627 (N_14627,N_6552,N_11544);
or U14628 (N_14628,N_9055,N_9580);
nor U14629 (N_14629,N_6640,N_12119);
nor U14630 (N_14630,N_11804,N_8325);
nor U14631 (N_14631,N_12023,N_12121);
nand U14632 (N_14632,N_8676,N_11400);
and U14633 (N_14633,N_9373,N_8403);
nor U14634 (N_14634,N_8412,N_9919);
and U14635 (N_14635,N_8911,N_11447);
and U14636 (N_14636,N_8823,N_12456);
nand U14637 (N_14637,N_9034,N_11101);
nand U14638 (N_14638,N_12047,N_10232);
nand U14639 (N_14639,N_12410,N_7558);
or U14640 (N_14640,N_11246,N_11667);
and U14641 (N_14641,N_8569,N_11191);
xor U14642 (N_14642,N_9624,N_10244);
and U14643 (N_14643,N_12061,N_8829);
or U14644 (N_14644,N_6448,N_11751);
xor U14645 (N_14645,N_7901,N_10855);
and U14646 (N_14646,N_9694,N_11351);
and U14647 (N_14647,N_9390,N_8701);
nand U14648 (N_14648,N_10414,N_10501);
and U14649 (N_14649,N_11366,N_8757);
and U14650 (N_14650,N_9488,N_12232);
nor U14651 (N_14651,N_8195,N_8310);
nand U14652 (N_14652,N_11175,N_10047);
nor U14653 (N_14653,N_6940,N_10972);
and U14654 (N_14654,N_10516,N_7144);
nor U14655 (N_14655,N_6497,N_12158);
xnor U14656 (N_14656,N_9676,N_9054);
and U14657 (N_14657,N_7255,N_12105);
nand U14658 (N_14658,N_11286,N_8425);
nand U14659 (N_14659,N_9286,N_6563);
nand U14660 (N_14660,N_11852,N_9914);
nor U14661 (N_14661,N_6791,N_9216);
xnor U14662 (N_14662,N_7115,N_8253);
or U14663 (N_14663,N_7280,N_10552);
and U14664 (N_14664,N_9108,N_10575);
nor U14665 (N_14665,N_11046,N_12213);
and U14666 (N_14666,N_12465,N_7004);
nand U14667 (N_14667,N_6911,N_7989);
or U14668 (N_14668,N_6325,N_8022);
and U14669 (N_14669,N_8321,N_8132);
or U14670 (N_14670,N_10973,N_12367);
and U14671 (N_14671,N_7366,N_10627);
and U14672 (N_14672,N_8060,N_8540);
or U14673 (N_14673,N_6610,N_7235);
and U14674 (N_14674,N_7405,N_7628);
nor U14675 (N_14675,N_8682,N_7874);
or U14676 (N_14676,N_9172,N_12020);
or U14677 (N_14677,N_11956,N_8234);
or U14678 (N_14678,N_11681,N_12396);
xor U14679 (N_14679,N_11532,N_6527);
nor U14680 (N_14680,N_10791,N_12055);
xor U14681 (N_14681,N_6729,N_9021);
or U14682 (N_14682,N_7365,N_9000);
and U14683 (N_14683,N_10034,N_10936);
or U14684 (N_14684,N_6635,N_11531);
nor U14685 (N_14685,N_7530,N_8397);
nand U14686 (N_14686,N_6675,N_6612);
nand U14687 (N_14687,N_10203,N_10191);
nand U14688 (N_14688,N_7408,N_7524);
xnor U14689 (N_14689,N_9354,N_7856);
nor U14690 (N_14690,N_8369,N_8910);
xor U14691 (N_14691,N_11263,N_9721);
nor U14692 (N_14692,N_8724,N_12284);
or U14693 (N_14693,N_11156,N_10987);
and U14694 (N_14694,N_10335,N_10532);
nand U14695 (N_14695,N_7457,N_12349);
and U14696 (N_14696,N_7470,N_6928);
nor U14697 (N_14697,N_12036,N_9397);
nor U14698 (N_14698,N_6365,N_9730);
nor U14699 (N_14699,N_10497,N_12438);
and U14700 (N_14700,N_8608,N_8014);
or U14701 (N_14701,N_8519,N_10635);
nor U14702 (N_14702,N_8523,N_9808);
or U14703 (N_14703,N_11022,N_6439);
nand U14704 (N_14704,N_9960,N_8323);
and U14705 (N_14705,N_6838,N_6585);
nand U14706 (N_14706,N_7054,N_10294);
nor U14707 (N_14707,N_10670,N_9832);
nor U14708 (N_14708,N_11678,N_11160);
nand U14709 (N_14709,N_9625,N_12488);
or U14710 (N_14710,N_10985,N_12432);
and U14711 (N_14711,N_10425,N_9374);
xor U14712 (N_14712,N_6340,N_12474);
or U14713 (N_14713,N_9558,N_7469);
or U14714 (N_14714,N_9222,N_10468);
and U14715 (N_14715,N_7630,N_6364);
and U14716 (N_14716,N_10601,N_8057);
and U14717 (N_14717,N_6425,N_9922);
and U14718 (N_14718,N_9096,N_6510);
and U14719 (N_14719,N_10783,N_8298);
nor U14720 (N_14720,N_8662,N_12309);
or U14721 (N_14721,N_11898,N_12004);
and U14722 (N_14722,N_10290,N_11147);
nor U14723 (N_14723,N_9043,N_10133);
nor U14724 (N_14724,N_11068,N_7795);
nand U14725 (N_14725,N_9738,N_8181);
nand U14726 (N_14726,N_11249,N_9382);
and U14727 (N_14727,N_11062,N_6811);
or U14728 (N_14728,N_9516,N_10549);
and U14729 (N_14729,N_8105,N_11883);
or U14730 (N_14730,N_10056,N_10187);
or U14731 (N_14731,N_7016,N_8925);
nor U14732 (N_14732,N_7021,N_12043);
nor U14733 (N_14733,N_12341,N_10483);
nor U14734 (N_14734,N_7855,N_10890);
nand U14735 (N_14735,N_6467,N_8903);
nand U14736 (N_14736,N_12215,N_9073);
and U14737 (N_14737,N_10564,N_11765);
and U14738 (N_14738,N_9137,N_6950);
and U14739 (N_14739,N_7415,N_9274);
or U14740 (N_14740,N_9865,N_8611);
xnor U14741 (N_14741,N_10410,N_10014);
nand U14742 (N_14742,N_6698,N_11921);
nor U14743 (N_14743,N_10717,N_6857);
nor U14744 (N_14744,N_11128,N_11785);
nand U14745 (N_14745,N_11051,N_7949);
or U14746 (N_14746,N_8645,N_12083);
nor U14747 (N_14747,N_11036,N_8464);
nor U14748 (N_14748,N_11729,N_12277);
and U14749 (N_14749,N_11220,N_8497);
nand U14750 (N_14750,N_6620,N_8411);
or U14751 (N_14751,N_11843,N_11092);
nor U14752 (N_14752,N_12293,N_10746);
and U14753 (N_14753,N_10907,N_9174);
nand U14754 (N_14754,N_12205,N_9687);
and U14755 (N_14755,N_7109,N_10488);
and U14756 (N_14756,N_10769,N_12282);
nand U14757 (N_14757,N_8362,N_8782);
or U14758 (N_14758,N_11938,N_10375);
xnor U14759 (N_14759,N_9209,N_9486);
nor U14760 (N_14760,N_7214,N_8229);
nor U14761 (N_14761,N_11915,N_9644);
and U14762 (N_14762,N_11188,N_9755);
or U14763 (N_14763,N_9596,N_6954);
nand U14764 (N_14764,N_12217,N_11107);
or U14765 (N_14765,N_8703,N_10553);
and U14766 (N_14766,N_8677,N_11348);
nor U14767 (N_14767,N_10018,N_8865);
nand U14768 (N_14768,N_10730,N_11021);
nor U14769 (N_14769,N_12174,N_10507);
and U14770 (N_14770,N_12405,N_9456);
or U14771 (N_14771,N_7009,N_8287);
xor U14772 (N_14772,N_6279,N_11464);
or U14773 (N_14773,N_9825,N_9705);
and U14774 (N_14774,N_9450,N_11085);
or U14775 (N_14775,N_10707,N_7176);
and U14776 (N_14776,N_10279,N_10634);
and U14777 (N_14777,N_11663,N_8989);
nor U14778 (N_14778,N_12276,N_6262);
nor U14779 (N_14779,N_8869,N_6737);
nor U14780 (N_14780,N_11808,N_8471);
nor U14781 (N_14781,N_8237,N_6914);
or U14782 (N_14782,N_10082,N_7619);
nand U14783 (N_14783,N_11066,N_7677);
nand U14784 (N_14784,N_11374,N_8333);
or U14785 (N_14785,N_11031,N_12100);
nor U14786 (N_14786,N_8435,N_10977);
nor U14787 (N_14787,N_9605,N_7522);
nand U14788 (N_14788,N_12321,N_12436);
and U14789 (N_14789,N_9990,N_6669);
or U14790 (N_14790,N_8354,N_10651);
nor U14791 (N_14791,N_10976,N_6769);
nand U14792 (N_14792,N_11816,N_7785);
and U14793 (N_14793,N_9179,N_10259);
nand U14794 (N_14794,N_6540,N_10408);
or U14795 (N_14795,N_10299,N_12485);
and U14796 (N_14796,N_10669,N_9032);
or U14797 (N_14797,N_8673,N_9128);
and U14798 (N_14798,N_11262,N_6587);
nand U14799 (N_14799,N_8979,N_12491);
and U14800 (N_14800,N_11889,N_7463);
nand U14801 (N_14801,N_7018,N_11360);
and U14802 (N_14802,N_9310,N_10090);
and U14803 (N_14803,N_8807,N_10336);
nand U14804 (N_14804,N_7443,N_10638);
nand U14805 (N_14805,N_10563,N_9894);
nor U14806 (N_14806,N_11195,N_7669);
or U14807 (N_14807,N_7050,N_9044);
nand U14808 (N_14808,N_7501,N_11917);
nand U14809 (N_14809,N_12454,N_6593);
nor U14810 (N_14810,N_6355,N_10250);
and U14811 (N_14811,N_6566,N_10211);
nand U14812 (N_14812,N_8239,N_10311);
or U14813 (N_14813,N_8296,N_7294);
nor U14814 (N_14814,N_8991,N_12494);
xnor U14815 (N_14815,N_8506,N_12328);
xor U14816 (N_14816,N_10301,N_10260);
nor U14817 (N_14817,N_11503,N_11754);
nand U14818 (N_14818,N_12462,N_7799);
nand U14819 (N_14819,N_8582,N_8400);
or U14820 (N_14820,N_10275,N_7979);
or U14821 (N_14821,N_8580,N_9637);
and U14822 (N_14822,N_12060,N_8748);
and U14823 (N_14823,N_7747,N_9980);
nand U14824 (N_14824,N_7215,N_10802);
nor U14825 (N_14825,N_9997,N_6834);
and U14826 (N_14826,N_6800,N_10998);
or U14827 (N_14827,N_10764,N_12231);
and U14828 (N_14828,N_8494,N_9027);
or U14829 (N_14829,N_9669,N_11421);
or U14830 (N_14830,N_7727,N_9728);
and U14831 (N_14831,N_11042,N_10193);
nand U14832 (N_14832,N_9935,N_8429);
and U14833 (N_14833,N_11657,N_9683);
nand U14834 (N_14834,N_9616,N_7954);
or U14835 (N_14835,N_7318,N_10334);
nand U14836 (N_14836,N_6740,N_9201);
and U14837 (N_14837,N_9889,N_9014);
nor U14838 (N_14838,N_8810,N_8171);
or U14839 (N_14839,N_7542,N_7779);
and U14840 (N_14840,N_7834,N_9647);
and U14841 (N_14841,N_9437,N_7614);
nand U14842 (N_14842,N_11847,N_7107);
nand U14843 (N_14843,N_9662,N_11210);
nand U14844 (N_14844,N_12414,N_7400);
and U14845 (N_14845,N_11899,N_11393);
nor U14846 (N_14846,N_11935,N_6495);
and U14847 (N_14847,N_7207,N_12012);
and U14848 (N_14848,N_6719,N_10368);
nor U14849 (N_14849,N_10535,N_6590);
xnor U14850 (N_14850,N_11493,N_11607);
and U14851 (N_14851,N_12446,N_7853);
or U14852 (N_14852,N_10013,N_11199);
nor U14853 (N_14853,N_9458,N_9840);
or U14854 (N_14854,N_10008,N_12226);
or U14855 (N_14855,N_6989,N_11289);
or U14856 (N_14856,N_9859,N_6648);
nand U14857 (N_14857,N_7938,N_7968);
nor U14858 (N_14858,N_12198,N_9386);
or U14859 (N_14859,N_11505,N_12220);
or U14860 (N_14860,N_12114,N_9731);
and U14861 (N_14861,N_12180,N_6753);
or U14862 (N_14862,N_8574,N_6854);
nor U14863 (N_14863,N_10878,N_8697);
nor U14864 (N_14864,N_11748,N_9191);
nor U14865 (N_14865,N_6586,N_10340);
and U14866 (N_14866,N_8220,N_8621);
or U14867 (N_14867,N_9194,N_9629);
nand U14868 (N_14868,N_8154,N_9257);
nand U14869 (N_14869,N_12286,N_11978);
and U14870 (N_14870,N_11355,N_8089);
nand U14871 (N_14871,N_6758,N_8912);
nand U14872 (N_14872,N_7239,N_7340);
and U14873 (N_14873,N_11265,N_6486);
or U14874 (N_14874,N_11149,N_7858);
and U14875 (N_14875,N_9850,N_8185);
or U14876 (N_14876,N_11019,N_9420);
nand U14877 (N_14877,N_9560,N_8837);
nor U14878 (N_14878,N_9991,N_10297);
nor U14879 (N_14879,N_12333,N_8801);
nand U14880 (N_14880,N_9231,N_10445);
or U14881 (N_14881,N_10693,N_8390);
nor U14882 (N_14882,N_12375,N_7787);
and U14883 (N_14883,N_11827,N_7426);
or U14884 (N_14884,N_11677,N_12492);
and U14885 (N_14885,N_10543,N_6487);
nor U14886 (N_14886,N_10555,N_9164);
and U14887 (N_14887,N_6603,N_6469);
or U14888 (N_14888,N_11602,N_8808);
or U14889 (N_14889,N_11495,N_11805);
nor U14890 (N_14890,N_10748,N_9425);
nor U14891 (N_14891,N_6881,N_7761);
xnor U14892 (N_14892,N_9112,N_6684);
or U14893 (N_14893,N_9853,N_11323);
xnor U14894 (N_14894,N_10181,N_10566);
nor U14895 (N_14895,N_6969,N_7571);
and U14896 (N_14896,N_9040,N_12452);
xor U14897 (N_14897,N_7615,N_10132);
nor U14898 (N_14898,N_9444,N_11310);
nand U14899 (N_14899,N_7755,N_8338);
xor U14900 (N_14900,N_9431,N_9401);
nor U14901 (N_14901,N_7097,N_8563);
nor U14902 (N_14902,N_8597,N_9849);
nor U14903 (N_14903,N_6326,N_6252);
nor U14904 (N_14904,N_6360,N_9723);
xnor U14905 (N_14905,N_7367,N_12272);
xor U14906 (N_14906,N_10136,N_8341);
or U14907 (N_14907,N_11964,N_9833);
and U14908 (N_14908,N_11626,N_7612);
or U14909 (N_14909,N_8416,N_12109);
nand U14910 (N_14910,N_10446,N_10702);
nor U14911 (N_14911,N_10562,N_10537);
and U14912 (N_14912,N_10565,N_11067);
and U14913 (N_14913,N_9173,N_6601);
nor U14914 (N_14914,N_11009,N_10380);
and U14915 (N_14915,N_8348,N_8512);
or U14916 (N_14916,N_9351,N_12175);
and U14917 (N_14917,N_11203,N_11402);
xor U14918 (N_14918,N_7844,N_10716);
and U14919 (N_14919,N_9831,N_10022);
nand U14920 (N_14920,N_12089,N_10840);
nor U14921 (N_14921,N_9787,N_11902);
nand U14922 (N_14922,N_9270,N_6858);
and U14923 (N_14923,N_8671,N_7729);
or U14924 (N_14924,N_10687,N_8792);
or U14925 (N_14925,N_12359,N_9321);
xor U14926 (N_14926,N_6395,N_10514);
nand U14927 (N_14927,N_9398,N_11079);
nand U14928 (N_14928,N_8102,N_6458);
nand U14929 (N_14929,N_11820,N_11381);
and U14930 (N_14930,N_8804,N_10138);
nor U14931 (N_14931,N_8061,N_6286);
xor U14932 (N_14932,N_8427,N_8828);
nand U14933 (N_14933,N_7835,N_10521);
nor U14934 (N_14934,N_11241,N_9189);
or U14935 (N_14935,N_12092,N_6409);
nand U14936 (N_14936,N_12201,N_8194);
nor U14937 (N_14937,N_8019,N_6573);
or U14938 (N_14938,N_6311,N_12395);
or U14939 (N_14939,N_9557,N_11597);
nor U14940 (N_14940,N_9052,N_10667);
and U14941 (N_14941,N_7651,N_6988);
and U14942 (N_14942,N_10568,N_7058);
nor U14943 (N_14943,N_9029,N_9798);
and U14944 (N_14944,N_8059,N_11407);
nor U14945 (N_14945,N_7864,N_9277);
nand U14946 (N_14946,N_9001,N_9989);
nor U14947 (N_14947,N_9106,N_10186);
nand U14948 (N_14948,N_8200,N_11171);
nand U14949 (N_14949,N_10571,N_10364);
nor U14950 (N_14950,N_11512,N_11910);
or U14951 (N_14951,N_8462,N_11780);
nor U14952 (N_14952,N_10015,N_8216);
and U14953 (N_14953,N_7328,N_10527);
nand U14954 (N_14954,N_11133,N_7876);
nor U14955 (N_14955,N_12419,N_8544);
nand U14956 (N_14956,N_7059,N_9311);
and U14957 (N_14957,N_10583,N_10856);
xor U14958 (N_14958,N_12477,N_7386);
nor U14959 (N_14959,N_9821,N_12424);
xnor U14960 (N_14960,N_6708,N_11654);
or U14961 (N_14961,N_7064,N_9086);
or U14962 (N_14962,N_9328,N_9300);
and U14963 (N_14963,N_10877,N_10650);
or U14964 (N_14964,N_7663,N_7659);
nand U14965 (N_14965,N_10005,N_7753);
or U14966 (N_14966,N_7827,N_11481);
nand U14967 (N_14967,N_9298,N_9170);
xor U14968 (N_14968,N_9684,N_9967);
or U14969 (N_14969,N_7174,N_11891);
xnor U14970 (N_14970,N_12449,N_12434);
nand U14971 (N_14971,N_6961,N_11976);
and U14972 (N_14972,N_7822,N_9707);
or U14973 (N_14973,N_11004,N_12392);
or U14974 (N_14974,N_12159,N_10809);
nor U14975 (N_14975,N_9036,N_11295);
nor U14976 (N_14976,N_9145,N_11387);
nand U14977 (N_14977,N_10066,N_11981);
and U14978 (N_14978,N_9410,N_12250);
or U14979 (N_14979,N_11029,N_8535);
nand U14980 (N_14980,N_7943,N_11094);
nor U14981 (N_14981,N_10481,N_6631);
or U14982 (N_14982,N_9528,N_8034);
xnor U14983 (N_14983,N_9693,N_10837);
or U14984 (N_14984,N_10736,N_6662);
or U14985 (N_14985,N_10473,N_10202);
nor U14986 (N_14986,N_10784,N_6726);
or U14987 (N_14987,N_7359,N_11410);
nor U14988 (N_14988,N_12490,N_6498);
and U14989 (N_14989,N_6384,N_7945);
or U14990 (N_14990,N_12469,N_10598);
nor U14991 (N_14991,N_12335,N_8575);
nor U14992 (N_14992,N_8351,N_11084);
and U14993 (N_14993,N_7027,N_9233);
or U14994 (N_14994,N_12268,N_11106);
and U14995 (N_14995,N_7578,N_11484);
nor U14996 (N_14996,N_8073,N_10648);
or U14997 (N_14997,N_7001,N_7374);
and U14998 (N_14998,N_11541,N_9101);
nor U14999 (N_14999,N_10763,N_8889);
nand U15000 (N_15000,N_11204,N_7244);
nor U15001 (N_15001,N_9657,N_8334);
or U15002 (N_15002,N_9121,N_8172);
and U15003 (N_15003,N_7602,N_8420);
nor U15004 (N_15004,N_10238,N_11675);
xor U15005 (N_15005,N_6745,N_8159);
and U15006 (N_15006,N_8960,N_6889);
nand U15007 (N_15007,N_8590,N_10988);
or U15008 (N_15008,N_12164,N_9567);
xnor U15009 (N_15009,N_9800,N_9881);
and U15010 (N_15010,N_11132,N_10712);
xnor U15011 (N_15011,N_11966,N_7748);
xnor U15012 (N_15012,N_8927,N_11794);
or U15013 (N_15013,N_9255,N_9823);
or U15014 (N_15014,N_12178,N_8393);
nand U15015 (N_15015,N_8766,N_6700);
and U15016 (N_15016,N_6765,N_6865);
and U15017 (N_15017,N_8028,N_8246);
or U15018 (N_15018,N_9573,N_11123);
nand U15019 (N_15019,N_10190,N_10918);
nand U15020 (N_15020,N_8700,N_9080);
nand U15021 (N_15021,N_7192,N_6541);
nor U15022 (N_15022,N_6502,N_11946);
xnor U15023 (N_15023,N_8138,N_11618);
or U15024 (N_15024,N_10394,N_8097);
xor U15025 (N_15025,N_8678,N_8607);
and U15026 (N_15026,N_6259,N_11730);
and U15027 (N_15027,N_8272,N_9077);
and U15028 (N_15028,N_9047,N_9700);
nand U15029 (N_15029,N_7570,N_8725);
nand U15030 (N_15030,N_10623,N_11078);
xor U15031 (N_15031,N_9931,N_12133);
or U15032 (N_15032,N_9810,N_11273);
and U15033 (N_15033,N_7320,N_6481);
and U15034 (N_15034,N_10396,N_9608);
xor U15035 (N_15035,N_8928,N_10496);
and U15036 (N_15036,N_9474,N_9236);
nor U15037 (N_15037,N_11086,N_6902);
and U15038 (N_15038,N_8958,N_9380);
and U15039 (N_15039,N_6430,N_9603);
nand U15040 (N_15040,N_7581,N_7985);
nand U15041 (N_15041,N_7633,N_7256);
and U15042 (N_15042,N_8706,N_8855);
or U15043 (N_15043,N_6963,N_9778);
nand U15044 (N_15044,N_8248,N_7777);
or U15045 (N_15045,N_6822,N_8213);
xor U15046 (N_15046,N_10946,N_8249);
nor U15047 (N_15047,N_9663,N_8349);
or U15048 (N_15048,N_11373,N_11179);
or U15049 (N_15049,N_9265,N_8933);
and U15050 (N_15050,N_10229,N_10912);
or U15051 (N_15051,N_8789,N_11682);
and U15052 (N_15052,N_6632,N_9679);
nand U15053 (N_15053,N_8492,N_6893);
and U15054 (N_15054,N_9870,N_12408);
nand U15055 (N_15055,N_9392,N_6878);
or U15056 (N_15056,N_8769,N_12051);
nand U15057 (N_15057,N_12104,N_6866);
and U15058 (N_15058,N_10739,N_11093);
nor U15059 (N_15059,N_11181,N_6288);
and U15060 (N_15060,N_7480,N_10493);
xor U15061 (N_15061,N_10164,N_6396);
xor U15062 (N_15062,N_6879,N_12237);
or U15063 (N_15063,N_11918,N_12444);
nand U15064 (N_15064,N_8146,N_8983);
nand U15065 (N_15065,N_9551,N_7511);
or U15066 (N_15066,N_9593,N_8176);
xnor U15067 (N_15067,N_12478,N_8268);
nand U15068 (N_15068,N_6967,N_10775);
or U15069 (N_15069,N_7947,N_11430);
nor U15070 (N_15070,N_9664,N_7329);
or U15071 (N_15071,N_11193,N_10852);
or U15072 (N_15072,N_6829,N_10596);
or U15073 (N_15073,N_7142,N_12398);
or U15074 (N_15074,N_10024,N_10577);
nand U15075 (N_15075,N_10726,N_10893);
nand U15076 (N_15076,N_8980,N_11842);
xor U15077 (N_15077,N_11944,N_7029);
nor U15078 (N_15078,N_11958,N_8964);
nor U15079 (N_15079,N_7698,N_6307);
and U15080 (N_15080,N_8279,N_10897);
nor U15081 (N_15081,N_11266,N_9520);
and U15082 (N_15082,N_8503,N_9020);
nor U15083 (N_15083,N_7601,N_10880);
nor U15084 (N_15084,N_12142,N_12307);
or U15085 (N_15085,N_7277,N_7010);
xor U15086 (N_15086,N_9717,N_8261);
nor U15087 (N_15087,N_11621,N_12382);
nand U15088 (N_15088,N_6551,N_12496);
or U15089 (N_15089,N_9002,N_10542);
or U15090 (N_15090,N_8197,N_9866);
nor U15091 (N_15091,N_9876,N_7442);
nor U15092 (N_15092,N_11873,N_6550);
nor U15093 (N_15093,N_10839,N_11637);
and U15094 (N_15094,N_12368,N_11030);
nand U15095 (N_15095,N_8632,N_11538);
nand U15096 (N_15096,N_8842,N_6431);
nand U15097 (N_15097,N_10570,N_7216);
nand U15098 (N_15098,N_10955,N_9353);
nor U15099 (N_15099,N_7708,N_8969);
xnor U15100 (N_15100,N_7681,N_9485);
nor U15101 (N_15101,N_11750,N_12086);
nand U15102 (N_15102,N_6756,N_10698);
nand U15103 (N_15103,N_9726,N_8173);
nand U15104 (N_15104,N_10291,N_9868);
nor U15105 (N_15105,N_9708,N_11596);
nand U15106 (N_15106,N_6987,N_7896);
nand U15107 (N_15107,N_10879,N_8273);
nor U15108 (N_15108,N_8651,N_12149);
nand U15109 (N_15109,N_11714,N_11100);
xnor U15110 (N_15110,N_8555,N_11671);
nor U15111 (N_15111,N_9860,N_8672);
or U15112 (N_15112,N_7994,N_6253);
nand U15113 (N_15113,N_11492,N_10767);
or U15114 (N_15114,N_7875,N_9171);
xnor U15115 (N_15115,N_7952,N_7546);
or U15116 (N_15116,N_9329,N_11540);
nand U15117 (N_15117,N_11993,N_11429);
nor U15118 (N_15118,N_9053,N_10028);
nand U15119 (N_15119,N_7842,N_8256);
nor U15120 (N_15120,N_8840,N_8916);
xnor U15121 (N_15121,N_8819,N_12132);
nor U15122 (N_15122,N_10999,N_12340);
or U15123 (N_15123,N_6976,N_9913);
or U15124 (N_15124,N_10561,N_12450);
or U15125 (N_15125,N_9317,N_10374);
nand U15126 (N_15126,N_7993,N_6894);
and U15127 (N_15127,N_11971,N_9544);
nand U15128 (N_15128,N_11112,N_11403);
or U15129 (N_15129,N_8062,N_6715);
and U15130 (N_15130,N_11326,N_8900);
nand U15131 (N_15131,N_6611,N_7249);
xnor U15132 (N_15132,N_11734,N_11652);
xnor U15133 (N_15133,N_6713,N_7582);
nor U15134 (N_15134,N_11604,N_11236);
or U15135 (N_15135,N_11325,N_8794);
nand U15136 (N_15136,N_7154,N_10860);
nand U15137 (N_15137,N_10541,N_11831);
nor U15138 (N_15138,N_9187,N_10592);
and U15139 (N_15139,N_10666,N_7155);
and U15140 (N_15140,N_9430,N_12135);
nor U15141 (N_15141,N_10607,N_8674);
and U15142 (N_15142,N_9531,N_7552);
and U15143 (N_15143,N_7505,N_7030);
nand U15144 (N_15144,N_7758,N_7605);
and U15145 (N_15145,N_11020,N_7624);
nor U15146 (N_15146,N_6545,N_9383);
and U15147 (N_15147,N_9753,N_10804);
and U15148 (N_15148,N_9154,N_10934);
and U15149 (N_15149,N_8430,N_9190);
and U15150 (N_15150,N_11422,N_10116);
or U15151 (N_15151,N_11546,N_7643);
and U15152 (N_15152,N_10824,N_9126);
nor U15153 (N_15153,N_11370,N_8669);
nand U15154 (N_15154,N_7780,N_7723);
nor U15155 (N_15155,N_11328,N_10160);
nand U15156 (N_15156,N_9066,N_7655);
and U15157 (N_15157,N_7807,N_8300);
and U15158 (N_15158,N_11766,N_11624);
nor U15159 (N_15159,N_12406,N_6900);
or U15160 (N_15160,N_6619,N_10016);
nor U15161 (N_15161,N_8929,N_7726);
nor U15162 (N_15162,N_10032,N_10104);
or U15163 (N_15163,N_8474,N_9855);
or U15164 (N_15164,N_6389,N_8401);
xnor U15165 (N_15165,N_11849,N_12265);
nand U15166 (N_15166,N_7257,N_6779);
or U15167 (N_15167,N_9941,N_8628);
and U15168 (N_15168,N_7031,N_6598);
nor U15169 (N_15169,N_11556,N_8040);
and U15170 (N_15170,N_6503,N_11669);
or U15171 (N_15171,N_12140,N_12212);
and U15172 (N_15172,N_9272,N_9533);
nand U15173 (N_15173,N_7243,N_10039);
nand U15174 (N_15174,N_8843,N_11548);
and U15175 (N_15175,N_10011,N_8612);
and U15176 (N_15176,N_12181,N_11810);
nor U15177 (N_15177,N_7811,N_11857);
or U15178 (N_15178,N_8413,N_11863);
nand U15179 (N_15179,N_8921,N_6689);
or U15180 (N_15180,N_12224,N_6741);
and U15181 (N_15181,N_7646,N_8116);
and U15182 (N_15182,N_12458,N_8930);
or U15183 (N_15183,N_8006,N_10691);
xnor U15184 (N_15184,N_11811,N_9974);
nor U15185 (N_15185,N_11287,N_8455);
nor U15186 (N_15186,N_10515,N_7487);
or U15187 (N_15187,N_11919,N_9577);
or U15188 (N_15188,N_6474,N_9547);
or U15189 (N_15189,N_10844,N_6977);
nor U15190 (N_15190,N_12029,N_11727);
nor U15191 (N_15191,N_11679,N_10600);
or U15192 (N_15192,N_10938,N_8680);
or U15193 (N_15193,N_7485,N_6653);
nor U15194 (N_15194,N_9847,N_6604);
nand U15195 (N_15195,N_8884,N_8913);
or U15196 (N_15196,N_7441,N_9740);
or U15197 (N_15197,N_7891,N_12101);
nand U15198 (N_15198,N_8183,N_8618);
or U15199 (N_15199,N_6994,N_9950);
and U15200 (N_15200,N_12471,N_10422);
and U15201 (N_15201,N_12482,N_10919);
and U15202 (N_15202,N_12314,N_8280);
and U15203 (N_15203,N_8141,N_10992);
and U15204 (N_15204,N_8366,N_6835);
and U15205 (N_15205,N_7897,N_8774);
or U15206 (N_15206,N_7976,N_8533);
or U15207 (N_15207,N_10728,N_11229);
and U15208 (N_15208,N_10683,N_7259);
nor U15209 (N_15209,N_11016,N_11312);
or U15210 (N_15210,N_8432,N_9051);
or U15211 (N_15211,N_8761,N_7489);
nor U15212 (N_15212,N_8001,N_11672);
or U15213 (N_15213,N_8361,N_7860);
nor U15214 (N_15214,N_9063,N_9784);
nand U15215 (N_15215,N_8122,N_10235);
and U15216 (N_15216,N_10308,N_8339);
and U15217 (N_15217,N_8352,N_11903);
nand U15218 (N_15218,N_8863,N_6805);
nand U15219 (N_15219,N_7814,N_11048);
nand U15220 (N_15220,N_8224,N_11833);
or U15221 (N_15221,N_9115,N_11167);
nand U15222 (N_15222,N_6477,N_11573);
nor U15223 (N_15223,N_11320,N_9330);
or U15224 (N_15224,N_8058,N_8294);
and U15225 (N_15225,N_12269,N_10102);
nor U15226 (N_15226,N_9476,N_11549);
xor U15227 (N_15227,N_6520,N_12376);
nand U15228 (N_15228,N_11459,N_8071);
nand U15229 (N_15229,N_6864,N_10891);
and U15230 (N_15230,N_7700,N_11039);
and U15231 (N_15231,N_6322,N_8557);
and U15232 (N_15232,N_11806,N_11396);
nand U15233 (N_15233,N_10920,N_6926);
or U15234 (N_15234,N_9899,N_8877);
nor U15235 (N_15235,N_7909,N_9016);
nand U15236 (N_15236,N_12481,N_8027);
nand U15237 (N_15237,N_6983,N_11023);
or U15238 (N_15238,N_6547,N_7704);
nor U15239 (N_15239,N_11931,N_7596);
xor U15240 (N_15240,N_7653,N_6885);
nor U15241 (N_15241,N_10341,N_7977);
or U15242 (N_15242,N_10961,N_12275);
xnor U15243 (N_15243,N_6875,N_12460);
or U15244 (N_15244,N_8008,N_8644);
nor U15245 (N_15245,N_11834,N_9651);
or U15246 (N_15246,N_8667,N_9399);
nor U15247 (N_15247,N_11040,N_11117);
or U15248 (N_15248,N_10248,N_7229);
nand U15249 (N_15249,N_11533,N_11145);
and U15250 (N_15250,N_11615,N_12421);
nor U15251 (N_15251,N_9506,N_7129);
xor U15252 (N_15252,N_6250,N_7309);
nor U15253 (N_15253,N_7840,N_8633);
or U15254 (N_15254,N_9863,N_11412);
nand U15255 (N_15255,N_7285,N_9048);
xor U15256 (N_15256,N_12206,N_6417);
nand U15257 (N_15257,N_8655,N_8439);
or U15258 (N_15258,N_10694,N_7291);
nand U15259 (N_15259,N_10777,N_8803);
nor U15260 (N_15260,N_8642,N_7707);
or U15261 (N_15261,N_7711,N_11879);
nand U15262 (N_15262,N_11157,N_6849);
and U15263 (N_15263,N_7015,N_7462);
nand U15264 (N_15264,N_12431,N_12202);
xnor U15265 (N_15265,N_9157,N_7420);
nand U15266 (N_15266,N_8318,N_7972);
and U15267 (N_15267,N_11823,N_11629);
xor U15268 (N_15268,N_6369,N_11006);
nor U15269 (N_15269,N_11995,N_8212);
or U15270 (N_15270,N_11244,N_11111);
nor U15271 (N_15271,N_11054,N_8052);
or U15272 (N_15272,N_7978,N_9013);
nor U15273 (N_15273,N_9575,N_6488);
nor U15274 (N_15274,N_11979,N_12312);
and U15275 (N_15275,N_7298,N_11630);
nand U15276 (N_15276,N_7986,N_9661);
nand U15277 (N_15277,N_8196,N_11390);
and U15278 (N_15278,N_9674,N_7428);
or U15279 (N_15279,N_10935,N_9902);
or U15280 (N_15280,N_11327,N_7686);
and U15281 (N_15281,N_6935,N_7573);
and U15282 (N_15282,N_9093,N_12153);
nand U15283 (N_15283,N_11208,N_11623);
xnor U15284 (N_15284,N_9192,N_6291);
nand U15285 (N_15285,N_8963,N_7961);
nor U15286 (N_15286,N_7421,N_8167);
nor U15287 (N_15287,N_11703,N_12459);
or U15288 (N_15288,N_6509,N_7370);
nor U15289 (N_15289,N_6531,N_6251);
or U15290 (N_15290,N_9136,N_7345);
or U15291 (N_15291,N_11380,N_10697);
nor U15292 (N_15292,N_9113,N_9176);
xnor U15293 (N_15293,N_7620,N_10451);
or U15294 (N_15294,N_8549,N_9025);
or U15295 (N_15295,N_6615,N_10452);
nand U15296 (N_15296,N_7205,N_8547);
or U15297 (N_15297,N_7454,N_9388);
nor U15298 (N_15298,N_11527,N_9094);
nor U15299 (N_15299,N_7908,N_11870);
and U15300 (N_15300,N_7278,N_7085);
nor U15301 (N_15301,N_12077,N_9448);
and U15302 (N_15302,N_10652,N_11121);
nand U15303 (N_15303,N_8157,N_9467);
nor U15304 (N_15304,N_6273,N_10019);
xor U15305 (N_15305,N_8515,N_11776);
nor U15306 (N_15306,N_7088,N_9841);
nor U15307 (N_15307,N_11925,N_8223);
nor U15308 (N_15308,N_11796,N_7114);
nand U15309 (N_15309,N_9457,N_9590);
and U15310 (N_15310,N_9871,N_8373);
nand U15311 (N_15311,N_9623,N_8016);
or U15312 (N_15312,N_9911,N_6444);
nand U15313 (N_15313,N_8776,N_7002);
nor U15314 (N_15314,N_11584,N_12099);
and U15315 (N_15315,N_6808,N_8545);
nand U15316 (N_15316,N_8120,N_11223);
nand U15317 (N_15317,N_8454,N_11974);
nand U15318 (N_15318,N_10742,N_10476);
and U15319 (N_15319,N_7063,N_8530);
xor U15320 (N_15320,N_8125,N_7044);
and U15321 (N_15321,N_10172,N_7168);
or U15322 (N_15322,N_12466,N_9463);
nand U15323 (N_15323,N_8649,N_11508);
nor U15324 (N_15324,N_10419,N_7884);
nand U15325 (N_15325,N_9141,N_6492);
nor U15326 (N_15326,N_6363,N_11943);
or U15327 (N_15327,N_12156,N_10283);
or U15328 (N_15328,N_6688,N_6394);
and U15329 (N_15329,N_6564,N_10594);
xor U15330 (N_15330,N_12017,N_7579);
or U15331 (N_15331,N_11561,N_7691);
nand U15332 (N_15332,N_9904,N_9501);
and U15333 (N_15333,N_8595,N_8024);
nor U15334 (N_15334,N_11443,N_9829);
and U15335 (N_15335,N_10550,N_6293);
xor U15336 (N_15336,N_11047,N_12002);
nor U15337 (N_15337,N_9011,N_7539);
or U15338 (N_15338,N_11405,N_10581);
nor U15339 (N_15339,N_10118,N_9635);
or U15340 (N_15340,N_6398,N_8299);
nand U15341 (N_15341,N_10886,N_10115);
or U15342 (N_15342,N_11788,N_10035);
and U15343 (N_15343,N_10484,N_6974);
nor U15344 (N_15344,N_12071,N_11343);
nand U15345 (N_15345,N_8143,N_9620);
and U15346 (N_15346,N_9219,N_7111);
nor U15347 (N_15347,N_7923,N_10125);
and U15348 (N_15348,N_11494,N_10910);
xnor U15349 (N_15349,N_11603,N_9759);
and U15350 (N_15350,N_7468,N_10243);
nand U15351 (N_15351,N_9384,N_7014);
nand U15352 (N_15352,N_9103,N_8950);
and U15353 (N_15353,N_9327,N_7668);
and U15354 (N_15354,N_12182,N_9549);
nand U15355 (N_15355,N_11997,N_10296);
nand U15356 (N_15356,N_6621,N_7486);
nor U15357 (N_15357,N_9774,N_9650);
and U15358 (N_15358,N_10091,N_11904);
or U15359 (N_15359,N_10779,N_7051);
nand U15360 (N_15360,N_10286,N_8704);
and U15361 (N_15361,N_7543,N_11498);
nor U15362 (N_15362,N_10358,N_9326);
xnor U15363 (N_15363,N_12422,N_9737);
nand U15364 (N_15364,N_10355,N_11283);
and U15365 (N_15365,N_6392,N_10225);
or U15366 (N_15366,N_9613,N_9727);
and U15367 (N_15367,N_8622,N_6943);
nand U15368 (N_15368,N_10883,N_10665);
and U15369 (N_15369,N_6500,N_12336);
nand U15370 (N_15370,N_9792,N_10829);
and U15371 (N_15371,N_10448,N_11465);
xnor U15372 (N_15372,N_8717,N_8905);
nor U15373 (N_15373,N_11859,N_8043);
and U15374 (N_15374,N_7509,N_9280);
nand U15375 (N_15375,N_8209,N_11190);
or U15376 (N_15376,N_8235,N_9581);
nand U15377 (N_15377,N_10462,N_10979);
nand U15378 (N_15378,N_9510,N_11547);
nor U15379 (N_15379,N_6682,N_11658);
nor U15380 (N_15380,N_10719,N_10612);
and U15381 (N_15381,N_6290,N_6390);
nor U15382 (N_15382,N_11994,N_12295);
xor U15383 (N_15383,N_7157,N_9748);
and U15384 (N_15384,N_10720,N_12204);
nand U15385 (N_15385,N_10757,N_9918);
and U15386 (N_15386,N_12354,N_11509);
xnor U15387 (N_15387,N_12355,N_10618);
nor U15388 (N_15388,N_10911,N_8897);
and U15389 (N_15389,N_9147,N_8326);
nand U15390 (N_15390,N_6583,N_6912);
nor U15391 (N_15391,N_9492,N_12302);
and U15392 (N_15392,N_6491,N_11141);
nor U15393 (N_15393,N_10708,N_6464);
and U15394 (N_15394,N_9155,N_10904);
and U15395 (N_15395,N_8156,N_7203);
nor U15396 (N_15396,N_7036,N_11530);
xnor U15397 (N_15397,N_10696,N_6300);
and U15398 (N_15398,N_7595,N_7231);
nor U15399 (N_15399,N_11953,N_8214);
or U15400 (N_15400,N_9445,N_8760);
nor U15401 (N_15401,N_10858,N_10964);
xnor U15402 (N_15402,N_8773,N_11739);
nor U15403 (N_15403,N_7551,N_6721);
and U15404 (N_15404,N_11217,N_9619);
nor U15405 (N_15405,N_10790,N_6992);
and U15406 (N_15406,N_8011,N_12429);
nor U15407 (N_15407,N_11648,N_12373);
and U15408 (N_15408,N_9295,N_12150);
xnor U15409 (N_15409,N_10586,N_12425);
and U15410 (N_15410,N_11913,N_10438);
nor U15411 (N_15411,N_10950,N_9874);
nor U15412 (N_15412,N_7905,N_11920);
and U15413 (N_15413,N_11202,N_8846);
nor U15414 (N_15414,N_8816,N_6597);
and U15415 (N_15415,N_11900,N_9254);
nor U15416 (N_15416,N_11260,N_9230);
nor U15417 (N_15417,N_8666,N_10672);
or U15418 (N_15418,N_7790,N_10184);
and U15419 (N_15419,N_10688,N_7112);
and U15420 (N_15420,N_9953,N_8314);
nand U15421 (N_15421,N_10442,N_10168);
nand U15422 (N_15422,N_11341,N_7302);
xnor U15423 (N_15423,N_10088,N_9898);
nand U15424 (N_15424,N_6792,N_11710);
and U15425 (N_15425,N_8036,N_7446);
nand U15426 (N_15426,N_6595,N_8461);
and U15427 (N_15427,N_12289,N_7465);
and U15428 (N_15428,N_10048,N_12472);
and U15429 (N_15429,N_8440,N_7106);
nand U15430 (N_15430,N_8727,N_10131);
and U15431 (N_15431,N_7327,N_7241);
nand U15432 (N_15432,N_9568,N_7099);
and U15433 (N_15433,N_9741,N_7599);
nor U15434 (N_15434,N_10392,N_8163);
and U15435 (N_15435,N_11371,N_6608);
and U15436 (N_15436,N_11418,N_11129);
xnor U15437 (N_15437,N_11840,N_7236);
and U15438 (N_15438,N_10423,N_9507);
nand U15439 (N_15439,N_10148,N_12407);
or U15440 (N_15440,N_12115,N_12402);
and U15441 (N_15441,N_12118,N_7068);
and U15442 (N_15442,N_10525,N_10544);
xnor U15443 (N_15443,N_9611,N_10021);
nor U15444 (N_15444,N_8251,N_11382);
or U15445 (N_15445,N_8308,N_10069);
nor U15446 (N_15446,N_7866,N_8255);
xnor U15447 (N_15447,N_9776,N_11059);
nor U15448 (N_15448,N_11579,N_10970);
nor U15449 (N_15449,N_10490,N_7342);
and U15450 (N_15450,N_10631,N_9830);
or U15451 (N_15451,N_6651,N_7966);
nor U15452 (N_15452,N_6472,N_7296);
nor U15453 (N_15453,N_10494,N_7534);
or U15454 (N_15454,N_8852,N_6315);
nand U15455 (N_15455,N_10906,N_7924);
or U15456 (N_15456,N_9537,N_12028);
nand U15457 (N_15457,N_6411,N_12350);
or U15458 (N_15458,N_9046,N_12337);
nor U15459 (N_15459,N_9699,N_9308);
or U15460 (N_15460,N_10778,N_7057);
and U15461 (N_15461,N_6937,N_12018);
or U15462 (N_15462,N_12357,N_7629);
and U15463 (N_15463,N_9224,N_6999);
nand U15464 (N_15464,N_12412,N_8311);
nand U15465 (N_15465,N_10385,N_12499);
and U15466 (N_15466,N_8050,N_7527);
nand U15467 (N_15467,N_8593,N_10547);
nor U15468 (N_15468,N_9256,N_6397);
nand U15469 (N_15469,N_11911,N_10216);
nand U15470 (N_15470,N_6735,N_12245);
nand U15471 (N_15471,N_10302,N_10901);
and U15472 (N_15472,N_12166,N_8169);
nor U15473 (N_15473,N_8112,N_9817);
nor U15474 (N_15474,N_12468,N_11359);
xnor U15475 (N_15475,N_7999,N_6596);
and U15476 (N_15476,N_7225,N_7110);
and U15477 (N_15477,N_9193,N_6814);
and U15478 (N_15478,N_11211,N_11628);
or U15479 (N_15479,N_6405,N_6840);
nor U15480 (N_15480,N_9161,N_9336);
and U15481 (N_15481,N_7337,N_7922);
and U15482 (N_15482,N_9470,N_11425);
or U15483 (N_15483,N_8820,N_9939);
nand U15484 (N_15484,N_10073,N_7268);
nor U15485 (N_15485,N_9548,N_6981);
and U15486 (N_15486,N_7763,N_11206);
nand U15487 (N_15487,N_9639,N_10655);
or U15488 (N_15488,N_7461,N_10559);
or U15489 (N_15489,N_8723,N_6660);
xnor U15490 (N_15490,N_12439,N_6922);
nor U15491 (N_15491,N_10695,N_9591);
or U15492 (N_15492,N_8295,N_12059);
nand U15493 (N_15493,N_10740,N_11034);
and U15494 (N_15494,N_8552,N_9948);
nand U15495 (N_15495,N_8441,N_10894);
nor U15496 (N_15496,N_10182,N_6637);
nor U15497 (N_15497,N_11952,N_7737);
nor U15498 (N_15498,N_11774,N_9642);
nand U15499 (N_15499,N_6812,N_7325);
nor U15500 (N_15500,N_8834,N_12091);
and U15501 (N_15501,N_7600,N_6898);
nor U15502 (N_15502,N_12300,N_9475);
or U15503 (N_15503,N_6558,N_8312);
and U15504 (N_15504,N_7349,N_9400);
nand U15505 (N_15505,N_7209,N_8421);
or U15506 (N_15506,N_6308,N_8114);
nor U15507 (N_15507,N_8047,N_12399);
or U15508 (N_15508,N_12141,N_12107);
and U15509 (N_15509,N_10926,N_6289);
and U15510 (N_15510,N_10673,N_8696);
nand U15511 (N_15511,N_9848,N_12052);
nand U15512 (N_15512,N_9797,N_6882);
nor U15513 (N_15513,N_11130,N_11939);
nor U15514 (N_15514,N_8203,N_12390);
nand U15515 (N_15515,N_11528,N_11861);
xnor U15516 (N_15516,N_9827,N_11033);
or U15517 (N_15517,N_9854,N_8355);
xnor U15518 (N_15518,N_10233,N_8654);
nor U15519 (N_15519,N_8586,N_7117);
xnor U15520 (N_15520,N_12057,N_7299);
xnor U15521 (N_15521,N_9118,N_6574);
nor U15522 (N_15522,N_12195,N_6335);
and U15523 (N_15523,N_11008,N_7246);
or U15524 (N_15524,N_12370,N_12377);
or U15525 (N_15525,N_7123,N_6995);
or U15526 (N_15526,N_10399,N_9091);
and U15527 (N_15527,N_9129,N_12325);
nor U15528 (N_15528,N_7504,N_9364);
nand U15529 (N_15529,N_10436,N_7564);
and U15530 (N_15530,N_7565,N_9836);
or U15531 (N_15531,N_11896,N_6732);
nand U15532 (N_15532,N_7019,N_9003);
and U15533 (N_15533,N_11468,N_7331);
nor U15534 (N_15534,N_10256,N_11526);
or U15535 (N_15535,N_12041,N_9033);
nand U15536 (N_15536,N_7792,N_9890);
nand U15537 (N_15537,N_9434,N_8670);
nor U15538 (N_15538,N_10126,N_6258);
xnor U15539 (N_15539,N_6691,N_7991);
and U15540 (N_15540,N_6568,N_7120);
nor U15541 (N_15541,N_9407,N_9238);
nand U15542 (N_15542,N_7410,N_7560);
nor U15543 (N_15543,N_12221,N_10272);
nand U15544 (N_15544,N_10000,N_9134);
nor U15545 (N_15545,N_11826,N_7586);
and U15546 (N_15546,N_6260,N_7171);
nand U15547 (N_15547,N_8999,N_12241);
and U15548 (N_15548,N_9621,N_11436);
nand U15549 (N_15549,N_11480,N_9588);
or U15550 (N_15550,N_11927,N_10352);
and U15551 (N_15551,N_7071,N_10915);
or U15552 (N_15552,N_6771,N_6599);
nor U15553 (N_15553,N_9304,N_11267);
xnor U15554 (N_15554,N_11395,N_7143);
or U15555 (N_15555,N_10621,N_12493);
xnor U15556 (N_15556,N_12489,N_12199);
xor U15557 (N_15557,N_9585,N_7496);
or U15558 (N_15558,N_8000,N_6855);
xnor U15559 (N_15559,N_8987,N_10214);
nor U15560 (N_15560,N_11166,N_8599);
nand U15561 (N_15561,N_7078,N_9166);
nor U15562 (N_15562,N_8520,N_7759);
nor U15563 (N_15563,N_7052,N_7275);
nand U15564 (N_15564,N_6455,N_6670);
and U15565 (N_15565,N_6275,N_8409);
or U15566 (N_15566,N_7886,N_6681);
nand U15567 (N_15567,N_9416,N_9057);
nor U15568 (N_15568,N_8153,N_11258);
or U15569 (N_15569,N_12227,N_9856);
and U15570 (N_15570,N_6254,N_7635);
and U15571 (N_15571,N_11731,N_7731);
nand U15572 (N_15572,N_10199,N_10836);
and U15573 (N_15573,N_10967,N_7813);
nand U15574 (N_15574,N_9489,N_11102);
or U15575 (N_15575,N_7208,N_6594);
nand U15576 (N_15576,N_9371,N_7576);
or U15577 (N_15577,N_11000,N_11239);
nor U15578 (N_15578,N_6772,N_8093);
and U15579 (N_15579,N_7034,N_11115);
nand U15580 (N_15580,N_10959,N_7053);
nor U15581 (N_15581,N_6910,N_9843);
or U15582 (N_15582,N_8695,N_6744);
or U15583 (N_15583,N_11991,N_11024);
and U15584 (N_15584,N_10609,N_10144);
and U15585 (N_15585,N_9930,N_12157);
nor U15586 (N_15586,N_10731,N_8066);
or U15587 (N_15587,N_11990,N_8496);
or U15588 (N_15588,N_6301,N_7693);
xnor U15589 (N_15589,N_6494,N_6742);
nand U15590 (N_15590,N_8219,N_8119);
and U15591 (N_15591,N_11466,N_7245);
nor U15592 (N_15592,N_6528,N_11143);
or U15593 (N_15593,N_10502,N_6457);
and U15594 (N_15594,N_8074,N_7695);
and U15595 (N_15595,N_6663,N_11970);
or U15596 (N_15596,N_8955,N_10923);
nor U15597 (N_15597,N_7846,N_9396);
or U15598 (N_15598,N_6869,N_10096);
and U15599 (N_15599,N_12093,N_6915);
nor U15600 (N_15600,N_9337,N_9009);
and U15601 (N_15601,N_11519,N_7191);
nor U15602 (N_15602,N_6556,N_11301);
nand U15603 (N_15603,N_8763,N_8168);
xor U15604 (N_15604,N_9169,N_8527);
or U15605 (N_15605,N_8956,N_7902);
or U15606 (N_15606,N_7569,N_10952);
xor U15607 (N_15607,N_6701,N_6368);
xnor U15608 (N_15608,N_11110,N_12261);
or U15609 (N_15609,N_8045,N_7478);
or U15610 (N_15610,N_11963,N_10456);
or U15611 (N_15611,N_10857,N_6445);
or U15612 (N_15612,N_11674,N_11518);
nand U15613 (N_15613,N_11850,N_6538);
or U15614 (N_15614,N_6607,N_7308);
xor U15615 (N_15615,N_11317,N_11688);
and U15616 (N_15616,N_11485,N_7035);
or U15617 (N_15617,N_8616,N_8858);
nor U15618 (N_15618,N_6886,N_7160);
nand U15619 (N_15619,N_10825,N_8899);
xnor U15620 (N_15620,N_8570,N_8292);
and U15621 (N_15621,N_8405,N_12188);
or U15622 (N_15622,N_7149,N_9656);
or U15623 (N_15623,N_6848,N_8603);
xnor U15624 (N_15624,N_7817,N_8814);
and U15625 (N_15625,N_9797,N_6698);
nand U15626 (N_15626,N_8926,N_10257);
or U15627 (N_15627,N_8825,N_8187);
or U15628 (N_15628,N_12487,N_12486);
and U15629 (N_15629,N_6478,N_10756);
and U15630 (N_15630,N_9508,N_11878);
and U15631 (N_15631,N_10417,N_9683);
nand U15632 (N_15632,N_9077,N_10538);
xnor U15633 (N_15633,N_7612,N_6930);
nor U15634 (N_15634,N_8055,N_7226);
nor U15635 (N_15635,N_6284,N_9301);
and U15636 (N_15636,N_10510,N_9168);
and U15637 (N_15637,N_11127,N_7438);
or U15638 (N_15638,N_10483,N_9351);
and U15639 (N_15639,N_7328,N_7932);
nor U15640 (N_15640,N_8892,N_10704);
xor U15641 (N_15641,N_9148,N_6936);
or U15642 (N_15642,N_12025,N_9974);
nand U15643 (N_15643,N_9480,N_7187);
and U15644 (N_15644,N_6496,N_9571);
nor U15645 (N_15645,N_8463,N_9868);
and U15646 (N_15646,N_10346,N_9420);
and U15647 (N_15647,N_11376,N_6651);
nor U15648 (N_15648,N_7881,N_9821);
nand U15649 (N_15649,N_8781,N_8209);
nand U15650 (N_15650,N_7755,N_12314);
or U15651 (N_15651,N_7001,N_8636);
or U15652 (N_15652,N_9945,N_9798);
nand U15653 (N_15653,N_8892,N_11590);
nand U15654 (N_15654,N_8532,N_8101);
nand U15655 (N_15655,N_8118,N_8622);
nand U15656 (N_15656,N_6621,N_7340);
and U15657 (N_15657,N_10741,N_9168);
or U15658 (N_15658,N_10833,N_9807);
nand U15659 (N_15659,N_9865,N_6553);
or U15660 (N_15660,N_9405,N_11374);
nor U15661 (N_15661,N_9500,N_8698);
nand U15662 (N_15662,N_10107,N_7234);
nand U15663 (N_15663,N_9394,N_8932);
or U15664 (N_15664,N_7655,N_11052);
and U15665 (N_15665,N_12300,N_11118);
xnor U15666 (N_15666,N_12237,N_12329);
or U15667 (N_15667,N_10790,N_9529);
nand U15668 (N_15668,N_6731,N_11989);
or U15669 (N_15669,N_10955,N_9141);
nand U15670 (N_15670,N_9521,N_6386);
and U15671 (N_15671,N_8518,N_7233);
nor U15672 (N_15672,N_10135,N_11901);
nand U15673 (N_15673,N_7774,N_10592);
xnor U15674 (N_15674,N_9710,N_8898);
or U15675 (N_15675,N_11694,N_7378);
xor U15676 (N_15676,N_9794,N_10862);
or U15677 (N_15677,N_9343,N_10925);
and U15678 (N_15678,N_7194,N_7883);
and U15679 (N_15679,N_8832,N_7486);
nand U15680 (N_15680,N_6856,N_8224);
nor U15681 (N_15681,N_6283,N_12106);
nor U15682 (N_15682,N_6933,N_9951);
nor U15683 (N_15683,N_12206,N_10140);
or U15684 (N_15684,N_12006,N_10694);
nor U15685 (N_15685,N_6846,N_11709);
nor U15686 (N_15686,N_9575,N_9101);
or U15687 (N_15687,N_9557,N_11500);
and U15688 (N_15688,N_6824,N_10456);
nand U15689 (N_15689,N_10372,N_6279);
nor U15690 (N_15690,N_7814,N_7930);
and U15691 (N_15691,N_12097,N_7962);
nand U15692 (N_15692,N_10505,N_6459);
or U15693 (N_15693,N_12310,N_11396);
and U15694 (N_15694,N_10812,N_7312);
or U15695 (N_15695,N_10612,N_6655);
and U15696 (N_15696,N_8535,N_10984);
and U15697 (N_15697,N_7889,N_11389);
nand U15698 (N_15698,N_12143,N_11125);
or U15699 (N_15699,N_7355,N_10571);
or U15700 (N_15700,N_6509,N_8453);
xor U15701 (N_15701,N_12224,N_10439);
and U15702 (N_15702,N_9722,N_8982);
or U15703 (N_15703,N_9771,N_9982);
and U15704 (N_15704,N_11985,N_8220);
xnor U15705 (N_15705,N_10287,N_6728);
nor U15706 (N_15706,N_10468,N_7265);
or U15707 (N_15707,N_9765,N_11264);
or U15708 (N_15708,N_8871,N_9368);
nand U15709 (N_15709,N_10891,N_8474);
nor U15710 (N_15710,N_10435,N_7878);
or U15711 (N_15711,N_8118,N_11897);
and U15712 (N_15712,N_11563,N_10867);
or U15713 (N_15713,N_11538,N_10302);
or U15714 (N_15714,N_7323,N_10401);
or U15715 (N_15715,N_10881,N_8214);
nor U15716 (N_15716,N_8102,N_6706);
nand U15717 (N_15717,N_9325,N_8300);
xor U15718 (N_15718,N_6960,N_9784);
nor U15719 (N_15719,N_9697,N_6268);
or U15720 (N_15720,N_8313,N_9663);
and U15721 (N_15721,N_10073,N_6763);
nand U15722 (N_15722,N_6813,N_10502);
nand U15723 (N_15723,N_11765,N_12362);
nor U15724 (N_15724,N_12271,N_9323);
and U15725 (N_15725,N_10104,N_6988);
nand U15726 (N_15726,N_9192,N_9071);
xor U15727 (N_15727,N_12259,N_12137);
nor U15728 (N_15728,N_7044,N_8505);
nand U15729 (N_15729,N_10779,N_11280);
nor U15730 (N_15730,N_7388,N_10464);
nand U15731 (N_15731,N_11098,N_10361);
or U15732 (N_15732,N_12238,N_10944);
and U15733 (N_15733,N_7534,N_11321);
or U15734 (N_15734,N_10851,N_11170);
or U15735 (N_15735,N_6724,N_7134);
and U15736 (N_15736,N_9428,N_8896);
xor U15737 (N_15737,N_9520,N_11755);
xnor U15738 (N_15738,N_9544,N_7322);
nand U15739 (N_15739,N_7856,N_9669);
and U15740 (N_15740,N_8929,N_9330);
nor U15741 (N_15741,N_8182,N_10058);
nand U15742 (N_15742,N_6386,N_9683);
or U15743 (N_15743,N_7088,N_11869);
xnor U15744 (N_15744,N_7793,N_8382);
nand U15745 (N_15745,N_11931,N_9239);
nor U15746 (N_15746,N_10418,N_11224);
nand U15747 (N_15747,N_7678,N_11846);
and U15748 (N_15748,N_11836,N_6650);
nor U15749 (N_15749,N_8227,N_8158);
xor U15750 (N_15750,N_11867,N_10031);
nor U15751 (N_15751,N_10451,N_11172);
nand U15752 (N_15752,N_10068,N_11619);
nand U15753 (N_15753,N_8888,N_7874);
nand U15754 (N_15754,N_6612,N_9632);
nor U15755 (N_15755,N_6720,N_11462);
or U15756 (N_15756,N_8891,N_7909);
nor U15757 (N_15757,N_10112,N_8017);
nand U15758 (N_15758,N_9351,N_9394);
or U15759 (N_15759,N_11775,N_7766);
nand U15760 (N_15760,N_8200,N_10812);
nand U15761 (N_15761,N_12480,N_8148);
or U15762 (N_15762,N_6557,N_10569);
or U15763 (N_15763,N_10060,N_11079);
or U15764 (N_15764,N_12416,N_10503);
xnor U15765 (N_15765,N_8048,N_8908);
nand U15766 (N_15766,N_7284,N_10966);
nor U15767 (N_15767,N_8090,N_8888);
and U15768 (N_15768,N_7406,N_11387);
and U15769 (N_15769,N_11855,N_9688);
nor U15770 (N_15770,N_7824,N_7510);
nor U15771 (N_15771,N_9740,N_8128);
or U15772 (N_15772,N_12330,N_7288);
nand U15773 (N_15773,N_8338,N_12021);
nand U15774 (N_15774,N_7793,N_8921);
xnor U15775 (N_15775,N_11082,N_8419);
nand U15776 (N_15776,N_11987,N_10621);
nand U15777 (N_15777,N_11590,N_8751);
and U15778 (N_15778,N_10086,N_9868);
and U15779 (N_15779,N_12218,N_11837);
nor U15780 (N_15780,N_11537,N_11389);
or U15781 (N_15781,N_7483,N_9587);
nand U15782 (N_15782,N_11236,N_9227);
nor U15783 (N_15783,N_6299,N_8644);
xor U15784 (N_15784,N_11213,N_8201);
nor U15785 (N_15785,N_9461,N_9194);
nor U15786 (N_15786,N_6904,N_11604);
or U15787 (N_15787,N_12466,N_7403);
nand U15788 (N_15788,N_9589,N_6964);
nand U15789 (N_15789,N_11051,N_9049);
nand U15790 (N_15790,N_12493,N_7762);
nor U15791 (N_15791,N_9248,N_7796);
xnor U15792 (N_15792,N_9099,N_8504);
nand U15793 (N_15793,N_11975,N_11008);
or U15794 (N_15794,N_10390,N_10146);
nor U15795 (N_15795,N_9669,N_9491);
or U15796 (N_15796,N_9367,N_9477);
or U15797 (N_15797,N_7290,N_12277);
nand U15798 (N_15798,N_7545,N_6388);
nand U15799 (N_15799,N_8543,N_11993);
and U15800 (N_15800,N_10816,N_10934);
nand U15801 (N_15801,N_11201,N_11158);
xnor U15802 (N_15802,N_6672,N_10259);
xnor U15803 (N_15803,N_6522,N_7557);
and U15804 (N_15804,N_8294,N_6329);
xor U15805 (N_15805,N_8298,N_7828);
and U15806 (N_15806,N_10924,N_6663);
nor U15807 (N_15807,N_10607,N_6511);
or U15808 (N_15808,N_6902,N_6948);
nor U15809 (N_15809,N_11488,N_9870);
xnor U15810 (N_15810,N_7187,N_7017);
nand U15811 (N_15811,N_8611,N_9971);
or U15812 (N_15812,N_7121,N_6588);
nand U15813 (N_15813,N_12442,N_10279);
nor U15814 (N_15814,N_11894,N_7399);
nor U15815 (N_15815,N_8112,N_8415);
nand U15816 (N_15816,N_6407,N_8520);
and U15817 (N_15817,N_10338,N_11920);
and U15818 (N_15818,N_7110,N_11616);
and U15819 (N_15819,N_12376,N_8823);
xnor U15820 (N_15820,N_11046,N_10025);
nor U15821 (N_15821,N_9748,N_10046);
nor U15822 (N_15822,N_10978,N_12024);
nand U15823 (N_15823,N_11777,N_7679);
nand U15824 (N_15824,N_7783,N_8368);
nor U15825 (N_15825,N_11804,N_9505);
xnor U15826 (N_15826,N_9104,N_9376);
or U15827 (N_15827,N_7323,N_10793);
or U15828 (N_15828,N_7930,N_6734);
and U15829 (N_15829,N_9899,N_10163);
nor U15830 (N_15830,N_6974,N_10308);
nand U15831 (N_15831,N_7783,N_10535);
and U15832 (N_15832,N_11981,N_8008);
nor U15833 (N_15833,N_6620,N_7917);
nand U15834 (N_15834,N_9948,N_11738);
or U15835 (N_15835,N_8937,N_9656);
xor U15836 (N_15836,N_8605,N_11520);
or U15837 (N_15837,N_8774,N_6257);
xnor U15838 (N_15838,N_11982,N_8949);
and U15839 (N_15839,N_6548,N_11807);
nor U15840 (N_15840,N_11011,N_12335);
nor U15841 (N_15841,N_9798,N_6483);
or U15842 (N_15842,N_8793,N_7601);
nand U15843 (N_15843,N_8795,N_10915);
nand U15844 (N_15844,N_11728,N_11015);
xnor U15845 (N_15845,N_11536,N_10568);
nor U15846 (N_15846,N_9635,N_10186);
nor U15847 (N_15847,N_7011,N_9130);
or U15848 (N_15848,N_10687,N_7403);
nand U15849 (N_15849,N_11336,N_8248);
nand U15850 (N_15850,N_10846,N_11880);
nand U15851 (N_15851,N_10540,N_9224);
xnor U15852 (N_15852,N_10165,N_10120);
nor U15853 (N_15853,N_11670,N_11130);
nor U15854 (N_15854,N_12063,N_7513);
or U15855 (N_15855,N_10587,N_11884);
nand U15856 (N_15856,N_12478,N_8535);
or U15857 (N_15857,N_9012,N_10442);
nor U15858 (N_15858,N_6744,N_12371);
and U15859 (N_15859,N_7023,N_8358);
or U15860 (N_15860,N_6758,N_9875);
nor U15861 (N_15861,N_8835,N_6383);
nand U15862 (N_15862,N_7132,N_8792);
nor U15863 (N_15863,N_7027,N_11118);
or U15864 (N_15864,N_7653,N_8697);
and U15865 (N_15865,N_9592,N_8239);
nand U15866 (N_15866,N_9440,N_8844);
or U15867 (N_15867,N_6283,N_11429);
or U15868 (N_15868,N_8926,N_10605);
xor U15869 (N_15869,N_9282,N_7589);
and U15870 (N_15870,N_7481,N_8782);
or U15871 (N_15871,N_6517,N_8546);
nor U15872 (N_15872,N_7524,N_7412);
nand U15873 (N_15873,N_9152,N_10588);
and U15874 (N_15874,N_10006,N_7372);
nand U15875 (N_15875,N_8471,N_7969);
nand U15876 (N_15876,N_6965,N_6937);
nor U15877 (N_15877,N_9018,N_10247);
and U15878 (N_15878,N_7965,N_10325);
and U15879 (N_15879,N_9919,N_7674);
and U15880 (N_15880,N_11110,N_12101);
or U15881 (N_15881,N_10305,N_9738);
nor U15882 (N_15882,N_6995,N_10943);
nand U15883 (N_15883,N_10378,N_6714);
nand U15884 (N_15884,N_7619,N_10780);
and U15885 (N_15885,N_11644,N_8410);
and U15886 (N_15886,N_11847,N_11506);
or U15887 (N_15887,N_9469,N_11144);
nor U15888 (N_15888,N_10964,N_11017);
nand U15889 (N_15889,N_11009,N_7230);
or U15890 (N_15890,N_10590,N_6637);
or U15891 (N_15891,N_10637,N_12082);
nor U15892 (N_15892,N_8397,N_8900);
nor U15893 (N_15893,N_12361,N_9328);
nor U15894 (N_15894,N_7262,N_11547);
xnor U15895 (N_15895,N_11103,N_10670);
and U15896 (N_15896,N_8558,N_10201);
and U15897 (N_15897,N_9370,N_9160);
and U15898 (N_15898,N_12154,N_8271);
nand U15899 (N_15899,N_11746,N_6935);
and U15900 (N_15900,N_7725,N_9046);
nor U15901 (N_15901,N_11969,N_9840);
or U15902 (N_15902,N_11357,N_10785);
and U15903 (N_15903,N_9100,N_8672);
nor U15904 (N_15904,N_12444,N_6564);
nor U15905 (N_15905,N_7071,N_12433);
or U15906 (N_15906,N_7024,N_6621);
nand U15907 (N_15907,N_12019,N_9296);
or U15908 (N_15908,N_11670,N_8563);
and U15909 (N_15909,N_7884,N_11429);
and U15910 (N_15910,N_10192,N_9751);
and U15911 (N_15911,N_7407,N_10558);
and U15912 (N_15912,N_9794,N_8230);
and U15913 (N_15913,N_8114,N_11342);
nor U15914 (N_15914,N_12181,N_8304);
nand U15915 (N_15915,N_6617,N_10385);
nand U15916 (N_15916,N_6785,N_11748);
and U15917 (N_15917,N_6748,N_10993);
xor U15918 (N_15918,N_10650,N_6863);
nand U15919 (N_15919,N_10382,N_9132);
nand U15920 (N_15920,N_7757,N_7164);
or U15921 (N_15921,N_10884,N_12277);
or U15922 (N_15922,N_11524,N_12410);
and U15923 (N_15923,N_9479,N_6922);
nand U15924 (N_15924,N_7215,N_7218);
and U15925 (N_15925,N_8279,N_6580);
or U15926 (N_15926,N_8650,N_11834);
nor U15927 (N_15927,N_12237,N_10944);
nand U15928 (N_15928,N_7001,N_12092);
nand U15929 (N_15929,N_12033,N_9070);
nand U15930 (N_15930,N_10445,N_7774);
nand U15931 (N_15931,N_9139,N_8941);
nor U15932 (N_15932,N_11913,N_11522);
and U15933 (N_15933,N_10639,N_7370);
nand U15934 (N_15934,N_8985,N_7569);
nand U15935 (N_15935,N_7434,N_8383);
and U15936 (N_15936,N_10421,N_10948);
and U15937 (N_15937,N_6370,N_11240);
nand U15938 (N_15938,N_8408,N_9546);
nand U15939 (N_15939,N_9843,N_8871);
xor U15940 (N_15940,N_11337,N_8707);
nor U15941 (N_15941,N_8161,N_9090);
nor U15942 (N_15942,N_12074,N_6705);
or U15943 (N_15943,N_8516,N_9981);
or U15944 (N_15944,N_6939,N_11829);
nor U15945 (N_15945,N_7214,N_11658);
and U15946 (N_15946,N_9609,N_7010);
nor U15947 (N_15947,N_10653,N_7444);
or U15948 (N_15948,N_10689,N_10854);
or U15949 (N_15949,N_9285,N_10876);
or U15950 (N_15950,N_10188,N_8281);
xor U15951 (N_15951,N_11397,N_6584);
nand U15952 (N_15952,N_6802,N_6402);
nor U15953 (N_15953,N_6630,N_8148);
xnor U15954 (N_15954,N_11019,N_8036);
nor U15955 (N_15955,N_6377,N_9548);
nand U15956 (N_15956,N_9577,N_12436);
nor U15957 (N_15957,N_10539,N_10954);
nor U15958 (N_15958,N_7263,N_10528);
or U15959 (N_15959,N_12129,N_6916);
and U15960 (N_15960,N_11489,N_8224);
and U15961 (N_15961,N_7116,N_9225);
xnor U15962 (N_15962,N_7185,N_8336);
and U15963 (N_15963,N_8413,N_9413);
and U15964 (N_15964,N_10674,N_12218);
or U15965 (N_15965,N_8765,N_9252);
and U15966 (N_15966,N_10622,N_7955);
or U15967 (N_15967,N_8121,N_7387);
or U15968 (N_15968,N_10460,N_6524);
nand U15969 (N_15969,N_11654,N_7213);
nor U15970 (N_15970,N_12440,N_12066);
xnor U15971 (N_15971,N_7441,N_10121);
nand U15972 (N_15972,N_7356,N_10512);
or U15973 (N_15973,N_8468,N_8961);
or U15974 (N_15974,N_9840,N_8376);
xnor U15975 (N_15975,N_10312,N_9332);
or U15976 (N_15976,N_8168,N_10071);
nor U15977 (N_15977,N_8787,N_10449);
nor U15978 (N_15978,N_10289,N_9878);
nor U15979 (N_15979,N_9222,N_9527);
nand U15980 (N_15980,N_7162,N_11154);
nor U15981 (N_15981,N_9574,N_7560);
or U15982 (N_15982,N_10291,N_6745);
or U15983 (N_15983,N_12161,N_11989);
xor U15984 (N_15984,N_8900,N_7211);
nand U15985 (N_15985,N_9932,N_12423);
or U15986 (N_15986,N_6730,N_9354);
nand U15987 (N_15987,N_11792,N_10118);
nand U15988 (N_15988,N_11433,N_12293);
nor U15989 (N_15989,N_6883,N_9984);
nand U15990 (N_15990,N_11107,N_11637);
and U15991 (N_15991,N_6893,N_11895);
and U15992 (N_15992,N_9427,N_6251);
nand U15993 (N_15993,N_9869,N_10758);
nor U15994 (N_15994,N_7936,N_6933);
or U15995 (N_15995,N_10186,N_8574);
or U15996 (N_15996,N_6905,N_6514);
nor U15997 (N_15997,N_9575,N_7403);
nor U15998 (N_15998,N_7382,N_9464);
and U15999 (N_15999,N_9600,N_10146);
or U16000 (N_16000,N_10285,N_6746);
nor U16001 (N_16001,N_12105,N_12399);
and U16002 (N_16002,N_7984,N_7246);
or U16003 (N_16003,N_12294,N_7548);
or U16004 (N_16004,N_6593,N_11880);
nand U16005 (N_16005,N_6900,N_11395);
xor U16006 (N_16006,N_11613,N_7712);
nand U16007 (N_16007,N_11709,N_8195);
and U16008 (N_16008,N_8698,N_12494);
and U16009 (N_16009,N_9639,N_10488);
nor U16010 (N_16010,N_9602,N_10253);
xor U16011 (N_16011,N_7847,N_11967);
nor U16012 (N_16012,N_11012,N_12465);
and U16013 (N_16013,N_7322,N_9957);
or U16014 (N_16014,N_6645,N_10420);
nor U16015 (N_16015,N_12038,N_8873);
xor U16016 (N_16016,N_9402,N_8081);
nand U16017 (N_16017,N_8339,N_11369);
nand U16018 (N_16018,N_8490,N_11127);
nor U16019 (N_16019,N_11979,N_7054);
nor U16020 (N_16020,N_11689,N_12411);
and U16021 (N_16021,N_7245,N_9568);
nand U16022 (N_16022,N_8244,N_10362);
nor U16023 (N_16023,N_11615,N_11593);
nand U16024 (N_16024,N_10558,N_10135);
and U16025 (N_16025,N_7290,N_12494);
nor U16026 (N_16026,N_12360,N_6885);
xor U16027 (N_16027,N_8023,N_9436);
nand U16028 (N_16028,N_9337,N_9509);
xor U16029 (N_16029,N_6467,N_10003);
nand U16030 (N_16030,N_11591,N_8928);
and U16031 (N_16031,N_6770,N_12254);
nor U16032 (N_16032,N_7912,N_8503);
or U16033 (N_16033,N_12115,N_7727);
or U16034 (N_16034,N_8368,N_8268);
or U16035 (N_16035,N_7587,N_8495);
nor U16036 (N_16036,N_11960,N_12089);
or U16037 (N_16037,N_11573,N_7712);
or U16038 (N_16038,N_8701,N_7507);
nor U16039 (N_16039,N_10514,N_10460);
or U16040 (N_16040,N_7246,N_6324);
and U16041 (N_16041,N_7265,N_9143);
nor U16042 (N_16042,N_7024,N_9768);
nor U16043 (N_16043,N_11597,N_11185);
and U16044 (N_16044,N_11435,N_11259);
or U16045 (N_16045,N_10193,N_10299);
or U16046 (N_16046,N_9783,N_12316);
nand U16047 (N_16047,N_10565,N_6390);
and U16048 (N_16048,N_9315,N_10235);
and U16049 (N_16049,N_7220,N_7452);
nand U16050 (N_16050,N_10495,N_8392);
and U16051 (N_16051,N_11366,N_8862);
nor U16052 (N_16052,N_7364,N_7832);
nor U16053 (N_16053,N_10055,N_6778);
nand U16054 (N_16054,N_11023,N_7244);
and U16055 (N_16055,N_8453,N_8484);
nor U16056 (N_16056,N_10950,N_6289);
xor U16057 (N_16057,N_9964,N_6872);
nor U16058 (N_16058,N_7108,N_11190);
and U16059 (N_16059,N_7037,N_9468);
or U16060 (N_16060,N_6921,N_11336);
xor U16061 (N_16061,N_10318,N_9612);
or U16062 (N_16062,N_11544,N_6513);
nor U16063 (N_16063,N_6447,N_12208);
or U16064 (N_16064,N_11597,N_9934);
or U16065 (N_16065,N_8436,N_7906);
or U16066 (N_16066,N_11742,N_10433);
nand U16067 (N_16067,N_7251,N_12131);
and U16068 (N_16068,N_9354,N_11864);
and U16069 (N_16069,N_11461,N_12220);
and U16070 (N_16070,N_9935,N_8521);
nand U16071 (N_16071,N_10488,N_12409);
nand U16072 (N_16072,N_7228,N_7400);
nor U16073 (N_16073,N_9386,N_10423);
or U16074 (N_16074,N_11241,N_10680);
xor U16075 (N_16075,N_11125,N_12456);
and U16076 (N_16076,N_6628,N_9602);
or U16077 (N_16077,N_10621,N_7999);
nor U16078 (N_16078,N_7836,N_12096);
or U16079 (N_16079,N_11180,N_7541);
or U16080 (N_16080,N_7303,N_6382);
nor U16081 (N_16081,N_10481,N_8028);
nand U16082 (N_16082,N_11974,N_11645);
nand U16083 (N_16083,N_6671,N_11218);
nand U16084 (N_16084,N_9345,N_7680);
and U16085 (N_16085,N_7916,N_8381);
nand U16086 (N_16086,N_11564,N_9869);
nand U16087 (N_16087,N_6598,N_10553);
or U16088 (N_16088,N_9952,N_7196);
nand U16089 (N_16089,N_10322,N_6443);
nand U16090 (N_16090,N_9902,N_10401);
and U16091 (N_16091,N_8710,N_9139);
nand U16092 (N_16092,N_10285,N_10900);
nor U16093 (N_16093,N_10904,N_7939);
nor U16094 (N_16094,N_8819,N_8712);
or U16095 (N_16095,N_11527,N_12340);
or U16096 (N_16096,N_8280,N_8065);
nand U16097 (N_16097,N_9438,N_9015);
xor U16098 (N_16098,N_9809,N_7369);
nor U16099 (N_16099,N_8654,N_11426);
or U16100 (N_16100,N_10007,N_7753);
and U16101 (N_16101,N_11910,N_8276);
nor U16102 (N_16102,N_11618,N_10443);
xor U16103 (N_16103,N_10014,N_7655);
or U16104 (N_16104,N_12030,N_11142);
nand U16105 (N_16105,N_6324,N_6534);
nor U16106 (N_16106,N_10569,N_6506);
nand U16107 (N_16107,N_10492,N_10217);
nand U16108 (N_16108,N_6881,N_10630);
and U16109 (N_16109,N_6401,N_8146);
xor U16110 (N_16110,N_7375,N_12315);
and U16111 (N_16111,N_9248,N_7650);
xnor U16112 (N_16112,N_8814,N_9387);
and U16113 (N_16113,N_7181,N_9867);
nor U16114 (N_16114,N_6457,N_7498);
and U16115 (N_16115,N_8150,N_8571);
or U16116 (N_16116,N_9567,N_10446);
or U16117 (N_16117,N_12034,N_11033);
or U16118 (N_16118,N_7403,N_7612);
and U16119 (N_16119,N_9731,N_7548);
xnor U16120 (N_16120,N_8579,N_9727);
nand U16121 (N_16121,N_10490,N_8560);
nand U16122 (N_16122,N_6610,N_7700);
nand U16123 (N_16123,N_7544,N_11520);
nand U16124 (N_16124,N_12297,N_11470);
xnor U16125 (N_16125,N_10835,N_7241);
nor U16126 (N_16126,N_11114,N_11595);
and U16127 (N_16127,N_6789,N_9893);
and U16128 (N_16128,N_9620,N_7439);
nor U16129 (N_16129,N_7527,N_8461);
nand U16130 (N_16130,N_7155,N_12239);
nand U16131 (N_16131,N_11396,N_7039);
nor U16132 (N_16132,N_7508,N_9744);
nand U16133 (N_16133,N_12086,N_10717);
and U16134 (N_16134,N_7159,N_8380);
nor U16135 (N_16135,N_11993,N_6431);
nor U16136 (N_16136,N_8877,N_8550);
nand U16137 (N_16137,N_10683,N_7313);
and U16138 (N_16138,N_7615,N_6649);
xnor U16139 (N_16139,N_7277,N_8551);
nor U16140 (N_16140,N_7955,N_11448);
nand U16141 (N_16141,N_11143,N_9445);
or U16142 (N_16142,N_8829,N_6709);
nand U16143 (N_16143,N_8305,N_10685);
nand U16144 (N_16144,N_11965,N_10708);
and U16145 (N_16145,N_12296,N_9080);
and U16146 (N_16146,N_9070,N_12203);
and U16147 (N_16147,N_9459,N_11286);
or U16148 (N_16148,N_9139,N_8718);
or U16149 (N_16149,N_12307,N_6360);
and U16150 (N_16150,N_6580,N_11863);
and U16151 (N_16151,N_11587,N_9110);
and U16152 (N_16152,N_7772,N_7839);
nor U16153 (N_16153,N_10672,N_10857);
or U16154 (N_16154,N_11694,N_10319);
nor U16155 (N_16155,N_8588,N_7604);
nand U16156 (N_16156,N_6334,N_10604);
or U16157 (N_16157,N_11459,N_10954);
or U16158 (N_16158,N_11704,N_10987);
nor U16159 (N_16159,N_10078,N_10814);
nand U16160 (N_16160,N_10453,N_9497);
nand U16161 (N_16161,N_9749,N_8603);
nand U16162 (N_16162,N_8394,N_9731);
nor U16163 (N_16163,N_9281,N_6978);
nand U16164 (N_16164,N_12465,N_10979);
or U16165 (N_16165,N_6634,N_7995);
nand U16166 (N_16166,N_6696,N_8681);
nor U16167 (N_16167,N_11824,N_8317);
and U16168 (N_16168,N_8126,N_6504);
or U16169 (N_16169,N_7522,N_11259);
or U16170 (N_16170,N_6581,N_8358);
nand U16171 (N_16171,N_11368,N_9620);
and U16172 (N_16172,N_12152,N_8060);
nand U16173 (N_16173,N_11748,N_12041);
nand U16174 (N_16174,N_7864,N_8123);
nor U16175 (N_16175,N_12325,N_7251);
and U16176 (N_16176,N_7734,N_9373);
nand U16177 (N_16177,N_8905,N_8426);
xnor U16178 (N_16178,N_8675,N_11226);
xnor U16179 (N_16179,N_7179,N_7228);
nor U16180 (N_16180,N_7045,N_10487);
and U16181 (N_16181,N_7055,N_6450);
nand U16182 (N_16182,N_8016,N_12494);
and U16183 (N_16183,N_10163,N_8107);
or U16184 (N_16184,N_11531,N_7860);
nand U16185 (N_16185,N_11103,N_10850);
nor U16186 (N_16186,N_9939,N_10677);
xor U16187 (N_16187,N_11961,N_7275);
or U16188 (N_16188,N_9783,N_11811);
nand U16189 (N_16189,N_11633,N_8107);
nor U16190 (N_16190,N_6416,N_8322);
xor U16191 (N_16191,N_11059,N_11292);
and U16192 (N_16192,N_11951,N_7220);
nand U16193 (N_16193,N_7778,N_11770);
or U16194 (N_16194,N_10864,N_8576);
or U16195 (N_16195,N_7652,N_7564);
and U16196 (N_16196,N_10918,N_9477);
nor U16197 (N_16197,N_9577,N_11038);
nand U16198 (N_16198,N_7960,N_8445);
nand U16199 (N_16199,N_11104,N_9198);
xor U16200 (N_16200,N_7813,N_11631);
xnor U16201 (N_16201,N_8813,N_11000);
nand U16202 (N_16202,N_10847,N_12318);
or U16203 (N_16203,N_10763,N_9069);
and U16204 (N_16204,N_7160,N_11052);
or U16205 (N_16205,N_11014,N_8348);
or U16206 (N_16206,N_11642,N_11479);
and U16207 (N_16207,N_12279,N_8532);
nor U16208 (N_16208,N_11127,N_9079);
or U16209 (N_16209,N_11000,N_11352);
xnor U16210 (N_16210,N_9452,N_9242);
nor U16211 (N_16211,N_8764,N_8589);
nand U16212 (N_16212,N_10019,N_11880);
nand U16213 (N_16213,N_10731,N_9526);
or U16214 (N_16214,N_9939,N_11158);
xor U16215 (N_16215,N_9447,N_12453);
or U16216 (N_16216,N_7204,N_10771);
xnor U16217 (N_16217,N_12234,N_10583);
nor U16218 (N_16218,N_7339,N_7070);
and U16219 (N_16219,N_7176,N_9955);
or U16220 (N_16220,N_7239,N_7467);
or U16221 (N_16221,N_11272,N_8175);
or U16222 (N_16222,N_6256,N_6959);
nor U16223 (N_16223,N_11106,N_9334);
nand U16224 (N_16224,N_8867,N_8862);
nor U16225 (N_16225,N_10977,N_9564);
and U16226 (N_16226,N_12186,N_6323);
nand U16227 (N_16227,N_6903,N_7928);
or U16228 (N_16228,N_7331,N_9683);
and U16229 (N_16229,N_9076,N_6620);
nand U16230 (N_16230,N_11929,N_6606);
nand U16231 (N_16231,N_12262,N_10764);
nor U16232 (N_16232,N_11901,N_7230);
and U16233 (N_16233,N_8390,N_11219);
nor U16234 (N_16234,N_12018,N_6774);
or U16235 (N_16235,N_6531,N_8344);
or U16236 (N_16236,N_10251,N_9400);
nor U16237 (N_16237,N_8001,N_8920);
or U16238 (N_16238,N_8991,N_9974);
nand U16239 (N_16239,N_11863,N_10210);
and U16240 (N_16240,N_10077,N_11768);
or U16241 (N_16241,N_11249,N_10472);
nor U16242 (N_16242,N_8636,N_7757);
and U16243 (N_16243,N_7325,N_7637);
nand U16244 (N_16244,N_6847,N_6882);
nand U16245 (N_16245,N_9313,N_10133);
and U16246 (N_16246,N_9206,N_8253);
or U16247 (N_16247,N_9800,N_11879);
or U16248 (N_16248,N_9793,N_10483);
and U16249 (N_16249,N_6920,N_11515);
nor U16250 (N_16250,N_11306,N_7604);
or U16251 (N_16251,N_12350,N_12111);
or U16252 (N_16252,N_12116,N_11877);
nand U16253 (N_16253,N_7480,N_10288);
xor U16254 (N_16254,N_11286,N_11504);
or U16255 (N_16255,N_10550,N_11655);
or U16256 (N_16256,N_12493,N_10663);
or U16257 (N_16257,N_7071,N_10475);
nand U16258 (N_16258,N_11884,N_10855);
nor U16259 (N_16259,N_7684,N_9708);
or U16260 (N_16260,N_10968,N_10693);
xor U16261 (N_16261,N_11573,N_8631);
nor U16262 (N_16262,N_12185,N_6560);
and U16263 (N_16263,N_11485,N_11333);
and U16264 (N_16264,N_10982,N_12394);
nor U16265 (N_16265,N_6902,N_7483);
or U16266 (N_16266,N_11811,N_10947);
and U16267 (N_16267,N_6775,N_10142);
and U16268 (N_16268,N_8145,N_12231);
nor U16269 (N_16269,N_10468,N_8535);
and U16270 (N_16270,N_12159,N_7201);
and U16271 (N_16271,N_10557,N_10597);
nand U16272 (N_16272,N_7012,N_9255);
xnor U16273 (N_16273,N_11332,N_8433);
nand U16274 (N_16274,N_7447,N_10524);
nand U16275 (N_16275,N_8688,N_12480);
nor U16276 (N_16276,N_8462,N_8159);
nand U16277 (N_16277,N_6326,N_6455);
xnor U16278 (N_16278,N_10622,N_11608);
or U16279 (N_16279,N_8554,N_12117);
and U16280 (N_16280,N_8890,N_7645);
and U16281 (N_16281,N_12047,N_9704);
xor U16282 (N_16282,N_11447,N_10661);
nor U16283 (N_16283,N_8807,N_8981);
nand U16284 (N_16284,N_6791,N_11488);
nor U16285 (N_16285,N_12185,N_9002);
xnor U16286 (N_16286,N_6755,N_11593);
and U16287 (N_16287,N_8121,N_8409);
nor U16288 (N_16288,N_8439,N_7795);
or U16289 (N_16289,N_6758,N_10735);
and U16290 (N_16290,N_8267,N_9394);
or U16291 (N_16291,N_8392,N_8371);
nand U16292 (N_16292,N_9118,N_11098);
and U16293 (N_16293,N_12151,N_7612);
nor U16294 (N_16294,N_10733,N_10972);
and U16295 (N_16295,N_12429,N_7051);
and U16296 (N_16296,N_10349,N_9486);
xnor U16297 (N_16297,N_11434,N_11189);
nand U16298 (N_16298,N_9657,N_11274);
nand U16299 (N_16299,N_9040,N_6631);
and U16300 (N_16300,N_11998,N_8718);
or U16301 (N_16301,N_6936,N_6773);
or U16302 (N_16302,N_10375,N_7755);
nor U16303 (N_16303,N_9074,N_10099);
nand U16304 (N_16304,N_10193,N_11615);
nor U16305 (N_16305,N_8845,N_10168);
or U16306 (N_16306,N_8049,N_7388);
or U16307 (N_16307,N_6267,N_6360);
and U16308 (N_16308,N_9293,N_10750);
xnor U16309 (N_16309,N_12459,N_7536);
nand U16310 (N_16310,N_12297,N_6280);
nor U16311 (N_16311,N_9567,N_10277);
nand U16312 (N_16312,N_8012,N_11017);
nor U16313 (N_16313,N_7292,N_6669);
nand U16314 (N_16314,N_9303,N_7892);
or U16315 (N_16315,N_7359,N_10294);
or U16316 (N_16316,N_9248,N_10307);
nand U16317 (N_16317,N_11982,N_6987);
and U16318 (N_16318,N_12319,N_10543);
nand U16319 (N_16319,N_9157,N_8746);
nand U16320 (N_16320,N_7310,N_7036);
and U16321 (N_16321,N_6903,N_11201);
nor U16322 (N_16322,N_10235,N_7204);
or U16323 (N_16323,N_9655,N_10685);
nand U16324 (N_16324,N_9554,N_9235);
or U16325 (N_16325,N_6318,N_8280);
nand U16326 (N_16326,N_11148,N_10591);
or U16327 (N_16327,N_9829,N_8103);
nor U16328 (N_16328,N_7024,N_9950);
and U16329 (N_16329,N_7434,N_7312);
or U16330 (N_16330,N_6360,N_10094);
nand U16331 (N_16331,N_7781,N_7046);
and U16332 (N_16332,N_9928,N_8607);
nor U16333 (N_16333,N_7615,N_9727);
or U16334 (N_16334,N_12385,N_9572);
nand U16335 (N_16335,N_7743,N_8408);
nand U16336 (N_16336,N_10596,N_9693);
and U16337 (N_16337,N_9050,N_9490);
xor U16338 (N_16338,N_7814,N_9085);
and U16339 (N_16339,N_12259,N_9101);
xnor U16340 (N_16340,N_10146,N_6910);
or U16341 (N_16341,N_6459,N_6270);
nand U16342 (N_16342,N_10086,N_10500);
nand U16343 (N_16343,N_10191,N_7722);
or U16344 (N_16344,N_11002,N_6722);
and U16345 (N_16345,N_6345,N_10732);
nand U16346 (N_16346,N_6576,N_6738);
nand U16347 (N_16347,N_8205,N_7351);
nor U16348 (N_16348,N_10164,N_7019);
xnor U16349 (N_16349,N_8742,N_9493);
nand U16350 (N_16350,N_8285,N_7284);
and U16351 (N_16351,N_7785,N_11631);
nand U16352 (N_16352,N_10904,N_10035);
or U16353 (N_16353,N_11653,N_6267);
xor U16354 (N_16354,N_11047,N_6407);
and U16355 (N_16355,N_9818,N_9473);
nor U16356 (N_16356,N_7193,N_9772);
xnor U16357 (N_16357,N_10397,N_11396);
nor U16358 (N_16358,N_6820,N_12495);
and U16359 (N_16359,N_11397,N_10853);
or U16360 (N_16360,N_6657,N_9390);
and U16361 (N_16361,N_9990,N_6780);
nor U16362 (N_16362,N_9686,N_11819);
nor U16363 (N_16363,N_10643,N_7410);
and U16364 (N_16364,N_8730,N_7645);
and U16365 (N_16365,N_12307,N_11069);
nor U16366 (N_16366,N_8770,N_7371);
or U16367 (N_16367,N_11657,N_8575);
or U16368 (N_16368,N_10513,N_8717);
and U16369 (N_16369,N_6494,N_9675);
or U16370 (N_16370,N_6579,N_8690);
and U16371 (N_16371,N_7759,N_11033);
and U16372 (N_16372,N_10200,N_9851);
nand U16373 (N_16373,N_12157,N_7030);
nor U16374 (N_16374,N_11897,N_7609);
xnor U16375 (N_16375,N_10644,N_7125);
nand U16376 (N_16376,N_9587,N_9236);
xor U16377 (N_16377,N_7395,N_9012);
nand U16378 (N_16378,N_12091,N_7579);
nand U16379 (N_16379,N_7226,N_6541);
or U16380 (N_16380,N_9887,N_8150);
nor U16381 (N_16381,N_9391,N_9307);
or U16382 (N_16382,N_11993,N_8283);
and U16383 (N_16383,N_9305,N_12223);
nor U16384 (N_16384,N_7884,N_6796);
and U16385 (N_16385,N_6523,N_10527);
nor U16386 (N_16386,N_10047,N_6580);
or U16387 (N_16387,N_10561,N_8247);
nor U16388 (N_16388,N_7241,N_11969);
and U16389 (N_16389,N_7108,N_9333);
or U16390 (N_16390,N_11277,N_7681);
or U16391 (N_16391,N_7907,N_8162);
nand U16392 (N_16392,N_10986,N_7056);
nor U16393 (N_16393,N_8863,N_11299);
nor U16394 (N_16394,N_8088,N_8578);
nand U16395 (N_16395,N_6430,N_9394);
nand U16396 (N_16396,N_9797,N_9939);
nand U16397 (N_16397,N_12466,N_7571);
and U16398 (N_16398,N_12097,N_10656);
nor U16399 (N_16399,N_7130,N_12290);
nor U16400 (N_16400,N_8416,N_9455);
and U16401 (N_16401,N_6369,N_7447);
nor U16402 (N_16402,N_10949,N_10102);
nor U16403 (N_16403,N_6383,N_6814);
or U16404 (N_16404,N_10116,N_10619);
or U16405 (N_16405,N_8543,N_7401);
or U16406 (N_16406,N_6483,N_6484);
or U16407 (N_16407,N_12353,N_7972);
nor U16408 (N_16408,N_7926,N_8134);
nor U16409 (N_16409,N_9605,N_6705);
nor U16410 (N_16410,N_6587,N_9433);
nor U16411 (N_16411,N_9907,N_9117);
nor U16412 (N_16412,N_9441,N_7583);
nand U16413 (N_16413,N_8671,N_7190);
and U16414 (N_16414,N_7596,N_6916);
or U16415 (N_16415,N_7500,N_10104);
or U16416 (N_16416,N_9360,N_10989);
and U16417 (N_16417,N_8884,N_12485);
nand U16418 (N_16418,N_8052,N_9144);
nand U16419 (N_16419,N_8928,N_10453);
or U16420 (N_16420,N_12176,N_11887);
nand U16421 (N_16421,N_10979,N_6888);
nor U16422 (N_16422,N_10706,N_10872);
nand U16423 (N_16423,N_10612,N_7516);
nand U16424 (N_16424,N_7712,N_9442);
nor U16425 (N_16425,N_11799,N_6563);
xor U16426 (N_16426,N_10397,N_10109);
nand U16427 (N_16427,N_11500,N_7191);
nor U16428 (N_16428,N_11817,N_8631);
nor U16429 (N_16429,N_11214,N_11045);
xor U16430 (N_16430,N_6631,N_8455);
nand U16431 (N_16431,N_9891,N_8433);
nand U16432 (N_16432,N_12421,N_12331);
and U16433 (N_16433,N_9538,N_8444);
xnor U16434 (N_16434,N_9215,N_7375);
nor U16435 (N_16435,N_6779,N_6251);
and U16436 (N_16436,N_10607,N_8617);
nand U16437 (N_16437,N_7527,N_10163);
and U16438 (N_16438,N_12111,N_7431);
or U16439 (N_16439,N_8341,N_9844);
or U16440 (N_16440,N_8611,N_7994);
nand U16441 (N_16441,N_7156,N_10641);
and U16442 (N_16442,N_11684,N_9939);
nor U16443 (N_16443,N_12325,N_7921);
and U16444 (N_16444,N_7946,N_9382);
nand U16445 (N_16445,N_6411,N_7666);
and U16446 (N_16446,N_12494,N_8847);
nor U16447 (N_16447,N_8553,N_12419);
nand U16448 (N_16448,N_10029,N_7906);
nor U16449 (N_16449,N_7783,N_7892);
and U16450 (N_16450,N_9570,N_6285);
nand U16451 (N_16451,N_8950,N_7396);
xor U16452 (N_16452,N_10370,N_7562);
and U16453 (N_16453,N_6310,N_8658);
xnor U16454 (N_16454,N_10774,N_7447);
and U16455 (N_16455,N_8303,N_10677);
nand U16456 (N_16456,N_8728,N_12181);
and U16457 (N_16457,N_11607,N_12173);
or U16458 (N_16458,N_11942,N_7025);
and U16459 (N_16459,N_9601,N_6802);
and U16460 (N_16460,N_10912,N_12488);
and U16461 (N_16461,N_12026,N_10902);
and U16462 (N_16462,N_10546,N_12155);
nand U16463 (N_16463,N_6795,N_8734);
nand U16464 (N_16464,N_9146,N_8469);
nor U16465 (N_16465,N_8804,N_9772);
and U16466 (N_16466,N_11865,N_8098);
and U16467 (N_16467,N_11102,N_11220);
or U16468 (N_16468,N_9689,N_6881);
or U16469 (N_16469,N_9014,N_8626);
or U16470 (N_16470,N_12394,N_7576);
and U16471 (N_16471,N_10827,N_11136);
nand U16472 (N_16472,N_8701,N_8230);
nor U16473 (N_16473,N_8125,N_10071);
and U16474 (N_16474,N_11532,N_10587);
and U16475 (N_16475,N_8863,N_11704);
and U16476 (N_16476,N_9380,N_10849);
and U16477 (N_16477,N_11919,N_9582);
nand U16478 (N_16478,N_11859,N_6307);
nand U16479 (N_16479,N_10872,N_10125);
nand U16480 (N_16480,N_9577,N_11000);
and U16481 (N_16481,N_10808,N_9674);
nand U16482 (N_16482,N_10457,N_7770);
nor U16483 (N_16483,N_12391,N_8748);
or U16484 (N_16484,N_12097,N_8591);
and U16485 (N_16485,N_10165,N_12137);
or U16486 (N_16486,N_8096,N_11271);
or U16487 (N_16487,N_8654,N_6869);
and U16488 (N_16488,N_9308,N_9757);
or U16489 (N_16489,N_6576,N_9265);
nor U16490 (N_16490,N_8891,N_10638);
and U16491 (N_16491,N_7212,N_9594);
and U16492 (N_16492,N_7600,N_11460);
nor U16493 (N_16493,N_12043,N_9998);
and U16494 (N_16494,N_12355,N_10774);
or U16495 (N_16495,N_6654,N_10513);
nor U16496 (N_16496,N_9230,N_11786);
nor U16497 (N_16497,N_10150,N_11561);
nand U16498 (N_16498,N_9622,N_9944);
nand U16499 (N_16499,N_11697,N_8757);
nand U16500 (N_16500,N_6901,N_7229);
or U16501 (N_16501,N_9207,N_10454);
nor U16502 (N_16502,N_7291,N_7308);
xor U16503 (N_16503,N_7250,N_10992);
xor U16504 (N_16504,N_11781,N_9801);
or U16505 (N_16505,N_10739,N_12268);
nand U16506 (N_16506,N_8014,N_7963);
and U16507 (N_16507,N_11347,N_11991);
xor U16508 (N_16508,N_6915,N_12413);
nor U16509 (N_16509,N_8686,N_6652);
nand U16510 (N_16510,N_7854,N_9993);
and U16511 (N_16511,N_12154,N_11989);
or U16512 (N_16512,N_7580,N_7805);
or U16513 (N_16513,N_8303,N_11539);
and U16514 (N_16514,N_9208,N_11076);
or U16515 (N_16515,N_12264,N_11106);
or U16516 (N_16516,N_12224,N_7985);
or U16517 (N_16517,N_9922,N_8696);
nor U16518 (N_16518,N_8708,N_12238);
xnor U16519 (N_16519,N_9488,N_9392);
nor U16520 (N_16520,N_7698,N_7502);
nand U16521 (N_16521,N_6938,N_10773);
nand U16522 (N_16522,N_7350,N_11978);
xnor U16523 (N_16523,N_9320,N_7266);
nor U16524 (N_16524,N_10644,N_10515);
xor U16525 (N_16525,N_6519,N_7918);
or U16526 (N_16526,N_7033,N_12439);
and U16527 (N_16527,N_6906,N_9093);
xnor U16528 (N_16528,N_7590,N_7596);
nand U16529 (N_16529,N_7968,N_12268);
or U16530 (N_16530,N_11148,N_9730);
or U16531 (N_16531,N_10405,N_6902);
nor U16532 (N_16532,N_9498,N_10507);
and U16533 (N_16533,N_8407,N_6720);
nor U16534 (N_16534,N_10335,N_6721);
and U16535 (N_16535,N_9558,N_6969);
and U16536 (N_16536,N_11189,N_11386);
nand U16537 (N_16537,N_11095,N_9759);
or U16538 (N_16538,N_7983,N_11518);
nor U16539 (N_16539,N_12337,N_6912);
nand U16540 (N_16540,N_10506,N_9131);
nor U16541 (N_16541,N_8239,N_10361);
nand U16542 (N_16542,N_11393,N_7594);
and U16543 (N_16543,N_9399,N_10948);
or U16544 (N_16544,N_7060,N_6252);
nand U16545 (N_16545,N_9463,N_8014);
nand U16546 (N_16546,N_10790,N_10824);
and U16547 (N_16547,N_7408,N_9955);
nand U16548 (N_16548,N_10637,N_7658);
nand U16549 (N_16549,N_6897,N_9624);
xnor U16550 (N_16550,N_7327,N_6901);
and U16551 (N_16551,N_7401,N_10035);
and U16552 (N_16552,N_10495,N_7972);
nand U16553 (N_16553,N_7492,N_9181);
xor U16554 (N_16554,N_7733,N_11689);
and U16555 (N_16555,N_7459,N_10739);
and U16556 (N_16556,N_9078,N_8636);
xnor U16557 (N_16557,N_7245,N_11072);
nor U16558 (N_16558,N_7259,N_10711);
and U16559 (N_16559,N_11471,N_6710);
nor U16560 (N_16560,N_11819,N_11190);
and U16561 (N_16561,N_7754,N_8921);
and U16562 (N_16562,N_11256,N_6866);
nand U16563 (N_16563,N_11716,N_11728);
and U16564 (N_16564,N_11623,N_6765);
nor U16565 (N_16565,N_12060,N_9209);
and U16566 (N_16566,N_11191,N_11681);
and U16567 (N_16567,N_9089,N_6494);
nand U16568 (N_16568,N_6613,N_10797);
and U16569 (N_16569,N_9876,N_8899);
nor U16570 (N_16570,N_11679,N_6760);
and U16571 (N_16571,N_9742,N_11094);
and U16572 (N_16572,N_9517,N_12110);
or U16573 (N_16573,N_8704,N_7002);
nand U16574 (N_16574,N_7903,N_9669);
nor U16575 (N_16575,N_8102,N_9475);
or U16576 (N_16576,N_11298,N_8716);
or U16577 (N_16577,N_7135,N_10119);
nor U16578 (N_16578,N_6371,N_8862);
nand U16579 (N_16579,N_6992,N_9569);
nor U16580 (N_16580,N_6508,N_7245);
nor U16581 (N_16581,N_11049,N_10825);
or U16582 (N_16582,N_7654,N_12325);
and U16583 (N_16583,N_7922,N_6795);
nand U16584 (N_16584,N_11742,N_12492);
or U16585 (N_16585,N_10914,N_11479);
nand U16586 (N_16586,N_11799,N_10245);
nand U16587 (N_16587,N_11735,N_9653);
and U16588 (N_16588,N_12110,N_7158);
and U16589 (N_16589,N_7386,N_12049);
nand U16590 (N_16590,N_10345,N_9192);
nor U16591 (N_16591,N_11103,N_9023);
nor U16592 (N_16592,N_12181,N_10060);
and U16593 (N_16593,N_11317,N_8889);
xnor U16594 (N_16594,N_11928,N_7075);
and U16595 (N_16595,N_11742,N_12279);
nand U16596 (N_16596,N_7954,N_8349);
nand U16597 (N_16597,N_7216,N_7025);
nor U16598 (N_16598,N_9789,N_10541);
nor U16599 (N_16599,N_7355,N_6273);
nand U16600 (N_16600,N_9528,N_10474);
nand U16601 (N_16601,N_7640,N_6907);
or U16602 (N_16602,N_11430,N_7395);
and U16603 (N_16603,N_11419,N_9900);
nor U16604 (N_16604,N_10741,N_12000);
xor U16605 (N_16605,N_6735,N_9273);
nor U16606 (N_16606,N_9593,N_12153);
and U16607 (N_16607,N_10913,N_12471);
and U16608 (N_16608,N_9306,N_11130);
nor U16609 (N_16609,N_9701,N_8460);
nand U16610 (N_16610,N_8427,N_8892);
nor U16611 (N_16611,N_10614,N_7112);
or U16612 (N_16612,N_11688,N_11682);
nand U16613 (N_16613,N_9464,N_6608);
nor U16614 (N_16614,N_6459,N_6357);
xor U16615 (N_16615,N_6486,N_6551);
xnor U16616 (N_16616,N_6895,N_11257);
and U16617 (N_16617,N_7738,N_10880);
and U16618 (N_16618,N_12027,N_11797);
and U16619 (N_16619,N_9632,N_10965);
and U16620 (N_16620,N_12402,N_9644);
nor U16621 (N_16621,N_10016,N_7391);
or U16622 (N_16622,N_8024,N_12371);
or U16623 (N_16623,N_9592,N_11347);
nand U16624 (N_16624,N_6475,N_11328);
or U16625 (N_16625,N_6415,N_12474);
and U16626 (N_16626,N_8211,N_7096);
and U16627 (N_16627,N_6954,N_8965);
nor U16628 (N_16628,N_11541,N_12312);
nor U16629 (N_16629,N_9662,N_10765);
or U16630 (N_16630,N_10645,N_10380);
xnor U16631 (N_16631,N_8953,N_9661);
nand U16632 (N_16632,N_8202,N_8473);
xor U16633 (N_16633,N_8550,N_12152);
nor U16634 (N_16634,N_10341,N_6993);
and U16635 (N_16635,N_10485,N_7602);
or U16636 (N_16636,N_7158,N_7352);
and U16637 (N_16637,N_10478,N_12153);
nand U16638 (N_16638,N_6987,N_6580);
or U16639 (N_16639,N_11136,N_11993);
and U16640 (N_16640,N_11783,N_10063);
or U16641 (N_16641,N_11542,N_9086);
nand U16642 (N_16642,N_10634,N_8562);
nor U16643 (N_16643,N_7774,N_9277);
or U16644 (N_16644,N_8387,N_7564);
or U16645 (N_16645,N_10675,N_8946);
and U16646 (N_16646,N_10112,N_7235);
nor U16647 (N_16647,N_7252,N_7840);
and U16648 (N_16648,N_11331,N_7393);
and U16649 (N_16649,N_8143,N_10670);
and U16650 (N_16650,N_12400,N_9505);
or U16651 (N_16651,N_8975,N_10624);
nor U16652 (N_16652,N_8253,N_9615);
nor U16653 (N_16653,N_11729,N_10004);
or U16654 (N_16654,N_8561,N_7281);
or U16655 (N_16655,N_10090,N_12426);
or U16656 (N_16656,N_8396,N_10359);
or U16657 (N_16657,N_9014,N_11962);
nand U16658 (N_16658,N_11752,N_7183);
and U16659 (N_16659,N_12315,N_6828);
xnor U16660 (N_16660,N_8170,N_12374);
xor U16661 (N_16661,N_9081,N_11668);
and U16662 (N_16662,N_8362,N_7132);
or U16663 (N_16663,N_11235,N_11887);
or U16664 (N_16664,N_9718,N_11465);
nand U16665 (N_16665,N_6595,N_8648);
or U16666 (N_16666,N_7792,N_11388);
xor U16667 (N_16667,N_7747,N_11007);
or U16668 (N_16668,N_10793,N_9461);
and U16669 (N_16669,N_6421,N_11140);
nor U16670 (N_16670,N_12251,N_6596);
or U16671 (N_16671,N_6662,N_6382);
nor U16672 (N_16672,N_8425,N_7847);
and U16673 (N_16673,N_10139,N_11841);
nand U16674 (N_16674,N_8530,N_7166);
nor U16675 (N_16675,N_12386,N_7461);
or U16676 (N_16676,N_7261,N_12167);
nand U16677 (N_16677,N_9871,N_10405);
or U16678 (N_16678,N_8190,N_10794);
nand U16679 (N_16679,N_11298,N_8163);
xor U16680 (N_16680,N_7668,N_12308);
or U16681 (N_16681,N_7811,N_6901);
and U16682 (N_16682,N_12182,N_8210);
and U16683 (N_16683,N_6471,N_9436);
nor U16684 (N_16684,N_6860,N_7406);
or U16685 (N_16685,N_8840,N_11686);
and U16686 (N_16686,N_8429,N_8984);
and U16687 (N_16687,N_8602,N_11624);
and U16688 (N_16688,N_8572,N_8850);
nand U16689 (N_16689,N_11594,N_12063);
xor U16690 (N_16690,N_10233,N_10940);
and U16691 (N_16691,N_7484,N_8041);
or U16692 (N_16692,N_11399,N_8606);
and U16693 (N_16693,N_7718,N_7008);
nand U16694 (N_16694,N_9255,N_8190);
nor U16695 (N_16695,N_12269,N_10151);
xnor U16696 (N_16696,N_7149,N_6951);
and U16697 (N_16697,N_12172,N_9778);
nand U16698 (N_16698,N_7142,N_10195);
nor U16699 (N_16699,N_6256,N_7928);
nand U16700 (N_16700,N_8644,N_8256);
and U16701 (N_16701,N_11111,N_9420);
nand U16702 (N_16702,N_7180,N_10867);
xor U16703 (N_16703,N_9091,N_10799);
xor U16704 (N_16704,N_6891,N_11681);
xor U16705 (N_16705,N_10053,N_7821);
and U16706 (N_16706,N_6345,N_7458);
and U16707 (N_16707,N_9295,N_8043);
or U16708 (N_16708,N_7021,N_7692);
nor U16709 (N_16709,N_12472,N_9480);
and U16710 (N_16710,N_6898,N_9559);
nand U16711 (N_16711,N_8317,N_7715);
nor U16712 (N_16712,N_11086,N_6432);
nor U16713 (N_16713,N_11593,N_12032);
nand U16714 (N_16714,N_12027,N_11666);
nand U16715 (N_16715,N_9232,N_9087);
nor U16716 (N_16716,N_12444,N_7431);
nand U16717 (N_16717,N_8845,N_12248);
and U16718 (N_16718,N_10698,N_11137);
and U16719 (N_16719,N_8140,N_12334);
and U16720 (N_16720,N_8858,N_9363);
and U16721 (N_16721,N_6735,N_12086);
nand U16722 (N_16722,N_8661,N_12156);
nor U16723 (N_16723,N_9152,N_7529);
nand U16724 (N_16724,N_11609,N_8327);
or U16725 (N_16725,N_7335,N_8532);
and U16726 (N_16726,N_8761,N_12184);
nor U16727 (N_16727,N_9542,N_12329);
or U16728 (N_16728,N_11856,N_12481);
nand U16729 (N_16729,N_7510,N_10308);
nand U16730 (N_16730,N_7222,N_10335);
xor U16731 (N_16731,N_10768,N_7557);
xor U16732 (N_16732,N_12475,N_11703);
or U16733 (N_16733,N_9739,N_6739);
and U16734 (N_16734,N_10061,N_12232);
nor U16735 (N_16735,N_7526,N_11950);
and U16736 (N_16736,N_8308,N_11540);
or U16737 (N_16737,N_8474,N_11339);
xor U16738 (N_16738,N_7234,N_8768);
and U16739 (N_16739,N_8638,N_9297);
and U16740 (N_16740,N_6326,N_11816);
and U16741 (N_16741,N_7862,N_10979);
xnor U16742 (N_16742,N_10130,N_11163);
nor U16743 (N_16743,N_10181,N_7549);
nand U16744 (N_16744,N_9955,N_9612);
and U16745 (N_16745,N_10385,N_10164);
nand U16746 (N_16746,N_7480,N_10620);
nand U16747 (N_16747,N_11360,N_11977);
nand U16748 (N_16748,N_10592,N_6370);
nor U16749 (N_16749,N_7949,N_6572);
or U16750 (N_16750,N_6668,N_10891);
and U16751 (N_16751,N_7995,N_12147);
nor U16752 (N_16752,N_7648,N_12084);
nor U16753 (N_16753,N_11379,N_8937);
nor U16754 (N_16754,N_10966,N_7492);
xor U16755 (N_16755,N_11933,N_9148);
or U16756 (N_16756,N_12277,N_9126);
and U16757 (N_16757,N_11419,N_12320);
nor U16758 (N_16758,N_6465,N_10841);
nand U16759 (N_16759,N_7477,N_10953);
and U16760 (N_16760,N_6672,N_8578);
or U16761 (N_16761,N_12411,N_9267);
and U16762 (N_16762,N_9446,N_11577);
or U16763 (N_16763,N_7553,N_6822);
nor U16764 (N_16764,N_9848,N_6729);
nor U16765 (N_16765,N_8414,N_7804);
and U16766 (N_16766,N_8817,N_10933);
nand U16767 (N_16767,N_9433,N_12422);
or U16768 (N_16768,N_12395,N_6733);
nor U16769 (N_16769,N_11963,N_10062);
or U16770 (N_16770,N_6475,N_6313);
and U16771 (N_16771,N_11669,N_9453);
or U16772 (N_16772,N_12078,N_7692);
nand U16773 (N_16773,N_11305,N_11035);
or U16774 (N_16774,N_12267,N_9756);
xor U16775 (N_16775,N_11424,N_10135);
nand U16776 (N_16776,N_11323,N_9029);
nor U16777 (N_16777,N_7629,N_12161);
or U16778 (N_16778,N_10320,N_11443);
or U16779 (N_16779,N_8075,N_7985);
and U16780 (N_16780,N_7610,N_9069);
and U16781 (N_16781,N_7602,N_11634);
nor U16782 (N_16782,N_10716,N_10056);
nand U16783 (N_16783,N_10882,N_6622);
and U16784 (N_16784,N_12342,N_10430);
nor U16785 (N_16785,N_11808,N_8523);
nand U16786 (N_16786,N_8248,N_10195);
nor U16787 (N_16787,N_9343,N_6279);
nor U16788 (N_16788,N_9069,N_8117);
and U16789 (N_16789,N_7097,N_10237);
nor U16790 (N_16790,N_11735,N_7593);
nand U16791 (N_16791,N_10962,N_6686);
or U16792 (N_16792,N_9062,N_8362);
nand U16793 (N_16793,N_6460,N_9577);
or U16794 (N_16794,N_8625,N_9198);
nand U16795 (N_16795,N_9387,N_6930);
and U16796 (N_16796,N_8823,N_7504);
and U16797 (N_16797,N_6626,N_10536);
or U16798 (N_16798,N_7271,N_9478);
and U16799 (N_16799,N_10553,N_7093);
nor U16800 (N_16800,N_11647,N_12488);
xnor U16801 (N_16801,N_10373,N_6653);
or U16802 (N_16802,N_9779,N_6594);
nor U16803 (N_16803,N_8416,N_7806);
nand U16804 (N_16804,N_7553,N_11360);
nor U16805 (N_16805,N_6435,N_8245);
nand U16806 (N_16806,N_12095,N_9362);
and U16807 (N_16807,N_11506,N_9671);
or U16808 (N_16808,N_11060,N_6888);
nand U16809 (N_16809,N_11339,N_9656);
and U16810 (N_16810,N_11414,N_10631);
nor U16811 (N_16811,N_10478,N_8329);
and U16812 (N_16812,N_11810,N_11251);
nand U16813 (N_16813,N_7190,N_9431);
and U16814 (N_16814,N_12457,N_11517);
nand U16815 (N_16815,N_7339,N_10747);
xnor U16816 (N_16816,N_7642,N_6670);
xnor U16817 (N_16817,N_7225,N_11855);
xnor U16818 (N_16818,N_11368,N_6476);
nand U16819 (N_16819,N_11911,N_8076);
xnor U16820 (N_16820,N_10532,N_7558);
or U16821 (N_16821,N_10509,N_9730);
nor U16822 (N_16822,N_8806,N_10782);
nand U16823 (N_16823,N_11471,N_11055);
nand U16824 (N_16824,N_11476,N_9796);
nand U16825 (N_16825,N_10111,N_11210);
nand U16826 (N_16826,N_11068,N_7967);
or U16827 (N_16827,N_9452,N_7984);
or U16828 (N_16828,N_11731,N_9240);
and U16829 (N_16829,N_10618,N_11280);
and U16830 (N_16830,N_9326,N_6655);
nor U16831 (N_16831,N_9535,N_8028);
or U16832 (N_16832,N_6855,N_8434);
xnor U16833 (N_16833,N_10973,N_7930);
nor U16834 (N_16834,N_7901,N_10749);
nor U16835 (N_16835,N_8549,N_12164);
nor U16836 (N_16836,N_10236,N_8199);
nor U16837 (N_16837,N_7021,N_12465);
nor U16838 (N_16838,N_6447,N_10149);
or U16839 (N_16839,N_10954,N_12187);
nor U16840 (N_16840,N_9522,N_11742);
and U16841 (N_16841,N_6596,N_7257);
or U16842 (N_16842,N_9545,N_6657);
and U16843 (N_16843,N_7709,N_9148);
nand U16844 (N_16844,N_6724,N_7068);
nand U16845 (N_16845,N_11723,N_9302);
nand U16846 (N_16846,N_7130,N_6254);
nand U16847 (N_16847,N_10595,N_6948);
and U16848 (N_16848,N_8240,N_8192);
and U16849 (N_16849,N_9128,N_10336);
or U16850 (N_16850,N_9425,N_7076);
and U16851 (N_16851,N_8352,N_8851);
xnor U16852 (N_16852,N_11912,N_6727);
nor U16853 (N_16853,N_10308,N_12295);
nand U16854 (N_16854,N_9929,N_10869);
xor U16855 (N_16855,N_9187,N_9102);
nand U16856 (N_16856,N_7678,N_6714);
xnor U16857 (N_16857,N_7407,N_10711);
and U16858 (N_16858,N_10034,N_7812);
or U16859 (N_16859,N_10979,N_6361);
and U16860 (N_16860,N_12193,N_6651);
nor U16861 (N_16861,N_7923,N_7228);
and U16862 (N_16862,N_8120,N_9092);
nor U16863 (N_16863,N_12062,N_8026);
nand U16864 (N_16864,N_7330,N_7362);
nand U16865 (N_16865,N_10469,N_9830);
nor U16866 (N_16866,N_7420,N_8464);
or U16867 (N_16867,N_6379,N_8098);
nor U16868 (N_16868,N_8227,N_9582);
or U16869 (N_16869,N_11363,N_12385);
nand U16870 (N_16870,N_12211,N_10167);
and U16871 (N_16871,N_10656,N_6835);
nor U16872 (N_16872,N_7908,N_11809);
nand U16873 (N_16873,N_11806,N_10275);
and U16874 (N_16874,N_7779,N_8615);
nand U16875 (N_16875,N_10664,N_11196);
nor U16876 (N_16876,N_10060,N_10241);
or U16877 (N_16877,N_11912,N_7858);
and U16878 (N_16878,N_9091,N_10798);
and U16879 (N_16879,N_12379,N_7301);
or U16880 (N_16880,N_8844,N_6382);
xnor U16881 (N_16881,N_12341,N_7345);
xnor U16882 (N_16882,N_8001,N_9712);
and U16883 (N_16883,N_9665,N_9876);
nor U16884 (N_16884,N_8483,N_10259);
or U16885 (N_16885,N_11116,N_9193);
and U16886 (N_16886,N_9431,N_7656);
or U16887 (N_16887,N_11337,N_6510);
nor U16888 (N_16888,N_11531,N_11343);
xnor U16889 (N_16889,N_10422,N_10315);
and U16890 (N_16890,N_11684,N_8931);
nor U16891 (N_16891,N_7917,N_7620);
nor U16892 (N_16892,N_9765,N_7861);
nor U16893 (N_16893,N_10598,N_10143);
or U16894 (N_16894,N_11580,N_9519);
nand U16895 (N_16895,N_6903,N_11096);
nand U16896 (N_16896,N_12272,N_6772);
xor U16897 (N_16897,N_8763,N_9344);
xor U16898 (N_16898,N_9798,N_10206);
nand U16899 (N_16899,N_9757,N_9171);
xnor U16900 (N_16900,N_8264,N_12295);
nand U16901 (N_16901,N_11411,N_6880);
and U16902 (N_16902,N_11119,N_9570);
and U16903 (N_16903,N_6772,N_11710);
nand U16904 (N_16904,N_7526,N_7950);
and U16905 (N_16905,N_12027,N_10087);
nor U16906 (N_16906,N_12243,N_11890);
nor U16907 (N_16907,N_7793,N_8296);
or U16908 (N_16908,N_11764,N_12280);
nor U16909 (N_16909,N_12028,N_11029);
and U16910 (N_16910,N_8151,N_12078);
nand U16911 (N_16911,N_6656,N_9210);
and U16912 (N_16912,N_6292,N_11336);
or U16913 (N_16913,N_7235,N_10214);
nand U16914 (N_16914,N_8731,N_9638);
or U16915 (N_16915,N_7426,N_11129);
or U16916 (N_16916,N_10595,N_9531);
and U16917 (N_16917,N_11866,N_6378);
xnor U16918 (N_16918,N_7545,N_10916);
and U16919 (N_16919,N_10017,N_6347);
nor U16920 (N_16920,N_10207,N_11940);
nor U16921 (N_16921,N_7629,N_6437);
or U16922 (N_16922,N_11774,N_10181);
nand U16923 (N_16923,N_6526,N_8003);
nand U16924 (N_16924,N_7964,N_10674);
and U16925 (N_16925,N_8485,N_12110);
or U16926 (N_16926,N_8598,N_10857);
nand U16927 (N_16927,N_8830,N_8999);
xnor U16928 (N_16928,N_7500,N_8484);
nand U16929 (N_16929,N_7976,N_10799);
and U16930 (N_16930,N_10282,N_12206);
and U16931 (N_16931,N_11342,N_11330);
nand U16932 (N_16932,N_11822,N_9089);
and U16933 (N_16933,N_10031,N_10468);
nand U16934 (N_16934,N_7148,N_9790);
and U16935 (N_16935,N_10414,N_10027);
or U16936 (N_16936,N_8908,N_10778);
xor U16937 (N_16937,N_12296,N_9044);
nor U16938 (N_16938,N_9939,N_6393);
and U16939 (N_16939,N_9231,N_10555);
and U16940 (N_16940,N_8618,N_6575);
or U16941 (N_16941,N_9757,N_7128);
nand U16942 (N_16942,N_11171,N_10585);
and U16943 (N_16943,N_9450,N_9699);
xor U16944 (N_16944,N_8435,N_8869);
nor U16945 (N_16945,N_11145,N_6832);
or U16946 (N_16946,N_7523,N_8279);
nand U16947 (N_16947,N_8456,N_11145);
nor U16948 (N_16948,N_10387,N_9149);
and U16949 (N_16949,N_11932,N_9755);
nor U16950 (N_16950,N_11805,N_11266);
and U16951 (N_16951,N_9111,N_10339);
and U16952 (N_16952,N_9765,N_7770);
xnor U16953 (N_16953,N_8496,N_9590);
or U16954 (N_16954,N_8832,N_12424);
nor U16955 (N_16955,N_7092,N_12117);
xnor U16956 (N_16956,N_12300,N_10676);
nor U16957 (N_16957,N_12103,N_11371);
xor U16958 (N_16958,N_7379,N_6497);
xor U16959 (N_16959,N_8042,N_10380);
and U16960 (N_16960,N_8030,N_6440);
and U16961 (N_16961,N_11285,N_10502);
xor U16962 (N_16962,N_9095,N_9477);
or U16963 (N_16963,N_9947,N_11447);
xnor U16964 (N_16964,N_9964,N_11288);
nand U16965 (N_16965,N_9801,N_11231);
or U16966 (N_16966,N_9530,N_11231);
nand U16967 (N_16967,N_8483,N_10361);
or U16968 (N_16968,N_7620,N_7864);
nor U16969 (N_16969,N_6812,N_11692);
nor U16970 (N_16970,N_12112,N_11211);
nor U16971 (N_16971,N_9523,N_8660);
nand U16972 (N_16972,N_11567,N_8877);
nand U16973 (N_16973,N_6276,N_9780);
and U16974 (N_16974,N_8542,N_11121);
or U16975 (N_16975,N_6592,N_7430);
and U16976 (N_16976,N_11365,N_7846);
xnor U16977 (N_16977,N_10306,N_10576);
and U16978 (N_16978,N_9044,N_12064);
and U16979 (N_16979,N_10666,N_7356);
nor U16980 (N_16980,N_6880,N_7379);
and U16981 (N_16981,N_6687,N_8692);
nor U16982 (N_16982,N_6634,N_6632);
and U16983 (N_16983,N_10323,N_9374);
and U16984 (N_16984,N_12291,N_7479);
nor U16985 (N_16985,N_9673,N_7996);
nand U16986 (N_16986,N_10727,N_7812);
and U16987 (N_16987,N_11958,N_7133);
nor U16988 (N_16988,N_9763,N_10613);
and U16989 (N_16989,N_9680,N_10451);
nand U16990 (N_16990,N_9221,N_7358);
xor U16991 (N_16991,N_8421,N_9715);
and U16992 (N_16992,N_11851,N_11771);
nand U16993 (N_16993,N_8376,N_8909);
xnor U16994 (N_16994,N_7087,N_12332);
or U16995 (N_16995,N_10109,N_10083);
xnor U16996 (N_16996,N_11622,N_12087);
and U16997 (N_16997,N_9527,N_12056);
or U16998 (N_16998,N_6669,N_11238);
and U16999 (N_16999,N_11137,N_10906);
nand U17000 (N_17000,N_11685,N_12382);
and U17001 (N_17001,N_12244,N_12018);
and U17002 (N_17002,N_12069,N_10978);
or U17003 (N_17003,N_9359,N_10427);
nor U17004 (N_17004,N_9129,N_8533);
xnor U17005 (N_17005,N_7994,N_7691);
xnor U17006 (N_17006,N_6643,N_12385);
and U17007 (N_17007,N_7360,N_11464);
xnor U17008 (N_17008,N_9737,N_10547);
nand U17009 (N_17009,N_7981,N_6598);
and U17010 (N_17010,N_10477,N_9880);
xor U17011 (N_17011,N_10318,N_12014);
xnor U17012 (N_17012,N_7592,N_12335);
or U17013 (N_17013,N_7859,N_8933);
nor U17014 (N_17014,N_11439,N_12031);
nand U17015 (N_17015,N_12452,N_11899);
nor U17016 (N_17016,N_8741,N_7056);
nor U17017 (N_17017,N_9729,N_9910);
and U17018 (N_17018,N_10598,N_12165);
nor U17019 (N_17019,N_10461,N_7493);
and U17020 (N_17020,N_9826,N_7451);
nor U17021 (N_17021,N_7135,N_10453);
or U17022 (N_17022,N_8285,N_8379);
nor U17023 (N_17023,N_10959,N_8823);
and U17024 (N_17024,N_9218,N_9593);
or U17025 (N_17025,N_11239,N_10946);
or U17026 (N_17026,N_10838,N_9348);
and U17027 (N_17027,N_8711,N_9425);
nor U17028 (N_17028,N_11596,N_7346);
and U17029 (N_17029,N_8670,N_8135);
nand U17030 (N_17030,N_11115,N_10658);
and U17031 (N_17031,N_6722,N_6474);
and U17032 (N_17032,N_11097,N_11988);
nor U17033 (N_17033,N_11325,N_6397);
or U17034 (N_17034,N_9306,N_7374);
nand U17035 (N_17035,N_7651,N_9707);
or U17036 (N_17036,N_8565,N_6571);
nor U17037 (N_17037,N_12377,N_9761);
nand U17038 (N_17038,N_11544,N_8965);
nand U17039 (N_17039,N_8241,N_12035);
or U17040 (N_17040,N_7800,N_7352);
nand U17041 (N_17041,N_7194,N_10420);
nand U17042 (N_17042,N_10353,N_8467);
xor U17043 (N_17043,N_6416,N_9468);
or U17044 (N_17044,N_7361,N_10637);
or U17045 (N_17045,N_12133,N_12006);
nand U17046 (N_17046,N_7734,N_12135);
and U17047 (N_17047,N_9952,N_10060);
nand U17048 (N_17048,N_11211,N_10621);
xnor U17049 (N_17049,N_10993,N_7643);
or U17050 (N_17050,N_10580,N_8303);
or U17051 (N_17051,N_11817,N_9814);
nand U17052 (N_17052,N_8070,N_6697);
or U17053 (N_17053,N_11720,N_7971);
nand U17054 (N_17054,N_9064,N_7775);
nand U17055 (N_17055,N_7480,N_10281);
nor U17056 (N_17056,N_12357,N_7873);
nor U17057 (N_17057,N_8347,N_6357);
nor U17058 (N_17058,N_6250,N_10465);
nand U17059 (N_17059,N_7363,N_11409);
nand U17060 (N_17060,N_6660,N_10999);
or U17061 (N_17061,N_11092,N_6767);
and U17062 (N_17062,N_7891,N_11884);
nor U17063 (N_17063,N_7667,N_6258);
and U17064 (N_17064,N_11492,N_12236);
xnor U17065 (N_17065,N_8920,N_9860);
and U17066 (N_17066,N_10039,N_9559);
or U17067 (N_17067,N_6308,N_7708);
and U17068 (N_17068,N_11998,N_7540);
nand U17069 (N_17069,N_9669,N_8133);
nand U17070 (N_17070,N_9632,N_12024);
xnor U17071 (N_17071,N_10927,N_6658);
nand U17072 (N_17072,N_10582,N_6853);
and U17073 (N_17073,N_11988,N_9961);
nor U17074 (N_17074,N_12377,N_8907);
or U17075 (N_17075,N_11043,N_11329);
nor U17076 (N_17076,N_7263,N_10526);
nand U17077 (N_17077,N_6362,N_9000);
nand U17078 (N_17078,N_11695,N_9566);
or U17079 (N_17079,N_7068,N_10922);
nand U17080 (N_17080,N_11007,N_8330);
nand U17081 (N_17081,N_12030,N_9336);
nor U17082 (N_17082,N_7920,N_11559);
xor U17083 (N_17083,N_7738,N_10700);
and U17084 (N_17084,N_12114,N_11367);
nor U17085 (N_17085,N_7660,N_9772);
and U17086 (N_17086,N_7178,N_9065);
xnor U17087 (N_17087,N_11034,N_10422);
and U17088 (N_17088,N_7921,N_7638);
nor U17089 (N_17089,N_11112,N_6449);
xor U17090 (N_17090,N_7535,N_12371);
or U17091 (N_17091,N_8315,N_8224);
nand U17092 (N_17092,N_8664,N_8439);
xor U17093 (N_17093,N_6836,N_10060);
or U17094 (N_17094,N_7500,N_7197);
nor U17095 (N_17095,N_7622,N_10069);
or U17096 (N_17096,N_10781,N_8780);
nor U17097 (N_17097,N_10045,N_6758);
xor U17098 (N_17098,N_10279,N_6328);
nand U17099 (N_17099,N_7619,N_11394);
nand U17100 (N_17100,N_11964,N_6701);
and U17101 (N_17101,N_8930,N_12011);
xor U17102 (N_17102,N_11141,N_10195);
and U17103 (N_17103,N_10903,N_10919);
nand U17104 (N_17104,N_11431,N_8636);
nand U17105 (N_17105,N_8258,N_9458);
nand U17106 (N_17106,N_11113,N_10219);
xor U17107 (N_17107,N_10820,N_6286);
xnor U17108 (N_17108,N_6511,N_7024);
nor U17109 (N_17109,N_7261,N_7192);
nor U17110 (N_17110,N_11030,N_11510);
xnor U17111 (N_17111,N_7377,N_8578);
nand U17112 (N_17112,N_10305,N_12479);
nand U17113 (N_17113,N_11253,N_11345);
nor U17114 (N_17114,N_9933,N_11429);
nor U17115 (N_17115,N_6436,N_8100);
or U17116 (N_17116,N_10172,N_11346);
nand U17117 (N_17117,N_8041,N_10374);
nand U17118 (N_17118,N_8671,N_11322);
nor U17119 (N_17119,N_11104,N_12175);
nand U17120 (N_17120,N_7180,N_8879);
nor U17121 (N_17121,N_6541,N_7336);
and U17122 (N_17122,N_6749,N_6626);
nor U17123 (N_17123,N_7755,N_6342);
or U17124 (N_17124,N_9967,N_8635);
nor U17125 (N_17125,N_8600,N_12240);
nor U17126 (N_17126,N_12394,N_11969);
nand U17127 (N_17127,N_10261,N_11846);
xor U17128 (N_17128,N_7355,N_6486);
nand U17129 (N_17129,N_10586,N_7991);
and U17130 (N_17130,N_10688,N_12176);
nand U17131 (N_17131,N_8535,N_9931);
or U17132 (N_17132,N_6362,N_9756);
nor U17133 (N_17133,N_8527,N_8643);
xnor U17134 (N_17134,N_6250,N_7649);
nor U17135 (N_17135,N_12473,N_9191);
nand U17136 (N_17136,N_12487,N_8468);
nand U17137 (N_17137,N_9883,N_10396);
nor U17138 (N_17138,N_12499,N_10225);
nand U17139 (N_17139,N_8814,N_6542);
nand U17140 (N_17140,N_11950,N_10055);
and U17141 (N_17141,N_9434,N_7121);
and U17142 (N_17142,N_12046,N_11759);
and U17143 (N_17143,N_8196,N_6765);
nand U17144 (N_17144,N_7747,N_11213);
or U17145 (N_17145,N_9944,N_8525);
and U17146 (N_17146,N_8105,N_7758);
or U17147 (N_17147,N_9529,N_8559);
xnor U17148 (N_17148,N_7596,N_7020);
or U17149 (N_17149,N_9321,N_10673);
and U17150 (N_17150,N_6931,N_8255);
or U17151 (N_17151,N_7615,N_11005);
or U17152 (N_17152,N_10380,N_11834);
nand U17153 (N_17153,N_9190,N_10174);
or U17154 (N_17154,N_11158,N_12038);
or U17155 (N_17155,N_6906,N_11207);
or U17156 (N_17156,N_12461,N_11734);
or U17157 (N_17157,N_6650,N_11256);
nor U17158 (N_17158,N_11282,N_9903);
nand U17159 (N_17159,N_9348,N_7260);
and U17160 (N_17160,N_12078,N_9086);
nor U17161 (N_17161,N_8957,N_10457);
nor U17162 (N_17162,N_12055,N_11321);
nand U17163 (N_17163,N_8020,N_10905);
or U17164 (N_17164,N_10065,N_7820);
nor U17165 (N_17165,N_8034,N_9350);
nand U17166 (N_17166,N_11844,N_9654);
or U17167 (N_17167,N_9622,N_6559);
nor U17168 (N_17168,N_11783,N_7991);
or U17169 (N_17169,N_10255,N_11709);
or U17170 (N_17170,N_11728,N_9756);
nor U17171 (N_17171,N_6472,N_7423);
nor U17172 (N_17172,N_9983,N_9134);
nor U17173 (N_17173,N_9584,N_8456);
and U17174 (N_17174,N_9332,N_8965);
and U17175 (N_17175,N_12445,N_10891);
nor U17176 (N_17176,N_8952,N_6748);
nor U17177 (N_17177,N_11889,N_12056);
and U17178 (N_17178,N_8679,N_9815);
xnor U17179 (N_17179,N_10254,N_9128);
nor U17180 (N_17180,N_7874,N_6799);
and U17181 (N_17181,N_6886,N_9358);
and U17182 (N_17182,N_12463,N_11483);
nor U17183 (N_17183,N_9656,N_6737);
nand U17184 (N_17184,N_12019,N_7516);
and U17185 (N_17185,N_7415,N_12399);
or U17186 (N_17186,N_9154,N_12126);
nor U17187 (N_17187,N_11010,N_8977);
nor U17188 (N_17188,N_8136,N_12254);
nor U17189 (N_17189,N_11472,N_7578);
or U17190 (N_17190,N_6563,N_8559);
and U17191 (N_17191,N_12433,N_12116);
nor U17192 (N_17192,N_11761,N_11907);
nand U17193 (N_17193,N_8538,N_11778);
xnor U17194 (N_17194,N_10861,N_10388);
xor U17195 (N_17195,N_9032,N_12486);
nor U17196 (N_17196,N_9054,N_8219);
xor U17197 (N_17197,N_8635,N_7586);
or U17198 (N_17198,N_6388,N_8684);
nand U17199 (N_17199,N_12243,N_9913);
nor U17200 (N_17200,N_9069,N_6329);
nand U17201 (N_17201,N_10809,N_12154);
or U17202 (N_17202,N_10075,N_10306);
nand U17203 (N_17203,N_9276,N_12487);
nor U17204 (N_17204,N_8438,N_10870);
or U17205 (N_17205,N_8824,N_7904);
and U17206 (N_17206,N_6498,N_8601);
nand U17207 (N_17207,N_9805,N_6720);
xor U17208 (N_17208,N_7334,N_10695);
or U17209 (N_17209,N_9944,N_8967);
or U17210 (N_17210,N_9626,N_8685);
and U17211 (N_17211,N_9636,N_10173);
nand U17212 (N_17212,N_7883,N_7206);
nor U17213 (N_17213,N_7272,N_11193);
and U17214 (N_17214,N_12465,N_8973);
nor U17215 (N_17215,N_11045,N_7294);
or U17216 (N_17216,N_10992,N_9117);
or U17217 (N_17217,N_9426,N_9742);
xnor U17218 (N_17218,N_7817,N_10282);
nor U17219 (N_17219,N_11380,N_11571);
or U17220 (N_17220,N_10651,N_11732);
or U17221 (N_17221,N_11518,N_10968);
or U17222 (N_17222,N_7524,N_11202);
or U17223 (N_17223,N_11774,N_6314);
or U17224 (N_17224,N_7058,N_11780);
or U17225 (N_17225,N_10380,N_10920);
nor U17226 (N_17226,N_7847,N_12405);
xnor U17227 (N_17227,N_9665,N_8066);
xor U17228 (N_17228,N_8744,N_12002);
nor U17229 (N_17229,N_7872,N_8001);
nor U17230 (N_17230,N_7643,N_11112);
and U17231 (N_17231,N_9854,N_7682);
nor U17232 (N_17232,N_12379,N_7072);
nor U17233 (N_17233,N_8830,N_9972);
or U17234 (N_17234,N_7989,N_8764);
nand U17235 (N_17235,N_8900,N_11775);
nand U17236 (N_17236,N_9273,N_9668);
nor U17237 (N_17237,N_11064,N_10826);
nor U17238 (N_17238,N_9522,N_10078);
nor U17239 (N_17239,N_10849,N_8264);
or U17240 (N_17240,N_11534,N_8559);
nor U17241 (N_17241,N_11006,N_12410);
nor U17242 (N_17242,N_10529,N_8671);
nand U17243 (N_17243,N_9266,N_6965);
xnor U17244 (N_17244,N_9175,N_11690);
or U17245 (N_17245,N_12488,N_6517);
nand U17246 (N_17246,N_9004,N_9065);
xnor U17247 (N_17247,N_6846,N_12233);
nand U17248 (N_17248,N_7191,N_10833);
or U17249 (N_17249,N_6652,N_12282);
and U17250 (N_17250,N_11834,N_11894);
nor U17251 (N_17251,N_9118,N_7365);
or U17252 (N_17252,N_10107,N_6795);
nor U17253 (N_17253,N_8012,N_7250);
nor U17254 (N_17254,N_9768,N_7598);
or U17255 (N_17255,N_12467,N_8585);
nor U17256 (N_17256,N_7558,N_10820);
or U17257 (N_17257,N_8168,N_10929);
nor U17258 (N_17258,N_10668,N_7603);
or U17259 (N_17259,N_6897,N_7526);
nand U17260 (N_17260,N_7335,N_9225);
nor U17261 (N_17261,N_7974,N_10771);
nand U17262 (N_17262,N_8118,N_8988);
nor U17263 (N_17263,N_6831,N_7230);
and U17264 (N_17264,N_12455,N_10674);
nor U17265 (N_17265,N_6287,N_6530);
nor U17266 (N_17266,N_9684,N_9543);
and U17267 (N_17267,N_12192,N_9052);
and U17268 (N_17268,N_6384,N_10242);
and U17269 (N_17269,N_9297,N_10330);
nand U17270 (N_17270,N_9660,N_8965);
and U17271 (N_17271,N_9142,N_7180);
or U17272 (N_17272,N_8306,N_6912);
nand U17273 (N_17273,N_8659,N_9465);
nor U17274 (N_17274,N_6734,N_11563);
xor U17275 (N_17275,N_7920,N_8626);
nand U17276 (N_17276,N_6480,N_7334);
nand U17277 (N_17277,N_8319,N_9173);
nor U17278 (N_17278,N_6464,N_6421);
and U17279 (N_17279,N_6452,N_10401);
nand U17280 (N_17280,N_6987,N_9806);
nand U17281 (N_17281,N_10419,N_8908);
and U17282 (N_17282,N_8653,N_9339);
nor U17283 (N_17283,N_9365,N_10209);
and U17284 (N_17284,N_8733,N_11841);
nor U17285 (N_17285,N_12290,N_10865);
nand U17286 (N_17286,N_9748,N_6266);
xnor U17287 (N_17287,N_9886,N_10170);
nand U17288 (N_17288,N_10708,N_12208);
or U17289 (N_17289,N_12286,N_8928);
nor U17290 (N_17290,N_10585,N_11428);
nand U17291 (N_17291,N_6292,N_11716);
and U17292 (N_17292,N_12037,N_12358);
nor U17293 (N_17293,N_7303,N_8101);
nor U17294 (N_17294,N_9516,N_9661);
and U17295 (N_17295,N_11392,N_7349);
nor U17296 (N_17296,N_11362,N_10201);
or U17297 (N_17297,N_9277,N_6657);
or U17298 (N_17298,N_8710,N_12292);
and U17299 (N_17299,N_8660,N_6361);
and U17300 (N_17300,N_7095,N_10610);
xor U17301 (N_17301,N_11507,N_7136);
or U17302 (N_17302,N_8332,N_8718);
nand U17303 (N_17303,N_10902,N_10179);
nand U17304 (N_17304,N_9268,N_8081);
and U17305 (N_17305,N_9871,N_10424);
and U17306 (N_17306,N_7283,N_10924);
or U17307 (N_17307,N_12412,N_6825);
and U17308 (N_17308,N_6523,N_6953);
or U17309 (N_17309,N_9798,N_9283);
or U17310 (N_17310,N_7446,N_10235);
xor U17311 (N_17311,N_7356,N_8495);
and U17312 (N_17312,N_8090,N_7725);
and U17313 (N_17313,N_6684,N_9067);
or U17314 (N_17314,N_6487,N_7104);
and U17315 (N_17315,N_8498,N_7593);
and U17316 (N_17316,N_11647,N_9339);
and U17317 (N_17317,N_9711,N_10730);
or U17318 (N_17318,N_9180,N_6416);
or U17319 (N_17319,N_8231,N_7715);
nand U17320 (N_17320,N_10463,N_10370);
nand U17321 (N_17321,N_12286,N_10709);
xor U17322 (N_17322,N_8625,N_7028);
or U17323 (N_17323,N_7085,N_10909);
and U17324 (N_17324,N_11821,N_12373);
or U17325 (N_17325,N_9444,N_9368);
and U17326 (N_17326,N_12190,N_6932);
nor U17327 (N_17327,N_10639,N_9081);
xnor U17328 (N_17328,N_6576,N_10676);
and U17329 (N_17329,N_10032,N_7228);
nor U17330 (N_17330,N_7938,N_7372);
nand U17331 (N_17331,N_7275,N_8936);
nor U17332 (N_17332,N_6944,N_11351);
and U17333 (N_17333,N_11055,N_10963);
nor U17334 (N_17334,N_7730,N_11627);
nor U17335 (N_17335,N_11049,N_11299);
or U17336 (N_17336,N_11408,N_8679);
nand U17337 (N_17337,N_10993,N_10744);
or U17338 (N_17338,N_11834,N_6621);
nor U17339 (N_17339,N_6883,N_9936);
and U17340 (N_17340,N_10787,N_10301);
and U17341 (N_17341,N_6541,N_12059);
nand U17342 (N_17342,N_6653,N_8614);
xnor U17343 (N_17343,N_10302,N_8857);
or U17344 (N_17344,N_6722,N_11814);
nor U17345 (N_17345,N_11458,N_9677);
or U17346 (N_17346,N_8260,N_8931);
or U17347 (N_17347,N_10568,N_12387);
nor U17348 (N_17348,N_7236,N_8624);
nor U17349 (N_17349,N_7382,N_10266);
and U17350 (N_17350,N_10571,N_8747);
nor U17351 (N_17351,N_9732,N_11473);
and U17352 (N_17352,N_9652,N_9963);
nand U17353 (N_17353,N_10366,N_8455);
nand U17354 (N_17354,N_9006,N_12428);
and U17355 (N_17355,N_6564,N_8786);
nor U17356 (N_17356,N_9781,N_8477);
nand U17357 (N_17357,N_12099,N_7024);
nand U17358 (N_17358,N_9327,N_7591);
nor U17359 (N_17359,N_8070,N_10098);
nor U17360 (N_17360,N_6643,N_11943);
nor U17361 (N_17361,N_8854,N_11002);
nand U17362 (N_17362,N_9697,N_11934);
and U17363 (N_17363,N_6703,N_9134);
nand U17364 (N_17364,N_8528,N_7853);
xnor U17365 (N_17365,N_10440,N_11811);
nor U17366 (N_17366,N_8581,N_9888);
or U17367 (N_17367,N_9093,N_6763);
nand U17368 (N_17368,N_10437,N_10904);
nand U17369 (N_17369,N_6934,N_6688);
nor U17370 (N_17370,N_10925,N_10120);
and U17371 (N_17371,N_10859,N_11834);
and U17372 (N_17372,N_8145,N_12491);
nand U17373 (N_17373,N_10759,N_8985);
xor U17374 (N_17374,N_7427,N_9795);
or U17375 (N_17375,N_11125,N_10561);
nor U17376 (N_17376,N_7282,N_8726);
or U17377 (N_17377,N_12360,N_8490);
and U17378 (N_17378,N_7359,N_12471);
nor U17379 (N_17379,N_9580,N_7715);
or U17380 (N_17380,N_7636,N_11205);
nor U17381 (N_17381,N_9834,N_10973);
or U17382 (N_17382,N_9503,N_12030);
or U17383 (N_17383,N_8525,N_8182);
nand U17384 (N_17384,N_7769,N_7637);
nor U17385 (N_17385,N_9656,N_6949);
xor U17386 (N_17386,N_6465,N_11413);
nor U17387 (N_17387,N_10206,N_10116);
and U17388 (N_17388,N_11463,N_12081);
nor U17389 (N_17389,N_9605,N_10039);
and U17390 (N_17390,N_10362,N_10037);
and U17391 (N_17391,N_9403,N_11071);
and U17392 (N_17392,N_7414,N_7212);
nor U17393 (N_17393,N_6902,N_9627);
xnor U17394 (N_17394,N_9905,N_12313);
nand U17395 (N_17395,N_6621,N_11801);
nand U17396 (N_17396,N_10655,N_7930);
nor U17397 (N_17397,N_8734,N_8202);
and U17398 (N_17398,N_9898,N_8521);
nor U17399 (N_17399,N_11457,N_11496);
or U17400 (N_17400,N_6852,N_9271);
xor U17401 (N_17401,N_7887,N_9401);
nor U17402 (N_17402,N_12026,N_6307);
or U17403 (N_17403,N_8956,N_11226);
and U17404 (N_17404,N_6372,N_7460);
nor U17405 (N_17405,N_6937,N_7780);
nand U17406 (N_17406,N_11519,N_9921);
nand U17407 (N_17407,N_8664,N_10818);
and U17408 (N_17408,N_9686,N_7646);
and U17409 (N_17409,N_10379,N_8161);
nand U17410 (N_17410,N_9625,N_8710);
xnor U17411 (N_17411,N_7749,N_12467);
nand U17412 (N_17412,N_10391,N_8870);
and U17413 (N_17413,N_9492,N_9094);
and U17414 (N_17414,N_10661,N_8590);
or U17415 (N_17415,N_7579,N_11306);
nor U17416 (N_17416,N_6439,N_11669);
nand U17417 (N_17417,N_7037,N_8284);
or U17418 (N_17418,N_8507,N_6787);
or U17419 (N_17419,N_10217,N_11153);
nor U17420 (N_17420,N_7950,N_11343);
and U17421 (N_17421,N_10060,N_10553);
and U17422 (N_17422,N_11773,N_9418);
and U17423 (N_17423,N_10259,N_10674);
nor U17424 (N_17424,N_9657,N_11845);
nor U17425 (N_17425,N_6799,N_6290);
and U17426 (N_17426,N_9788,N_7201);
nor U17427 (N_17427,N_9758,N_12436);
and U17428 (N_17428,N_9616,N_8424);
nand U17429 (N_17429,N_6971,N_10110);
nand U17430 (N_17430,N_7084,N_8729);
nand U17431 (N_17431,N_7070,N_7523);
nand U17432 (N_17432,N_12099,N_9120);
xnor U17433 (N_17433,N_8563,N_11610);
nand U17434 (N_17434,N_11258,N_8399);
nor U17435 (N_17435,N_7527,N_9187);
or U17436 (N_17436,N_7064,N_8218);
nand U17437 (N_17437,N_11258,N_8317);
xor U17438 (N_17438,N_7391,N_11251);
nand U17439 (N_17439,N_8970,N_8110);
nor U17440 (N_17440,N_12386,N_9412);
and U17441 (N_17441,N_9367,N_8260);
and U17442 (N_17442,N_11680,N_8711);
xor U17443 (N_17443,N_10706,N_11734);
nand U17444 (N_17444,N_7400,N_8112);
nor U17445 (N_17445,N_8628,N_9718);
and U17446 (N_17446,N_6505,N_10276);
or U17447 (N_17447,N_6546,N_7771);
and U17448 (N_17448,N_8324,N_11834);
nand U17449 (N_17449,N_6298,N_12412);
or U17450 (N_17450,N_11727,N_10161);
or U17451 (N_17451,N_12377,N_11747);
or U17452 (N_17452,N_10227,N_8840);
and U17453 (N_17453,N_7590,N_10290);
and U17454 (N_17454,N_6889,N_9653);
or U17455 (N_17455,N_12422,N_6614);
or U17456 (N_17456,N_6740,N_8995);
and U17457 (N_17457,N_10976,N_7803);
nand U17458 (N_17458,N_6767,N_11382);
nand U17459 (N_17459,N_12469,N_10981);
nand U17460 (N_17460,N_9231,N_10679);
or U17461 (N_17461,N_6624,N_7652);
nand U17462 (N_17462,N_10501,N_6548);
nand U17463 (N_17463,N_7751,N_8746);
xor U17464 (N_17464,N_10599,N_11079);
and U17465 (N_17465,N_7405,N_7913);
and U17466 (N_17466,N_7276,N_8439);
and U17467 (N_17467,N_6950,N_8509);
or U17468 (N_17468,N_7928,N_9558);
nor U17469 (N_17469,N_8852,N_7008);
and U17470 (N_17470,N_8756,N_7727);
xor U17471 (N_17471,N_8605,N_9476);
xor U17472 (N_17472,N_7362,N_11394);
and U17473 (N_17473,N_11608,N_9140);
nand U17474 (N_17474,N_6421,N_8403);
xor U17475 (N_17475,N_9071,N_7114);
or U17476 (N_17476,N_9664,N_6906);
or U17477 (N_17477,N_10634,N_6780);
or U17478 (N_17478,N_9630,N_11827);
or U17479 (N_17479,N_7163,N_8293);
or U17480 (N_17480,N_8858,N_7920);
nand U17481 (N_17481,N_10097,N_7366);
or U17482 (N_17482,N_12172,N_9324);
or U17483 (N_17483,N_9812,N_7594);
nor U17484 (N_17484,N_10571,N_7900);
nor U17485 (N_17485,N_8908,N_6662);
nand U17486 (N_17486,N_11005,N_9874);
nor U17487 (N_17487,N_9914,N_6477);
and U17488 (N_17488,N_6399,N_10356);
or U17489 (N_17489,N_6573,N_8783);
and U17490 (N_17490,N_6354,N_11484);
and U17491 (N_17491,N_7366,N_12333);
nand U17492 (N_17492,N_7308,N_10395);
nor U17493 (N_17493,N_11459,N_9326);
xor U17494 (N_17494,N_8616,N_8567);
and U17495 (N_17495,N_10222,N_8873);
or U17496 (N_17496,N_9304,N_10994);
and U17497 (N_17497,N_8126,N_10804);
nor U17498 (N_17498,N_8284,N_11972);
nand U17499 (N_17499,N_10802,N_9845);
nor U17500 (N_17500,N_8273,N_9523);
and U17501 (N_17501,N_8832,N_7769);
nor U17502 (N_17502,N_10629,N_7719);
or U17503 (N_17503,N_6494,N_8089);
or U17504 (N_17504,N_8854,N_9743);
or U17505 (N_17505,N_8062,N_12405);
or U17506 (N_17506,N_6441,N_9982);
nand U17507 (N_17507,N_9401,N_10061);
nor U17508 (N_17508,N_12084,N_8924);
xnor U17509 (N_17509,N_11880,N_6807);
nand U17510 (N_17510,N_9864,N_9386);
nand U17511 (N_17511,N_6686,N_6350);
or U17512 (N_17512,N_11421,N_7540);
or U17513 (N_17513,N_12463,N_7070);
nand U17514 (N_17514,N_7012,N_9025);
nor U17515 (N_17515,N_11023,N_11789);
nand U17516 (N_17516,N_6726,N_6457);
or U17517 (N_17517,N_10075,N_7446);
nand U17518 (N_17518,N_10670,N_6863);
or U17519 (N_17519,N_8504,N_12167);
and U17520 (N_17520,N_10328,N_9661);
and U17521 (N_17521,N_10196,N_11264);
or U17522 (N_17522,N_8001,N_8194);
and U17523 (N_17523,N_7528,N_6737);
nor U17524 (N_17524,N_10920,N_10402);
or U17525 (N_17525,N_8785,N_10863);
or U17526 (N_17526,N_9613,N_6733);
nor U17527 (N_17527,N_7670,N_11100);
or U17528 (N_17528,N_11573,N_7911);
nor U17529 (N_17529,N_9407,N_7607);
nor U17530 (N_17530,N_12436,N_7361);
nand U17531 (N_17531,N_11471,N_10746);
nor U17532 (N_17532,N_10812,N_8356);
nor U17533 (N_17533,N_7641,N_6779);
or U17534 (N_17534,N_8925,N_7239);
nor U17535 (N_17535,N_12262,N_12456);
nor U17536 (N_17536,N_6386,N_6760);
nor U17537 (N_17537,N_8743,N_6644);
or U17538 (N_17538,N_8379,N_9375);
and U17539 (N_17539,N_8711,N_6690);
or U17540 (N_17540,N_10006,N_10445);
or U17541 (N_17541,N_12338,N_7232);
and U17542 (N_17542,N_8380,N_9569);
nor U17543 (N_17543,N_8777,N_9705);
and U17544 (N_17544,N_12277,N_7799);
nand U17545 (N_17545,N_10965,N_6935);
nand U17546 (N_17546,N_7836,N_8185);
nor U17547 (N_17547,N_7100,N_7551);
or U17548 (N_17548,N_7958,N_8802);
or U17549 (N_17549,N_6557,N_11331);
nor U17550 (N_17550,N_7009,N_11641);
and U17551 (N_17551,N_6394,N_10673);
nand U17552 (N_17552,N_12069,N_8596);
or U17553 (N_17553,N_7530,N_10674);
nor U17554 (N_17554,N_10873,N_11919);
nand U17555 (N_17555,N_9056,N_9156);
nor U17556 (N_17556,N_11667,N_11158);
nor U17557 (N_17557,N_9852,N_11185);
or U17558 (N_17558,N_7341,N_8980);
and U17559 (N_17559,N_12354,N_9875);
or U17560 (N_17560,N_9486,N_9580);
and U17561 (N_17561,N_10278,N_12484);
nand U17562 (N_17562,N_7362,N_7704);
or U17563 (N_17563,N_9199,N_12206);
nor U17564 (N_17564,N_10628,N_6655);
and U17565 (N_17565,N_9911,N_12475);
nor U17566 (N_17566,N_9675,N_8538);
xnor U17567 (N_17567,N_9369,N_11380);
and U17568 (N_17568,N_12110,N_6862);
nor U17569 (N_17569,N_8346,N_9924);
nor U17570 (N_17570,N_11402,N_12083);
nor U17571 (N_17571,N_9946,N_6717);
nand U17572 (N_17572,N_11296,N_7672);
nor U17573 (N_17573,N_9011,N_10457);
nand U17574 (N_17574,N_11814,N_7517);
or U17575 (N_17575,N_8952,N_7625);
or U17576 (N_17576,N_9160,N_6256);
or U17577 (N_17577,N_11333,N_10533);
or U17578 (N_17578,N_11511,N_9747);
or U17579 (N_17579,N_9345,N_11967);
nand U17580 (N_17580,N_11762,N_10939);
xnor U17581 (N_17581,N_11623,N_7887);
nor U17582 (N_17582,N_10882,N_11846);
nand U17583 (N_17583,N_11249,N_7754);
nand U17584 (N_17584,N_12221,N_12444);
nor U17585 (N_17585,N_7241,N_8283);
nor U17586 (N_17586,N_7516,N_8431);
or U17587 (N_17587,N_12295,N_8556);
nor U17588 (N_17588,N_11304,N_9383);
nand U17589 (N_17589,N_6616,N_8252);
nand U17590 (N_17590,N_7676,N_12476);
nand U17591 (N_17591,N_8071,N_7409);
and U17592 (N_17592,N_11508,N_7982);
nand U17593 (N_17593,N_11743,N_8085);
nand U17594 (N_17594,N_7533,N_9425);
or U17595 (N_17595,N_6629,N_11294);
or U17596 (N_17596,N_9187,N_6801);
or U17597 (N_17597,N_10534,N_8237);
nor U17598 (N_17598,N_7171,N_9867);
xnor U17599 (N_17599,N_7463,N_9351);
nor U17600 (N_17600,N_11740,N_8594);
or U17601 (N_17601,N_8575,N_11837);
or U17602 (N_17602,N_11032,N_9531);
or U17603 (N_17603,N_9817,N_8115);
or U17604 (N_17604,N_9333,N_9007);
xor U17605 (N_17605,N_11643,N_11691);
xor U17606 (N_17606,N_10917,N_7977);
nand U17607 (N_17607,N_10117,N_10757);
nor U17608 (N_17608,N_10443,N_10772);
and U17609 (N_17609,N_9700,N_7749);
nand U17610 (N_17610,N_7317,N_12469);
or U17611 (N_17611,N_7319,N_9355);
nand U17612 (N_17612,N_10012,N_11525);
xnor U17613 (N_17613,N_11664,N_9156);
nor U17614 (N_17614,N_11535,N_11706);
and U17615 (N_17615,N_8636,N_7346);
and U17616 (N_17616,N_10471,N_9632);
nor U17617 (N_17617,N_12153,N_8862);
nand U17618 (N_17618,N_8161,N_9577);
nand U17619 (N_17619,N_6420,N_7170);
nor U17620 (N_17620,N_11794,N_10824);
nand U17621 (N_17621,N_9474,N_10523);
nor U17622 (N_17622,N_9052,N_8679);
nand U17623 (N_17623,N_11152,N_12337);
nor U17624 (N_17624,N_11352,N_8856);
and U17625 (N_17625,N_11105,N_9788);
and U17626 (N_17626,N_10644,N_11894);
nand U17627 (N_17627,N_7238,N_10534);
nor U17628 (N_17628,N_10486,N_8108);
and U17629 (N_17629,N_7963,N_10341);
and U17630 (N_17630,N_10813,N_10505);
nand U17631 (N_17631,N_10329,N_8137);
and U17632 (N_17632,N_11672,N_12436);
nand U17633 (N_17633,N_11879,N_11952);
and U17634 (N_17634,N_11035,N_11307);
and U17635 (N_17635,N_7504,N_8031);
nor U17636 (N_17636,N_8858,N_9928);
and U17637 (N_17637,N_9971,N_10060);
and U17638 (N_17638,N_8424,N_7453);
nor U17639 (N_17639,N_6270,N_7100);
xor U17640 (N_17640,N_7416,N_9121);
nand U17641 (N_17641,N_12336,N_9022);
or U17642 (N_17642,N_9408,N_9300);
or U17643 (N_17643,N_12068,N_10783);
or U17644 (N_17644,N_11594,N_11944);
nand U17645 (N_17645,N_6516,N_12143);
xor U17646 (N_17646,N_8396,N_11311);
nor U17647 (N_17647,N_7150,N_10971);
nand U17648 (N_17648,N_12063,N_11085);
nand U17649 (N_17649,N_10923,N_6778);
nand U17650 (N_17650,N_9670,N_10853);
or U17651 (N_17651,N_11518,N_11569);
or U17652 (N_17652,N_9911,N_6868);
or U17653 (N_17653,N_11110,N_8209);
nand U17654 (N_17654,N_9810,N_9518);
nor U17655 (N_17655,N_12252,N_8243);
and U17656 (N_17656,N_8928,N_12325);
nor U17657 (N_17657,N_8015,N_7089);
xor U17658 (N_17658,N_9106,N_6532);
or U17659 (N_17659,N_9226,N_6382);
and U17660 (N_17660,N_8937,N_10284);
xor U17661 (N_17661,N_10964,N_11396);
nand U17662 (N_17662,N_10855,N_12156);
and U17663 (N_17663,N_8615,N_7399);
nand U17664 (N_17664,N_11983,N_7306);
nand U17665 (N_17665,N_6764,N_8960);
nor U17666 (N_17666,N_8181,N_7398);
nand U17667 (N_17667,N_11711,N_8875);
nand U17668 (N_17668,N_6283,N_7544);
and U17669 (N_17669,N_8034,N_9279);
nand U17670 (N_17670,N_10032,N_9555);
and U17671 (N_17671,N_9944,N_7822);
or U17672 (N_17672,N_8881,N_11991);
nand U17673 (N_17673,N_11125,N_11824);
nor U17674 (N_17674,N_9597,N_8142);
or U17675 (N_17675,N_9538,N_9322);
nor U17676 (N_17676,N_11598,N_8739);
or U17677 (N_17677,N_9971,N_9099);
xor U17678 (N_17678,N_6893,N_7175);
nor U17679 (N_17679,N_10224,N_7978);
nand U17680 (N_17680,N_11257,N_7636);
nand U17681 (N_17681,N_8141,N_7719);
or U17682 (N_17682,N_9336,N_7760);
nand U17683 (N_17683,N_10791,N_8413);
and U17684 (N_17684,N_10149,N_11298);
xnor U17685 (N_17685,N_8032,N_9997);
nor U17686 (N_17686,N_7272,N_9189);
and U17687 (N_17687,N_10135,N_11924);
and U17688 (N_17688,N_8061,N_12472);
and U17689 (N_17689,N_7837,N_7883);
and U17690 (N_17690,N_10382,N_6783);
nor U17691 (N_17691,N_7697,N_9938);
nor U17692 (N_17692,N_10954,N_7330);
nand U17693 (N_17693,N_7327,N_9921);
and U17694 (N_17694,N_9488,N_12101);
nor U17695 (N_17695,N_10970,N_12223);
or U17696 (N_17696,N_8237,N_9887);
nand U17697 (N_17697,N_8520,N_8833);
and U17698 (N_17698,N_10411,N_8754);
and U17699 (N_17699,N_9891,N_7481);
nand U17700 (N_17700,N_12455,N_7546);
and U17701 (N_17701,N_11247,N_7490);
nor U17702 (N_17702,N_12405,N_9377);
nand U17703 (N_17703,N_8505,N_9349);
xor U17704 (N_17704,N_11968,N_6862);
or U17705 (N_17705,N_10584,N_8291);
nand U17706 (N_17706,N_11756,N_6850);
or U17707 (N_17707,N_8706,N_12256);
and U17708 (N_17708,N_7343,N_11950);
and U17709 (N_17709,N_11925,N_8126);
or U17710 (N_17710,N_8405,N_6544);
and U17711 (N_17711,N_7238,N_7182);
nor U17712 (N_17712,N_11380,N_7909);
and U17713 (N_17713,N_10861,N_8399);
nor U17714 (N_17714,N_10971,N_11614);
and U17715 (N_17715,N_10940,N_10399);
nand U17716 (N_17716,N_6795,N_11568);
nor U17717 (N_17717,N_6844,N_11575);
and U17718 (N_17718,N_9763,N_10276);
and U17719 (N_17719,N_11594,N_9608);
and U17720 (N_17720,N_12329,N_6490);
and U17721 (N_17721,N_11977,N_11575);
nor U17722 (N_17722,N_9929,N_9803);
or U17723 (N_17723,N_8349,N_6734);
nor U17724 (N_17724,N_10654,N_6825);
or U17725 (N_17725,N_9341,N_6976);
xor U17726 (N_17726,N_8195,N_9421);
or U17727 (N_17727,N_6916,N_7665);
or U17728 (N_17728,N_7783,N_8305);
and U17729 (N_17729,N_12339,N_8420);
or U17730 (N_17730,N_12269,N_12031);
nor U17731 (N_17731,N_8789,N_10473);
nand U17732 (N_17732,N_11754,N_10760);
or U17733 (N_17733,N_6584,N_11296);
nand U17734 (N_17734,N_6648,N_9112);
or U17735 (N_17735,N_10223,N_6606);
nor U17736 (N_17736,N_10686,N_9311);
and U17737 (N_17737,N_9000,N_9588);
nand U17738 (N_17738,N_10849,N_8844);
nor U17739 (N_17739,N_7759,N_8958);
nand U17740 (N_17740,N_8423,N_11108);
nand U17741 (N_17741,N_9796,N_10900);
and U17742 (N_17742,N_9306,N_10387);
or U17743 (N_17743,N_12344,N_10750);
xnor U17744 (N_17744,N_11895,N_12390);
and U17745 (N_17745,N_12470,N_12232);
and U17746 (N_17746,N_9489,N_6812);
nor U17747 (N_17747,N_10779,N_7542);
nand U17748 (N_17748,N_9729,N_7421);
xor U17749 (N_17749,N_7831,N_12291);
xor U17750 (N_17750,N_11684,N_11566);
nand U17751 (N_17751,N_8280,N_7205);
or U17752 (N_17752,N_10987,N_8809);
or U17753 (N_17753,N_6398,N_8872);
nand U17754 (N_17754,N_9137,N_7593);
nor U17755 (N_17755,N_6750,N_11870);
and U17756 (N_17756,N_12235,N_10131);
and U17757 (N_17757,N_8657,N_12484);
nand U17758 (N_17758,N_9762,N_7718);
nor U17759 (N_17759,N_10804,N_10990);
or U17760 (N_17760,N_8508,N_7033);
or U17761 (N_17761,N_6313,N_11437);
nand U17762 (N_17762,N_10467,N_12228);
or U17763 (N_17763,N_11685,N_6808);
nor U17764 (N_17764,N_7912,N_8309);
and U17765 (N_17765,N_9601,N_6664);
nand U17766 (N_17766,N_9830,N_6966);
nand U17767 (N_17767,N_9725,N_9632);
nand U17768 (N_17768,N_8445,N_7995);
and U17769 (N_17769,N_10740,N_7806);
or U17770 (N_17770,N_10890,N_10482);
nand U17771 (N_17771,N_11981,N_8350);
nor U17772 (N_17772,N_8184,N_9047);
or U17773 (N_17773,N_11001,N_12187);
or U17774 (N_17774,N_10915,N_9399);
nor U17775 (N_17775,N_10945,N_11983);
or U17776 (N_17776,N_9473,N_12394);
nor U17777 (N_17777,N_6784,N_10095);
or U17778 (N_17778,N_9469,N_11993);
nor U17779 (N_17779,N_8148,N_7737);
nor U17780 (N_17780,N_10795,N_7234);
xnor U17781 (N_17781,N_9960,N_6401);
and U17782 (N_17782,N_11957,N_11326);
nor U17783 (N_17783,N_12213,N_6519);
or U17784 (N_17784,N_12240,N_10640);
xor U17785 (N_17785,N_9992,N_10017);
nand U17786 (N_17786,N_9486,N_10491);
xnor U17787 (N_17787,N_6471,N_11593);
nor U17788 (N_17788,N_10323,N_8541);
xnor U17789 (N_17789,N_6274,N_10869);
nor U17790 (N_17790,N_11097,N_11846);
xor U17791 (N_17791,N_9235,N_10822);
and U17792 (N_17792,N_9030,N_8871);
or U17793 (N_17793,N_7827,N_7994);
or U17794 (N_17794,N_11659,N_7317);
or U17795 (N_17795,N_11180,N_11736);
and U17796 (N_17796,N_6943,N_12174);
nand U17797 (N_17797,N_9688,N_11693);
or U17798 (N_17798,N_8999,N_10628);
nor U17799 (N_17799,N_9487,N_11379);
nand U17800 (N_17800,N_12038,N_12384);
xor U17801 (N_17801,N_11177,N_7985);
and U17802 (N_17802,N_6613,N_12024);
nand U17803 (N_17803,N_10043,N_6723);
xor U17804 (N_17804,N_11714,N_7054);
nor U17805 (N_17805,N_11309,N_9634);
nand U17806 (N_17806,N_6634,N_6421);
or U17807 (N_17807,N_7001,N_9474);
nor U17808 (N_17808,N_9294,N_10505);
xor U17809 (N_17809,N_10534,N_10518);
xor U17810 (N_17810,N_7034,N_9333);
and U17811 (N_17811,N_7430,N_9055);
nand U17812 (N_17812,N_12120,N_9451);
nor U17813 (N_17813,N_9031,N_7980);
and U17814 (N_17814,N_8680,N_7348);
nor U17815 (N_17815,N_9083,N_8800);
nor U17816 (N_17816,N_11860,N_9153);
and U17817 (N_17817,N_9053,N_11589);
or U17818 (N_17818,N_8812,N_7957);
or U17819 (N_17819,N_8042,N_6298);
nor U17820 (N_17820,N_8160,N_6964);
and U17821 (N_17821,N_11302,N_10961);
nor U17822 (N_17822,N_10875,N_11959);
or U17823 (N_17823,N_7202,N_9880);
and U17824 (N_17824,N_10997,N_11416);
nand U17825 (N_17825,N_8583,N_12235);
and U17826 (N_17826,N_8558,N_9348);
nor U17827 (N_17827,N_6433,N_11801);
nand U17828 (N_17828,N_8190,N_11334);
nand U17829 (N_17829,N_9087,N_7996);
or U17830 (N_17830,N_12331,N_10328);
or U17831 (N_17831,N_6999,N_9858);
nand U17832 (N_17832,N_6675,N_6640);
and U17833 (N_17833,N_8490,N_11170);
nor U17834 (N_17834,N_10339,N_6494);
nand U17835 (N_17835,N_9717,N_11569);
or U17836 (N_17836,N_9843,N_6629);
nor U17837 (N_17837,N_10983,N_7974);
nor U17838 (N_17838,N_9072,N_11814);
nor U17839 (N_17839,N_10213,N_12090);
nor U17840 (N_17840,N_6699,N_7088);
or U17841 (N_17841,N_7195,N_10852);
nand U17842 (N_17842,N_9348,N_11325);
and U17843 (N_17843,N_10196,N_8458);
nor U17844 (N_17844,N_7194,N_10157);
xnor U17845 (N_17845,N_9686,N_6493);
nor U17846 (N_17846,N_9809,N_6531);
or U17847 (N_17847,N_10522,N_8906);
or U17848 (N_17848,N_10926,N_7546);
nand U17849 (N_17849,N_9712,N_11280);
or U17850 (N_17850,N_9665,N_11486);
or U17851 (N_17851,N_6545,N_9281);
and U17852 (N_17852,N_7809,N_8477);
or U17853 (N_17853,N_9660,N_10782);
and U17854 (N_17854,N_9922,N_9496);
nor U17855 (N_17855,N_6714,N_9365);
xnor U17856 (N_17856,N_10686,N_7056);
and U17857 (N_17857,N_9095,N_9831);
or U17858 (N_17858,N_10573,N_11850);
nand U17859 (N_17859,N_8629,N_9035);
nand U17860 (N_17860,N_10504,N_9139);
and U17861 (N_17861,N_11816,N_12261);
or U17862 (N_17862,N_10093,N_11171);
and U17863 (N_17863,N_10186,N_8605);
or U17864 (N_17864,N_6769,N_6695);
and U17865 (N_17865,N_9479,N_8201);
and U17866 (N_17866,N_8591,N_12296);
xnor U17867 (N_17867,N_10762,N_11656);
nor U17868 (N_17868,N_12087,N_8813);
or U17869 (N_17869,N_7955,N_6318);
and U17870 (N_17870,N_8859,N_9445);
nor U17871 (N_17871,N_8607,N_7931);
and U17872 (N_17872,N_7773,N_9633);
nand U17873 (N_17873,N_9953,N_12386);
or U17874 (N_17874,N_9765,N_8732);
or U17875 (N_17875,N_10002,N_11484);
and U17876 (N_17876,N_9628,N_10641);
nor U17877 (N_17877,N_7674,N_11167);
xnor U17878 (N_17878,N_8357,N_7480);
nor U17879 (N_17879,N_7400,N_7504);
or U17880 (N_17880,N_7435,N_7883);
nor U17881 (N_17881,N_8435,N_7696);
nor U17882 (N_17882,N_6865,N_11031);
nand U17883 (N_17883,N_10796,N_12038);
nand U17884 (N_17884,N_6741,N_9828);
or U17885 (N_17885,N_8030,N_10327);
xnor U17886 (N_17886,N_9966,N_11337);
nor U17887 (N_17887,N_9112,N_8763);
nor U17888 (N_17888,N_6757,N_8038);
xor U17889 (N_17889,N_11052,N_7507);
xnor U17890 (N_17890,N_9871,N_7860);
and U17891 (N_17891,N_7021,N_7629);
nand U17892 (N_17892,N_7416,N_6432);
nand U17893 (N_17893,N_9873,N_11354);
and U17894 (N_17894,N_11950,N_7410);
and U17895 (N_17895,N_11432,N_7849);
nor U17896 (N_17896,N_7781,N_8399);
nand U17897 (N_17897,N_9329,N_8459);
xor U17898 (N_17898,N_8687,N_12465);
nand U17899 (N_17899,N_8687,N_8698);
and U17900 (N_17900,N_8993,N_6693);
or U17901 (N_17901,N_6778,N_11765);
nand U17902 (N_17902,N_7407,N_8459);
or U17903 (N_17903,N_8620,N_11786);
and U17904 (N_17904,N_11803,N_9220);
nand U17905 (N_17905,N_11944,N_8355);
nor U17906 (N_17906,N_11302,N_7794);
nor U17907 (N_17907,N_6768,N_10782);
nor U17908 (N_17908,N_8077,N_11336);
and U17909 (N_17909,N_8112,N_8990);
nor U17910 (N_17910,N_9322,N_7222);
nand U17911 (N_17911,N_8573,N_8335);
nor U17912 (N_17912,N_8581,N_10895);
nand U17913 (N_17913,N_10893,N_12413);
nor U17914 (N_17914,N_8200,N_11141);
nand U17915 (N_17915,N_6631,N_10918);
nor U17916 (N_17916,N_6585,N_6870);
nand U17917 (N_17917,N_11118,N_11910);
nor U17918 (N_17918,N_6437,N_10987);
nand U17919 (N_17919,N_9899,N_7673);
nor U17920 (N_17920,N_10329,N_9292);
and U17921 (N_17921,N_7377,N_9658);
nand U17922 (N_17922,N_7357,N_9667);
nor U17923 (N_17923,N_6374,N_11223);
or U17924 (N_17924,N_12478,N_7749);
or U17925 (N_17925,N_12184,N_7254);
xnor U17926 (N_17926,N_11948,N_7010);
nand U17927 (N_17927,N_11485,N_7007);
and U17928 (N_17928,N_9021,N_9539);
and U17929 (N_17929,N_10735,N_11197);
and U17930 (N_17930,N_11223,N_8082);
or U17931 (N_17931,N_6534,N_11701);
nand U17932 (N_17932,N_9721,N_7579);
xor U17933 (N_17933,N_9266,N_9867);
nand U17934 (N_17934,N_11263,N_9492);
nand U17935 (N_17935,N_8225,N_7096);
and U17936 (N_17936,N_8331,N_7831);
nor U17937 (N_17937,N_12063,N_9919);
and U17938 (N_17938,N_9764,N_10102);
nand U17939 (N_17939,N_8881,N_9927);
and U17940 (N_17940,N_8920,N_8222);
and U17941 (N_17941,N_6925,N_11386);
and U17942 (N_17942,N_7220,N_6369);
nor U17943 (N_17943,N_9827,N_10349);
nand U17944 (N_17944,N_7958,N_10852);
and U17945 (N_17945,N_9281,N_8973);
nor U17946 (N_17946,N_10891,N_12152);
nand U17947 (N_17947,N_7525,N_7506);
or U17948 (N_17948,N_7857,N_8206);
and U17949 (N_17949,N_11947,N_11726);
nand U17950 (N_17950,N_10421,N_8694);
nand U17951 (N_17951,N_9180,N_12106);
nor U17952 (N_17952,N_8238,N_9079);
and U17953 (N_17953,N_11167,N_11414);
nor U17954 (N_17954,N_10214,N_12278);
nand U17955 (N_17955,N_6815,N_8333);
and U17956 (N_17956,N_10845,N_8425);
and U17957 (N_17957,N_7249,N_7350);
nor U17958 (N_17958,N_8421,N_9802);
nor U17959 (N_17959,N_12376,N_12470);
nor U17960 (N_17960,N_11262,N_10497);
or U17961 (N_17961,N_7137,N_9009);
xor U17962 (N_17962,N_9171,N_9797);
nand U17963 (N_17963,N_11286,N_8738);
nand U17964 (N_17964,N_11870,N_7296);
nor U17965 (N_17965,N_7902,N_6271);
nor U17966 (N_17966,N_11603,N_7333);
and U17967 (N_17967,N_7336,N_7776);
or U17968 (N_17968,N_11541,N_10648);
xnor U17969 (N_17969,N_7430,N_8243);
nand U17970 (N_17970,N_10478,N_11591);
nand U17971 (N_17971,N_12387,N_6584);
nor U17972 (N_17972,N_10732,N_10597);
and U17973 (N_17973,N_9480,N_11916);
or U17974 (N_17974,N_9724,N_12302);
or U17975 (N_17975,N_10781,N_8305);
and U17976 (N_17976,N_7107,N_9927);
xor U17977 (N_17977,N_7774,N_7187);
or U17978 (N_17978,N_7889,N_7811);
and U17979 (N_17979,N_9676,N_10400);
or U17980 (N_17980,N_10329,N_11718);
and U17981 (N_17981,N_9105,N_9497);
nor U17982 (N_17982,N_11235,N_10867);
nor U17983 (N_17983,N_6347,N_10567);
xnor U17984 (N_17984,N_8188,N_9992);
nand U17985 (N_17985,N_8530,N_6607);
or U17986 (N_17986,N_11636,N_7821);
nor U17987 (N_17987,N_12005,N_6503);
nor U17988 (N_17988,N_12345,N_11284);
nor U17989 (N_17989,N_7046,N_7565);
nor U17990 (N_17990,N_9697,N_9386);
nand U17991 (N_17991,N_10020,N_6901);
xor U17992 (N_17992,N_10176,N_8543);
or U17993 (N_17993,N_9234,N_10362);
nand U17994 (N_17994,N_9480,N_6671);
nor U17995 (N_17995,N_11877,N_10156);
or U17996 (N_17996,N_11785,N_12183);
and U17997 (N_17997,N_7781,N_8085);
nor U17998 (N_17998,N_9147,N_10332);
or U17999 (N_17999,N_10131,N_11097);
nand U18000 (N_18000,N_7595,N_7699);
or U18001 (N_18001,N_9097,N_11360);
nor U18002 (N_18002,N_7346,N_11341);
and U18003 (N_18003,N_8991,N_10206);
or U18004 (N_18004,N_9940,N_11403);
nor U18005 (N_18005,N_8316,N_9893);
nor U18006 (N_18006,N_9642,N_9497);
and U18007 (N_18007,N_6337,N_7592);
nor U18008 (N_18008,N_6851,N_7732);
nand U18009 (N_18009,N_7925,N_11126);
nand U18010 (N_18010,N_9600,N_11154);
nor U18011 (N_18011,N_7643,N_10691);
nand U18012 (N_18012,N_8939,N_6509);
or U18013 (N_18013,N_6789,N_11784);
nand U18014 (N_18014,N_9900,N_12432);
nand U18015 (N_18015,N_10471,N_11986);
or U18016 (N_18016,N_10875,N_10160);
nor U18017 (N_18017,N_12313,N_12283);
and U18018 (N_18018,N_10354,N_7572);
xor U18019 (N_18019,N_10536,N_8960);
or U18020 (N_18020,N_7911,N_7206);
and U18021 (N_18021,N_10065,N_10921);
nor U18022 (N_18022,N_12240,N_6875);
or U18023 (N_18023,N_7558,N_8531);
nor U18024 (N_18024,N_9696,N_8809);
nor U18025 (N_18025,N_9045,N_10641);
xnor U18026 (N_18026,N_11212,N_8359);
and U18027 (N_18027,N_12212,N_6919);
or U18028 (N_18028,N_9399,N_7579);
or U18029 (N_18029,N_10337,N_8879);
nand U18030 (N_18030,N_11242,N_6290);
or U18031 (N_18031,N_10967,N_9346);
and U18032 (N_18032,N_7914,N_8897);
and U18033 (N_18033,N_7646,N_10358);
or U18034 (N_18034,N_12173,N_9146);
and U18035 (N_18035,N_10336,N_10849);
nand U18036 (N_18036,N_7535,N_10304);
nor U18037 (N_18037,N_11229,N_9690);
nor U18038 (N_18038,N_10228,N_8754);
nor U18039 (N_18039,N_10442,N_8322);
nand U18040 (N_18040,N_12098,N_12449);
nand U18041 (N_18041,N_9292,N_11642);
nand U18042 (N_18042,N_8068,N_10670);
nor U18043 (N_18043,N_8403,N_8226);
nand U18044 (N_18044,N_10768,N_8290);
or U18045 (N_18045,N_11981,N_10144);
or U18046 (N_18046,N_10260,N_7004);
nor U18047 (N_18047,N_10718,N_11709);
nor U18048 (N_18048,N_6626,N_12037);
nand U18049 (N_18049,N_8741,N_10306);
nand U18050 (N_18050,N_8324,N_12028);
nand U18051 (N_18051,N_10240,N_9212);
or U18052 (N_18052,N_7927,N_10284);
xor U18053 (N_18053,N_6713,N_9718);
and U18054 (N_18054,N_8006,N_11275);
or U18055 (N_18055,N_9185,N_8197);
xor U18056 (N_18056,N_10377,N_9980);
or U18057 (N_18057,N_10154,N_8248);
and U18058 (N_18058,N_6386,N_9000);
or U18059 (N_18059,N_6682,N_6799);
nor U18060 (N_18060,N_9777,N_10561);
or U18061 (N_18061,N_8098,N_10561);
and U18062 (N_18062,N_10998,N_7768);
or U18063 (N_18063,N_11139,N_6609);
nand U18064 (N_18064,N_7066,N_8706);
and U18065 (N_18065,N_11198,N_6841);
nand U18066 (N_18066,N_8844,N_11720);
and U18067 (N_18067,N_10502,N_10426);
nand U18068 (N_18068,N_11586,N_8251);
xnor U18069 (N_18069,N_10927,N_6865);
nand U18070 (N_18070,N_7377,N_12368);
xor U18071 (N_18071,N_11050,N_7175);
nand U18072 (N_18072,N_8842,N_12420);
and U18073 (N_18073,N_7545,N_12331);
or U18074 (N_18074,N_10870,N_10607);
xor U18075 (N_18075,N_10060,N_6466);
or U18076 (N_18076,N_6705,N_9151);
nor U18077 (N_18077,N_9471,N_12212);
and U18078 (N_18078,N_11383,N_9699);
or U18079 (N_18079,N_9903,N_10832);
xnor U18080 (N_18080,N_8616,N_11338);
xnor U18081 (N_18081,N_9975,N_9625);
or U18082 (N_18082,N_6731,N_9609);
and U18083 (N_18083,N_10390,N_11072);
and U18084 (N_18084,N_7121,N_7907);
nor U18085 (N_18085,N_9520,N_11540);
and U18086 (N_18086,N_12415,N_8733);
or U18087 (N_18087,N_11122,N_12283);
or U18088 (N_18088,N_8194,N_7689);
nor U18089 (N_18089,N_9022,N_12451);
and U18090 (N_18090,N_8595,N_11459);
nand U18091 (N_18091,N_9788,N_11306);
nor U18092 (N_18092,N_9217,N_11832);
nand U18093 (N_18093,N_11427,N_7727);
or U18094 (N_18094,N_8332,N_9312);
and U18095 (N_18095,N_6259,N_11073);
nand U18096 (N_18096,N_7846,N_9608);
nor U18097 (N_18097,N_9123,N_7703);
xnor U18098 (N_18098,N_7376,N_7419);
nand U18099 (N_18099,N_9970,N_8757);
nor U18100 (N_18100,N_7746,N_6396);
nor U18101 (N_18101,N_6849,N_10435);
nand U18102 (N_18102,N_10949,N_11241);
nand U18103 (N_18103,N_11392,N_8527);
or U18104 (N_18104,N_7425,N_7028);
nor U18105 (N_18105,N_11258,N_8749);
or U18106 (N_18106,N_6475,N_9686);
nand U18107 (N_18107,N_11752,N_8241);
and U18108 (N_18108,N_7842,N_6404);
xnor U18109 (N_18109,N_6926,N_9249);
and U18110 (N_18110,N_12317,N_8410);
xnor U18111 (N_18111,N_11666,N_9172);
xor U18112 (N_18112,N_9167,N_6643);
xnor U18113 (N_18113,N_6744,N_9920);
or U18114 (N_18114,N_10434,N_7373);
or U18115 (N_18115,N_9935,N_8808);
nand U18116 (N_18116,N_6488,N_11100);
and U18117 (N_18117,N_7094,N_6412);
nand U18118 (N_18118,N_9033,N_7683);
and U18119 (N_18119,N_11753,N_8011);
nor U18120 (N_18120,N_9220,N_11540);
or U18121 (N_18121,N_8838,N_7154);
or U18122 (N_18122,N_10607,N_11205);
nand U18123 (N_18123,N_10453,N_6796);
or U18124 (N_18124,N_8992,N_12321);
or U18125 (N_18125,N_12355,N_6542);
nor U18126 (N_18126,N_11558,N_6657);
and U18127 (N_18127,N_7409,N_10837);
or U18128 (N_18128,N_7355,N_6644);
nor U18129 (N_18129,N_11620,N_12154);
xor U18130 (N_18130,N_10343,N_8777);
and U18131 (N_18131,N_12119,N_9421);
and U18132 (N_18132,N_7780,N_11802);
xnor U18133 (N_18133,N_8963,N_8161);
nand U18134 (N_18134,N_8448,N_6478);
and U18135 (N_18135,N_11771,N_6694);
nand U18136 (N_18136,N_12032,N_11329);
nand U18137 (N_18137,N_8748,N_12248);
nand U18138 (N_18138,N_7189,N_12044);
or U18139 (N_18139,N_11834,N_12461);
nand U18140 (N_18140,N_7728,N_8431);
xnor U18141 (N_18141,N_7254,N_9576);
nand U18142 (N_18142,N_10281,N_11817);
nand U18143 (N_18143,N_9024,N_9506);
xnor U18144 (N_18144,N_11454,N_7612);
xor U18145 (N_18145,N_9765,N_10791);
nand U18146 (N_18146,N_6468,N_9556);
or U18147 (N_18147,N_10486,N_7976);
nor U18148 (N_18148,N_8706,N_9269);
nor U18149 (N_18149,N_9251,N_7146);
xnor U18150 (N_18150,N_10043,N_12430);
and U18151 (N_18151,N_11799,N_12418);
or U18152 (N_18152,N_6302,N_7239);
xor U18153 (N_18153,N_7046,N_8774);
nand U18154 (N_18154,N_9645,N_8147);
xor U18155 (N_18155,N_8476,N_11936);
or U18156 (N_18156,N_8481,N_8212);
nand U18157 (N_18157,N_12187,N_7215);
and U18158 (N_18158,N_8294,N_9590);
xor U18159 (N_18159,N_9819,N_9498);
nor U18160 (N_18160,N_12185,N_9596);
xnor U18161 (N_18161,N_8223,N_8789);
nand U18162 (N_18162,N_7672,N_9156);
xor U18163 (N_18163,N_9527,N_7138);
and U18164 (N_18164,N_8547,N_12414);
nor U18165 (N_18165,N_7638,N_9160);
or U18166 (N_18166,N_11004,N_10297);
nor U18167 (N_18167,N_10945,N_11725);
nor U18168 (N_18168,N_7623,N_11264);
nor U18169 (N_18169,N_7892,N_7925);
or U18170 (N_18170,N_11541,N_11538);
nand U18171 (N_18171,N_6663,N_6840);
or U18172 (N_18172,N_8212,N_11493);
xor U18173 (N_18173,N_10034,N_6515);
or U18174 (N_18174,N_9404,N_10229);
and U18175 (N_18175,N_11740,N_10099);
and U18176 (N_18176,N_8615,N_8099);
xor U18177 (N_18177,N_6791,N_11649);
nand U18178 (N_18178,N_8580,N_7796);
or U18179 (N_18179,N_11558,N_11928);
nor U18180 (N_18180,N_11777,N_9416);
nand U18181 (N_18181,N_10554,N_8100);
nor U18182 (N_18182,N_10441,N_6510);
or U18183 (N_18183,N_7813,N_8589);
nor U18184 (N_18184,N_9513,N_9141);
and U18185 (N_18185,N_10413,N_8767);
and U18186 (N_18186,N_11757,N_9386);
nor U18187 (N_18187,N_7834,N_6471);
nand U18188 (N_18188,N_8344,N_9914);
or U18189 (N_18189,N_6311,N_9155);
nor U18190 (N_18190,N_6981,N_11647);
or U18191 (N_18191,N_11227,N_8111);
nor U18192 (N_18192,N_12164,N_8105);
nand U18193 (N_18193,N_12253,N_9846);
or U18194 (N_18194,N_10824,N_8300);
or U18195 (N_18195,N_7652,N_8226);
or U18196 (N_18196,N_7766,N_11502);
and U18197 (N_18197,N_8020,N_11759);
and U18198 (N_18198,N_10397,N_11820);
xnor U18199 (N_18199,N_6734,N_6620);
and U18200 (N_18200,N_10228,N_9971);
nor U18201 (N_18201,N_12160,N_6710);
or U18202 (N_18202,N_7689,N_9183);
nand U18203 (N_18203,N_10618,N_6484);
or U18204 (N_18204,N_10610,N_7636);
xnor U18205 (N_18205,N_7432,N_9068);
nor U18206 (N_18206,N_8743,N_10576);
or U18207 (N_18207,N_8250,N_10456);
nor U18208 (N_18208,N_7465,N_11098);
and U18209 (N_18209,N_8336,N_11513);
xnor U18210 (N_18210,N_6587,N_11859);
nor U18211 (N_18211,N_12395,N_8918);
or U18212 (N_18212,N_6623,N_9914);
or U18213 (N_18213,N_10565,N_9221);
or U18214 (N_18214,N_11548,N_12325);
nor U18215 (N_18215,N_8694,N_8262);
and U18216 (N_18216,N_6649,N_8676);
nand U18217 (N_18217,N_7982,N_9095);
nand U18218 (N_18218,N_9495,N_10161);
or U18219 (N_18219,N_10124,N_9755);
nand U18220 (N_18220,N_11141,N_12316);
nand U18221 (N_18221,N_10448,N_9200);
nor U18222 (N_18222,N_6611,N_10513);
xnor U18223 (N_18223,N_9027,N_7263);
or U18224 (N_18224,N_8734,N_6273);
nor U18225 (N_18225,N_10144,N_8172);
and U18226 (N_18226,N_11525,N_11825);
nor U18227 (N_18227,N_6576,N_11622);
nand U18228 (N_18228,N_7860,N_6480);
or U18229 (N_18229,N_10793,N_9508);
or U18230 (N_18230,N_8074,N_9687);
nand U18231 (N_18231,N_7902,N_11481);
or U18232 (N_18232,N_7521,N_8169);
nand U18233 (N_18233,N_7454,N_11607);
or U18234 (N_18234,N_7135,N_11698);
and U18235 (N_18235,N_9303,N_9885);
nand U18236 (N_18236,N_9789,N_11333);
or U18237 (N_18237,N_7247,N_11038);
and U18238 (N_18238,N_11369,N_6832);
nand U18239 (N_18239,N_9331,N_9207);
or U18240 (N_18240,N_11005,N_9426);
nor U18241 (N_18241,N_7230,N_6638);
or U18242 (N_18242,N_7185,N_7044);
nor U18243 (N_18243,N_12483,N_7695);
nand U18244 (N_18244,N_9961,N_6346);
or U18245 (N_18245,N_7600,N_12420);
nand U18246 (N_18246,N_11921,N_10424);
or U18247 (N_18247,N_11478,N_9220);
xnor U18248 (N_18248,N_9331,N_6432);
nand U18249 (N_18249,N_6267,N_12435);
nand U18250 (N_18250,N_8617,N_9857);
nand U18251 (N_18251,N_7124,N_6672);
xor U18252 (N_18252,N_9218,N_7939);
nor U18253 (N_18253,N_9117,N_9502);
nand U18254 (N_18254,N_10155,N_7348);
or U18255 (N_18255,N_9918,N_12174);
and U18256 (N_18256,N_8948,N_6799);
nor U18257 (N_18257,N_6254,N_7309);
and U18258 (N_18258,N_10551,N_9748);
and U18259 (N_18259,N_9888,N_9869);
and U18260 (N_18260,N_10445,N_6735);
or U18261 (N_18261,N_6453,N_9859);
nor U18262 (N_18262,N_8219,N_9750);
and U18263 (N_18263,N_7021,N_11336);
nor U18264 (N_18264,N_9891,N_11189);
nor U18265 (N_18265,N_10564,N_10235);
or U18266 (N_18266,N_10577,N_7373);
nor U18267 (N_18267,N_12075,N_11791);
or U18268 (N_18268,N_9359,N_8378);
and U18269 (N_18269,N_6556,N_7334);
nor U18270 (N_18270,N_12419,N_9691);
and U18271 (N_18271,N_11906,N_9478);
nor U18272 (N_18272,N_6408,N_8992);
or U18273 (N_18273,N_12289,N_9225);
or U18274 (N_18274,N_7090,N_6637);
and U18275 (N_18275,N_8769,N_7231);
and U18276 (N_18276,N_8760,N_9339);
and U18277 (N_18277,N_7731,N_9612);
or U18278 (N_18278,N_10669,N_11941);
xnor U18279 (N_18279,N_7711,N_8173);
or U18280 (N_18280,N_7269,N_11217);
nand U18281 (N_18281,N_11558,N_11256);
and U18282 (N_18282,N_9838,N_11197);
nand U18283 (N_18283,N_6523,N_7079);
or U18284 (N_18284,N_6869,N_6369);
or U18285 (N_18285,N_7008,N_9207);
or U18286 (N_18286,N_9773,N_8646);
nand U18287 (N_18287,N_8514,N_9870);
nor U18288 (N_18288,N_9505,N_11523);
nor U18289 (N_18289,N_10956,N_8925);
xor U18290 (N_18290,N_10618,N_11668);
or U18291 (N_18291,N_10815,N_8548);
nand U18292 (N_18292,N_7717,N_9884);
and U18293 (N_18293,N_9049,N_9549);
and U18294 (N_18294,N_10362,N_11498);
and U18295 (N_18295,N_9766,N_7346);
nor U18296 (N_18296,N_9293,N_11380);
or U18297 (N_18297,N_7329,N_11118);
or U18298 (N_18298,N_9116,N_10652);
or U18299 (N_18299,N_9289,N_7040);
nor U18300 (N_18300,N_7976,N_6767);
nor U18301 (N_18301,N_11429,N_7374);
nor U18302 (N_18302,N_11161,N_9867);
nor U18303 (N_18303,N_12147,N_12187);
nor U18304 (N_18304,N_9857,N_12336);
nor U18305 (N_18305,N_10941,N_9117);
or U18306 (N_18306,N_8592,N_10078);
nand U18307 (N_18307,N_10453,N_8911);
or U18308 (N_18308,N_7747,N_9995);
nand U18309 (N_18309,N_7613,N_7222);
and U18310 (N_18310,N_9727,N_7279);
nor U18311 (N_18311,N_8994,N_9698);
xnor U18312 (N_18312,N_12154,N_9322);
xor U18313 (N_18313,N_9351,N_10766);
xnor U18314 (N_18314,N_11491,N_10962);
and U18315 (N_18315,N_6624,N_8204);
or U18316 (N_18316,N_6595,N_8776);
and U18317 (N_18317,N_9999,N_8156);
nand U18318 (N_18318,N_10198,N_10880);
nand U18319 (N_18319,N_9492,N_10432);
or U18320 (N_18320,N_11518,N_6907);
nor U18321 (N_18321,N_9204,N_7040);
or U18322 (N_18322,N_6528,N_6901);
or U18323 (N_18323,N_7731,N_9178);
nor U18324 (N_18324,N_6575,N_8593);
or U18325 (N_18325,N_6376,N_6784);
and U18326 (N_18326,N_10740,N_6325);
and U18327 (N_18327,N_12203,N_8335);
or U18328 (N_18328,N_9837,N_6449);
nand U18329 (N_18329,N_12217,N_10348);
and U18330 (N_18330,N_10828,N_9990);
xor U18331 (N_18331,N_7025,N_12029);
nor U18332 (N_18332,N_11792,N_7783);
nor U18333 (N_18333,N_6629,N_9675);
nand U18334 (N_18334,N_10569,N_11585);
nand U18335 (N_18335,N_9657,N_9991);
nor U18336 (N_18336,N_9817,N_11530);
nor U18337 (N_18337,N_7554,N_10489);
or U18338 (N_18338,N_7779,N_8330);
and U18339 (N_18339,N_7403,N_10441);
and U18340 (N_18340,N_6712,N_8174);
nor U18341 (N_18341,N_6378,N_8346);
and U18342 (N_18342,N_6716,N_9497);
nor U18343 (N_18343,N_12232,N_8747);
nand U18344 (N_18344,N_9424,N_8904);
nand U18345 (N_18345,N_7749,N_6484);
or U18346 (N_18346,N_12366,N_9340);
nand U18347 (N_18347,N_6744,N_8848);
nor U18348 (N_18348,N_10026,N_8213);
nor U18349 (N_18349,N_8697,N_11208);
and U18350 (N_18350,N_7135,N_10776);
nand U18351 (N_18351,N_11175,N_10663);
or U18352 (N_18352,N_6733,N_9332);
nand U18353 (N_18353,N_8926,N_8209);
xnor U18354 (N_18354,N_12441,N_10124);
nand U18355 (N_18355,N_7427,N_9169);
or U18356 (N_18356,N_11565,N_9413);
or U18357 (N_18357,N_8522,N_6584);
and U18358 (N_18358,N_12203,N_9489);
nor U18359 (N_18359,N_6818,N_9042);
nand U18360 (N_18360,N_11081,N_10311);
and U18361 (N_18361,N_7414,N_11845);
or U18362 (N_18362,N_7148,N_10196);
or U18363 (N_18363,N_9747,N_7757);
and U18364 (N_18364,N_8018,N_11091);
xor U18365 (N_18365,N_7030,N_11023);
or U18366 (N_18366,N_6836,N_8661);
or U18367 (N_18367,N_7991,N_8708);
and U18368 (N_18368,N_6873,N_6899);
or U18369 (N_18369,N_12095,N_7724);
or U18370 (N_18370,N_8917,N_11186);
and U18371 (N_18371,N_8382,N_8550);
nor U18372 (N_18372,N_11744,N_9852);
nor U18373 (N_18373,N_11055,N_7086);
xnor U18374 (N_18374,N_6583,N_11374);
or U18375 (N_18375,N_11721,N_12008);
nor U18376 (N_18376,N_9251,N_8809);
xor U18377 (N_18377,N_9184,N_10661);
or U18378 (N_18378,N_9220,N_7375);
nor U18379 (N_18379,N_7898,N_7185);
and U18380 (N_18380,N_9350,N_10601);
nand U18381 (N_18381,N_9139,N_6468);
and U18382 (N_18382,N_8532,N_8071);
nor U18383 (N_18383,N_7685,N_6849);
nor U18384 (N_18384,N_9908,N_6615);
nand U18385 (N_18385,N_9525,N_8440);
or U18386 (N_18386,N_6781,N_8815);
nand U18387 (N_18387,N_8647,N_10941);
nand U18388 (N_18388,N_7050,N_9095);
or U18389 (N_18389,N_7020,N_11179);
nand U18390 (N_18390,N_9032,N_10269);
nor U18391 (N_18391,N_10943,N_9281);
or U18392 (N_18392,N_10696,N_12350);
and U18393 (N_18393,N_12008,N_7844);
nand U18394 (N_18394,N_8234,N_10068);
or U18395 (N_18395,N_6511,N_7175);
nor U18396 (N_18396,N_10449,N_9131);
nand U18397 (N_18397,N_7788,N_8061);
nand U18398 (N_18398,N_10905,N_7233);
and U18399 (N_18399,N_10606,N_9942);
nor U18400 (N_18400,N_8299,N_10943);
or U18401 (N_18401,N_11790,N_9513);
nor U18402 (N_18402,N_9831,N_7399);
or U18403 (N_18403,N_7405,N_7767);
nor U18404 (N_18404,N_10883,N_11266);
nand U18405 (N_18405,N_8431,N_11877);
nand U18406 (N_18406,N_11598,N_6684);
nand U18407 (N_18407,N_11483,N_7957);
xor U18408 (N_18408,N_9942,N_10862);
nor U18409 (N_18409,N_11105,N_11477);
or U18410 (N_18410,N_9800,N_7586);
and U18411 (N_18411,N_7951,N_11443);
nand U18412 (N_18412,N_10284,N_11833);
nand U18413 (N_18413,N_6632,N_10400);
nor U18414 (N_18414,N_11652,N_11138);
nand U18415 (N_18415,N_9772,N_7435);
xor U18416 (N_18416,N_8295,N_9028);
or U18417 (N_18417,N_11696,N_12134);
and U18418 (N_18418,N_6592,N_9023);
nand U18419 (N_18419,N_10093,N_11905);
and U18420 (N_18420,N_7048,N_10397);
nand U18421 (N_18421,N_7059,N_7309);
and U18422 (N_18422,N_7370,N_8923);
nor U18423 (N_18423,N_10672,N_9052);
xor U18424 (N_18424,N_9757,N_7801);
nor U18425 (N_18425,N_7575,N_10506);
nand U18426 (N_18426,N_9487,N_10073);
or U18427 (N_18427,N_7475,N_6679);
nand U18428 (N_18428,N_8622,N_11458);
and U18429 (N_18429,N_11826,N_11117);
nand U18430 (N_18430,N_7149,N_7633);
nor U18431 (N_18431,N_6394,N_10636);
and U18432 (N_18432,N_6743,N_7916);
nor U18433 (N_18433,N_9916,N_7657);
nand U18434 (N_18434,N_10005,N_9946);
and U18435 (N_18435,N_10559,N_8946);
or U18436 (N_18436,N_10758,N_7494);
nand U18437 (N_18437,N_9487,N_8273);
or U18438 (N_18438,N_10498,N_10173);
or U18439 (N_18439,N_9833,N_7137);
and U18440 (N_18440,N_12024,N_8778);
xor U18441 (N_18441,N_10319,N_7071);
and U18442 (N_18442,N_9688,N_11450);
and U18443 (N_18443,N_6375,N_9126);
and U18444 (N_18444,N_10413,N_9581);
and U18445 (N_18445,N_11731,N_10445);
and U18446 (N_18446,N_11989,N_10658);
and U18447 (N_18447,N_9054,N_9112);
and U18448 (N_18448,N_7134,N_11264);
xnor U18449 (N_18449,N_11406,N_6647);
nor U18450 (N_18450,N_8888,N_8878);
or U18451 (N_18451,N_11719,N_7808);
or U18452 (N_18452,N_11495,N_7159);
and U18453 (N_18453,N_11842,N_10333);
xor U18454 (N_18454,N_10930,N_7419);
or U18455 (N_18455,N_12451,N_10646);
nand U18456 (N_18456,N_12049,N_9162);
nor U18457 (N_18457,N_7728,N_9319);
and U18458 (N_18458,N_6442,N_6684);
or U18459 (N_18459,N_8206,N_8243);
xor U18460 (N_18460,N_7733,N_7999);
and U18461 (N_18461,N_8783,N_8209);
nand U18462 (N_18462,N_9431,N_6646);
and U18463 (N_18463,N_6361,N_8549);
or U18464 (N_18464,N_7711,N_6497);
or U18465 (N_18465,N_9191,N_9178);
and U18466 (N_18466,N_8578,N_8265);
and U18467 (N_18467,N_8315,N_6391);
nor U18468 (N_18468,N_11387,N_7962);
and U18469 (N_18469,N_11469,N_9246);
and U18470 (N_18470,N_8593,N_10261);
nand U18471 (N_18471,N_6916,N_6284);
nor U18472 (N_18472,N_9998,N_11420);
and U18473 (N_18473,N_12436,N_7079);
and U18474 (N_18474,N_11641,N_9719);
nand U18475 (N_18475,N_7139,N_6947);
nand U18476 (N_18476,N_11679,N_10084);
nand U18477 (N_18477,N_9095,N_6598);
nor U18478 (N_18478,N_6684,N_11278);
nor U18479 (N_18479,N_11973,N_8250);
xnor U18480 (N_18480,N_7850,N_10350);
and U18481 (N_18481,N_10431,N_10615);
nand U18482 (N_18482,N_11720,N_11686);
or U18483 (N_18483,N_8036,N_10315);
xor U18484 (N_18484,N_7760,N_7382);
or U18485 (N_18485,N_6868,N_11042);
nand U18486 (N_18486,N_9874,N_12092);
nor U18487 (N_18487,N_12099,N_11908);
nand U18488 (N_18488,N_7487,N_7745);
and U18489 (N_18489,N_6435,N_7016);
or U18490 (N_18490,N_6813,N_12136);
or U18491 (N_18491,N_7634,N_8912);
nor U18492 (N_18492,N_6790,N_10049);
nand U18493 (N_18493,N_8062,N_7080);
and U18494 (N_18494,N_11557,N_8417);
or U18495 (N_18495,N_9754,N_8829);
and U18496 (N_18496,N_9901,N_9850);
or U18497 (N_18497,N_8870,N_9133);
nor U18498 (N_18498,N_10372,N_8359);
nand U18499 (N_18499,N_6256,N_8921);
nand U18500 (N_18500,N_11983,N_12282);
nand U18501 (N_18501,N_11403,N_11905);
or U18502 (N_18502,N_9329,N_11339);
and U18503 (N_18503,N_9217,N_11386);
and U18504 (N_18504,N_12041,N_9615);
nand U18505 (N_18505,N_6849,N_10310);
or U18506 (N_18506,N_11078,N_11408);
and U18507 (N_18507,N_9474,N_8745);
nor U18508 (N_18508,N_8720,N_8616);
xor U18509 (N_18509,N_10932,N_10730);
and U18510 (N_18510,N_10498,N_6639);
nand U18511 (N_18511,N_10184,N_11991);
or U18512 (N_18512,N_8103,N_8702);
or U18513 (N_18513,N_10380,N_8771);
nand U18514 (N_18514,N_11234,N_7317);
xor U18515 (N_18515,N_11956,N_11924);
and U18516 (N_18516,N_8724,N_10735);
nand U18517 (N_18517,N_10245,N_8016);
or U18518 (N_18518,N_7353,N_6838);
and U18519 (N_18519,N_7192,N_9720);
nor U18520 (N_18520,N_8855,N_12295);
and U18521 (N_18521,N_10189,N_7673);
nor U18522 (N_18522,N_6956,N_6688);
xnor U18523 (N_18523,N_7830,N_12188);
or U18524 (N_18524,N_11275,N_9624);
xor U18525 (N_18525,N_8762,N_6421);
or U18526 (N_18526,N_8546,N_9018);
or U18527 (N_18527,N_6468,N_8601);
nor U18528 (N_18528,N_11042,N_12309);
nor U18529 (N_18529,N_8754,N_6654);
nand U18530 (N_18530,N_10565,N_6626);
nand U18531 (N_18531,N_6436,N_11276);
and U18532 (N_18532,N_8501,N_12047);
and U18533 (N_18533,N_7715,N_8720);
xnor U18534 (N_18534,N_9946,N_8730);
or U18535 (N_18535,N_9107,N_8686);
and U18536 (N_18536,N_8463,N_10006);
nor U18537 (N_18537,N_8311,N_10610);
nor U18538 (N_18538,N_6402,N_12146);
and U18539 (N_18539,N_6532,N_6999);
or U18540 (N_18540,N_11942,N_12241);
and U18541 (N_18541,N_6347,N_10937);
and U18542 (N_18542,N_6291,N_12398);
nand U18543 (N_18543,N_9116,N_6748);
and U18544 (N_18544,N_9356,N_7316);
and U18545 (N_18545,N_9802,N_6974);
or U18546 (N_18546,N_7435,N_7896);
nand U18547 (N_18547,N_9674,N_6539);
and U18548 (N_18548,N_12315,N_6586);
or U18549 (N_18549,N_11770,N_7830);
nor U18550 (N_18550,N_8955,N_7014);
nand U18551 (N_18551,N_6686,N_6357);
nor U18552 (N_18552,N_7225,N_8272);
nand U18553 (N_18553,N_6428,N_9500);
or U18554 (N_18554,N_7850,N_7578);
nand U18555 (N_18555,N_7890,N_11347);
nand U18556 (N_18556,N_10688,N_11751);
nor U18557 (N_18557,N_9238,N_6902);
and U18558 (N_18558,N_7173,N_7215);
nor U18559 (N_18559,N_11163,N_9369);
nand U18560 (N_18560,N_10571,N_10013);
xnor U18561 (N_18561,N_10804,N_6332);
or U18562 (N_18562,N_10186,N_6490);
and U18563 (N_18563,N_9891,N_7510);
and U18564 (N_18564,N_9385,N_11349);
nand U18565 (N_18565,N_7923,N_7595);
and U18566 (N_18566,N_8396,N_8934);
nand U18567 (N_18567,N_6786,N_6713);
nand U18568 (N_18568,N_8136,N_11172);
nor U18569 (N_18569,N_10018,N_10327);
and U18570 (N_18570,N_10639,N_8029);
nand U18571 (N_18571,N_7468,N_6962);
or U18572 (N_18572,N_12324,N_12466);
or U18573 (N_18573,N_7154,N_7639);
or U18574 (N_18574,N_8713,N_6453);
and U18575 (N_18575,N_6666,N_9780);
xor U18576 (N_18576,N_9905,N_7681);
nand U18577 (N_18577,N_6897,N_11240);
nor U18578 (N_18578,N_8619,N_6518);
nor U18579 (N_18579,N_10519,N_10308);
xnor U18580 (N_18580,N_7142,N_8014);
nand U18581 (N_18581,N_7682,N_11014);
nor U18582 (N_18582,N_9981,N_12124);
nand U18583 (N_18583,N_7108,N_10036);
or U18584 (N_18584,N_6964,N_9477);
xnor U18585 (N_18585,N_6461,N_11318);
xor U18586 (N_18586,N_10556,N_11786);
nand U18587 (N_18587,N_7805,N_8684);
nor U18588 (N_18588,N_8124,N_12084);
nand U18589 (N_18589,N_9969,N_10676);
nor U18590 (N_18590,N_10298,N_10102);
nand U18591 (N_18591,N_10988,N_7615);
nand U18592 (N_18592,N_11090,N_12076);
or U18593 (N_18593,N_7796,N_8836);
and U18594 (N_18594,N_9196,N_7994);
nor U18595 (N_18595,N_10327,N_9218);
or U18596 (N_18596,N_10937,N_6295);
xor U18597 (N_18597,N_7042,N_7940);
xnor U18598 (N_18598,N_8568,N_9264);
and U18599 (N_18599,N_11940,N_9662);
and U18600 (N_18600,N_8983,N_7104);
nand U18601 (N_18601,N_9001,N_10065);
nor U18602 (N_18602,N_7007,N_12201);
or U18603 (N_18603,N_10549,N_9981);
or U18604 (N_18604,N_6328,N_9017);
nand U18605 (N_18605,N_8810,N_6740);
or U18606 (N_18606,N_6895,N_11614);
and U18607 (N_18607,N_8755,N_11421);
nand U18608 (N_18608,N_11313,N_10009);
nand U18609 (N_18609,N_12327,N_9873);
and U18610 (N_18610,N_9221,N_7973);
nor U18611 (N_18611,N_10567,N_11039);
xnor U18612 (N_18612,N_9273,N_11777);
nor U18613 (N_18613,N_7401,N_12498);
and U18614 (N_18614,N_12188,N_9661);
and U18615 (N_18615,N_9401,N_7787);
nand U18616 (N_18616,N_11810,N_7542);
or U18617 (N_18617,N_6444,N_12074);
nand U18618 (N_18618,N_8589,N_7587);
xor U18619 (N_18619,N_11902,N_11261);
nor U18620 (N_18620,N_9765,N_10291);
or U18621 (N_18621,N_8174,N_11043);
or U18622 (N_18622,N_6976,N_11324);
or U18623 (N_18623,N_11335,N_12361);
and U18624 (N_18624,N_9913,N_7155);
and U18625 (N_18625,N_12384,N_11779);
xnor U18626 (N_18626,N_7909,N_10452);
and U18627 (N_18627,N_9350,N_8366);
and U18628 (N_18628,N_7879,N_8965);
and U18629 (N_18629,N_11555,N_7310);
or U18630 (N_18630,N_9901,N_11288);
xor U18631 (N_18631,N_11603,N_9360);
nor U18632 (N_18632,N_11272,N_9725);
or U18633 (N_18633,N_9512,N_6938);
or U18634 (N_18634,N_9963,N_6629);
and U18635 (N_18635,N_10180,N_11799);
nand U18636 (N_18636,N_6784,N_6464);
nor U18637 (N_18637,N_8274,N_8245);
or U18638 (N_18638,N_6717,N_8639);
nor U18639 (N_18639,N_12401,N_9709);
or U18640 (N_18640,N_7844,N_10550);
nor U18641 (N_18641,N_6935,N_6622);
nand U18642 (N_18642,N_12198,N_9764);
or U18643 (N_18643,N_7604,N_11334);
nand U18644 (N_18644,N_11470,N_9341);
xnor U18645 (N_18645,N_7202,N_11758);
nand U18646 (N_18646,N_10514,N_10923);
xor U18647 (N_18647,N_12014,N_8299);
nand U18648 (N_18648,N_10835,N_10855);
xnor U18649 (N_18649,N_10347,N_6742);
nor U18650 (N_18650,N_7735,N_7385);
nor U18651 (N_18651,N_6672,N_10880);
nor U18652 (N_18652,N_11690,N_6738);
or U18653 (N_18653,N_6755,N_10873);
nor U18654 (N_18654,N_9985,N_6763);
nand U18655 (N_18655,N_7282,N_8383);
and U18656 (N_18656,N_6756,N_11413);
or U18657 (N_18657,N_9116,N_7378);
nand U18658 (N_18658,N_9083,N_9433);
and U18659 (N_18659,N_6276,N_6394);
or U18660 (N_18660,N_7413,N_9981);
nor U18661 (N_18661,N_10067,N_8487);
nor U18662 (N_18662,N_8575,N_7766);
and U18663 (N_18663,N_12108,N_10111);
xnor U18664 (N_18664,N_9843,N_11726);
xor U18665 (N_18665,N_11857,N_11654);
nand U18666 (N_18666,N_11963,N_9688);
xor U18667 (N_18667,N_8166,N_8904);
and U18668 (N_18668,N_8804,N_12359);
and U18669 (N_18669,N_11950,N_9142);
nor U18670 (N_18670,N_12460,N_12261);
or U18671 (N_18671,N_11913,N_7186);
or U18672 (N_18672,N_12130,N_7799);
nor U18673 (N_18673,N_6660,N_12088);
and U18674 (N_18674,N_9677,N_12229);
xnor U18675 (N_18675,N_11997,N_10815);
and U18676 (N_18676,N_9448,N_11020);
nor U18677 (N_18677,N_9724,N_8769);
and U18678 (N_18678,N_8671,N_10166);
and U18679 (N_18679,N_10963,N_11916);
xnor U18680 (N_18680,N_10146,N_7280);
nor U18681 (N_18681,N_8594,N_7240);
nand U18682 (N_18682,N_8542,N_7720);
and U18683 (N_18683,N_11257,N_11467);
nor U18684 (N_18684,N_9674,N_10829);
xor U18685 (N_18685,N_12400,N_7120);
or U18686 (N_18686,N_11023,N_12439);
and U18687 (N_18687,N_7977,N_11716);
nor U18688 (N_18688,N_11301,N_10092);
and U18689 (N_18689,N_7928,N_12211);
nor U18690 (N_18690,N_8118,N_11772);
nor U18691 (N_18691,N_8612,N_11769);
nand U18692 (N_18692,N_9574,N_9683);
xor U18693 (N_18693,N_7391,N_9527);
nor U18694 (N_18694,N_7722,N_6336);
and U18695 (N_18695,N_7117,N_10233);
nand U18696 (N_18696,N_10831,N_9387);
or U18697 (N_18697,N_6424,N_10044);
nand U18698 (N_18698,N_12029,N_6339);
and U18699 (N_18699,N_9458,N_9199);
or U18700 (N_18700,N_9986,N_11241);
and U18701 (N_18701,N_7576,N_10145);
xor U18702 (N_18702,N_6350,N_8523);
or U18703 (N_18703,N_12251,N_7459);
or U18704 (N_18704,N_9790,N_10472);
nor U18705 (N_18705,N_7897,N_8712);
and U18706 (N_18706,N_9135,N_10575);
and U18707 (N_18707,N_6377,N_10984);
xnor U18708 (N_18708,N_8913,N_11950);
nor U18709 (N_18709,N_7415,N_11325);
and U18710 (N_18710,N_11789,N_12289);
nand U18711 (N_18711,N_10307,N_9394);
nand U18712 (N_18712,N_7041,N_7081);
nor U18713 (N_18713,N_9163,N_12056);
and U18714 (N_18714,N_6480,N_7956);
and U18715 (N_18715,N_9796,N_6701);
and U18716 (N_18716,N_7418,N_8558);
nor U18717 (N_18717,N_9490,N_10050);
xor U18718 (N_18718,N_12236,N_7074);
or U18719 (N_18719,N_12418,N_9602);
and U18720 (N_18720,N_10597,N_12072);
or U18721 (N_18721,N_6553,N_9210);
nand U18722 (N_18722,N_11673,N_8148);
nand U18723 (N_18723,N_8207,N_6586);
and U18724 (N_18724,N_11556,N_8220);
nor U18725 (N_18725,N_6353,N_11865);
nand U18726 (N_18726,N_12396,N_7688);
nor U18727 (N_18727,N_8767,N_6689);
and U18728 (N_18728,N_8851,N_9979);
or U18729 (N_18729,N_7005,N_11865);
or U18730 (N_18730,N_10493,N_11197);
nand U18731 (N_18731,N_6716,N_7466);
nand U18732 (N_18732,N_8754,N_6553);
and U18733 (N_18733,N_12223,N_10920);
nand U18734 (N_18734,N_6596,N_6617);
and U18735 (N_18735,N_7892,N_7847);
nand U18736 (N_18736,N_11633,N_7046);
nand U18737 (N_18737,N_11730,N_11045);
nand U18738 (N_18738,N_7417,N_7463);
nand U18739 (N_18739,N_9759,N_8396);
nor U18740 (N_18740,N_11524,N_8554);
or U18741 (N_18741,N_12445,N_10651);
nor U18742 (N_18742,N_9492,N_8689);
or U18743 (N_18743,N_12280,N_9521);
nand U18744 (N_18744,N_9688,N_8460);
and U18745 (N_18745,N_10378,N_9821);
and U18746 (N_18746,N_7244,N_9638);
or U18747 (N_18747,N_10498,N_10006);
and U18748 (N_18748,N_10509,N_11657);
nor U18749 (N_18749,N_9188,N_10961);
nor U18750 (N_18750,N_15508,N_15623);
or U18751 (N_18751,N_13743,N_18556);
nor U18752 (N_18752,N_17150,N_15885);
or U18753 (N_18753,N_18127,N_17286);
xnor U18754 (N_18754,N_13575,N_17282);
and U18755 (N_18755,N_16631,N_14757);
and U18756 (N_18756,N_13860,N_13132);
or U18757 (N_18757,N_14028,N_13447);
nand U18758 (N_18758,N_13476,N_13044);
nand U18759 (N_18759,N_15230,N_15617);
xor U18760 (N_18760,N_13140,N_14384);
and U18761 (N_18761,N_15234,N_13244);
nand U18762 (N_18762,N_14686,N_14188);
or U18763 (N_18763,N_15828,N_16951);
or U18764 (N_18764,N_16344,N_15942);
or U18765 (N_18765,N_14192,N_15320);
or U18766 (N_18766,N_16908,N_18230);
nand U18767 (N_18767,N_13961,N_13848);
nor U18768 (N_18768,N_15066,N_16143);
nand U18769 (N_18769,N_17367,N_18680);
nor U18770 (N_18770,N_15010,N_12904);
or U18771 (N_18771,N_12665,N_14595);
nor U18772 (N_18772,N_16216,N_16297);
and U18773 (N_18773,N_15439,N_17226);
nand U18774 (N_18774,N_12797,N_18667);
xnor U18775 (N_18775,N_18412,N_17340);
or U18776 (N_18776,N_14756,N_14526);
nor U18777 (N_18777,N_16357,N_14607);
and U18778 (N_18778,N_14973,N_13464);
or U18779 (N_18779,N_15161,N_13789);
or U18780 (N_18780,N_14452,N_13274);
and U18781 (N_18781,N_15824,N_18078);
nor U18782 (N_18782,N_17982,N_12616);
or U18783 (N_18783,N_14136,N_12833);
nor U18784 (N_18784,N_13703,N_17347);
or U18785 (N_18785,N_15476,N_14509);
nor U18786 (N_18786,N_13059,N_16615);
and U18787 (N_18787,N_16140,N_13290);
nand U18788 (N_18788,N_16762,N_18338);
and U18789 (N_18789,N_14948,N_16236);
or U18790 (N_18790,N_16442,N_15354);
nor U18791 (N_18791,N_16607,N_15856);
nand U18792 (N_18792,N_14097,N_12610);
nor U18793 (N_18793,N_15091,N_15886);
nor U18794 (N_18794,N_15125,N_18345);
and U18795 (N_18795,N_14524,N_15314);
and U18796 (N_18796,N_18578,N_14959);
nor U18797 (N_18797,N_12935,N_13495);
nand U18798 (N_18798,N_13395,N_16658);
and U18799 (N_18799,N_18298,N_14742);
nor U18800 (N_18800,N_18673,N_14781);
nor U18801 (N_18801,N_15352,N_14634);
nand U18802 (N_18802,N_15548,N_16982);
nand U18803 (N_18803,N_15945,N_13298);
nand U18804 (N_18804,N_18214,N_13824);
xor U18805 (N_18805,N_17195,N_13317);
nor U18806 (N_18806,N_17970,N_15844);
xnor U18807 (N_18807,N_17214,N_16926);
and U18808 (N_18808,N_13436,N_15065);
nor U18809 (N_18809,N_15495,N_15387);
or U18810 (N_18810,N_15690,N_14465);
and U18811 (N_18811,N_15843,N_17866);
xor U18812 (N_18812,N_15076,N_17089);
nand U18813 (N_18813,N_16057,N_17619);
nand U18814 (N_18814,N_17622,N_14897);
nand U18815 (N_18815,N_18456,N_17243);
and U18816 (N_18816,N_16989,N_18146);
xor U18817 (N_18817,N_13027,N_13911);
or U18818 (N_18818,N_14515,N_14852);
nand U18819 (N_18819,N_15121,N_17879);
nor U18820 (N_18820,N_16688,N_14484);
and U18821 (N_18821,N_16376,N_17287);
or U18822 (N_18822,N_16849,N_18051);
or U18823 (N_18823,N_12880,N_15277);
xor U18824 (N_18824,N_15849,N_14287);
and U18825 (N_18825,N_16068,N_18421);
or U18826 (N_18826,N_13401,N_17071);
and U18827 (N_18827,N_17918,N_13407);
nand U18828 (N_18828,N_12513,N_16099);
xor U18829 (N_18829,N_15009,N_17810);
nor U18830 (N_18830,N_18734,N_14712);
or U18831 (N_18831,N_15745,N_17821);
nand U18832 (N_18832,N_13029,N_14992);
nor U18833 (N_18833,N_16605,N_16977);
or U18834 (N_18834,N_14132,N_16269);
nand U18835 (N_18835,N_17635,N_16756);
nor U18836 (N_18836,N_16327,N_15041);
nor U18837 (N_18837,N_13483,N_14870);
nor U18838 (N_18838,N_15131,N_12932);
nand U18839 (N_18839,N_18687,N_18396);
or U18840 (N_18840,N_14886,N_17670);
nor U18841 (N_18841,N_14049,N_13385);
and U18842 (N_18842,N_13942,N_13580);
nand U18843 (N_18843,N_18703,N_15530);
nand U18844 (N_18844,N_16034,N_14464);
xnor U18845 (N_18845,N_13758,N_14373);
or U18846 (N_18846,N_15363,N_14473);
nand U18847 (N_18847,N_17310,N_12678);
and U18848 (N_18848,N_16538,N_16023);
and U18849 (N_18849,N_15500,N_16905);
or U18850 (N_18850,N_14692,N_18130);
nand U18851 (N_18851,N_18503,N_16222);
nand U18852 (N_18852,N_17319,N_18087);
nor U18853 (N_18853,N_13172,N_16828);
nor U18854 (N_18854,N_16548,N_17080);
nand U18855 (N_18855,N_17379,N_13466);
nor U18856 (N_18856,N_17435,N_14525);
and U18857 (N_18857,N_16571,N_14985);
xnor U18858 (N_18858,N_17415,N_17536);
xor U18859 (N_18859,N_18458,N_13135);
or U18860 (N_18860,N_18304,N_18611);
nor U18861 (N_18861,N_13035,N_17634);
and U18862 (N_18862,N_18589,N_17646);
or U18863 (N_18863,N_18061,N_12819);
nor U18864 (N_18864,N_14153,N_14416);
and U18865 (N_18865,N_18093,N_15517);
and U18866 (N_18866,N_15164,N_18662);
or U18867 (N_18867,N_16561,N_16271);
or U18868 (N_18868,N_13171,N_16799);
nand U18869 (N_18869,N_14297,N_12743);
nor U18870 (N_18870,N_14654,N_14547);
nor U18871 (N_18871,N_12754,N_17992);
and U18872 (N_18872,N_13562,N_14288);
nand U18873 (N_18873,N_15589,N_12906);
nand U18874 (N_18874,N_15829,N_14655);
nor U18875 (N_18875,N_16659,N_14989);
nor U18876 (N_18876,N_12648,N_17855);
or U18877 (N_18877,N_17601,N_13754);
nor U18878 (N_18878,N_15715,N_14885);
or U18879 (N_18879,N_14353,N_14414);
nor U18880 (N_18880,N_16932,N_16501);
nor U18881 (N_18881,N_14089,N_15022);
or U18882 (N_18882,N_17489,N_12722);
and U18883 (N_18883,N_18402,N_12840);
xnor U18884 (N_18884,N_16698,N_14573);
nand U18885 (N_18885,N_12632,N_17370);
and U18886 (N_18886,N_14128,N_14862);
or U18887 (N_18887,N_16856,N_14859);
or U18888 (N_18888,N_12786,N_13262);
and U18889 (N_18889,N_12962,N_16809);
xnor U18890 (N_18890,N_14081,N_15101);
nor U18891 (N_18891,N_17180,N_12866);
and U18892 (N_18892,N_13057,N_13790);
nor U18893 (N_18893,N_14449,N_15126);
nor U18894 (N_18894,N_12690,N_16875);
nor U18895 (N_18895,N_14226,N_14344);
nor U18896 (N_18896,N_18222,N_12612);
nor U18897 (N_18897,N_15964,N_16305);
nor U18898 (N_18898,N_13305,N_12631);
or U18899 (N_18899,N_16946,N_12776);
nand U18900 (N_18900,N_15763,N_18710);
nand U18901 (N_18901,N_17207,N_17767);
and U18902 (N_18902,N_18097,N_16554);
nand U18903 (N_18903,N_17575,N_17822);
nand U18904 (N_18904,N_15380,N_17562);
nand U18905 (N_18905,N_17225,N_16781);
xor U18906 (N_18906,N_18475,N_17981);
or U18907 (N_18907,N_16287,N_17338);
nor U18908 (N_18908,N_16628,N_14938);
xor U18909 (N_18909,N_15540,N_17936);
nor U18910 (N_18910,N_15104,N_18606);
xnor U18911 (N_18911,N_17306,N_18018);
and U18912 (N_18912,N_14699,N_15420);
or U18913 (N_18913,N_17045,N_14102);
nor U18914 (N_18914,N_18508,N_12970);
and U18915 (N_18915,N_15701,N_14813);
or U18916 (N_18916,N_14844,N_13312);
and U18917 (N_18917,N_18356,N_18208);
xnor U18918 (N_18918,N_15328,N_16007);
nor U18919 (N_18919,N_15952,N_15923);
nand U18920 (N_18920,N_14808,N_15096);
nand U18921 (N_18921,N_14235,N_17889);
xor U18922 (N_18922,N_13344,N_17757);
xnor U18923 (N_18923,N_18075,N_15193);
or U18924 (N_18924,N_14728,N_17247);
xor U18925 (N_18925,N_15562,N_16405);
nand U18926 (N_18926,N_12548,N_15310);
or U18927 (N_18927,N_13455,N_15696);
nor U18928 (N_18928,N_18332,N_18512);
and U18929 (N_18929,N_17327,N_14438);
and U18930 (N_18930,N_13153,N_17680);
nand U18931 (N_18931,N_14632,N_14935);
or U18932 (N_18932,N_15878,N_13705);
nand U18933 (N_18933,N_18015,N_15179);
nor U18934 (N_18934,N_13618,N_14325);
nor U18935 (N_18935,N_14502,N_17004);
nand U18936 (N_18936,N_13164,N_14977);
nand U18937 (N_18937,N_18228,N_17663);
nand U18938 (N_18938,N_16719,N_15598);
xnor U18939 (N_18939,N_16077,N_13460);
nand U18940 (N_18940,N_16382,N_18202);
or U18941 (N_18941,N_17104,N_13213);
nand U18942 (N_18942,N_18590,N_15266);
nor U18943 (N_18943,N_17668,N_15256);
nand U18944 (N_18944,N_12689,N_16508);
or U18945 (N_18945,N_17262,N_12567);
nand U18946 (N_18946,N_14854,N_15178);
nor U18947 (N_18947,N_12778,N_15231);
and U18948 (N_18948,N_14961,N_13877);
xnor U18949 (N_18949,N_13316,N_12658);
or U18950 (N_18950,N_16408,N_16331);
or U18951 (N_18951,N_18659,N_12719);
or U18952 (N_18952,N_14101,N_18420);
xnor U18953 (N_18953,N_17550,N_14806);
and U18954 (N_18954,N_18213,N_13334);
nand U18955 (N_18955,N_15628,N_13200);
nand U18956 (N_18956,N_12622,N_15515);
and U18957 (N_18957,N_16958,N_15583);
nand U18958 (N_18958,N_14881,N_13223);
nand U18959 (N_18959,N_14579,N_12793);
or U18960 (N_18960,N_13125,N_15211);
nor U18961 (N_18961,N_17795,N_12986);
and U18962 (N_18962,N_15894,N_17062);
and U18963 (N_18963,N_18206,N_17745);
nand U18964 (N_18964,N_14475,N_13040);
nor U18965 (N_18965,N_14779,N_16811);
and U18966 (N_18966,N_15019,N_15246);
nor U18967 (N_18967,N_13219,N_13878);
nor U18968 (N_18968,N_18566,N_14174);
nand U18969 (N_18969,N_13299,N_14154);
nand U18970 (N_18970,N_14534,N_13557);
nor U18971 (N_18971,N_18701,N_16858);
nor U18972 (N_18972,N_16701,N_13517);
nand U18973 (N_18973,N_16020,N_15846);
nor U18974 (N_18974,N_14307,N_13173);
and U18975 (N_18975,N_14394,N_17690);
and U18976 (N_18976,N_17197,N_16087);
nand U18977 (N_18977,N_12582,N_18696);
xor U18978 (N_18978,N_13480,N_15316);
or U18979 (N_18979,N_14248,N_14903);
nand U18980 (N_18980,N_14251,N_16380);
and U18981 (N_18981,N_15912,N_16539);
xor U18982 (N_18982,N_18628,N_13018);
or U18983 (N_18983,N_18722,N_17912);
nor U18984 (N_18984,N_16448,N_12640);
nor U18985 (N_18985,N_18273,N_16993);
xor U18986 (N_18986,N_12521,N_13991);
xnor U18987 (N_18987,N_16521,N_14166);
nand U18988 (N_18988,N_18650,N_14802);
or U18989 (N_18989,N_17657,N_18244);
and U18990 (N_18990,N_14604,N_18585);
and U18991 (N_18991,N_13440,N_17436);
and U18992 (N_18992,N_15272,N_16915);
or U18993 (N_18993,N_17812,N_14921);
nor U18994 (N_18994,N_17136,N_16675);
and U18995 (N_18995,N_16687,N_12684);
nand U18996 (N_18996,N_14074,N_15522);
or U18997 (N_18997,N_14633,N_12895);
or U18998 (N_18998,N_18594,N_16436);
nor U18999 (N_18999,N_14617,N_15271);
or U19000 (N_19000,N_12977,N_15177);
xnor U19001 (N_19001,N_17541,N_15307);
and U19002 (N_19002,N_17824,N_14837);
or U19003 (N_19003,N_13257,N_13893);
or U19004 (N_19004,N_12604,N_16909);
xor U19005 (N_19005,N_16552,N_15326);
or U19006 (N_19006,N_17922,N_14593);
nor U19007 (N_19007,N_17701,N_17940);
nand U19008 (N_19008,N_16999,N_13356);
nor U19009 (N_19009,N_15214,N_15007);
or U19010 (N_19010,N_17205,N_12509);
and U19011 (N_19011,N_14066,N_14974);
xor U19012 (N_19012,N_13386,N_16558);
and U19013 (N_19013,N_15641,N_14126);
and U19014 (N_19014,N_13937,N_17244);
nand U19015 (N_19015,N_14706,N_13046);
nor U19016 (N_19016,N_12586,N_16527);
and U19017 (N_19017,N_13746,N_18597);
nor U19018 (N_19018,N_15809,N_15005);
and U19019 (N_19019,N_14422,N_14011);
and U19020 (N_19020,N_16243,N_18540);
or U19021 (N_19021,N_18248,N_13183);
or U19022 (N_19022,N_13062,N_14163);
and U19023 (N_19023,N_18110,N_17395);
or U19024 (N_19024,N_15248,N_14406);
and U19025 (N_19025,N_13413,N_13740);
nand U19026 (N_19026,N_12900,N_18415);
nor U19027 (N_19027,N_15336,N_12940);
and U19028 (N_19028,N_15804,N_13446);
or U19029 (N_19029,N_15513,N_16280);
nand U19030 (N_19030,N_16172,N_13103);
nand U19031 (N_19031,N_18299,N_18197);
and U19032 (N_19032,N_16472,N_18587);
nor U19033 (N_19033,N_13851,N_13639);
xor U19034 (N_19034,N_17784,N_12738);
and U19035 (N_19035,N_13988,N_16107);
nand U19036 (N_19036,N_14214,N_16174);
nand U19037 (N_19037,N_15581,N_18677);
or U19038 (N_19038,N_13060,N_15822);
and U19039 (N_19039,N_13134,N_14912);
and U19040 (N_19040,N_17148,N_13782);
xor U19041 (N_19041,N_13028,N_16772);
and U19042 (N_19042,N_15864,N_17764);
xnor U19043 (N_19043,N_14545,N_14819);
nand U19044 (N_19044,N_14486,N_16559);
nor U19045 (N_19045,N_14062,N_14130);
nor U19046 (N_19046,N_18252,N_15511);
nand U19047 (N_19047,N_13362,N_17255);
nand U19048 (N_19048,N_17762,N_14342);
and U19049 (N_19049,N_17772,N_14853);
nor U19050 (N_19050,N_18275,N_15728);
xor U19051 (N_19051,N_16544,N_12881);
nor U19052 (N_19052,N_17744,N_16292);
or U19053 (N_19053,N_13972,N_15134);
or U19054 (N_19054,N_14663,N_13017);
and U19055 (N_19055,N_15660,N_17869);
and U19056 (N_19056,N_16202,N_18143);
xor U19057 (N_19057,N_15603,N_12893);
nor U19058 (N_19058,N_18315,N_12818);
nor U19059 (N_19059,N_17689,N_18454);
xnor U19060 (N_19060,N_17109,N_14976);
nand U19061 (N_19061,N_17857,N_15772);
or U19062 (N_19062,N_17002,N_15213);
xnor U19063 (N_19063,N_17280,N_12966);
nor U19064 (N_19064,N_17705,N_16830);
nand U19065 (N_19065,N_16689,N_16429);
or U19066 (N_19066,N_12644,N_17307);
nor U19067 (N_19067,N_13025,N_15327);
or U19068 (N_19068,N_17376,N_17697);
xnor U19069 (N_19069,N_14405,N_16991);
nor U19070 (N_19070,N_16748,N_14334);
nor U19071 (N_19071,N_15280,N_13950);
nor U19072 (N_19072,N_17427,N_18283);
or U19073 (N_19073,N_18414,N_17488);
and U19074 (N_19074,N_16633,N_16332);
nor U19075 (N_19075,N_14095,N_15305);
nor U19076 (N_19076,N_13596,N_15329);
nor U19077 (N_19077,N_16976,N_14237);
nor U19078 (N_19078,N_14937,N_13658);
or U19079 (N_19079,N_16677,N_13646);
nand U19080 (N_19080,N_12523,N_16081);
or U19081 (N_19081,N_14072,N_16874);
xor U19082 (N_19082,N_15494,N_15863);
or U19083 (N_19083,N_14477,N_17237);
nand U19084 (N_19084,N_14058,N_16250);
or U19085 (N_19085,N_17946,N_17907);
xnor U19086 (N_19086,N_18221,N_18306);
nor U19087 (N_19087,N_17653,N_13537);
or U19088 (N_19088,N_17994,N_13787);
nor U19089 (N_19089,N_15176,N_14627);
nand U19090 (N_19090,N_13817,N_15204);
and U19091 (N_19091,N_15723,N_14258);
nor U19092 (N_19092,N_14093,N_12968);
nor U19093 (N_19093,N_14548,N_16136);
nor U19094 (N_19094,N_13648,N_15874);
and U19095 (N_19095,N_17369,N_14759);
or U19096 (N_19096,N_17266,N_15974);
and U19097 (N_19097,N_17892,N_18249);
xnor U19098 (N_19098,N_14086,N_17563);
xor U19099 (N_19099,N_12815,N_17532);
nor U19100 (N_19100,N_14556,N_14120);
nor U19101 (N_19101,N_12967,N_15401);
or U19102 (N_19102,N_15845,N_17441);
nor U19103 (N_19103,N_17654,N_16647);
or U19104 (N_19104,N_17194,N_13513);
nor U19105 (N_19105,N_15854,N_12855);
and U19106 (N_19106,N_14114,N_18325);
xor U19107 (N_19107,N_15985,N_13124);
nand U19108 (N_19108,N_16914,N_14087);
nand U19109 (N_19109,N_18101,N_14221);
and U19110 (N_19110,N_16597,N_15276);
or U19111 (N_19111,N_16740,N_16211);
and U19112 (N_19112,N_12989,N_17919);
nand U19113 (N_19113,N_14263,N_16003);
or U19114 (N_19114,N_13276,N_12988);
and U19115 (N_19115,N_14277,N_16208);
nand U19116 (N_19116,N_14669,N_15529);
and U19117 (N_19117,N_14708,N_13050);
nor U19118 (N_19118,N_14978,N_17937);
and U19119 (N_19119,N_14158,N_18341);
and U19120 (N_19120,N_12985,N_14563);
nand U19121 (N_19121,N_13081,N_16308);
and U19122 (N_19122,N_18425,N_12923);
nor U19123 (N_19123,N_14319,N_16090);
or U19124 (N_19124,N_14091,N_15170);
or U19125 (N_19125,N_16386,N_14879);
or U19126 (N_19126,N_14027,N_12804);
nand U19127 (N_19127,N_15639,N_15760);
xor U19128 (N_19128,N_13019,N_16589);
nand U19129 (N_19129,N_16489,N_14882);
or U19130 (N_19130,N_17829,N_18698);
nand U19131 (N_19131,N_14581,N_13948);
xor U19132 (N_19132,N_16520,N_16457);
nor U19133 (N_19133,N_15151,N_16666);
nand U19134 (N_19134,N_14433,N_16346);
or U19135 (N_19135,N_16741,N_15223);
or U19136 (N_19136,N_14138,N_18541);
nand U19137 (N_19137,N_18121,N_15789);
xnor U19138 (N_19138,N_14271,N_14164);
nor U19139 (N_19139,N_13031,N_15459);
or U19140 (N_19140,N_16636,N_14644);
or U19141 (N_19141,N_14343,N_18564);
or U19142 (N_19142,N_17951,N_15827);
nand U19143 (N_19143,N_15069,N_17093);
and U19144 (N_19144,N_13524,N_13829);
nor U19145 (N_19145,N_13692,N_17743);
and U19146 (N_19146,N_18358,N_15813);
or U19147 (N_19147,N_13642,N_16795);
and U19148 (N_19148,N_17468,N_12891);
nand U19149 (N_19149,N_13635,N_13956);
and U19150 (N_19150,N_15454,N_14127);
nor U19151 (N_19151,N_18518,N_14615);
nand U19152 (N_19152,N_13306,N_18226);
xor U19153 (N_19153,N_16549,N_12823);
nor U19154 (N_19154,N_13729,N_18607);
xor U19155 (N_19155,N_14872,N_12905);
nor U19156 (N_19156,N_15877,N_13636);
or U19157 (N_19157,N_16818,N_17135);
nand U19158 (N_19158,N_15503,N_15646);
or U19159 (N_19159,N_15222,N_18272);
nor U19160 (N_19160,N_13641,N_16700);
nand U19161 (N_19161,N_18003,N_18666);
or U19162 (N_19162,N_14594,N_12590);
nor U19163 (N_19163,N_18613,N_15203);
nor U19164 (N_19164,N_17979,N_14971);
nand U19165 (N_19165,N_13565,N_17811);
nor U19166 (N_19166,N_15528,N_15818);
nor U19167 (N_19167,N_16540,N_17437);
and U19168 (N_19168,N_13560,N_18162);
nand U19169 (N_19169,N_13655,N_16012);
or U19170 (N_19170,N_18581,N_18547);
or U19171 (N_19171,N_18343,N_18140);
xnor U19172 (N_19172,N_17193,N_16956);
nand U19173 (N_19173,N_14677,N_17787);
and U19174 (N_19174,N_17948,N_13421);
and U19175 (N_19175,N_17048,N_13249);
nor U19176 (N_19176,N_14429,N_13041);
nor U19177 (N_19177,N_13958,N_16779);
and U19178 (N_19178,N_14659,N_18023);
or U19179 (N_19179,N_17322,N_16345);
or U19180 (N_19180,N_17371,N_17598);
nor U19181 (N_19181,N_18282,N_14415);
nor U19182 (N_19182,N_14245,N_15649);
nand U19183 (N_19183,N_17304,N_13204);
or U19184 (N_19184,N_14690,N_16312);
nor U19185 (N_19185,N_13732,N_16319);
and U19186 (N_19186,N_13576,N_15106);
xnor U19187 (N_19187,N_17449,N_18237);
and U19188 (N_19188,N_16560,N_13611);
nor U19189 (N_19189,N_13070,N_15457);
or U19190 (N_19190,N_16347,N_14898);
xor U19191 (N_19191,N_12697,N_16102);
xnor U19192 (N_19192,N_13825,N_15676);
nand U19193 (N_19193,N_14570,N_17259);
xor U19194 (N_19194,N_18120,N_12959);
nand U19195 (N_19195,N_14362,N_14740);
nor U19196 (N_19196,N_14358,N_13764);
nand U19197 (N_19197,N_13903,N_17260);
or U19198 (N_19198,N_15502,N_13426);
or U19199 (N_19199,N_18133,N_18626);
nand U19200 (N_19200,N_13706,N_15062);
xnor U19201 (N_19201,N_13023,N_15133);
and U19202 (N_19202,N_15183,N_18484);
nor U19203 (N_19203,N_17715,N_13731);
and U19204 (N_19204,N_13485,N_14889);
or U19205 (N_19205,N_16138,N_18570);
and U19206 (N_19206,N_14378,N_16998);
and U19207 (N_19207,N_13788,N_14636);
nor U19208 (N_19208,N_18647,N_15774);
and U19209 (N_19209,N_14159,N_15718);
nor U19210 (N_19210,N_13906,N_17236);
and U19211 (N_19211,N_14048,N_13331);
and U19212 (N_19212,N_15880,N_16227);
or U19213 (N_19213,N_12767,N_16248);
nor U19214 (N_19214,N_16485,N_17599);
and U19215 (N_19215,N_17311,N_17530);
nor U19216 (N_19216,N_17816,N_14666);
nor U19217 (N_19217,N_15933,N_17731);
and U19218 (N_19218,N_16255,N_17916);
or U19219 (N_19219,N_16646,N_16703);
or U19220 (N_19220,N_12723,N_16969);
nand U19221 (N_19221,N_14206,N_15677);
nor U19222 (N_19222,N_16133,N_18164);
nand U19223 (N_19223,N_13767,N_14283);
xor U19224 (N_19224,N_18600,N_18410);
and U19225 (N_19225,N_17451,N_13669);
nand U19226 (N_19226,N_17667,N_14281);
and U19227 (N_19227,N_12558,N_16746);
nand U19228 (N_19228,N_17538,N_16066);
or U19229 (N_19229,N_13619,N_16887);
nor U19230 (N_19230,N_16826,N_17897);
or U19231 (N_19231,N_16446,N_14914);
nand U19232 (N_19232,N_16445,N_14233);
and U19233 (N_19233,N_12515,N_15250);
or U19234 (N_19234,N_12530,N_14268);
nor U19235 (N_19235,N_14688,N_17399);
nor U19236 (N_19236,N_13924,N_14957);
xor U19237 (N_19237,N_17524,N_17021);
nor U19238 (N_19238,N_13071,N_14832);
and U19239 (N_19239,N_13377,N_13253);
nor U19240 (N_19240,N_13075,N_15590);
and U19241 (N_19241,N_13841,N_15642);
nor U19242 (N_19242,N_17250,N_15750);
nor U19243 (N_19243,N_15883,N_18220);
nor U19244 (N_19244,N_14784,N_13228);
and U19245 (N_19245,N_17173,N_12563);
and U19246 (N_19246,N_16710,N_13994);
nor U19247 (N_19247,N_13925,N_13854);
or U19248 (N_19248,N_16643,N_17057);
nand U19249 (N_19249,N_13954,N_13320);
nor U19250 (N_19250,N_13520,N_14939);
nor U19251 (N_19251,N_12976,N_17377);
or U19252 (N_19252,N_16722,N_15785);
or U19253 (N_19253,N_15644,N_13497);
nor U19254 (N_19254,N_17878,N_13008);
nand U19255 (N_19255,N_15770,N_16718);
or U19256 (N_19256,N_14625,N_15673);
nor U19257 (N_19257,N_13637,N_12583);
nor U19258 (N_19258,N_13727,N_16141);
or U19259 (N_19259,N_14064,N_18353);
and U19260 (N_19260,N_14302,N_12843);
and U19261 (N_19261,N_14046,N_14349);
and U19262 (N_19262,N_16266,N_18138);
and U19263 (N_19263,N_14367,N_18223);
or U19264 (N_19264,N_13496,N_16812);
nor U19265 (N_19265,N_15403,N_14493);
nand U19266 (N_19266,N_18324,N_17580);
and U19267 (N_19267,N_13021,N_12756);
nor U19268 (N_19268,N_13327,N_14732);
xnor U19269 (N_19269,N_15306,N_17125);
xor U19270 (N_19270,N_16859,N_14363);
nand U19271 (N_19271,N_15340,N_14902);
nor U19272 (N_19272,N_14803,N_17658);
nand U19273 (N_19273,N_13273,N_12836);
xor U19274 (N_19274,N_14037,N_17746);
xor U19275 (N_19275,N_16857,N_17028);
and U19276 (N_19276,N_14584,N_13811);
nand U19277 (N_19277,N_18102,N_16434);
and U19278 (N_19278,N_13365,N_13112);
nor U19279 (N_19279,N_14043,N_14476);
nor U19280 (N_19280,N_13490,N_14958);
nor U19281 (N_19281,N_15499,N_18403);
and U19282 (N_19282,N_16717,N_15593);
or U19283 (N_19283,N_15421,N_13128);
and U19284 (N_19284,N_13295,N_14150);
or U19285 (N_19285,N_17790,N_17792);
nand U19286 (N_19286,N_15285,N_17941);
nor U19287 (N_19287,N_14915,N_17722);
nor U19288 (N_19288,N_14665,N_16578);
nor U19289 (N_19289,N_13268,N_15379);
nor U19290 (N_19290,N_14498,N_17184);
and U19291 (N_19291,N_15756,N_17181);
nor U19292 (N_19292,N_12742,N_16103);
nand U19293 (N_19293,N_13738,N_12536);
nor U19294 (N_19294,N_17886,N_15901);
nand U19295 (N_19295,N_16054,N_14892);
or U19296 (N_19296,N_18572,N_13250);
or U19297 (N_19297,N_15269,N_14275);
and U19298 (N_19298,N_14021,N_14168);
or U19299 (N_19299,N_14739,N_18106);
or U19300 (N_19300,N_13503,N_17224);
and U19301 (N_19301,N_12633,N_13303);
nor U19302 (N_19302,N_17210,N_18467);
nor U19303 (N_19303,N_16567,N_13235);
nor U19304 (N_19304,N_18695,N_16363);
nor U19305 (N_19305,N_13332,N_17407);
and U19306 (N_19306,N_17138,N_12746);
and U19307 (N_19307,N_14117,N_16423);
nor U19308 (N_19308,N_15228,N_16058);
or U19309 (N_19309,N_18636,N_15708);
xor U19310 (N_19310,N_18339,N_17358);
nand U19311 (N_19311,N_12516,N_14664);
nand U19312 (N_19312,N_13345,N_17393);
nand U19313 (N_19313,N_14485,N_14259);
or U19314 (N_19314,N_17042,N_18046);
xnor U19315 (N_19315,N_14927,N_15796);
xnor U19316 (N_19316,N_13484,N_13607);
xnor U19317 (N_19317,N_17628,N_13572);
nor U19318 (N_19318,N_14161,N_17142);
and U19319 (N_19319,N_16449,N_18741);
xor U19320 (N_19320,N_15695,N_13237);
and U19321 (N_19321,N_15702,N_17461);
or U19322 (N_19322,N_13267,N_15468);
and U19323 (N_19323,N_14050,N_16458);
and U19324 (N_19324,N_13117,N_16361);
nand U19325 (N_19325,N_17206,N_18715);
and U19326 (N_19326,N_13967,N_13939);
nor U19327 (N_19327,N_16794,N_18638);
or U19328 (N_19328,N_15820,N_15569);
nor U19329 (N_19329,N_12889,N_16681);
and U19330 (N_19330,N_16004,N_15445);
and U19331 (N_19331,N_16639,N_16025);
and U19332 (N_19332,N_18435,N_14273);
nor U19333 (N_19333,N_16247,N_13077);
nor U19334 (N_19334,N_18502,N_15006);
nand U19335 (N_19335,N_16881,N_16062);
xor U19336 (N_19336,N_15795,N_13379);
nor U19337 (N_19337,N_16039,N_15705);
nor U19338 (N_19338,N_16483,N_14599);
and U19339 (N_19339,N_14614,N_14376);
xor U19340 (N_19340,N_15903,N_17666);
nor U19341 (N_19341,N_18416,N_18655);
or U19342 (N_19342,N_13283,N_13030);
nand U19343 (N_19343,N_18039,N_15663);
nand U19344 (N_19344,N_18187,N_16640);
nand U19345 (N_19345,N_14612,N_14023);
nor U19346 (N_19346,N_17157,N_18105);
and U19347 (N_19347,N_16793,N_16109);
nor U19348 (N_19348,N_14750,N_15165);
nor U19349 (N_19349,N_13186,N_15274);
nand U19350 (N_19350,N_18692,N_17880);
and U19351 (N_19351,N_17607,N_16845);
and U19352 (N_19352,N_14098,N_16215);
and U19353 (N_19353,N_12687,N_15037);
or U19354 (N_19354,N_15312,N_18083);
nor U19355 (N_19355,N_15323,N_12641);
nor U19356 (N_19356,N_15984,N_15664);
and U19357 (N_19357,N_18705,N_18464);
and U19358 (N_19358,N_17345,N_13941);
nand U19359 (N_19359,N_13766,N_14842);
and U19360 (N_19360,N_16671,N_15549);
and U19361 (N_19361,N_12748,N_17526);
or U19362 (N_19362,N_14328,N_15599);
or U19363 (N_19363,N_14054,N_16026);
nand U19364 (N_19364,N_17613,N_18417);
nand U19365 (N_19365,N_16426,N_12745);
nand U19366 (N_19366,N_18509,N_13867);
xor U19367 (N_19367,N_18129,N_12514);
nand U19368 (N_19368,N_17699,N_13552);
and U19369 (N_19369,N_18082,N_15751);
and U19370 (N_19370,N_13522,N_13026);
and U19371 (N_19371,N_16656,N_15948);
xnor U19372 (N_19372,N_17504,N_17771);
or U19373 (N_19373,N_14182,N_18658);
or U19374 (N_19374,N_16275,N_12614);
nand U19375 (N_19375,N_12553,N_18525);
nand U19376 (N_19376,N_18259,N_16239);
nand U19377 (N_19377,N_16805,N_13900);
or U19378 (N_19378,N_12806,N_12579);
xnor U19379 (N_19379,N_18555,N_14309);
or U19380 (N_19380,N_18406,N_16091);
nor U19381 (N_19381,N_12808,N_15220);
or U19382 (N_19382,N_14990,N_13561);
nor U19383 (N_19383,N_14847,N_13510);
nand U19384 (N_19384,N_12755,N_14061);
nand U19385 (N_19385,N_16529,N_17245);
and U19386 (N_19386,N_14234,N_13979);
nand U19387 (N_19387,N_18371,N_15981);
nor U19388 (N_19388,N_15504,N_17510);
nand U19389 (N_19389,N_15890,N_14825);
or U19390 (N_19390,N_18285,N_15095);
nand U19391 (N_19391,N_14016,N_16821);
nor U19392 (N_19392,N_13794,N_18177);
nor U19393 (N_19393,N_17299,N_18233);
nand U19394 (N_19394,N_13833,N_13009);
or U19395 (N_19395,N_13151,N_16177);
and U19396 (N_19396,N_13240,N_13473);
or U19397 (N_19397,N_17052,N_13653);
and U19398 (N_19398,N_17807,N_15103);
or U19399 (N_19399,N_15814,N_17398);
or U19400 (N_19400,N_15392,N_15426);
nor U19401 (N_19401,N_16630,N_17198);
nand U19402 (N_19402,N_16726,N_15585);
nor U19403 (N_19403,N_17788,N_13489);
or U19404 (N_19404,N_16231,N_15163);
nand U19405 (N_19405,N_14350,N_17894);
or U19406 (N_19406,N_14170,N_13987);
nor U19407 (N_19407,N_18468,N_17196);
xnor U19408 (N_19408,N_16317,N_17442);
nand U19409 (N_19409,N_16660,N_16205);
and U19410 (N_19410,N_14942,N_13184);
and U19411 (N_19411,N_15949,N_18496);
nand U19412 (N_19412,N_12653,N_14679);
nand U19413 (N_19413,N_18193,N_14843);
nand U19414 (N_19414,N_17846,N_13801);
and U19415 (N_19415,N_17323,N_18149);
and U19416 (N_19416,N_14907,N_18660);
or U19417 (N_19417,N_17600,N_14147);
nor U19418 (N_19418,N_17497,N_12956);
and U19419 (N_19419,N_15265,N_15734);
nor U19420 (N_19420,N_18480,N_18398);
and U19421 (N_19421,N_14834,N_18577);
nor U19422 (N_19422,N_14348,N_13033);
nor U19423 (N_19423,N_17665,N_16920);
nor U19424 (N_19424,N_17611,N_17543);
and U19425 (N_19425,N_13374,N_17302);
nor U19426 (N_19426,N_13462,N_13749);
nand U19427 (N_19427,N_14077,N_12885);
nor U19428 (N_19428,N_16955,N_16966);
nand U19429 (N_19429,N_13786,N_14734);
and U19430 (N_19430,N_15000,N_14603);
nor U19431 (N_19431,N_13804,N_13842);
nand U19432 (N_19432,N_16067,N_15629);
nand U19433 (N_19433,N_17014,N_14705);
and U19434 (N_19434,N_16988,N_14754);
nand U19435 (N_19435,N_16083,N_18035);
xor U19436 (N_19436,N_18179,N_17566);
and U19437 (N_19437,N_13238,N_13680);
or U19438 (N_19438,N_14339,N_17025);
and U19439 (N_19439,N_12953,N_16028);
and U19440 (N_19440,N_15205,N_17274);
nor U19441 (N_19441,N_12606,N_13177);
nor U19442 (N_19442,N_16262,N_14578);
nand U19443 (N_19443,N_18069,N_13187);
or U19444 (N_19444,N_16218,N_12878);
nand U19445 (N_19445,N_14673,N_14090);
and U19446 (N_19446,N_17440,N_16410);
nand U19447 (N_19447,N_16753,N_12869);
nor U19448 (N_19448,N_16632,N_17469);
xor U19449 (N_19449,N_16513,N_18423);
nor U19450 (N_19450,N_14103,N_18579);
or U19451 (N_19451,N_16356,N_12506);
nor U19452 (N_19452,N_16488,N_12731);
nand U19453 (N_19453,N_15159,N_17964);
nor U19454 (N_19454,N_13810,N_17130);
and U19455 (N_19455,N_15268,N_14505);
nor U19456 (N_19456,N_17815,N_16162);
xor U19457 (N_19457,N_16584,N_16749);
nand U19458 (N_19458,N_14356,N_15388);
xnor U19459 (N_19459,N_17209,N_18319);
nand U19460 (N_19460,N_17336,N_14238);
nor U19461 (N_19461,N_13944,N_14008);
nand U19462 (N_19462,N_17734,N_18654);
nor U19463 (N_19463,N_18088,N_12669);
nor U19464 (N_19464,N_16364,N_17276);
or U19465 (N_19465,N_12949,N_14590);
nand U19466 (N_19466,N_16819,N_15072);
and U19467 (N_19467,N_18131,N_13595);
or U19468 (N_19468,N_18378,N_13449);
and U19469 (N_19469,N_13501,N_13061);
or U19470 (N_19470,N_16616,N_16475);
nand U19471 (N_19471,N_14382,N_15397);
nor U19472 (N_19472,N_18592,N_15934);
or U19473 (N_19473,N_14398,N_12564);
or U19474 (N_19474,N_13161,N_12592);
and U19475 (N_19475,N_13254,N_14434);
nand U19476 (N_19476,N_13406,N_18314);
or U19477 (N_19477,N_12926,N_17284);
or U19478 (N_19478,N_13791,N_15994);
or U19479 (N_19479,N_13336,N_14208);
xor U19480 (N_19480,N_18348,N_14137);
and U19481 (N_19481,N_12624,N_14149);
or U19482 (N_19482,N_16574,N_12730);
and U19483 (N_19483,N_16572,N_15150);
or U19484 (N_19484,N_16088,N_14743);
nor U19485 (N_19485,N_17817,N_13159);
nand U19486 (N_19486,N_17949,N_15730);
nand U19487 (N_19487,N_16153,N_17717);
and U19488 (N_19488,N_15202,N_18168);
and U19489 (N_19489,N_18427,N_16115);
nand U19490 (N_19490,N_14560,N_18312);
nand U19491 (N_19491,N_17662,N_18501);
or U19492 (N_19492,N_18258,N_17839);
and U19493 (N_19493,N_16683,N_14056);
and U19494 (N_19494,N_13905,N_14777);
and U19495 (N_19495,N_15738,N_15028);
or U19496 (N_19496,N_15027,N_15724);
xnor U19497 (N_19497,N_15935,N_16581);
or U19498 (N_19498,N_15800,N_13022);
xnor U19499 (N_19499,N_13751,N_18738);
and U19500 (N_19500,N_13288,N_15758);
nand U19501 (N_19501,N_12546,N_13106);
and U19502 (N_19502,N_16506,N_15859);
and U19503 (N_19503,N_14207,N_13529);
nand U19504 (N_19504,N_18706,N_13175);
or U19505 (N_19505,N_18536,N_17267);
nor U19506 (N_19506,N_17523,N_16590);
xnor U19507 (N_19507,N_13393,N_16038);
nor U19508 (N_19508,N_14201,N_12873);
nand U19509 (N_19509,N_13291,N_18235);
nor U19510 (N_19510,N_15416,N_15914);
and U19511 (N_19511,N_12764,N_13042);
nand U19512 (N_19512,N_16124,N_14553);
nand U19513 (N_19513,N_17228,N_16203);
and U19514 (N_19514,N_14588,N_18400);
nand U19515 (N_19515,N_15749,N_14453);
nor U19516 (N_19516,N_15088,N_17609);
xnor U19517 (N_19517,N_13416,N_16949);
or U19518 (N_19518,N_18245,N_12568);
or U19519 (N_19519,N_15852,N_18517);
or U19520 (N_19520,N_18739,N_16478);
or U19521 (N_19521,N_18616,N_15697);
xor U19522 (N_19522,N_13211,N_17782);
nand U19523 (N_19523,N_16577,N_18707);
nand U19524 (N_19524,N_14219,N_16122);
nor U19525 (N_19525,N_13621,N_13352);
or U19526 (N_19526,N_14542,N_14946);
nand U19527 (N_19527,N_13359,N_15999);
nand U19528 (N_19528,N_12752,N_13468);
nand U19529 (N_19529,N_14890,N_12867);
nor U19530 (N_19530,N_15482,N_15922);
and U19531 (N_19531,N_15349,N_18013);
nand U19532 (N_19532,N_16902,N_14575);
and U19533 (N_19533,N_16713,N_17935);
nand U19534 (N_19534,N_13866,N_13323);
or U19535 (N_19535,N_17683,N_14122);
nor U19536 (N_19536,N_13045,N_17413);
nand U19537 (N_19537,N_14979,N_17603);
or U19538 (N_19538,N_14051,N_15656);
xnor U19539 (N_19539,N_16302,N_13425);
nor U19540 (N_19540,N_13222,N_14360);
nand U19541 (N_19541,N_13394,N_15498);
nor U19542 (N_19542,N_14587,N_17401);
xnor U19543 (N_19543,N_18580,N_18231);
nand U19544 (N_19544,N_18559,N_12862);
or U19545 (N_19545,N_14936,N_14185);
or U19546 (N_19546,N_14392,N_15413);
or U19547 (N_19547,N_13170,N_12561);
or U19548 (N_19548,N_15668,N_18210);
nand U19549 (N_19549,N_16186,N_16092);
and U19550 (N_19550,N_17841,N_14262);
or U19551 (N_19551,N_13616,N_15094);
xnor U19552 (N_19552,N_17200,N_15840);
or U19553 (N_19553,N_16188,N_15970);
nand U19554 (N_19554,N_12712,N_18439);
and U19555 (N_19555,N_15357,N_17027);
nor U19556 (N_19556,N_18669,N_18545);
and U19557 (N_19557,N_12569,N_17910);
nor U19558 (N_19558,N_17083,N_13055);
or U19559 (N_19559,N_13717,N_18612);
nand U19560 (N_19560,N_16052,N_15112);
or U19561 (N_19561,N_12736,N_17867);
xnor U19562 (N_19562,N_16525,N_13579);
or U19563 (N_19563,N_16246,N_15058);
and U19564 (N_19564,N_15294,N_18438);
or U19565 (N_19565,N_18326,N_15860);
or U19566 (N_19566,N_12657,N_16502);
nand U19567 (N_19567,N_14402,N_14256);
or U19568 (N_19568,N_15888,N_17796);
or U19569 (N_19569,N_18573,N_14229);
nor U19570 (N_19570,N_17137,N_17380);
xor U19571 (N_19571,N_17615,N_17968);
xnor U19572 (N_19572,N_16463,N_16395);
nor U19573 (N_19573,N_18551,N_18727);
nor U19574 (N_19574,N_14265,N_13367);
nand U19575 (N_19575,N_12987,N_14744);
or U19576 (N_19576,N_14204,N_18591);
nand U19577 (N_19577,N_17428,N_17433);
or U19578 (N_19578,N_16422,N_15471);
and U19579 (N_19579,N_16519,N_17186);
or U19580 (N_19580,N_16980,N_16085);
or U19581 (N_19581,N_12961,N_13836);
nor U19582 (N_19582,N_13534,N_18565);
and U19583 (N_19583,N_17904,N_13324);
or U19584 (N_19584,N_17363,N_18188);
nor U19585 (N_19585,N_18562,N_17314);
and U19586 (N_19586,N_15746,N_13998);
nand U19587 (N_19587,N_18553,N_14355);
nand U19588 (N_19588,N_14200,N_16759);
and U19589 (N_19589,N_18552,N_15386);
nand U19590 (N_19590,N_14855,N_18367);
nand U19591 (N_19591,N_13087,N_13000);
and U19592 (N_19592,N_13687,N_13671);
or U19593 (N_19593,N_14364,N_15462);
xnor U19594 (N_19594,N_12659,N_14657);
nor U19595 (N_19595,N_16168,N_17905);
or U19596 (N_19596,N_18429,N_17711);
and U19597 (N_19597,N_15118,N_13780);
or U19598 (N_19598,N_15146,N_13630);
nor U19599 (N_19599,N_16290,N_14129);
and U19600 (N_19600,N_15776,N_15525);
or U19601 (N_19601,N_14823,N_13964);
nand U19602 (N_19602,N_15152,N_17800);
nand U19603 (N_19603,N_18323,N_18567);
nor U19604 (N_19604,N_16876,N_12995);
nor U19605 (N_19605,N_18265,N_16661);
nand U19606 (N_19606,N_13971,N_18386);
and U19607 (N_19607,N_15608,N_16960);
nor U19608 (N_19608,N_14326,N_14932);
nand U19609 (N_19609,N_15967,N_18539);
nor U19610 (N_19610,N_13453,N_17106);
and U19611 (N_19611,N_13259,N_14304);
nor U19612 (N_19612,N_13960,N_13357);
nor U19613 (N_19613,N_15238,N_14232);
or U19614 (N_19614,N_16161,N_15737);
and U19615 (N_19615,N_14111,N_17724);
xnor U19616 (N_19616,N_13838,N_14773);
or U19617 (N_19617,N_14693,N_15570);
nand U19618 (N_19618,N_18002,N_13246);
and U19619 (N_19619,N_13844,N_12501);
and U19620 (N_19620,N_13197,N_13968);
nor U19621 (N_19621,N_17590,N_18290);
and U19622 (N_19622,N_18103,N_14601);
nand U19623 (N_19623,N_16055,N_16328);
and U19624 (N_19624,N_16295,N_13230);
nand U19625 (N_19625,N_16604,N_16270);
and U19626 (N_19626,N_13512,N_16612);
or U19627 (N_19627,N_16072,N_17034);
or U19628 (N_19628,N_15682,N_12913);
or U19629 (N_19629,N_14012,N_14195);
nand U19630 (N_19630,N_17296,N_17364);
nand U19631 (N_19631,N_18465,N_15561);
and U19632 (N_19632,N_16968,N_15475);
nor U19633 (N_19633,N_15480,N_14134);
and U19634 (N_19634,N_18390,N_13897);
and U19635 (N_19635,N_16716,N_18198);
nor U19636 (N_19636,N_17517,N_13902);
or U19637 (N_19637,N_17119,N_17513);
or U19638 (N_19638,N_15070,N_15905);
or U19639 (N_19639,N_17623,N_15924);
or U19640 (N_19640,N_18697,N_14293);
nor U19641 (N_19641,N_15681,N_17639);
and U19642 (N_19642,N_14622,N_12710);
nor U19643 (N_19643,N_14381,N_13185);
nor U19644 (N_19644,N_12974,N_17661);
or U19645 (N_19645,N_16420,N_14546);
or U19646 (N_19646,N_14720,N_16961);
xnor U19647 (N_19647,N_17645,N_12852);
nor U19648 (N_19648,N_17636,N_12941);
nor U19649 (N_19649,N_17881,N_16371);
nor U19650 (N_19650,N_16706,N_14040);
nor U19651 (N_19651,N_18227,N_12928);
nand U19652 (N_19652,N_18716,N_17467);
nand U19653 (N_19653,N_14063,N_13670);
nor U19654 (N_19654,N_15286,N_14807);
and U19655 (N_19655,N_12825,N_12708);
nor U19656 (N_19656,N_18486,N_16642);
or U19657 (N_19657,N_15961,N_14672);
and U19658 (N_19658,N_13733,N_17594);
and U19659 (N_19659,N_13584,N_15064);
or U19660 (N_19660,N_16011,N_16444);
nor U19661 (N_19661,N_18135,N_17714);
nor U19662 (N_19662,N_13916,N_13896);
nand U19663 (N_19663,N_12503,N_12654);
nand U19664 (N_19664,N_13285,N_14270);
or U19665 (N_19665,N_13210,N_12599);
nand U19666 (N_19666,N_18074,N_14038);
nor U19667 (N_19667,N_16336,N_14084);
or U19668 (N_19668,N_13872,N_17429);
nor U19669 (N_19669,N_17024,N_14013);
xnor U19670 (N_19670,N_13591,N_18316);
nand U19671 (N_19671,N_18347,N_13430);
and U19672 (N_19672,N_16220,N_14115);
or U19673 (N_19673,N_18726,N_18713);
or U19674 (N_19674,N_16783,N_18243);
nor U19675 (N_19675,N_15717,N_16720);
nor U19676 (N_19676,N_13272,N_13602);
nor U19677 (N_19677,N_13207,N_15433);
and U19678 (N_19678,N_14876,N_15706);
nand U19679 (N_19679,N_12547,N_14146);
nor U19680 (N_19680,N_12721,N_16626);
nor U19681 (N_19681,N_17218,N_14497);
nor U19682 (N_19682,N_13467,N_15119);
and U19683 (N_19683,N_15747,N_18134);
and U19684 (N_19684,N_16402,N_15487);
or U19685 (N_19685,N_16106,N_17775);
xor U19686 (N_19686,N_14596,N_17858);
nor U19687 (N_19687,N_18189,N_17147);
and U19688 (N_19688,N_15531,N_18645);
and U19689 (N_19689,N_14749,N_17612);
nand U19690 (N_19690,N_17592,N_18391);
and U19691 (N_19691,N_18123,N_18250);
or U19692 (N_19692,N_16326,N_13957);
nor U19693 (N_19693,N_14794,N_18257);
or U19694 (N_19694,N_16145,N_18331);
nor U19695 (N_19695,N_17204,N_14471);
or U19696 (N_19696,N_12814,N_18279);
nand U19697 (N_19697,N_14900,N_16337);
xor U19698 (N_19698,N_13656,N_16784);
or U19699 (N_19699,N_13373,N_15650);
nand U19700 (N_19700,N_17234,N_16419);
nor U19701 (N_19701,N_15446,N_15679);
or U19702 (N_19702,N_14801,N_15982);
or U19703 (N_19703,N_16693,N_18062);
and U19704 (N_19704,N_12629,N_14082);
nor U19705 (N_19705,N_15395,N_17898);
nor U19706 (N_19706,N_12671,N_13378);
nor U19707 (N_19707,N_13776,N_15754);
or U19708 (N_19708,N_16110,N_16761);
and U19709 (N_19709,N_14067,N_15989);
or U19710 (N_19710,N_14763,N_13578);
nand U19711 (N_19711,N_17146,N_18229);
nor U19712 (N_19712,N_17281,N_17502);
xor U19713 (N_19713,N_14999,N_17980);
nor U19714 (N_19714,N_17955,N_15365);
nand U19715 (N_19715,N_12584,N_15242);
and U19716 (N_19716,N_18499,N_12571);
and U19717 (N_19717,N_16708,N_15210);
xor U19718 (N_19718,N_17160,N_17390);
nand U19719 (N_19719,N_16503,N_15198);
nand U19720 (N_19720,N_17264,N_16199);
xor U19721 (N_19721,N_13100,N_14753);
nor U19722 (N_19722,N_14828,N_13382);
nand U19723 (N_19723,N_17098,N_15128);
nor U19724 (N_19724,N_15099,N_16119);
and U19725 (N_19725,N_14736,N_16747);
or U19726 (N_19726,N_17548,N_15056);
xor U19727 (N_19727,N_14684,N_13149);
nor U19728 (N_19728,N_12813,N_14354);
and U19729 (N_19729,N_15309,N_16200);
nor U19730 (N_19730,N_16197,N_14592);
and U19731 (N_19731,N_18443,N_16031);
and U19732 (N_19732,N_17191,N_18107);
or U19733 (N_19733,N_16670,N_18641);
or U19734 (N_19734,N_16944,N_13507);
nor U19735 (N_19735,N_15342,N_12875);
or U19736 (N_19736,N_15461,N_12701);
nand U19737 (N_19737,N_16394,N_13221);
nand U19738 (N_19738,N_15568,N_15407);
or U19739 (N_19739,N_16839,N_17297);
xor U19740 (N_19740,N_13734,N_16848);
and U19741 (N_19741,N_13640,N_12796);
and U19742 (N_19742,N_15892,N_15465);
nand U19743 (N_19743,N_13452,N_15045);
nand U19744 (N_19744,N_14152,N_16070);
xnor U19745 (N_19745,N_15591,N_14320);
nor U19746 (N_19746,N_18058,N_12720);
or U19747 (N_19747,N_14267,N_14183);
nor U19748 (N_19748,N_14609,N_14361);
or U19749 (N_19749,N_18264,N_17261);
and U19750 (N_19750,N_17110,N_16635);
nand U19751 (N_19751,N_18674,N_15552);
nor U19752 (N_19752,N_15393,N_17350);
or U19753 (N_19753,N_16178,N_17679);
nand U19754 (N_19754,N_16921,N_16167);
or U19755 (N_19755,N_14156,N_16524);
nor U19756 (N_19756,N_16390,N_14875);
and U19757 (N_19757,N_12630,N_17584);
nand U19758 (N_19758,N_14566,N_15116);
nor U19759 (N_19759,N_17577,N_13862);
and U19760 (N_19760,N_14503,N_14909);
or U19761 (N_19761,N_15819,N_16595);
and U19762 (N_19762,N_15257,N_17602);
or U19763 (N_19763,N_13834,N_15474);
or U19764 (N_19764,N_16383,N_16368);
and U19765 (N_19765,N_17604,N_16264);
nand U19766 (N_19766,N_17954,N_17578);
nand U19767 (N_19767,N_15620,N_15296);
and U19768 (N_19768,N_13279,N_14899);
nor U19769 (N_19769,N_13115,N_14555);
nor U19770 (N_19770,N_14399,N_13157);
and U19771 (N_19771,N_15550,N_14867);
or U19772 (N_19772,N_13002,N_13992);
or U19773 (N_19773,N_16334,N_18364);
and U19774 (N_19774,N_16557,N_16546);
and U19775 (N_19775,N_14519,N_16017);
xnor U19776 (N_19776,N_14104,N_18098);
and U19777 (N_19777,N_17957,N_16806);
and U19778 (N_19778,N_16594,N_15559);
or U19779 (N_19779,N_17349,N_18055);
or U19780 (N_19780,N_13660,N_16791);
nor U19781 (N_19781,N_12999,N_12864);
xnor U19782 (N_19782,N_15408,N_18108);
nand U19783 (N_19783,N_17727,N_15424);
nand U19784 (N_19784,N_15700,N_12817);
or U19785 (N_19785,N_16492,N_17789);
nand U19786 (N_19786,N_18479,N_16692);
nor U19787 (N_19787,N_16916,N_12845);
nor U19788 (N_19788,N_18153,N_14606);
and U19789 (N_19789,N_12618,N_15129);
nor U19790 (N_19790,N_16664,N_13986);
nor U19791 (N_19791,N_13190,N_13975);
nand U19792 (N_19792,N_15434,N_13450);
nand U19793 (N_19793,N_15666,N_18505);
nand U19794 (N_19794,N_12609,N_17120);
nand U19795 (N_19795,N_12842,N_13546);
xor U19796 (N_19796,N_17675,N_15325);
xnor U19797 (N_19797,N_17412,N_17298);
or U19798 (N_19798,N_12693,N_16495);
and U19799 (N_19799,N_13005,N_17346);
nor U19800 (N_19800,N_12525,N_14479);
and U19801 (N_19801,N_16514,N_16733);
nor U19802 (N_19802,N_14236,N_13661);
nor U19803 (N_19803,N_12996,N_13855);
or U19804 (N_19804,N_13573,N_18387);
or U19805 (N_19805,N_17159,N_13494);
and U19806 (N_19806,N_16095,N_13707);
and U19807 (N_19807,N_13227,N_14930);
nor U19808 (N_19808,N_18059,N_12856);
or U19809 (N_19809,N_13090,N_15873);
or U19810 (N_19810,N_12838,N_14631);
nand U19811 (N_19811,N_15194,N_16553);
nand U19812 (N_19812,N_17381,N_12637);
or U19813 (N_19813,N_17165,N_15315);
nand U19814 (N_19814,N_15359,N_12874);
nor U19815 (N_19815,N_18563,N_16237);
nand U19816 (N_19816,N_12639,N_16732);
xnor U19817 (N_19817,N_15986,N_12925);
nor U19818 (N_19818,N_12802,N_16427);
nand U19819 (N_19819,N_16883,N_18274);
nor U19820 (N_19820,N_15683,N_13813);
and U19821 (N_19821,N_16482,N_13111);
nor U19822 (N_19822,N_17223,N_12747);
and U19823 (N_19823,N_17202,N_18079);
nand U19824 (N_19824,N_15545,N_13319);
or U19825 (N_19825,N_13989,N_15587);
or U19826 (N_19826,N_16673,N_14598);
nand U19827 (N_19827,N_14246,N_13800);
nor U19828 (N_19828,N_12625,N_13938);
or U19829 (N_19829,N_13949,N_17013);
nor U19830 (N_19830,N_18148,N_14840);
nand U19831 (N_19831,N_18494,N_15167);
nand U19832 (N_19832,N_17430,N_14691);
or U19833 (N_19833,N_18099,N_14397);
xnor U19834 (N_19834,N_14822,N_16547);
or U19835 (N_19835,N_15081,N_14697);
xor U19836 (N_19836,N_15369,N_18530);
nand U19837 (N_19837,N_14427,N_18196);
nand U19838 (N_19838,N_13581,N_13252);
nor U19839 (N_19839,N_16644,N_14923);
nand U19840 (N_19840,N_14995,N_13066);
nand U19841 (N_19841,N_16242,N_16810);
or U19842 (N_19842,N_16219,N_15444);
nand U19843 (N_19843,N_13098,N_17054);
or U19844 (N_19844,N_17009,N_17516);
nor U19845 (N_19845,N_18524,N_13651);
nand U19846 (N_19846,N_17595,N_15716);
and U19847 (N_19847,N_15940,N_17096);
and U19848 (N_19848,N_14006,N_14369);
nand U19849 (N_19849,N_14583,N_14108);
or U19850 (N_19850,N_17547,N_17169);
nand U19851 (N_19851,N_16100,N_16533);
nor U19852 (N_19852,N_18122,N_17344);
and U19853 (N_19853,N_14965,N_17094);
nor U19854 (N_19854,N_14718,N_13870);
nand U19855 (N_19855,N_12991,N_17443);
and U19856 (N_19856,N_13514,N_12559);
nor U19857 (N_19857,N_16550,N_16680);
and U19858 (N_19858,N_14983,N_16024);
nor U19859 (N_19859,N_13857,N_15488);
nor U19860 (N_19860,N_18280,N_16164);
nor U19861 (N_19861,N_18601,N_15122);
nor U19862 (N_19862,N_17542,N_14241);
or U19863 (N_19863,N_12688,N_14316);
xnor U19864 (N_19864,N_16263,N_17753);
or U19865 (N_19865,N_12512,N_15790);
xnor U19866 (N_19866,N_18445,N_17092);
and U19867 (N_19867,N_15534,N_15437);
or U19868 (N_19868,N_18520,N_12854);
xnor U19869 (N_19869,N_14695,N_18340);
nand U19870 (N_19870,N_14698,N_18746);
or U19871 (N_19871,N_15074,N_16459);
nor U19872 (N_19872,N_14851,N_13590);
and U19873 (N_19873,N_16479,N_18170);
and U19874 (N_19874,N_17718,N_17820);
or U19875 (N_19875,N_15338,N_14769);
nor U19876 (N_19876,N_12554,N_17466);
xnor U19877 (N_19877,N_13024,N_13914);
nand U19878 (N_19878,N_17742,N_13191);
nand U19879 (N_19879,N_16669,N_17553);
nor U19880 (N_19880,N_14145,N_18740);
or U19881 (N_19881,N_13681,N_15206);
and U19882 (N_19882,N_15973,N_16129);
or U19883 (N_19883,N_14637,N_16542);
and U19884 (N_19884,N_14512,N_17249);
nor U19885 (N_19885,N_16827,N_15402);
nand U19886 (N_19886,N_14463,N_18329);
or U19887 (N_19887,N_15875,N_14420);
nand U19888 (N_19888,N_17802,N_18292);
nand U19889 (N_19889,N_18382,N_15602);
xor U19890 (N_19890,N_13427,N_15344);
nor U19891 (N_19891,N_17961,N_17320);
nor U19892 (N_19892,N_15926,N_14878);
and U19893 (N_19893,N_15355,N_18038);
nor U19894 (N_19894,N_16135,N_14772);
nand U19895 (N_19895,N_13931,N_16768);
and U19896 (N_19896,N_12617,N_17172);
or U19897 (N_19897,N_15855,N_18732);
and U19898 (N_19898,N_18725,N_18717);
and U19899 (N_19899,N_17084,N_18711);
or U19900 (N_19900,N_15622,N_14910);
or U19901 (N_19901,N_16049,N_14727);
and U19902 (N_19902,N_13865,N_15588);
nor U19903 (N_19903,N_14715,N_14318);
and U19904 (N_19904,N_13419,N_17997);
and U19905 (N_19905,N_17156,N_15685);
or U19906 (N_19906,N_18749,N_15987);
nor U19907 (N_19907,N_15491,N_16516);
xnor U19908 (N_19908,N_14821,N_15906);
xnor U19909 (N_19909,N_18114,N_15147);
or U19910 (N_19910,N_14830,N_13470);
nand U19911 (N_19911,N_16787,N_17141);
nor U19912 (N_19912,N_13633,N_13886);
nor U19913 (N_19913,N_16033,N_17596);
and U19914 (N_19914,N_12627,N_13370);
and U19915 (N_19915,N_12850,N_17128);
nor U19916 (N_19916,N_15404,N_13147);
and U19917 (N_19917,N_13013,N_15802);
or U19918 (N_19918,N_16764,N_15811);
nor U19919 (N_19919,N_16776,N_14998);
nand U19920 (N_19920,N_14703,N_16304);
nor U19921 (N_19921,N_16375,N_14717);
or U19922 (N_19922,N_15083,N_13571);
and U19923 (N_19923,N_16562,N_15455);
nand U19924 (N_19924,N_16518,N_15033);
or U19925 (N_19925,N_14380,N_16229);
nor U19926 (N_19926,N_13620,N_18043);
nor U19927 (N_19927,N_15605,N_12857);
or U19928 (N_19928,N_16111,N_15002);
or U19929 (N_19929,N_16870,N_16499);
nand U19930 (N_19930,N_15497,N_15882);
or U19931 (N_19931,N_13712,N_12954);
or U19932 (N_19932,N_14767,N_13456);
nand U19933 (N_19933,N_15117,N_16665);
nor U19934 (N_19934,N_15604,N_14274);
and U19935 (N_19935,N_18544,N_16526);
or U19936 (N_19936,N_15943,N_14230);
xor U19937 (N_19937,N_17500,N_16466);
nor U19938 (N_19938,N_15087,N_16996);
nand U19939 (N_19939,N_15247,N_13708);
or U19940 (N_19940,N_18434,N_18158);
xor U19941 (N_19941,N_15792,N_12894);
or U19942 (N_19942,N_12772,N_16259);
and U19943 (N_19943,N_16313,N_18042);
nand U19944 (N_19944,N_15941,N_16112);
and U19945 (N_19945,N_12773,N_12964);
nand U19946 (N_19946,N_15832,N_17826);
xor U19947 (N_19947,N_17579,N_17383);
or U19948 (N_19948,N_18460,N_12694);
nor U19949 (N_19949,N_14205,N_17409);
nor U19950 (N_19950,N_12702,N_12882);
nor U19951 (N_19951,N_17208,N_17016);
xor U19952 (N_19952,N_18247,N_16997);
and U19953 (N_19953,N_12728,N_17416);
xor U19954 (N_19954,N_15781,N_18546);
nand U19955 (N_19955,N_12552,N_14956);
and U19956 (N_19956,N_17168,N_17035);
or U19957 (N_19957,N_17883,N_14052);
nor U19958 (N_19958,N_12805,N_14199);
and U19959 (N_19959,N_17158,N_15594);
nor U19960 (N_19960,N_18335,N_14142);
xnor U19961 (N_19961,N_18192,N_15635);
and U19962 (N_19962,N_16486,N_13675);
and U19963 (N_19963,N_13203,N_15613);
nand U19964 (N_19964,N_13360,N_16757);
and U19965 (N_19965,N_16930,N_12707);
nor U19966 (N_19966,N_15181,N_17631);
and U19967 (N_19967,N_12911,N_15962);
and U19968 (N_19968,N_17382,N_13154);
or U19969 (N_19969,N_13176,N_17633);
and U19970 (N_19970,N_17621,N_15721);
nand U19971 (N_19971,N_17331,N_13715);
and U19972 (N_19972,N_17453,N_13913);
or U19973 (N_19973,N_15267,N_18195);
nand U19974 (N_19974,N_13508,N_16570);
nand U19975 (N_19975,N_14552,N_17920);
and U19976 (N_19976,N_13830,N_16244);
or U19977 (N_19977,N_14829,N_13381);
or U19978 (N_19978,N_13683,N_17356);
nand U19979 (N_19979,N_16536,N_14668);
nor U19980 (N_19980,N_15258,N_14194);
nand U19981 (N_19981,N_17316,N_14469);
or U19982 (N_19982,N_17178,N_13770);
and U19983 (N_19983,N_16157,N_16919);
nor U19984 (N_19984,N_17567,N_14396);
or U19985 (N_19985,N_16293,N_18027);
nand U19986 (N_19986,N_13261,N_15390);
nor U19987 (N_19987,N_12709,N_14418);
or U19988 (N_19988,N_13544,N_16978);
and U19989 (N_19989,N_17512,N_16060);
and U19990 (N_19990,N_17908,N_15755);
nor U19991 (N_19991,N_12550,N_13909);
nor U19992 (N_19992,N_15687,N_16917);
and U19993 (N_19993,N_18681,N_14224);
nor U19994 (N_19994,N_13263,N_14482);
nand U19995 (N_19995,N_13769,N_18089);
nor U19996 (N_19996,N_13492,N_18437);
nand U19997 (N_19997,N_15848,N_12884);
nand U19998 (N_19998,N_17769,N_16891);
and U19999 (N_19999,N_18481,N_13236);
nor U20000 (N_20000,N_12799,N_13940);
or U20001 (N_20001,N_13631,N_13610);
or U20002 (N_20002,N_13724,N_12784);
nand U20003 (N_20003,N_16892,N_12718);
or U20004 (N_20004,N_13783,N_17385);
or U20005 (N_20005,N_18643,N_14094);
nor U20006 (N_20006,N_18418,N_15221);
and U20007 (N_20007,N_15505,N_15052);
or U20008 (N_20008,N_14250,N_18393);
nand U20009 (N_20009,N_12981,N_18708);
nor U20010 (N_20010,N_14704,N_14391);
or U20011 (N_20011,N_13920,N_16895);
xnor U20012 (N_20012,N_16193,N_15759);
and U20013 (N_20013,N_12868,N_17321);
xnor U20014 (N_20014,N_17127,N_17099);
nand U20015 (N_20015,N_13138,N_18702);
nor U20016 (N_20016,N_14180,N_13709);
nor U20017 (N_20017,N_18637,N_17438);
nand U20018 (N_20018,N_16555,N_16378);
nor U20019 (N_20019,N_14811,N_15823);
xor U20020 (N_20020,N_12522,N_14193);
or U20021 (N_20021,N_18608,N_14752);
xnor U20022 (N_20022,N_17696,N_14856);
nor U20023 (N_20023,N_18627,N_15732);
nor U20024 (N_20024,N_18067,N_14731);
or U20025 (N_20025,N_15950,N_17187);
nand U20026 (N_20026,N_16192,N_16184);
nor U20027 (N_20027,N_18266,N_12717);
nand U20028 (N_20028,N_17781,N_16306);
and U20029 (N_20029,N_14884,N_18115);
or U20030 (N_20030,N_18184,N_18575);
and U20031 (N_20031,N_13251,N_18743);
and U20032 (N_20032,N_14005,N_13012);
and U20033 (N_20033,N_12716,N_13383);
or U20034 (N_20034,N_15954,N_14678);
and U20035 (N_20035,N_16702,N_13689);
and U20036 (N_20036,N_14442,N_16268);
and U20037 (N_20037,N_13761,N_18165);
and U20038 (N_20038,N_14586,N_13638);
nand U20039 (N_20039,N_14791,N_13454);
nor U20040 (N_20040,N_13269,N_16841);
and U20041 (N_20041,N_12619,N_16569);
nand U20042 (N_20042,N_16752,N_15726);
or U20043 (N_20043,N_14106,N_13096);
and U20044 (N_20044,N_13114,N_18021);
nand U20045 (N_20045,N_16284,N_14849);
and U20046 (N_20046,N_17755,N_14947);
nand U20047 (N_20047,N_17357,N_16721);
or U20048 (N_20048,N_16369,N_18515);
nand U20049 (N_20049,N_13448,N_14187);
xnor U20050 (N_20050,N_16352,N_18699);
or U20051 (N_20051,N_14920,N_15375);
nor U20052 (N_20052,N_18277,N_15925);
nand U20053 (N_20053,N_12766,N_18225);
and U20054 (N_20054,N_13363,N_16583);
nand U20055 (N_20055,N_15626,N_18535);
nor U20056 (N_20056,N_16388,N_15753);
nor U20057 (N_20057,N_18022,N_17448);
nor U20058 (N_20058,N_16241,N_17122);
nand U20059 (N_20059,N_13212,N_16214);
nor U20060 (N_20060,N_16179,N_17278);
or U20061 (N_20061,N_15405,N_15951);
nor U20062 (N_20062,N_17015,N_14078);
and U20063 (N_20063,N_12927,N_16254);
nand U20064 (N_20064,N_17632,N_17694);
and U20065 (N_20065,N_14217,N_17642);
xor U20066 (N_20066,N_13915,N_14858);
nor U20067 (N_20067,N_16322,N_18271);
and U20068 (N_20068,N_14327,N_17426);
or U20069 (N_20069,N_14954,N_17219);
or U20070 (N_20070,N_15512,N_17403);
or U20071 (N_20071,N_15740,N_13074);
nor U20072 (N_20072,N_16739,N_16316);
or U20073 (N_20073,N_16450,N_12945);
and U20074 (N_20074,N_16873,N_18160);
or U20075 (N_20075,N_13927,N_14269);
or U20076 (N_20076,N_18742,N_13554);
and U20077 (N_20077,N_14189,N_12915);
and U20078 (N_20078,N_13672,N_12955);
and U20079 (N_20079,N_13716,N_13152);
nand U20080 (N_20080,N_16754,N_18683);
or U20081 (N_20081,N_16154,N_13063);
nor U20082 (N_20082,N_16430,N_17571);
and U20083 (N_20083,N_17794,N_14123);
nor U20084 (N_20084,N_15419,N_12860);
or U20085 (N_20085,N_16059,N_13779);
nor U20086 (N_20086,N_18533,N_15431);
and U20087 (N_20087,N_14848,N_16760);
or U20088 (N_20088,N_17454,N_12765);
and U20089 (N_20089,N_17763,N_18450);
and U20090 (N_20090,N_14160,N_16278);
and U20091 (N_20091,N_14211,N_13567);
or U20092 (N_20092,N_17026,N_17932);
nor U20093 (N_20093,N_17248,N_15544);
and U20094 (N_20094,N_15817,N_16785);
or U20095 (N_20095,N_18394,N_13412);
xor U20096 (N_20096,N_18366,N_17420);
nor U20097 (N_20097,N_14906,N_16065);
nor U20098 (N_20098,N_18147,N_18504);
and U20099 (N_20099,N_18407,N_15077);
or U20100 (N_20100,N_15443,N_13676);
nor U20101 (N_20101,N_15233,N_15839);
nor U20102 (N_20102,N_17856,N_16824);
and U20103 (N_20103,N_17337,N_17586);
nor U20104 (N_20104,N_14857,N_18278);
nand U20105 (N_20105,N_13891,N_16600);
or U20106 (N_20106,N_13392,N_12781);
nand U20107 (N_20107,N_18656,N_12936);
nand U20108 (N_20108,N_13739,N_15837);
nand U20109 (N_20109,N_17055,N_13995);
nor U20110 (N_20110,N_12621,N_17175);
or U20111 (N_20111,N_16225,N_17285);
nor U20112 (N_20112,N_16230,N_12539);
or U20113 (N_20113,N_17010,N_13504);
nor U20114 (N_20114,N_14922,N_17330);
and U20115 (N_20115,N_12595,N_13518);
nand U20116 (N_20116,N_17884,N_12835);
or U20117 (N_20117,N_12847,N_18154);
or U20118 (N_20118,N_18261,N_17515);
or U20119 (N_20119,N_16367,N_13714);
nand U20120 (N_20120,N_14306,N_18704);
nand U20121 (N_20121,N_15162,N_17664);
nor U20122 (N_20122,N_18053,N_15136);
and U20123 (N_20123,N_14611,N_17900);
nor U20124 (N_20124,N_17915,N_15139);
and U20125 (N_20125,N_14254,N_15130);
or U20126 (N_20126,N_15510,N_16504);
and U20127 (N_20127,N_17999,N_16453);
nor U20128 (N_20128,N_12783,N_12931);
and U20129 (N_20129,N_13181,N_17681);
nand U20130 (N_20130,N_18044,N_16086);
xnor U20131 (N_20131,N_13678,N_12549);
and U20132 (N_20132,N_14621,N_16907);
or U20133 (N_20133,N_18307,N_17389);
or U20134 (N_20134,N_14945,N_13215);
or U20135 (N_20135,N_14618,N_17559);
nand U20136 (N_20136,N_14496,N_14242);
nor U20137 (N_20137,N_17018,N_18011);
nand U20138 (N_20138,N_13634,N_15577);
or U20139 (N_20139,N_15201,N_13231);
xnor U20140 (N_20140,N_14404,N_14602);
and U20141 (N_20141,N_13123,N_12828);
nor U20142 (N_20142,N_18000,N_14835);
nand U20143 (N_20143,N_15135,N_17465);
nand U20144 (N_20144,N_15689,N_18295);
xor U20145 (N_20145,N_12587,N_17765);
or U20146 (N_20146,N_17047,N_12594);
and U20147 (N_20147,N_15669,N_14385);
nor U20148 (N_20148,N_15597,N_15647);
nand U20149 (N_20149,N_17059,N_12811);
nand U20150 (N_20150,N_12681,N_16765);
nor U20151 (N_20151,N_17031,N_16294);
nand U20152 (N_20152,N_13622,N_16010);
and U20153 (N_20153,N_13856,N_16137);
nor U20154 (N_20154,N_14919,N_15260);
xor U20155 (N_20155,N_16888,N_15331);
nor U20156 (N_20156,N_13472,N_17450);
or U20157 (N_20157,N_17740,N_18629);
nor U20158 (N_20158,N_15539,N_13946);
or U20159 (N_20159,N_15867,N_18090);
or U20160 (N_20160,N_17036,N_13803);
and U20161 (N_20161,N_13953,N_17927);
xor U20162 (N_20162,N_14118,N_16035);
nand U20163 (N_20163,N_13981,N_13307);
nand U20164 (N_20164,N_16362,N_16114);
and U20165 (N_20165,N_18328,N_18288);
or U20166 (N_20166,N_12897,N_14723);
or U20167 (N_20167,N_15110,N_13311);
or U20168 (N_20168,N_13277,N_12994);
nor U20169 (N_20169,N_18322,N_17928);
nand U20170 (N_20170,N_12596,N_17030);
nor U20171 (N_20171,N_13962,N_13375);
nand U20172 (N_20172,N_15538,N_17040);
or U20173 (N_20173,N_15175,N_13469);
or U20174 (N_20174,N_18646,N_17709);
or U20175 (N_20175,N_16288,N_15089);
xnor U20176 (N_20176,N_18631,N_17560);
nand U20177 (N_20177,N_14411,N_18346);
and U20178 (N_20178,N_15904,N_13058);
nor U20179 (N_20179,N_13598,N_15093);
nand U20180 (N_20180,N_17462,N_13965);
nor U20181 (N_20181,N_17038,N_14651);
xor U20182 (N_20182,N_14428,N_18392);
nand U20183 (N_20183,N_18623,N_16939);
or U20184 (N_20184,N_17851,N_12668);
or U20185 (N_20185,N_17097,N_14419);
or U20186 (N_20186,N_17108,N_15153);
and U20187 (N_20187,N_17490,N_17149);
nand U20188 (N_20188,N_17650,N_17638);
nand U20189 (N_20189,N_13673,N_16624);
nand U20190 (N_20190,N_15836,N_12556);
or U20191 (N_20191,N_12652,N_16606);
or U20192 (N_20192,N_16954,N_15251);
nand U20193 (N_20193,N_15812,N_17549);
nor U20194 (N_20194,N_18096,N_15637);
nand U20195 (N_20195,N_17671,N_13457);
nor U20196 (N_20196,N_15911,N_17539);
nor U20197 (N_20197,N_14057,N_17804);
or U20198 (N_20198,N_18690,N_12601);
nor U20199 (N_20199,N_18431,N_17326);
nand U20200 (N_20200,N_15592,N_16267);
or U20201 (N_20201,N_17809,N_13974);
nor U20202 (N_20202,N_16098,N_14366);
nand U20203 (N_20203,N_12504,N_17976);
and U20204 (N_20204,N_13193,N_17348);
or U20205 (N_20205,N_15341,N_15566);
xnor U20206 (N_20206,N_18268,N_15532);
nand U20207 (N_20207,N_15595,N_15831);
and U20208 (N_20208,N_13224,N_15897);
and U20209 (N_20209,N_16148,N_15624);
nand U20210 (N_20210,N_13966,N_17558);
and U20211 (N_20211,N_16084,N_16943);
nand U20212 (N_20212,N_18181,N_15526);
nand U20213 (N_20213,N_14616,N_18483);
or U20214 (N_20214,N_16071,N_18293);
nand U20215 (N_20215,N_18424,N_18092);
or U20216 (N_20216,N_13543,N_15229);
or U20217 (N_20217,N_16882,N_17960);
nand U20218 (N_20218,N_15658,N_13539);
nor U20219 (N_20219,N_12792,N_14809);
or U20220 (N_20220,N_17252,N_14068);
or U20221 (N_20221,N_15396,N_13541);
and U20222 (N_20222,N_18185,N_15547);
and U20223 (N_20223,N_16005,N_16807);
nor U20224 (N_20224,N_12816,N_14730);
and U20225 (N_20225,N_16884,N_15847);
xnor U20226 (N_20226,N_17317,N_13797);
nand U20227 (N_20227,N_17719,N_17917);
nand U20228 (N_20228,N_15891,N_12785);
or U20229 (N_20229,N_13202,N_15616);
and U20230 (N_20230,N_18297,N_16650);
or U20231 (N_20231,N_17967,N_13713);
and U20232 (N_20232,N_14792,N_17232);
nand U20233 (N_20233,N_13723,N_17989);
nand U20234 (N_20234,N_16690,N_16116);
xnor U20235 (N_20235,N_15343,N_14148);
nor U20236 (N_20236,N_14165,N_16942);
and U20237 (N_20237,N_18560,N_16209);
xor U20238 (N_20238,N_15507,N_16972);
nor U20239 (N_20239,N_16938,N_13569);
nor U20240 (N_20240,N_16773,N_17828);
or U20241 (N_20241,N_17456,N_17114);
and U20242 (N_20242,N_12635,N_15333);
xor U20243 (N_20243,N_15079,N_16963);
nand U20244 (N_20244,N_13617,N_16194);
or U20245 (N_20245,N_17134,N_13542);
nor U20246 (N_20246,N_17750,N_17085);
nand U20247 (N_20247,N_15394,N_17493);
nor U20248 (N_20248,N_12623,N_16625);
nand U20249 (N_20249,N_17644,N_17477);
or U20250 (N_20250,N_13049,N_15853);
and U20251 (N_20251,N_13284,N_14022);
or U20252 (N_20252,N_16893,N_18026);
and U20253 (N_20253,N_13195,N_14276);
and U20254 (N_20254,N_14812,N_18086);
or U20255 (N_20255,N_14774,N_18405);
nor U20256 (N_20256,N_12538,N_16166);
xnor U20257 (N_20257,N_12555,N_15358);
nand U20258 (N_20258,N_13693,N_16456);
nor U20259 (N_20259,N_14880,N_18337);
nand U20260 (N_20260,N_12574,N_12651);
or U20261 (N_20261,N_13568,N_17300);
nand U20262 (N_20262,N_13535,N_15470);
nor U20263 (N_20263,N_15798,N_13054);
nand U20264 (N_20264,N_14850,N_16089);
nand U20265 (N_20265,N_13519,N_17124);
nand U20266 (N_20266,N_13198,N_13006);
xor U20267 (N_20267,N_13566,N_18171);
nor U20268 (N_20268,N_13304,N_17480);
or U20269 (N_20269,N_13130,N_15671);
nand U20270 (N_20270,N_14055,N_18639);
nand U20271 (N_20271,N_17039,N_14647);
and U20272 (N_20272,N_16001,N_12903);
nor U20273 (N_20273,N_18462,N_13475);
nand U20274 (N_20274,N_15725,N_15634);
xor U20275 (N_20275,N_13921,N_14018);
nor U20276 (N_20276,N_15239,N_17741);
or U20277 (N_20277,N_13847,N_18619);
and U20278 (N_20278,N_14019,N_18651);
xnor U20279 (N_20279,N_13471,N_15172);
nor U20280 (N_20280,N_18745,N_12727);
nor U20281 (N_20281,N_17823,N_14780);
and U20282 (N_20282,N_13516,N_17164);
xor U20283 (N_20283,N_15609,N_17006);
or U20284 (N_20284,N_18305,N_16975);
or U20285 (N_20285,N_16281,N_17246);
nand U20286 (N_20286,N_16435,N_13281);
and U20287 (N_20287,N_14928,N_14533);
nor U20288 (N_20288,N_17251,N_15719);
xor U20289 (N_20289,N_18215,N_13343);
and U20290 (N_20290,N_12511,N_16603);
nand U20291 (N_20291,N_13389,N_12771);
or U20292 (N_20292,N_15290,N_16370);
and U20293 (N_20293,N_18052,N_15425);
or U20294 (N_20294,N_13613,N_17171);
nor U20295 (N_20295,N_18113,N_12774);
nor U20296 (N_20296,N_17060,N_18352);
or U20297 (N_20297,N_17876,N_17405);
or U20298 (N_20298,N_14481,N_14559);
or U20299 (N_20299,N_13282,N_17227);
xnor U20300 (N_20300,N_13463,N_12700);
nand U20301 (N_20301,N_13196,N_14386);
nand U20302 (N_20302,N_15612,N_17479);
or U20303 (N_20303,N_12980,N_13549);
nand U20304 (N_20304,N_17342,N_14042);
nand U20305 (N_20305,N_15889,N_14868);
or U20306 (N_20306,N_13999,N_16273);
or U20307 (N_20307,N_18661,N_17952);
nor U20308 (N_20308,N_16800,N_16543);
and U20309 (N_20309,N_17140,N_15808);
xor U20310 (N_20310,N_18510,N_16476);
nor U20311 (N_20311,N_13894,N_13521);
or U20312 (N_20312,N_16391,N_18379);
or U20313 (N_20313,N_17768,N_13827);
nand U20314 (N_20314,N_13350,N_15188);
nand U20315 (N_20315,N_14804,N_17827);
and U20316 (N_20316,N_17066,N_18583);
nand U20317 (N_20317,N_16496,N_14436);
nand U20318 (N_20318,N_17678,N_16272);
and U20319 (N_20319,N_14047,N_17651);
or U20320 (N_20320,N_12934,N_12779);
xnor U20321 (N_20321,N_15311,N_15582);
or U20322 (N_20322,N_13887,N_17283);
nand U20323 (N_20323,N_17525,N_17860);
xnor U20324 (N_20324,N_17288,N_12572);
nand U20325 (N_20325,N_18652,N_13113);
xor U20326 (N_20326,N_15729,N_15469);
nand U20327 (N_20327,N_15441,N_15428);
nor U20328 (N_20328,N_14294,N_12733);
and U20329 (N_20329,N_15189,N_15807);
and U20330 (N_20330,N_18375,N_13735);
nor U20331 (N_20331,N_16282,N_13122);
nand U20332 (N_20332,N_15881,N_16210);
nand U20333 (N_20333,N_12914,N_17366);
xor U20334 (N_20334,N_16321,N_16265);
nor U20335 (N_20335,N_16620,N_15435);
nand U20336 (N_20336,N_17263,N_14572);
and U20337 (N_20337,N_15160,N_13684);
nand U20338 (N_20338,N_13933,N_18595);
nor U20339 (N_20339,N_15409,N_16927);
nor U20340 (N_20340,N_15971,N_17446);
or U20341 (N_20341,N_12517,N_18137);
and U20342 (N_20342,N_17074,N_13318);
nand U20343 (N_20343,N_17312,N_16510);
and U20344 (N_20344,N_15565,N_16906);
and U20345 (N_20345,N_17583,N_17739);
or U20346 (N_20346,N_16043,N_17408);
nand U20347 (N_20347,N_18336,N_14060);
and U20348 (N_20348,N_14986,N_18550);
nor U20349 (N_20349,N_15080,N_12908);
nand U20350 (N_20350,N_18296,N_14751);
and U20351 (N_20351,N_13414,N_14216);
nand U20352 (N_20352,N_15451,N_16804);
xor U20353 (N_20353,N_16743,N_16651);
nand U20354 (N_20354,N_18161,N_17445);
and U20355 (N_20355,N_16144,N_12706);
nand U20356 (N_20356,N_16618,N_14827);
and U20357 (N_20357,N_16803,N_18497);
xor U20358 (N_20358,N_14395,N_16403);
nor U20359 (N_20359,N_13910,N_15640);
or U20360 (N_20360,N_13784,N_13095);
nor U20361 (N_20361,N_13220,N_18287);
and U20362 (N_20362,N_14991,N_14645);
and U20363 (N_20363,N_15572,N_14279);
xor U20364 (N_20364,N_18242,N_16473);
nor U20365 (N_20365,N_15596,N_14407);
or U20366 (N_20366,N_12902,N_15574);
or U20367 (N_20367,N_16861,N_18490);
xor U20368 (N_20368,N_14413,N_14775);
or U20369 (N_20369,N_12528,N_15422);
nor U20370 (N_20370,N_16289,N_15866);
or U20371 (N_20371,N_15182,N_13586);
xor U20372 (N_20372,N_18063,N_16285);
and U20373 (N_20373,N_15963,N_13728);
nor U20374 (N_20374,N_12800,N_17265);
nor U20375 (N_20375,N_14044,N_15584);
nor U20376 (N_20376,N_18554,N_12664);
nor U20377 (N_20377,N_12642,N_14755);
and U20378 (N_20378,N_12971,N_17495);
nand U20379 (N_20379,N_12540,N_18548);
or U20380 (N_20380,N_17660,N_14895);
xnor U20381 (N_20381,N_17503,N_15016);
nand U20382 (N_20382,N_16941,N_15464);
nand U20383 (N_20383,N_16097,N_14747);
nor U20384 (N_20384,N_13737,N_17131);
nand U20385 (N_20385,N_16207,N_18014);
xnor U20386 (N_20386,N_16728,N_16579);
nor U20387 (N_20387,N_18118,N_16831);
nand U20388 (N_20388,N_15633,N_15288);
and U20389 (N_20389,N_17877,N_17729);
nor U20390 (N_20390,N_14894,N_17360);
and U20391 (N_20391,N_17966,N_15793);
or U20392 (N_20392,N_13015,N_15319);
nor U20393 (N_20393,N_18363,N_18737);
nor U20394 (N_20394,N_17710,N_13816);
nor U20395 (N_20395,N_16817,N_13603);
or U20396 (N_20396,N_12909,N_17481);
and U20397 (N_20397,N_15743,N_15195);
or U20398 (N_20398,N_12620,N_12801);
nor U20399 (N_20399,N_14564,N_16608);
nand U20400 (N_20400,N_18355,N_17478);
xor U20401 (N_20401,N_15636,N_13889);
and U20402 (N_20402,N_13265,N_18209);
or U20403 (N_20403,N_12543,N_15236);
or U20404 (N_20404,N_17161,N_16040);
nand U20405 (N_20405,N_12939,N_16480);
and U20406 (N_20406,N_16256,N_14676);
and U20407 (N_20407,N_18571,N_18104);
xor U20408 (N_20408,N_15791,N_16415);
nor U20409 (N_20409,N_14635,N_15173);
and U20410 (N_20410,N_16213,N_14244);
or U20411 (N_20411,N_15227,N_14605);
nor U20412 (N_20412,N_12667,N_16096);
nor U20413 (N_20413,N_17531,N_15332);
nand U20414 (N_20414,N_13078,N_18150);
or U20415 (N_20415,N_16338,N_12822);
nand U20416 (N_20416,N_16027,N_16120);
nor U20417 (N_20417,N_13205,N_12585);
and U20418 (N_20418,N_17581,N_18144);
and U20419 (N_20419,N_14033,N_13020);
nand U20420 (N_20420,N_13973,N_17470);
nand U20421 (N_20421,N_15084,N_16431);
and U20422 (N_20422,N_13174,N_12901);
and U20423 (N_20423,N_17861,N_15415);
xor U20424 (N_20424,N_15932,N_17923);
or U20425 (N_20425,N_14403,N_16697);
and U20426 (N_20426,N_16952,N_16731);
nor U20427 (N_20427,N_14483,N_13435);
and U20428 (N_20428,N_15278,N_14962);
xnor U20429 (N_20429,N_13686,N_16676);
or U20430 (N_20430,N_18180,N_17439);
and U20431 (N_20431,N_12535,N_18404);
or U20432 (N_20432,N_17969,N_18263);
and U20433 (N_20433,N_13511,N_15063);
nor U20434 (N_20434,N_15123,N_18139);
nor U20435 (N_20435,N_12751,N_15031);
or U20436 (N_20436,N_15154,N_17167);
and U20437 (N_20437,N_13300,N_15140);
and U20438 (N_20438,N_14558,N_16763);
nor U20439 (N_20439,N_13884,N_13812);
and U20440 (N_20440,N_18207,N_15085);
xnor U20441 (N_20441,N_14024,N_15518);
nor U20442 (N_20442,N_17404,N_14778);
xor U20443 (N_20443,N_16484,N_16404);
and U20444 (N_20444,N_16053,N_12769);
or U20445 (N_20445,N_16169,N_18232);
and U20446 (N_20446,N_16774,N_13882);
nand U20447 (N_20447,N_16182,N_17335);
nand U20448 (N_20448,N_15190,N_17830);
nor U20449 (N_20449,N_16126,N_15322);
nand U20450 (N_20450,N_13806,N_18620);
nand U20451 (N_20451,N_17374,N_17386);
nand U20452 (N_20452,N_15614,N_17610);
or U20453 (N_20453,N_16301,N_15298);
nand U20454 (N_20454,N_16696,N_18446);
and U20455 (N_20455,N_12542,N_12832);
and U20456 (N_20456,N_16730,N_13730);
nand U20457 (N_20457,N_13720,N_15711);
nor U20458 (N_20458,N_17576,N_13901);
and U20459 (N_20459,N_15898,N_15661);
or U20460 (N_20460,N_16528,N_15975);
and U20461 (N_20461,N_16965,N_14371);
nand U20462 (N_20462,N_12729,N_14478);
nand U20463 (N_20463,N_15704,N_15372);
nor U20464 (N_20464,N_16623,N_17112);
nor U20465 (N_20465,N_13614,N_12662);
or U20466 (N_20466,N_15410,N_17626);
xor U20467 (N_20467,N_14648,N_18684);
or U20468 (N_20468,N_13846,N_14345);
nand U20469 (N_20469,N_17730,N_14597);
and U20470 (N_20470,N_18156,N_15779);
and U20471 (N_20471,N_13351,N_13798);
nand U20472 (N_20472,N_12510,N_17972);
nand U20473 (N_20473,N_17113,N_13126);
and U20474 (N_20474,N_13158,N_14222);
xor U20475 (N_20475,N_18218,N_18448);
and U20476 (N_20476,N_17836,N_16712);
nand U20477 (N_20477,N_14531,N_15712);
xor U20478 (N_20478,N_15991,N_18455);
nor U20479 (N_20479,N_14500,N_13104);
xor U20480 (N_20480,N_14039,N_14131);
and U20481 (N_20481,N_16611,N_15714);
or U20482 (N_20482,N_13338,N_13837);
nand U20483 (N_20483,N_14887,N_14988);
or U20484 (N_20484,N_13355,N_15187);
nor U20485 (N_20485,N_13201,N_18617);
and U20486 (N_20486,N_15440,N_14431);
nand U20487 (N_20487,N_17693,N_15479);
nand U20488 (N_20488,N_14975,N_13876);
nand U20489 (N_20489,N_16050,N_16454);
nor U20490 (N_20490,N_16046,N_17672);
or U20491 (N_20491,N_13458,N_17752);
or U20492 (N_20492,N_12859,N_16471);
and U20493 (N_20493,N_17256,N_18302);
or U20494 (N_20494,N_13431,N_14758);
or U20495 (N_20495,N_16407,N_17561);
nand U20496 (N_20496,N_12803,N_17988);
nor U20497 (N_20497,N_16339,N_17235);
nor U20498 (N_20498,N_17170,N_16872);
nor U20499 (N_20499,N_14532,N_17791);
or U20500 (N_20500,N_17017,N_13094);
nor U20501 (N_20501,N_14506,N_14994);
nor U20502 (N_20502,N_16865,N_13922);
xor U20503 (N_20503,N_17958,N_15449);
or U20504 (N_20504,N_13079,N_18238);
nor U20505 (N_20505,N_13310,N_13433);
nor U20506 (N_20506,N_16196,N_15969);
xnor U20507 (N_20507,N_17924,N_14454);
xor U20508 (N_20508,N_14643,N_17712);
nand U20509 (N_20509,N_16738,N_18300);
nor U20510 (N_20510,N_14913,N_16505);
and U20511 (N_20511,N_17648,N_16180);
nand U20512 (N_20512,N_13547,N_15458);
and U20513 (N_20513,N_12899,N_17616);
and U20514 (N_20514,N_14036,N_14144);
or U20515 (N_20515,N_16987,N_17001);
nor U20516 (N_20516,N_14996,N_15483);
nand U20517 (N_20517,N_15460,N_18397);
nor U20518 (N_20518,N_18538,N_13313);
and U20519 (N_20519,N_16766,N_16455);
or U20520 (N_20520,N_13131,N_13016);
xnor U20521 (N_20521,N_13477,N_17703);
and U20522 (N_20522,N_13984,N_17605);
nor U20523 (N_20523,N_16251,N_16030);
and U20524 (N_20524,N_17355,N_15490);
or U20525 (N_20525,N_16105,N_17618);
nand U20526 (N_20526,N_13768,N_16000);
nor U20527 (N_20527,N_12930,N_13488);
or U20528 (N_20528,N_14661,N_14351);
nand U20529 (N_20529,N_13309,N_13293);
nor U20530 (N_20530,N_17166,N_14333);
and U20531 (N_20531,N_18019,N_14667);
nor U20532 (N_20532,N_15158,N_17123);
or U20533 (N_20533,N_17508,N_18368);
nor U20534 (N_20534,N_18598,N_14967);
or U20535 (N_20535,N_15778,N_13585);
and U20536 (N_20536,N_17432,N_18151);
or U20537 (N_20537,N_18005,N_14100);
nand U20538 (N_20538,N_13434,N_13133);
or U20539 (N_20539,N_16981,N_18361);
xnor U20540 (N_20540,N_14788,N_13108);
nor U20541 (N_20541,N_13086,N_18720);
and U20542 (N_20542,N_16588,N_16325);
nor U20543 (N_20543,N_13548,N_14646);
xor U20544 (N_20544,N_13109,N_16591);
and U20545 (N_20545,N_15501,N_18111);
nor U20546 (N_20546,N_12677,N_15102);
and U20547 (N_20547,N_15192,N_16198);
and U20548 (N_20548,N_17557,N_13609);
and U20549 (N_20549,N_14490,N_12541);
and U20550 (N_20550,N_15218,N_13750);
or U20551 (N_20551,N_15021,N_13417);
and U20552 (N_20552,N_17837,N_17797);
or U20553 (N_20553,N_17075,N_16885);
nand U20554 (N_20554,N_18360,N_16384);
nor U20555 (N_20555,N_14943,N_15693);
or U20556 (N_20556,N_14714,N_16195);
xnor U20557 (N_20557,N_18718,N_15652);
nand U20558 (N_20558,N_16335,N_13119);
nand U20559 (N_20559,N_17212,N_16232);
or U20560 (N_20560,N_14383,N_14713);
and U20561 (N_20561,N_18219,N_14789);
or U20562 (N_20562,N_13428,N_17277);
nand U20563 (N_20563,N_16645,N_13437);
xor U20564 (N_20564,N_16412,N_17046);
or U20565 (N_20565,N_17230,N_14324);
nand U20566 (N_20566,N_14171,N_16855);
or U20567 (N_20567,N_17540,N_14368);
and U20568 (N_20568,N_13216,N_16079);
and U20569 (N_20569,N_18433,N_14298);
or U20570 (N_20570,N_17925,N_13612);
or U20571 (N_20571,N_14653,N_15068);
nor U20572 (N_20572,N_18471,N_12757);
and U20573 (N_20573,N_13649,N_13849);
nand U20574 (N_20574,N_13951,N_13545);
nor U20575 (N_20575,N_13482,N_13668);
or U20576 (N_20576,N_12938,N_14816);
or U20577 (N_20577,N_17079,N_14443);
nor U20578 (N_20578,N_17519,N_14323);
nor U20579 (N_20579,N_18294,N_18470);
and U20580 (N_20580,N_16413,N_15835);
or U20581 (N_20581,N_16113,N_13007);
or U20582 (N_20582,N_16820,N_16056);
xnor U20583 (N_20583,N_16714,N_12963);
and U20584 (N_20584,N_15186,N_16206);
nor U20585 (N_20585,N_14799,N_18719);
and U20586 (N_20586,N_15259,N_18709);
nor U20587 (N_20587,N_15287,N_14873);
nor U20588 (N_20588,N_13328,N_17521);
and U20589 (N_20589,N_17556,N_16032);
and U20590 (N_20590,N_14432,N_12876);
nand U20591 (N_20591,N_18362,N_15524);
nand U20592 (N_20592,N_14970,N_16191);
and U20593 (N_20593,N_16619,N_12692);
or U20594 (N_20594,N_12759,N_13722);
nor U20595 (N_20595,N_13597,N_13538);
nor U20596 (N_20596,N_18444,N_17163);
or U20597 (N_20597,N_12758,N_16132);
or U20598 (N_20598,N_15773,N_14517);
nand U20599 (N_20599,N_13654,N_17145);
or U20600 (N_20600,N_12870,N_16679);
and U20601 (N_20601,N_14521,N_17126);
nor U20602 (N_20602,N_18633,N_17572);
nor U20603 (N_20603,N_14585,N_14982);
and U20604 (N_20604,N_16847,N_15412);
nand U20605 (N_20605,N_16311,N_16314);
nor U20606 (N_20606,N_15553,N_14220);
nor U20607 (N_20607,N_14619,N_14696);
and U20608 (N_20608,N_17748,N_14514);
and U20609 (N_20609,N_18254,N_14504);
and U20610 (N_20610,N_18032,N_16613);
nor U20611 (N_20611,N_15803,N_16782);
nand U20612 (N_20612,N_14626,N_16276);
or U20613 (N_20613,N_17308,N_16481);
xor U20614 (N_20614,N_16715,N_13685);
nand U20615 (N_20615,N_16953,N_17179);
and U20616 (N_20616,N_17520,N_15348);
xor U20617 (N_20617,N_17893,N_18109);
or U20618 (N_20618,N_15929,N_15486);
and U20619 (N_20619,N_15020,N_16936);
xnor U20620 (N_20620,N_14001,N_14795);
xor U20621 (N_20621,N_12761,N_15263);
nor U20622 (N_20622,N_12851,N_18721);
or U20623 (N_20623,N_16397,N_16971);
or U20624 (N_20624,N_14457,N_15060);
nand U20625 (N_20625,N_18436,N_16349);
and U20626 (N_20626,N_14640,N_16467);
and U20627 (N_20627,N_16006,N_16964);
nand U20628 (N_20628,N_13823,N_12972);
and U20629 (N_20629,N_16576,N_13818);
or U20630 (N_20630,N_16493,N_17111);
xnor U20631 (N_20631,N_17934,N_13143);
nand U20632 (N_20632,N_17475,N_18049);
xor U20633 (N_20633,N_15615,N_12570);
nand U20634 (N_20634,N_16564,N_12982);
or U20635 (N_20635,N_16512,N_15558);
nor U20636 (N_20636,N_13853,N_14243);
and U20637 (N_20637,N_15353,N_18301);
or U20638 (N_20638,N_13478,N_14893);
or U20639 (N_20639,N_13232,N_16228);
nand U20640 (N_20640,N_17511,N_13881);
or U20641 (N_20641,N_14096,N_17033);
and U20642 (N_20642,N_13084,N_18344);
nor U20643 (N_20643,N_12647,N_18428);
or U20644 (N_20644,N_16320,N_14099);
or U20645 (N_20645,N_14656,N_16009);
or U20646 (N_20646,N_13904,N_17629);
and U20647 (N_20647,N_16816,N_15996);
and U20648 (N_20648,N_14488,N_14518);
or U20649 (N_20649,N_18012,N_13091);
or U20650 (N_20650,N_13315,N_15143);
and U20651 (N_20651,N_16134,N_14997);
and U20652 (N_20652,N_17095,N_15092);
and U20653 (N_20653,N_15057,N_17240);
nand U20654 (N_20654,N_15736,N_14311);
or U20655 (N_20655,N_18537,N_15448);
nand U20656 (N_20656,N_13418,N_12820);
and U20657 (N_20657,N_18634,N_15180);
nand U20658 (N_20658,N_16534,N_16986);
nor U20659 (N_20659,N_17061,N_15324);
and U20660 (N_20660,N_15373,N_16596);
nand U20661 (N_20661,N_15787,N_14257);
xor U20662 (N_20662,N_18234,N_16418);
nor U20663 (N_20663,N_13551,N_17144);
nand U20664 (N_20664,N_17906,N_17309);
nand U20665 (N_20665,N_15826,N_15196);
and U20666 (N_20666,N_14670,N_16868);
nand U20667 (N_20667,N_13879,N_16638);
and U20668 (N_20668,N_13928,N_15733);
or U20669 (N_20669,N_13399,N_12951);
nor U20670 (N_20670,N_14722,N_18688);
or U20671 (N_20671,N_17188,N_17818);
nor U20672 (N_20672,N_13657,N_18568);
nand U20673 (N_20673,N_15038,N_18186);
nor U20674 (N_20674,N_14523,N_16877);
and U20675 (N_20675,N_18095,N_14680);
nand U20676 (N_20676,N_18239,N_16258);
nand U20677 (N_20677,N_17545,N_18516);
and U20678 (N_20678,N_14184,N_13105);
nor U20679 (N_20679,N_18602,N_18519);
nor U20680 (N_20680,N_12984,N_18574);
or U20681 (N_20681,N_17995,N_16441);
and U20682 (N_20682,N_15947,N_14186);
nand U20683 (N_20683,N_16417,N_16257);
nand U20684 (N_20684,N_14212,N_16869);
nand U20685 (N_20685,N_13141,N_17305);
or U20686 (N_20686,N_14733,N_15990);
and U20687 (N_20687,N_17129,N_17702);
and U20688 (N_20688,N_15414,N_18357);
xor U20689 (N_20689,N_12724,N_17183);
or U20690 (N_20690,N_18532,N_14085);
or U20691 (N_20691,N_14507,N_14210);
xor U20692 (N_20692,N_13036,N_13429);
xor U20693 (N_20693,N_16260,N_16602);
nor U20694 (N_20694,N_13439,N_12957);
or U20695 (N_20695,N_17087,N_14073);
nand U20696 (N_20696,N_17105,N_12524);
and U20697 (N_20697,N_17546,N_14949);
nand U20698 (N_20698,N_14724,N_16163);
nand U20699 (N_20699,N_18459,N_16351);
xnor U20700 (N_20700,N_14860,N_13774);
or U20701 (N_20701,N_17835,N_17229);
nand U20702 (N_20702,N_12920,N_17930);
nand U20703 (N_20703,N_15930,N_14317);
and U20704 (N_20704,N_12794,N_17101);
and U20705 (N_20705,N_18376,N_12628);
and U20706 (N_20706,N_15899,N_13286);
nor U20707 (N_20707,N_17117,N_15920);
xnor U20708 (N_20708,N_12598,N_17238);
nor U20709 (N_20709,N_14824,N_12924);
nor U20710 (N_20710,N_14357,N_14796);
nor U20711 (N_20711,N_13652,N_12948);
or U20712 (N_20712,N_12831,N_12848);
nand U20713 (N_20713,N_17023,N_13892);
and U20714 (N_20714,N_16150,N_16042);
or U20715 (N_20715,N_13577,N_14255);
and U20716 (N_20716,N_17885,N_16147);
nor U20717 (N_20717,N_14388,N_13118);
nor U20718 (N_20718,N_18327,N_14642);
nor U20719 (N_20719,N_15302,N_15506);
nand U20720 (N_20720,N_15015,N_12611);
or U20721 (N_20721,N_16854,N_13593);
and U20722 (N_20722,N_16755,N_12780);
nand U20723 (N_20723,N_18648,N_12846);
or U20724 (N_20724,N_13698,N_15957);
or U20725 (N_20725,N_13778,N_18507);
xnor U20726 (N_20726,N_18640,N_17505);
and U20727 (N_20727,N_17185,N_14213);
or U20728 (N_20728,N_13863,N_17222);
and U20729 (N_20729,N_15270,N_15075);
or U20730 (N_20730,N_15907,N_15638);
xnor U20731 (N_20731,N_16742,N_17499);
or U20732 (N_20732,N_15301,N_13142);
nand U20733 (N_20733,N_16279,N_17088);
nand U20734 (N_20734,N_12675,N_14308);
xnor U20735 (N_20735,N_14076,N_12650);
or U20736 (N_20736,N_14197,N_13396);
nor U20737 (N_20737,N_12744,N_17962);
and U20738 (N_20738,N_13677,N_15918);
nor U20739 (N_20739,N_16379,N_18270);
and U20740 (N_20740,N_14387,N_14336);
or U20741 (N_20741,N_17786,N_12960);
or U20742 (N_20742,N_18668,N_14007);
nand U20743 (N_20743,N_16771,N_14785);
and U20744 (N_20744,N_16183,N_12519);
nand U20745 (N_20745,N_18495,N_17294);
nor U20746 (N_20746,N_16736,N_15958);
nor U20747 (N_20747,N_14805,N_14537);
and U20748 (N_20748,N_14441,N_15166);
nor U20749 (N_20749,N_18354,N_17254);
nand U20750 (N_20750,N_18388,N_15450);
nand U20751 (N_20751,N_15050,N_14550);
nand U20752 (N_20752,N_17151,N_16118);
nor U20753 (N_20753,N_12608,N_16871);
or U20754 (N_20754,N_16657,N_13990);
or U20755 (N_20755,N_16947,N_14674);
or U20756 (N_20756,N_17067,N_17459);
and U20757 (N_20757,N_13627,N_17460);
nand U20758 (N_20758,N_17333,N_14793);
or U20759 (N_20759,N_18675,N_17463);
nor U20760 (N_20760,N_15292,N_13038);
nand U20761 (N_20761,N_15900,N_18622);
and U20762 (N_20762,N_13339,N_14472);
or U20763 (N_20763,N_14941,N_15600);
or U20764 (N_20764,N_15382,N_16291);
or U20765 (N_20765,N_13068,N_17077);
or U20766 (N_20766,N_13461,N_13859);
or U20767 (N_20767,N_15477,N_12643);
and U20768 (N_20768,N_15048,N_13391);
nand U20769 (N_20769,N_15321,N_15769);
or U20770 (N_20770,N_17831,N_18072);
nor U20771 (N_20771,N_15966,N_15243);
nor U20772 (N_20772,N_15090,N_16424);
nor U20773 (N_20773,N_14017,N_17655);
and U20774 (N_20774,N_15521,N_14726);
nor U20775 (N_20775,N_12507,N_16678);
or U20776 (N_20776,N_17343,N_13819);
xor U20777 (N_20777,N_14196,N_13137);
nand U20778 (N_20778,N_13809,N_12696);
nand U20779 (N_20779,N_14782,N_18167);
xnor U20780 (N_20780,N_13912,N_17485);
xor U20781 (N_20781,N_17509,N_13398);
nor U20782 (N_20782,N_12760,N_13880);
and U20783 (N_20783,N_18240,N_14660);
xor U20784 (N_20784,N_12969,N_14010);
nand U20785 (N_20785,N_13828,N_17522);
and U20786 (N_20786,N_16593,N_15780);
xor U20787 (N_20787,N_18543,N_12740);
xnor U20788 (N_20788,N_16994,N_13048);
and U20789 (N_20789,N_15764,N_13752);
and U20790 (N_20790,N_17625,N_17153);
nor U20791 (N_20791,N_13696,N_15484);
or U20792 (N_20792,N_13505,N_15418);
and U20793 (N_20793,N_18342,N_13523);
or U20794 (N_20794,N_16750,N_14030);
nor U20795 (N_20795,N_14610,N_12888);
nand U20796 (N_20796,N_16142,N_15694);
nor U20797 (N_20797,N_13089,N_14765);
nor U20798 (N_20798,N_18624,N_14331);
and U20799 (N_20799,N_16074,N_15691);
and U20800 (N_20800,N_18330,N_17339);
nand U20801 (N_20801,N_15939,N_15833);
nand U20802 (N_20802,N_18733,N_14162);
or U20803 (N_20803,N_14458,N_17279);
nand U20804 (N_20804,N_17833,N_12983);
and U20805 (N_20805,N_17301,N_13899);
nor U20806 (N_20806,N_14409,N_15207);
nor U20807 (N_20807,N_13358,N_13264);
nor U20808 (N_20808,N_17295,N_13719);
and U20809 (N_20809,N_13600,N_17533);
and U20810 (N_20810,N_17073,N_18365);
or U20811 (N_20811,N_16522,N_18203);
or U20812 (N_20812,N_17554,N_18256);
and U20813 (N_20813,N_17203,N_17406);
xor U20814 (N_20814,N_15742,N_13559);
or U20815 (N_20815,N_15516,N_13947);
nand U20816 (N_20816,N_14445,N_14314);
and U20817 (N_20817,N_18472,N_14918);
nand U20818 (N_20818,N_17896,N_14285);
xnor U20819 (N_20819,N_14908,N_16990);
nand U20820 (N_20820,N_15953,N_16315);
xor U20821 (N_20821,N_17825,N_14075);
xor U20822 (N_20822,N_16416,N_12575);
or U20823 (N_20823,N_18267,N_14925);
xor U20824 (N_20824,N_17674,N_15496);
nand U20825 (N_20825,N_17738,N_15137);
or U20826 (N_20826,N_17873,N_13242);
nand U20827 (N_20827,N_13868,N_14707);
nor U20828 (N_20828,N_16121,N_16788);
nor U20829 (N_20829,N_17076,N_14425);
or U20830 (N_20830,N_17614,N_14652);
and U20831 (N_20831,N_13459,N_18593);
or U20832 (N_20832,N_16979,N_12713);
nor U20833 (N_20833,N_17707,N_16707);
and U20834 (N_20834,N_16155,N_13209);
nand U20835 (N_20835,N_16929,N_12849);
xnor U20836 (N_20836,N_16970,N_13890);
and U20837 (N_20837,N_12883,N_12557);
or U20838 (N_20838,N_14613,N_13555);
or U20839 (N_20839,N_17012,N_13726);
or U20840 (N_20840,N_15011,N_16737);
and U20841 (N_20841,N_15675,N_14240);
or U20842 (N_20842,N_17991,N_13550);
xor U20843 (N_20843,N_14107,N_16333);
and U20844 (N_20844,N_15543,N_13772);
and U20845 (N_20845,N_13163,N_17983);
nand U20846 (N_20846,N_14167,N_14577);
nand U20847 (N_20847,N_14340,N_16500);
nor U20848 (N_20848,N_14980,N_17996);
xor U20849 (N_20849,N_14571,N_17778);
and U20850 (N_20850,N_17000,N_12577);
or U20851 (N_20851,N_17365,N_18531);
and U20852 (N_20852,N_16509,N_16461);
nor U20853 (N_20853,N_16460,N_13690);
or U20854 (N_20854,N_18729,N_13741);
nand U20855 (N_20855,N_15115,N_17770);
and U20856 (N_20856,N_14624,N_17289);
nand U20857 (N_20857,N_14522,N_16156);
or U20858 (N_20858,N_18308,N_14456);
or U20859 (N_20859,N_15148,N_16318);
nor U20860 (N_20860,N_18369,N_17776);
or U20861 (N_20861,N_13917,N_15297);
nand U20862 (N_20862,N_17798,N_14689);
or U20863 (N_20863,N_17081,N_17853);
xor U20864 (N_20864,N_18142,N_14951);
nand U20865 (N_20865,N_14711,N_14771);
nor U20866 (N_20866,N_16468,N_17424);
xnor U20867 (N_20867,N_17573,N_14140);
or U20868 (N_20868,N_17216,N_16879);
and U20869 (N_20869,N_13700,N_14176);
or U20870 (N_20870,N_14014,N_12841);
and U20871 (N_20871,N_16889,N_16729);
nor U20872 (N_20872,N_18372,N_15902);
or U20873 (N_20873,N_14389,N_15879);
or U20874 (N_20874,N_15580,N_15944);
nand U20875 (N_20875,N_15887,N_16777);
or U20876 (N_20876,N_12646,N_13180);
nor U20877 (N_20877,N_14629,N_15481);
nand U20878 (N_20878,N_14215,N_13840);
and U20879 (N_20879,N_17761,N_17514);
or U20880 (N_20880,N_18065,N_14474);
and U20881 (N_20881,N_14953,N_16360);
and U20882 (N_20882,N_15752,N_15364);
xnor U20883 (N_20883,N_14177,N_12821);
xnor U20884 (N_20884,N_17043,N_14839);
or U20885 (N_20885,N_17998,N_16477);
xor U20886 (N_20886,N_16541,N_15370);
nor U20887 (N_20887,N_18389,N_17486);
nor U20888 (N_20888,N_17956,N_13099);
nor U20889 (N_20889,N_18463,N_14544);
or U20890 (N_20890,N_12589,N_15291);
xnor U20891 (N_20891,N_14926,N_13296);
nand U20892 (N_20892,N_13167,N_16330);
nor U20893 (N_20893,N_15377,N_17819);
nor U20894 (N_20894,N_13815,N_15519);
nor U20895 (N_20895,N_16494,N_13753);
nor U20896 (N_20896,N_18665,N_18534);
or U20897 (N_20897,N_18657,N_15264);
xor U20898 (N_20898,N_15910,N_15184);
nor U20899 (N_20899,N_16329,N_14000);
or U20900 (N_20900,N_14510,N_15051);
nand U20901 (N_20901,N_18432,N_15241);
or U20902 (N_20902,N_14620,N_15678);
nor U20903 (N_20903,N_13280,N_13587);
nor U20904 (N_20904,N_15199,N_14009);
nor U20905 (N_20905,N_12565,N_15289);
xor U20906 (N_20906,N_16080,N_16047);
or U20907 (N_20907,N_15542,N_16078);
nor U20908 (N_20908,N_14338,N_16019);
nor U20909 (N_20909,N_15362,N_16846);
nor U20910 (N_20910,N_13092,N_18033);
and U20911 (N_20911,N_14252,N_15872);
xor U20912 (N_20912,N_17291,N_17652);
and U20913 (N_20913,N_14143,N_14466);
or U20914 (N_20914,N_15215,N_13757);
or U20915 (N_20915,N_15997,N_14002);
xnor U20916 (N_20916,N_18333,N_17535);
or U20917 (N_20917,N_14459,N_13858);
nand U20918 (N_20918,N_13691,N_12749);
nand U20919 (N_20919,N_17421,N_16452);
nand U20920 (N_20920,N_14576,N_16769);
nor U20921 (N_20921,N_15851,N_14543);
nand U20922 (N_20922,N_15995,N_15346);
xor U20923 (N_20923,N_16663,N_17887);
and U20924 (N_20924,N_17534,N_12907);
and U20925 (N_20925,N_17659,N_14377);
or U20926 (N_20926,N_13907,N_15004);
or U20927 (N_20927,N_17215,N_16353);
nor U20928 (N_20928,N_16802,N_15862);
nor U20929 (N_20929,N_17392,N_14738);
nand U20930 (N_20930,N_17751,N_15145);
nor U20931 (N_20931,N_18451,N_13056);
nor U20932 (N_20932,N_17799,N_13643);
or U20933 (N_20933,N_13875,N_16146);
and U20934 (N_20934,N_14295,N_13438);
and U20935 (N_20935,N_15621,N_13873);
or U20936 (N_20936,N_17275,N_16217);
and U20937 (N_20937,N_16586,N_15919);
nand U20938 (N_20938,N_13932,N_14125);
xor U20939 (N_20939,N_13443,N_13945);
xnor U20940 (N_20940,N_15563,N_17354);
nand U20941 (N_20941,N_13083,N_16389);
nand U20942 (N_20942,N_14495,N_14460);
nand U20943 (N_20943,N_15631,N_17931);
or U20944 (N_20944,N_16860,N_16511);
nor U20945 (N_20945,N_17020,N_13745);
xor U20946 (N_20946,N_12714,N_17911);
nor U20947 (N_20947,N_16372,N_15399);
nand U20948 (N_20948,N_16786,N_13895);
nand U20949 (N_20949,N_13165,N_16901);
nor U20950 (N_20950,N_14641,N_16850);
or U20951 (N_20951,N_13218,N_14365);
and U20952 (N_20952,N_15643,N_18047);
or U20953 (N_20953,N_17864,N_18678);
or U20954 (N_20954,N_13839,N_18010);
nor U20955 (N_20955,N_18182,N_16898);
nand U20956 (N_20956,N_13850,N_12861);
or U20957 (N_20957,N_13588,N_14786);
or U20958 (N_20958,N_17987,N_13266);
or U20959 (N_20959,N_18395,N_14623);
nand U20960 (N_20960,N_14508,N_13808);
nor U20961 (N_20961,N_18216,N_18373);
or U20962 (N_20962,N_16992,N_14608);
xnor U20963 (N_20963,N_14253,N_16261);
or U20964 (N_20964,N_18712,N_15043);
xor U20965 (N_20965,N_17774,N_17359);
or U20966 (N_20966,N_17068,N_17397);
nand U20967 (N_20967,N_17843,N_12887);
nor U20968 (N_20968,N_14092,N_18284);
nand U20969 (N_20969,N_14529,N_15003);
and U20970 (N_20970,N_17929,N_12789);
nor U20971 (N_20971,N_16324,N_13536);
xor U20972 (N_20972,N_16758,N_16490);
and U20973 (N_20973,N_17473,N_14029);
nand U20974 (N_20974,N_12680,N_15946);
and U20975 (N_20975,N_16414,N_14461);
and U20976 (N_20976,N_15047,N_16125);
and U20977 (N_20977,N_12829,N_16566);
nand U20978 (N_20978,N_16127,N_14079);
and U20979 (N_20979,N_13935,N_13271);
nand U20980 (N_20980,N_13275,N_17953);
nand U20981 (N_20981,N_15226,N_16614);
and U20982 (N_20982,N_15535,N_14299);
nand U20983 (N_20983,N_14141,N_13615);
and U20984 (N_20984,N_14341,N_12580);
or U20985 (N_20985,N_14113,N_15727);
nand U20986 (N_20986,N_16437,N_17528);
and U20987 (N_20987,N_14228,N_12858);
and U20988 (N_20988,N_18119,N_15217);
nor U20989 (N_20989,N_16234,N_17850);
or U20990 (N_20990,N_13321,N_15630);
or U20991 (N_20991,N_15098,N_14139);
and U20992 (N_20992,N_13289,N_15086);
or U20993 (N_20993,N_17943,N_17691);
and U20994 (N_20994,N_14121,N_14198);
and U20995 (N_20995,N_17756,N_14209);
or U20996 (N_20996,N_16852,N_15335);
or U20997 (N_20997,N_16240,N_17947);
nor U20998 (N_20998,N_14181,N_15282);
nor U20999 (N_20999,N_17434,N_15607);
and U21000 (N_21000,N_13982,N_13179);
nor U21001 (N_21001,N_18028,N_18723);
nand U21002 (N_21002,N_17506,N_16815);
nand U21003 (N_21003,N_15692,N_12593);
xor U21004 (N_21004,N_18500,N_15858);
or U21005 (N_21005,N_18260,N_12753);
nor U21006 (N_21006,N_16711,N_15610);
nor U21007 (N_21007,N_18466,N_18262);
and U21008 (N_21008,N_16123,N_12990);
or U21009 (N_21009,N_15212,N_18747);
or U21010 (N_21010,N_13852,N_17239);
and U21011 (N_21011,N_15810,N_13674);
xnor U21012 (N_21012,N_18614,N_17913);
nand U21013 (N_21013,N_12526,N_13509);
and U21014 (N_21014,N_17990,N_15744);
xor U21015 (N_21015,N_16283,N_18309);
and U21016 (N_21016,N_12562,N_12602);
nand U21017 (N_21017,N_15114,N_13701);
and U21018 (N_21018,N_18041,N_14178);
nand U21019 (N_21019,N_15830,N_13725);
nand U21020 (N_21020,N_13444,N_17189);
or U21021 (N_21021,N_15869,N_14059);
nand U21022 (N_21022,N_17606,N_13234);
or U21023 (N_21023,N_17086,N_13380);
or U21024 (N_21024,N_16354,N_14820);
and U21025 (N_21025,N_13864,N_17692);
or U21026 (N_21026,N_17100,N_16392);
and U21027 (N_21027,N_12529,N_18599);
or U21028 (N_21028,N_15082,N_16948);
nand U21029 (N_21029,N_17713,N_15655);
nand U21030 (N_21030,N_16844,N_12998);
xor U21031 (N_21031,N_15825,N_14557);
and U21032 (N_21032,N_13663,N_16160);
nor U21033 (N_21033,N_15988,N_13697);
xnor U21034 (N_21034,N_17870,N_15536);
or U21035 (N_21035,N_15067,N_18735);
nor U21036 (N_21036,N_17152,N_17669);
and U21037 (N_21037,N_15557,N_17926);
nand U21038 (N_21038,N_12711,N_12768);
nor U21039 (N_21039,N_17324,N_14169);
nor U21040 (N_21040,N_13502,N_17190);
nor U21041 (N_21041,N_13985,N_13255);
nand U21042 (N_21042,N_16433,N_15303);
or U21043 (N_21043,N_17492,N_18125);
nor U21044 (N_21044,N_14300,N_12770);
nand U21045 (N_21045,N_17570,N_13182);
nor U21046 (N_21046,N_17103,N_17116);
xnor U21047 (N_21047,N_15564,N_17373);
nor U21048 (N_21048,N_16751,N_16498);
nor U21049 (N_21049,N_15225,N_15456);
or U21050 (N_21050,N_14447,N_18057);
nand U21051 (N_21051,N_14911,N_12682);
nor U21052 (N_21052,N_12879,N_15035);
or U21053 (N_21053,N_13102,N_14748);
and U21054 (N_21054,N_13831,N_16016);
and U21055 (N_21055,N_15417,N_16797);
and U21056 (N_21056,N_17630,N_13785);
and U21057 (N_21057,N_15132,N_18194);
and U21058 (N_21058,N_14455,N_17685);
or U21059 (N_21059,N_13759,N_17728);
or U21060 (N_21060,N_15611,N_13493);
xnor U21061 (N_21061,N_15149,N_14412);
nand U21062 (N_21062,N_17375,N_12613);
or U21063 (N_21063,N_14511,N_17617);
or U21064 (N_21064,N_14916,N_16037);
xnor U21065 (N_21065,N_16175,N_17241);
and U21066 (N_21066,N_17233,N_14516);
nand U21067 (N_21067,N_13558,N_14638);
or U21068 (N_21068,N_17458,N_12877);
and U21069 (N_21069,N_17425,N_18686);
xnor U21070 (N_21070,N_17587,N_13189);
or U21071 (N_21071,N_16641,N_15026);
and U21072 (N_21072,N_18349,N_14347);
nor U21073 (N_21073,N_12673,N_16587);
nand U21074 (N_21074,N_13664,N_15351);
or U21075 (N_21075,N_13245,N_12798);
nand U21076 (N_21076,N_18691,N_12588);
or U21077 (N_21077,N_14494,N_15509);
or U21078 (N_21078,N_14797,N_15815);
or U21079 (N_21079,N_15046,N_17293);
and U21080 (N_21080,N_16029,N_16359);
and U21081 (N_21081,N_13885,N_14539);
or U21082 (N_21082,N_16792,N_12826);
nand U21083 (N_21083,N_15978,N_12683);
or U21084 (N_21084,N_13532,N_16002);
or U21085 (N_21085,N_15127,N_18116);
nor U21086 (N_21086,N_14917,N_15360);
and U21087 (N_21087,N_15627,N_13898);
nand U21088 (N_21088,N_15097,N_18731);
or U21089 (N_21089,N_16686,N_14600);
xor U21090 (N_21090,N_12551,N_17849);
and U21091 (N_21091,N_12545,N_13805);
nand U21092 (N_21092,N_12997,N_13368);
or U21093 (N_21093,N_15654,N_18269);
and U21094 (N_21094,N_18442,N_13583);
and U21095 (N_21095,N_15662,N_17890);
nand U21096 (N_21096,N_15895,N_16051);
nor U21097 (N_21097,N_14764,N_13248);
and U21098 (N_21098,N_14080,N_13366);
nor U21099 (N_21099,N_15921,N_14179);
or U21100 (N_21100,N_13353,N_17882);
nor U21101 (N_21101,N_15249,N_13402);
nand U21102 (N_21102,N_14687,N_15979);
and U21103 (N_21103,N_14869,N_17041);
nor U21104 (N_21104,N_16935,N_18211);
nand U21105 (N_21105,N_18511,N_13665);
nor U21106 (N_21106,N_13923,N_13067);
nand U21107 (N_21107,N_13556,N_17003);
xor U21108 (N_21108,N_17574,N_13795);
xor U21109 (N_21109,N_18159,N_18080);
nand U21110 (N_21110,N_17942,N_13963);
xor U21111 (N_21111,N_13004,N_14883);
and U21112 (N_21112,N_17400,N_13871);
and U21113 (N_21113,N_16734,N_12508);
or U21114 (N_21114,N_15931,N_15279);
nor U21115 (N_21115,N_13424,N_15001);
nor U21116 (N_21116,N_18070,N_13072);
xnor U21117 (N_21117,N_13297,N_16967);
or U21118 (N_21118,N_15400,N_16896);
or U21119 (N_21119,N_14305,N_15345);
and U21120 (N_21120,N_12918,N_14451);
nor U21121 (N_21121,N_13694,N_15976);
nor U21122 (N_21122,N_14649,N_16224);
or U21123 (N_21123,N_16432,N_14286);
xor U21124 (N_21124,N_16487,N_14266);
and U21125 (N_21125,N_15308,N_14315);
or U21126 (N_21126,N_14562,N_15632);
xnor U21127 (N_21127,N_14448,N_13742);
xnor U21128 (N_21128,N_13335,N_17290);
or U21129 (N_21129,N_15968,N_13069);
nor U21130 (N_21130,N_17176,N_18584);
xor U21131 (N_21131,N_15797,N_18166);
or U21132 (N_21132,N_17431,N_17069);
nor U21133 (N_21133,N_14770,N_14520);
xnor U21134 (N_21134,N_12741,N_15896);
or U21135 (N_21135,N_12950,N_16537);
or U21136 (N_21136,N_13043,N_16253);
nand U21137 (N_21137,N_18621,N_15389);
nand U21138 (N_21138,N_18169,N_18064);
nor U21139 (N_21139,N_17555,N_15078);
nand U21140 (N_21140,N_13064,N_16451);
nor U21141 (N_21141,N_16443,N_17640);
and U21142 (N_21142,N_14964,N_15283);
or U21143 (N_21143,N_14535,N_13807);
nand U21144 (N_21144,N_15739,N_18145);
and U21145 (N_21145,N_18205,N_13756);
or U21146 (N_21146,N_16648,N_14877);
or U21147 (N_21147,N_15761,N_13384);
or U21148 (N_21148,N_16653,N_12763);
and U21149 (N_21149,N_14375,N_16008);
and U21150 (N_21150,N_16022,N_14934);
and U21151 (N_21151,N_14105,N_12603);
and U21152 (N_21152,N_13832,N_15571);
or U21153 (N_21153,N_12663,N_16685);
nand U21154 (N_21154,N_17682,N_16842);
nor U21155 (N_21155,N_17537,N_12518);
nand U21156 (N_21156,N_14289,N_13160);
nor U21157 (N_21157,N_17569,N_15262);
or U21158 (N_21158,N_16695,N_13843);
nand U21159 (N_21159,N_18630,N_17107);
nor U21160 (N_21160,N_14133,N_15191);
or U21161 (N_21161,N_15368,N_18649);
nand U21162 (N_21162,N_13410,N_14761);
or U21163 (N_21163,N_18523,N_14124);
nor U21164 (N_21164,N_17391,N_18582);
and U21165 (N_21165,N_13659,N_13405);
nand U21166 (N_21166,N_14569,N_12605);
nand U21167 (N_21167,N_13107,N_17977);
xnor U21168 (N_21168,N_15018,N_12533);
or U21169 (N_21169,N_18419,N_13076);
or U21170 (N_21170,N_15467,N_18694);
or U21171 (N_21171,N_12626,N_15575);
nand U21172 (N_21172,N_16439,N_17845);
nand U21173 (N_21173,N_14321,N_14468);
and U21174 (N_21174,N_18513,N_17974);
and U21175 (N_21175,N_13760,N_15029);
nor U21176 (N_21176,N_16061,N_14901);
and U21177 (N_21177,N_16385,N_18317);
nand U21178 (N_21178,N_13626,N_17852);
or U21179 (N_21179,N_17698,N_18124);
nor U21180 (N_21180,N_14260,N_13695);
nor U21181 (N_21181,N_13736,N_13037);
nor U21182 (N_21182,N_13599,N_18724);
or U21183 (N_21183,N_15299,N_13835);
xnor U21184 (N_21184,N_17844,N_12844);
nor U21185 (N_21185,N_16515,N_14071);
or U21186 (N_21186,N_16801,N_17091);
and U21187 (N_21187,N_17118,N_15667);
nand U21188 (N_21188,N_15366,N_18493);
nand U21189 (N_21189,N_17716,N_18048);
and U21190 (N_21190,N_14924,N_16303);
and U21191 (N_21191,N_18682,N_13397);
or U21192 (N_21192,N_15240,N_15254);
nand U21193 (N_21193,N_16438,N_14630);
or U21194 (N_21194,N_18054,N_16497);
nor U21195 (N_21195,N_15293,N_14322);
nor U21196 (N_21196,N_14332,N_15556);
nor U21197 (N_21197,N_18744,N_16015);
nand U21198 (N_21198,N_12787,N_16563);
nand U21199 (N_21199,N_17139,N_15909);
xnor U21200 (N_21200,N_13199,N_18557);
or U21201 (N_21201,N_13820,N_14440);
nor U21202 (N_21202,N_15391,N_15025);
or U21203 (N_21203,N_13129,N_16585);
or U21204 (N_21204,N_15124,N_15771);
or U21205 (N_21205,N_16044,N_18204);
nand U21206 (N_21206,N_13247,N_14280);
xor U21207 (N_21207,N_12872,N_16725);
nor U21208 (N_21208,N_16532,N_15533);
and U21209 (N_21209,N_16864,N_18440);
or U21210 (N_21210,N_13822,N_16832);
and U21211 (N_21211,N_14501,N_18173);
or U21212 (N_21212,N_17993,N_16637);
nor U21213 (N_21213,N_13156,N_14963);
xnor U21214 (N_21214,N_13605,N_16117);
or U21215 (N_21215,N_17939,N_12537);
nor U21216 (N_21216,N_13563,N_17162);
or U21217 (N_21217,N_18212,N_16189);
or U21218 (N_21218,N_12520,N_12735);
or U21219 (N_21219,N_13194,N_17708);
xor U21220 (N_21220,N_14675,N_17133);
or U21221 (N_21221,N_14031,N_13258);
and U21222 (N_21222,N_17754,N_16323);
or U21223 (N_21223,N_15036,N_15200);
nor U21224 (N_21224,N_13341,N_18384);
or U21225 (N_21225,N_17847,N_12916);
xor U21226 (N_21226,N_18001,N_13308);
nor U21227 (N_21227,N_16440,N_18311);
and U21228 (N_21228,N_16789,N_14112);
or U21229 (N_21229,N_16252,N_13208);
and U21230 (N_21230,N_13747,N_15313);
or U21231 (N_21231,N_13688,N_15371);
nor U21232 (N_21232,N_15834,N_18514);
or U21233 (N_21233,N_13388,N_16627);
nand U21234 (N_21234,N_12699,N_15703);
nor U21235 (N_21235,N_15436,N_13241);
nor U21236 (N_21236,N_15174,N_14487);
or U21237 (N_21237,N_15472,N_15244);
nor U21238 (N_21238,N_14004,N_13624);
and U21239 (N_21239,N_13645,N_14026);
or U21240 (N_21240,N_14681,N_14110);
and U21241 (N_21241,N_13781,N_13601);
nand U21242 (N_21242,N_18056,N_18401);
or U21243 (N_21243,N_16409,N_13256);
or U21244 (N_21244,N_15554,N_13744);
and U21245 (N_21245,N_14296,N_16173);
and U21246 (N_21246,N_17780,N_17457);
xnor U21247 (N_21247,N_14379,N_17686);
and U21248 (N_21248,N_16387,N_15142);
and U21249 (N_21249,N_17971,N_15601);
or U21250 (N_21250,N_17676,N_13499);
nor U21251 (N_21251,N_14944,N_17985);
or U21252 (N_21252,N_16447,N_15012);
nor U21253 (N_21253,N_17733,N_17588);
and U21254 (N_21254,N_14972,N_16863);
and U21255 (N_21255,N_13354,N_16165);
xor U21256 (N_21256,N_17591,N_18141);
and U21257 (N_21257,N_18596,N_14950);
and U21258 (N_21258,N_16867,N_16913);
nor U21259 (N_21259,N_14291,N_17396);
or U21260 (N_21260,N_16425,N_15514);
nor U21261 (N_21261,N_18126,N_16833);
nor U21262 (N_21262,N_15252,N_13411);
nor U21263 (N_21263,N_13908,N_13486);
xor U21264 (N_21264,N_18281,N_18644);
or U21265 (N_21265,N_15430,N_15648);
and U21266 (N_21266,N_12795,N_13491);
or U21267 (N_21267,N_14818,N_17447);
nand U21268 (N_21268,N_16365,N_13441);
xnor U21269 (N_21269,N_13442,N_15216);
xnor U21270 (N_21270,N_15670,N_14861);
nor U21271 (N_21271,N_13039,N_12978);
xnor U21272 (N_21272,N_16900,N_18603);
nand U21273 (N_21273,N_14846,N_16814);
nor U21274 (N_21274,N_17334,N_16545);
or U21275 (N_21275,N_18408,N_13718);
nand U21276 (N_21276,N_15014,N_16808);
nand U21277 (N_21277,N_16373,N_17529);
and U21278 (N_21278,N_12777,N_14863);
or U21279 (N_21279,N_12943,N_18588);
and U21280 (N_21280,N_12656,N_13292);
nand U21281 (N_21281,N_13604,N_14390);
nor U21282 (N_21282,N_17270,N_17115);
nor U21283 (N_21283,N_13052,N_15023);
nand U21284 (N_21284,N_13349,N_17854);
or U21285 (N_21285,N_15707,N_13445);
nand U21286 (N_21286,N_15275,N_18176);
or U21287 (N_21287,N_15959,N_12933);
and U21288 (N_21288,N_13777,N_14135);
nand U21289 (N_21289,N_14716,N_15378);
and U21290 (N_21290,N_15330,N_17760);
nor U21291 (N_21291,N_13206,N_14810);
and U21292 (N_21292,N_15735,N_18246);
nor U21293 (N_21293,N_13644,N_16796);
or U21294 (N_21294,N_17220,N_17482);
nor U21295 (N_21295,N_16837,N_16151);
nor U21296 (N_21296,N_14372,N_14574);
nand U21297 (N_21297,N_13342,N_13260);
or U21298 (N_21298,N_13667,N_17758);
nor U21299 (N_21299,N_16937,N_16245);
or U21300 (N_21300,N_18426,N_17773);
or U21301 (N_21301,N_13347,N_17840);
nand U21302 (N_21302,N_14462,N_14591);
nor U21303 (N_21303,N_15767,N_18474);
and U21304 (N_21304,N_18076,N_16507);
nor U21305 (N_21305,N_14710,N_13930);
or U21306 (N_21306,N_13978,N_14446);
and U21307 (N_21307,N_18473,N_12790);
xnor U21308 (N_21308,N_12695,N_12578);
and U21309 (N_21309,N_16310,N_16668);
or U21310 (N_21310,N_15155,N_17507);
nor U21311 (N_21311,N_18409,N_16101);
nand U21312 (N_21312,N_13762,N_18522);
xnor U21313 (N_21313,N_12691,N_18073);
nand U21314 (N_21314,N_13188,N_14845);
and U21315 (N_21315,N_13582,N_17620);
nor U21316 (N_21316,N_16705,N_13155);
nor U21317 (N_21317,N_13337,N_13540);
nand U21318 (N_21318,N_16013,N_14491);
xnor U21319 (N_21319,N_15537,N_14841);
nand U21320 (N_21320,N_12788,N_12992);
and U21321 (N_21321,N_16158,N_12896);
nor U21322 (N_21322,N_13775,N_17735);
nand U21323 (N_21323,N_17565,N_14313);
nor U21324 (N_21324,N_17496,N_16348);
or U21325 (N_21325,N_14172,N_15937);
nand U21326 (N_21326,N_17901,N_18447);
and U21327 (N_21327,N_13799,N_18172);
nand U21328 (N_21328,N_16104,N_17706);
and U21329 (N_21329,N_16853,N_16985);
nand U21330 (N_21330,N_16377,N_15111);
nor U21331 (N_21331,N_13145,N_12898);
and U21332 (N_21332,N_14833,N_17891);
nor U21333 (N_21333,N_17257,N_15857);
or U21334 (N_21334,N_15347,N_13704);
or U21335 (N_21335,N_13178,N_17551);
nand U21336 (N_21336,N_14155,N_16617);
and U21337 (N_21337,N_14536,N_16428);
and U21338 (N_21338,N_16928,N_18609);
nand U21339 (N_21339,N_15838,N_15684);
nor U21340 (N_21340,N_17268,N_13528);
and U21341 (N_21341,N_17213,N_14551);
nand U21342 (N_21342,N_16629,N_13088);
xor U21343 (N_21343,N_13422,N_16342);
xor U21344 (N_21344,N_17217,N_14865);
xor U21345 (N_21345,N_16491,N_17888);
nor U21346 (N_21346,N_16823,N_13792);
nand U21347 (N_21347,N_14682,N_12670);
nor U21348 (N_21348,N_13821,N_13371);
nand U21349 (N_21349,N_15674,N_16894);
or U21350 (N_21350,N_13034,N_13287);
xnor U21351 (N_21351,N_13192,N_15908);
xnor U21352 (N_21352,N_17005,N_17700);
nand U21353 (N_21353,N_16735,N_17102);
nand U21354 (N_21354,N_16212,N_16709);
nand U21355 (N_21355,N_13564,N_15799);
nand U21356 (N_21356,N_16374,N_14329);
nand U21357 (N_21357,N_18128,N_18030);
or U21358 (N_21358,N_17975,N_18610);
nand U21359 (N_21359,N_14437,N_17624);
and U21360 (N_21360,N_18191,N_14492);
nor U21361 (N_21361,N_18017,N_15913);
nor U21362 (N_21362,N_15606,N_13679);
or U21363 (N_21363,N_13162,N_15520);
nor U21364 (N_21364,N_15546,N_16634);
and U21365 (N_21365,N_14700,N_17037);
nor U21366 (N_21366,N_15983,N_16358);
nand U21367 (N_21367,N_17362,N_16983);
nand U21368 (N_21368,N_17552,N_12705);
nor U21369 (N_21369,N_17378,N_15762);
or U21370 (N_21370,N_17476,N_15463);
or U21371 (N_21371,N_18689,N_12560);
nor U21372 (N_21372,N_15757,N_17332);
nand U21373 (N_21373,N_12853,N_14231);
nand U21374 (N_21374,N_16575,N_12824);
and U21375 (N_21375,N_17785,N_16672);
xor U21376 (N_21376,N_13570,N_17419);
nor U21377 (N_21377,N_18334,N_13474);
nor U21378 (N_21378,N_16682,N_13748);
or U21379 (N_21379,N_17051,N_14335);
xnor U21380 (N_21380,N_17008,N_17875);
or U21381 (N_21381,N_18385,N_17695);
nor U21382 (N_21382,N_18381,N_18374);
nand U21383 (N_21383,N_15384,N_14776);
nand U21384 (N_21384,N_15956,N_17211);
and U21385 (N_21385,N_18491,N_13952);
nor U21386 (N_21386,N_13409,N_13763);
xnor U21387 (N_21387,N_15653,N_15805);
and U21388 (N_21388,N_17643,N_16139);
nor U21389 (N_21389,N_14045,N_12685);
nand U21390 (N_21390,N_18542,N_16277);
xnor U21391 (N_21391,N_18485,N_17806);
and U21392 (N_21392,N_17231,N_14346);
and U21393 (N_21393,N_15438,N_17973);
or U21394 (N_21394,N_18359,N_17011);
nor U21395 (N_21395,N_16411,N_17484);
xor U21396 (N_21396,N_18025,N_13553);
or U21397 (N_21397,N_18586,N_13166);
nand U21398 (N_21398,N_15998,N_15381);
nand U21399 (N_21399,N_15722,N_13608);
nor U21400 (N_21400,N_16131,N_17455);
and U21401 (N_21401,N_13148,N_17253);
and U21402 (N_21402,N_17328,N_16910);
nor U21403 (N_21403,N_16878,N_17950);
and U21404 (N_21404,N_13826,N_15485);
or U21405 (N_21405,N_14960,N_16835);
and U21406 (N_21406,N_14966,N_13623);
nor U21407 (N_21407,N_17464,N_16152);
or U21408 (N_21408,N_14766,N_16517);
xnor U21409 (N_21409,N_16286,N_13498);
xor U21410 (N_21410,N_12698,N_16465);
and U21411 (N_21411,N_14065,N_14650);
nand U21412 (N_21412,N_14424,N_18653);
nand U21413 (N_21413,N_18091,N_15071);
and U21414 (N_21414,N_12812,N_14800);
nor U21415 (N_21415,N_14513,N_16610);
nand U21416 (N_21416,N_16933,N_16775);
or U21417 (N_21417,N_13589,N_15573);
and U21418 (N_21418,N_15783,N_15478);
nand U21419 (N_21419,N_12958,N_12655);
and U21420 (N_21420,N_13329,N_18449);
or U21421 (N_21421,N_14203,N_17372);
nand U21422 (N_21422,N_16744,N_18350);
nor U21423 (N_21423,N_12674,N_18670);
or U21424 (N_21424,N_13625,N_16393);
nor U21425 (N_21425,N_18045,N_14746);
nand U21426 (N_21426,N_13085,N_16565);
nand U21427 (N_21427,N_13333,N_14467);
nor U21428 (N_21428,N_15960,N_15619);
xor U21429 (N_21429,N_16036,N_13926);
nand U21430 (N_21430,N_12739,N_18527);
or U21431 (N_21431,N_16918,N_15579);
and U21432 (N_21432,N_16840,N_13650);
or U21433 (N_21433,N_17759,N_13217);
nor U21434 (N_21434,N_17641,N_14278);
nor U21435 (N_21435,N_14393,N_14301);
nor U21436 (N_21436,N_13647,N_16149);
or U21437 (N_21437,N_16300,N_15261);
or U21438 (N_21438,N_14312,N_13996);
and U21439 (N_21439,N_18253,N_13980);
or U21440 (N_21440,N_17242,N_17070);
nand U21441 (N_21441,N_18461,N_16880);
or U21442 (N_21442,N_16601,N_18469);
or U21443 (N_21443,N_18241,N_12809);
nor U21444 (N_21444,N_12912,N_15972);
nor U21445 (N_21445,N_13404,N_17865);
or U21446 (N_21446,N_13225,N_13997);
or U21447 (N_21447,N_16021,N_13526);
nand U21448 (N_21448,N_13169,N_15113);
or U21449 (N_21449,N_18009,N_13606);
or U21450 (N_21450,N_18476,N_17518);
nor U21451 (N_21451,N_15680,N_17065);
nand U21452 (N_21452,N_14814,N_15698);
or U21453 (N_21453,N_12636,N_12600);
and U21454 (N_21454,N_14053,N_16662);
and U21455 (N_21455,N_12649,N_17568);
or U21456 (N_21456,N_14741,N_13390);
nand U21457 (N_21457,N_17201,N_17872);
nor U21458 (N_21458,N_14694,N_12638);
nor U21459 (N_21459,N_13080,N_16350);
nor U21460 (N_21460,N_16649,N_15560);
or U21461 (N_21461,N_12791,N_15618);
or U21462 (N_21462,N_17984,N_17199);
nor U21463 (N_21463,N_18452,N_18693);
and U21464 (N_21464,N_12834,N_12661);
and U21465 (N_21465,N_13531,N_17963);
and U21466 (N_21466,N_13423,N_18521);
or U21467 (N_21467,N_17673,N_12782);
nor U21468 (N_21468,N_14905,N_16406);
and U21469 (N_21469,N_14871,N_14561);
nor U21470 (N_21470,N_13711,N_14290);
nand U21471 (N_21471,N_14658,N_16274);
nor U21472 (N_21472,N_13364,N_12527);
nand U21473 (N_21473,N_14836,N_16185);
and U21474 (N_21474,N_13845,N_12734);
and U21475 (N_21475,N_16235,N_16745);
nor U21476 (N_21476,N_16829,N_13226);
or U21477 (N_21477,N_13533,N_17387);
nand U21478 (N_21478,N_16667,N_16573);
nand U21479 (N_21479,N_14034,N_16366);
and U21480 (N_21480,N_12910,N_16770);
nand U21481 (N_21481,N_13127,N_16530);
nor U21482 (N_21482,N_15185,N_18478);
nand U21483 (N_21483,N_13628,N_13993);
nor U21484 (N_21484,N_17132,N_16176);
nand U21485 (N_21485,N_13943,N_14787);
nor U21486 (N_21486,N_14683,N_15304);
and U21487 (N_21487,N_18004,N_15049);
and U21488 (N_21488,N_17064,N_18037);
or U21489 (N_21489,N_12810,N_15927);
and U21490 (N_21490,N_18576,N_12750);
xor U21491 (N_21491,N_16780,N_16249);
or U21492 (N_21492,N_17749,N_17221);
nor U21493 (N_21493,N_15709,N_16355);
nor U21494 (N_21494,N_17182,N_15659);
or U21495 (N_21495,N_18482,N_17805);
nand U21496 (N_21496,N_13243,N_14337);
nand U21497 (N_21497,N_15713,N_14760);
and U21498 (N_21498,N_16171,N_12942);
nor U21499 (N_21499,N_17589,N_14540);
or U21500 (N_21500,N_16523,N_13093);
nor U21501 (N_21501,N_18136,N_18163);
nor U21502 (N_21502,N_17315,N_14866);
and U21503 (N_21503,N_14831,N_17258);
and U21504 (N_21504,N_15748,N_17597);
or U21505 (N_21505,N_16899,N_17273);
nand U21506 (N_21506,N_18007,N_14628);
or U21507 (N_21507,N_14020,N_17341);
nand U21508 (N_21508,N_14762,N_18318);
and U21509 (N_21509,N_15350,N_18291);
nand U21510 (N_21510,N_12952,N_12505);
nor U21511 (N_21511,N_14003,N_16838);
and U21512 (N_21512,N_14955,N_18024);
and U21513 (N_21513,N_13116,N_17938);
or U21514 (N_21514,N_16931,N_16973);
or U21515 (N_21515,N_13233,N_12634);
xnor U21516 (N_21516,N_17747,N_14528);
or U21517 (N_21517,N_17269,N_12775);
nand U21518 (N_21518,N_16580,N_15318);
or U21519 (N_21519,N_14426,N_14041);
and U21520 (N_21520,N_14639,N_14929);
and U21521 (N_21521,N_13525,N_17072);
nor U21522 (N_21522,N_13110,N_12573);
or U21523 (N_21523,N_17472,N_16181);
or U21524 (N_21524,N_12544,N_18313);
nand U21525 (N_21525,N_14735,N_17394);
nor U21526 (N_21526,N_16464,N_16064);
or U21527 (N_21527,N_15109,N_18006);
nor U21528 (N_21528,N_16469,N_15144);
xnor U21529 (N_21529,N_14359,N_16822);
xor U21530 (N_21530,N_18016,N_17501);
nor U21531 (N_21531,N_17384,N_12726);
and U21532 (N_21532,N_16866,N_17944);
nor U21533 (N_21533,N_16959,N_18020);
nand U21534 (N_21534,N_18236,N_15893);
or U21535 (N_21535,N_14702,N_15053);
xnor U21536 (N_21536,N_17803,N_16421);
nor U21537 (N_21537,N_14157,N_13983);
nand U21538 (N_21538,N_14035,N_16340);
or U21539 (N_21539,N_16041,N_14940);
and U21540 (N_21540,N_14191,N_17909);
or U21541 (N_21541,N_14417,N_18036);
nor U21542 (N_21542,N_16654,N_18498);
or U21543 (N_21543,N_17608,N_17808);
or U21544 (N_21544,N_16130,N_13348);
nand U21545 (N_21545,N_15411,N_15219);
or U21546 (N_21546,N_15710,N_15406);
nand U21547 (N_21547,N_13662,N_13011);
nand U21548 (N_21548,N_18031,N_13869);
nand U21549 (N_21549,N_15527,N_18526);
xor U21550 (N_21550,N_18487,N_17871);
or U21551 (N_21551,N_17965,N_12922);
nor U21552 (N_21552,N_18377,N_12830);
nand U21553 (N_21553,N_16834,N_15447);
nor U21554 (N_21554,N_17842,N_16886);
and U21555 (N_21555,N_17720,N_17647);
or U21556 (N_21556,N_15427,N_14202);
nand U21557 (N_21557,N_16462,N_13302);
xnor U21558 (N_21558,N_12581,N_14116);
nor U21559 (N_21559,N_13755,N_18155);
and U21560 (N_21560,N_16851,N_17177);
or U21561 (N_21561,N_17914,N_15686);
or U21562 (N_21562,N_14783,N_15337);
nor U21563 (N_21563,N_15197,N_13010);
xnor U21564 (N_21564,N_16652,N_16582);
or U21565 (N_21565,N_14173,N_17725);
xor U21566 (N_21566,N_17368,N_16655);
nand U21567 (N_21567,N_18112,N_15466);
nand U21568 (N_21568,N_17959,N_14721);
nand U21569 (N_21569,N_15868,N_16551);
or U21570 (N_21570,N_15657,N_15731);
nor U21571 (N_21571,N_15055,N_14247);
nor U21572 (N_21572,N_14968,N_13346);
and U21573 (N_21573,N_16221,N_13032);
and U21574 (N_21574,N_17649,N_13278);
and U21575 (N_21575,N_15059,N_17684);
or U21576 (N_21576,N_17899,N_18679);
or U21577 (N_21577,N_15551,N_13970);
or U21578 (N_21578,N_17687,N_18671);
or U21579 (N_21579,N_16187,N_12965);
and U21580 (N_21580,N_15120,N_17903);
and U21581 (N_21581,N_14218,N_17313);
and U21582 (N_21582,N_12672,N_13481);
nor U21583 (N_21583,N_14874,N_13451);
nor U21584 (N_21584,N_13773,N_17121);
and U21585 (N_21585,N_15030,N_17814);
and U21586 (N_21586,N_12929,N_17732);
nor U21587 (N_21587,N_18174,N_15008);
nand U21588 (N_21588,N_14891,N_14582);
and U21589 (N_21589,N_12979,N_15356);
nand U21590 (N_21590,N_15367,N_17063);
nand U21591 (N_21591,N_12679,N_17986);
xnor U21592 (N_21592,N_16924,N_16699);
and U21593 (N_21593,N_13403,N_14401);
nor U21594 (N_21594,N_15374,N_18251);
nand U21595 (N_21595,N_16767,N_17272);
and U21596 (N_21596,N_12947,N_17292);
nor U21597 (N_21597,N_14530,N_15061);
or U21598 (N_21598,N_18071,N_16790);
and U21599 (N_21599,N_14798,N_13325);
nor U21600 (N_21600,N_14987,N_14549);
or U21601 (N_21601,N_17859,N_16048);
nand U21602 (N_21602,N_14838,N_14790);
and U21603 (N_21603,N_17721,N_17056);
xor U21604 (N_21604,N_13802,N_14025);
or U21605 (N_21605,N_15334,N_16170);
nand U21606 (N_21606,N_18632,N_15870);
nor U21607 (N_21607,N_18303,N_13918);
nor U21608 (N_21608,N_17271,N_13793);
nand U21609 (N_21609,N_16204,N_15794);
and U21610 (N_21610,N_17410,N_13053);
and U21611 (N_21611,N_17318,N_12946);
nor U21612 (N_21612,N_18152,N_15169);
and U21613 (N_21613,N_18642,N_18178);
and U21614 (N_21614,N_12919,N_17058);
or U21615 (N_21615,N_17656,N_15013);
and U21616 (N_21616,N_17779,N_15861);
nor U21617 (N_21617,N_15054,N_18199);
and U21618 (N_21618,N_16925,N_15917);
nand U21619 (N_21619,N_17736,N_18183);
and U21620 (N_21620,N_18413,N_13432);
xor U21621 (N_21621,N_17444,N_16609);
or U21622 (N_21622,N_15768,N_16798);
xor U21623 (N_21623,N_16381,N_15493);
and U21624 (N_21624,N_17978,N_16401);
nor U21625 (N_21625,N_16076,N_13270);
nor U21626 (N_21626,N_17417,N_14729);
nand U21627 (N_21627,N_14527,N_14284);
and U21628 (N_21628,N_18605,N_17483);
xnor U21629 (N_21629,N_14709,N_18635);
nand U21630 (N_21630,N_14662,N_16694);
nor U21631 (N_21631,N_14070,N_17704);
nand U21632 (N_21632,N_15567,N_16912);
nand U21633 (N_21633,N_15821,N_14410);
nor U21634 (N_21634,N_18201,N_14430);
nand U21635 (N_21635,N_17737,N_18506);
or U21636 (N_21636,N_16974,N_14444);
nor U21637 (N_21637,N_16621,N_13144);
or U21638 (N_21638,N_13047,N_16598);
nor U21639 (N_21639,N_12827,N_15980);
xor U21640 (N_21640,N_14227,N_15017);
and U21641 (N_21641,N_16341,N_13376);
nor U21642 (N_21642,N_18488,N_12975);
or U21643 (N_21643,N_18217,N_17801);
nand U21644 (N_21644,N_14470,N_14264);
xnor U21645 (N_21645,N_14580,N_15232);
nand U21646 (N_21646,N_14292,N_16299);
and U21647 (N_21647,N_12865,N_14370);
or U21648 (N_21648,N_13919,N_13796);
and U21649 (N_21649,N_17527,N_12890);
nor U21650 (N_21650,N_17688,N_15665);
or U21651 (N_21651,N_18117,N_16674);
nand U21652 (N_21652,N_16400,N_18453);
and U21653 (N_21653,N_18190,N_15993);
or U21654 (N_21654,N_15255,N_18528);
nor U21655 (N_21655,N_17487,N_14933);
or U21656 (N_21656,N_15720,N_18399);
nand U21657 (N_21657,N_16778,N_15876);
nor U21658 (N_21658,N_15171,N_16094);
nor U21659 (N_21659,N_13146,N_15034);
nand U21660 (N_21660,N_14119,N_16075);
nor U21661 (N_21661,N_14993,N_13699);
xnor U21662 (N_21662,N_16093,N_16069);
and U21663 (N_21663,N_18441,N_17053);
or U21664 (N_21664,N_17582,N_13888);
or U21665 (N_21665,N_13861,N_17723);
nand U21666 (N_21666,N_15766,N_14109);
nor U21667 (N_21667,N_16226,N_17082);
xnor U21668 (N_21668,N_17933,N_18492);
nand U21669 (N_21669,N_17895,N_17361);
and U21670 (N_21670,N_13369,N_16128);
or U21671 (N_21671,N_14745,N_16704);
nor U21672 (N_21672,N_17677,N_18430);
and U21673 (N_21673,N_12704,N_18728);
and U21674 (N_21674,N_17838,N_17090);
and U21675 (N_21675,N_13955,N_18422);
and U21676 (N_21676,N_14952,N_13465);
nor U21677 (N_21677,N_14088,N_15625);
nor U21678 (N_21678,N_18370,N_17862);
or U21679 (N_21679,N_14151,N_17414);
nor U21680 (N_21680,N_15850,N_14421);
xor U21681 (N_21681,N_16296,N_13415);
or U21682 (N_21682,N_17044,N_14400);
and U21683 (N_21683,N_17564,N_15916);
or U21684 (N_21684,N_18310,N_18100);
nor U21685 (N_21685,N_15235,N_18676);
or U21686 (N_21686,N_14408,N_18008);
xor U21687 (N_21687,N_14261,N_12725);
nand U21688 (N_21688,N_13361,N_14815);
or U21689 (N_21689,N_16190,N_13051);
nor U21690 (N_21690,N_16684,N_17192);
nand U21691 (N_21691,N_14480,N_17491);
and U21692 (N_21692,N_13969,N_15281);
xnor U21693 (N_21693,N_13340,N_14554);
nand U21694 (N_21694,N_13120,N_15453);
nor U21695 (N_21695,N_13101,N_13765);
nand U21696 (N_21696,N_17351,N_14725);
nor U21697 (N_21697,N_12762,N_15672);
nand U21698 (N_21698,N_16108,N_16298);
and U21699 (N_21699,N_12566,N_13710);
or U21700 (N_21700,N_13929,N_13594);
and U21701 (N_21701,N_12863,N_12686);
and U21702 (N_21702,N_17637,N_18411);
and U21703 (N_21703,N_15108,N_13771);
nor U21704 (N_21704,N_17154,N_18736);
nor U21705 (N_21705,N_14671,N_17813);
and U21706 (N_21706,N_12597,N_13121);
and U21707 (N_21707,N_17143,N_17474);
nand U21708 (N_21708,N_13387,N_15775);
nor U21709 (N_21709,N_18029,N_16691);
nor U21710 (N_21710,N_12500,N_12615);
xnor U21711 (N_21711,N_17874,N_12807);
nand U21712 (N_21712,N_18529,N_15651);
or U21713 (N_21713,N_17155,N_15936);
and U21714 (N_21714,N_18081,N_16238);
nand U21715 (N_21715,N_17303,N_15100);
nand U21716 (N_21716,N_13721,N_12732);
xor U21717 (N_21717,N_13097,N_13702);
xor U21718 (N_21718,N_15044,N_16082);
or U21719 (N_21719,N_13082,N_18085);
or U21720 (N_21720,N_16923,N_13294);
nor U21721 (N_21721,N_15273,N_17777);
nand U21722 (N_21722,N_14701,N_13326);
and U21723 (N_21723,N_15865,N_15376);
xnor U21724 (N_21724,N_17049,N_17329);
nor U21725 (N_21725,N_16903,N_12892);
nor U21726 (N_21726,N_13592,N_16014);
nor U21727 (N_21727,N_15168,N_15473);
or U21728 (N_21728,N_12703,N_12917);
nor U21729 (N_21729,N_14435,N_15786);
nand U21730 (N_21730,N_13003,N_15523);
xnor U21731 (N_21731,N_14310,N_12937);
or U21732 (N_21732,N_14015,N_18060);
and U21733 (N_21733,N_14896,N_18289);
nand U21734 (N_21734,N_18157,N_14352);
nor U21735 (N_21735,N_17945,N_14083);
xnor U21736 (N_21736,N_16159,N_17834);
and U21737 (N_21737,N_14864,N_17029);
or U21738 (N_21738,N_16836,N_18286);
nand U21739 (N_21739,N_18380,N_15806);
nand U21740 (N_21740,N_16474,N_12645);
or U21741 (N_21741,N_17863,N_14904);
or U21742 (N_21742,N_17471,N_13322);
and U21743 (N_21743,N_18050,N_14568);
and U21744 (N_21744,N_13530,N_15042);
xnor U21745 (N_21745,N_13959,N_16343);
nor U21746 (N_21746,N_12607,N_16843);
nand U21747 (N_21747,N_18321,N_18200);
or U21748 (N_21748,N_13229,N_12921);
nor U21749 (N_21749,N_17007,N_18625);
or U21750 (N_21750,N_17793,N_12591);
and U21751 (N_21751,N_18618,N_15442);
xnor U21752 (N_21752,N_12886,N_12676);
nor U21753 (N_21753,N_16897,N_15965);
nor U21754 (N_21754,N_18224,N_17388);
and U21755 (N_21755,N_16727,N_18549);
nor U21756 (N_21756,N_15039,N_18457);
nor U21757 (N_21757,N_13301,N_14374);
and U21758 (N_21758,N_12944,N_13400);
nor U21759 (N_21759,N_16950,N_18077);
and U21760 (N_21760,N_15699,N_18175);
or U21761 (N_21761,N_16724,N_15423);
or U21762 (N_21762,N_16723,N_13814);
or U21763 (N_21763,N_15928,N_13515);
or U21764 (N_21764,N_12837,N_15541);
and U21765 (N_21765,N_15398,N_14175);
xor U21766 (N_21766,N_14190,N_13883);
or U21767 (N_21767,N_14499,N_18320);
and U21768 (N_21768,N_13506,N_17452);
or U21769 (N_21769,N_17174,N_12871);
nor U21770 (N_21770,N_13001,N_17868);
nand U21771 (N_21771,N_14423,N_16556);
xnor U21772 (N_21772,N_14225,N_16223);
and U21773 (N_21773,N_15317,N_16825);
nor U21774 (N_21774,N_15765,N_14223);
or U21775 (N_21775,N_17585,N_17902);
xor U21776 (N_21776,N_15138,N_13065);
or U21777 (N_21777,N_16904,N_14330);
and U21778 (N_21778,N_13632,N_14685);
or U21779 (N_21779,N_15253,N_15032);
and U21780 (N_21780,N_15300,N_13168);
and U21781 (N_21781,N_15040,N_16862);
nand U21782 (N_21782,N_13574,N_14984);
xnor U21783 (N_21783,N_16535,N_16962);
or U21784 (N_21784,N_14931,N_17022);
nand U21785 (N_21785,N_15237,N_16201);
nor U21786 (N_21786,N_16599,N_12715);
nand U21787 (N_21787,N_14303,N_17593);
and U21788 (N_21788,N_18569,N_15073);
nor U21789 (N_21789,N_16307,N_14768);
nand U21790 (N_21790,N_13479,N_15992);
xnor U21791 (N_21791,N_18383,N_15842);
nand U21792 (N_21792,N_17921,N_13934);
nor U21793 (N_21793,N_13874,N_17418);
xnor U21794 (N_21794,N_14450,N_15024);
nand U21795 (N_21795,N_12502,N_16622);
nand U21796 (N_21796,N_15938,N_18068);
and U21797 (N_21797,N_12531,N_18672);
and U21798 (N_21798,N_14969,N_17783);
and U21799 (N_21799,N_16945,N_18615);
and U21800 (N_21800,N_15383,N_15977);
and U21801 (N_21801,N_15245,N_18094);
or U21802 (N_21802,N_12737,N_14239);
and U21803 (N_21803,N_12576,N_13682);
nor U21804 (N_21804,N_14489,N_18255);
and U21805 (N_21805,N_13150,N_14719);
and U21806 (N_21806,N_15361,N_18558);
and U21807 (N_21807,N_18561,N_15801);
and U21808 (N_21808,N_14282,N_16399);
or U21809 (N_21809,N_15208,N_13214);
nor U21810 (N_21810,N_12993,N_13976);
and U21811 (N_21811,N_16995,N_16957);
nand U21812 (N_21812,N_16813,N_18714);
or U21813 (N_21813,N_15224,N_15578);
nor U21814 (N_21814,N_15107,N_15955);
and U21815 (N_21815,N_15209,N_13014);
nand U21816 (N_21816,N_18685,N_18040);
and U21817 (N_21817,N_14817,N_13073);
nor U21818 (N_21818,N_13420,N_13239);
nand U21819 (N_21819,N_12534,N_18034);
nand U21820 (N_21820,N_18730,N_15489);
and U21821 (N_21821,N_18489,N_16063);
nand U21822 (N_21822,N_16045,N_18604);
nand U21823 (N_21823,N_16940,N_13629);
nor U21824 (N_21824,N_17544,N_12666);
nor U21825 (N_21825,N_13666,N_18084);
nor U21826 (N_21826,N_18663,N_17422);
nor U21827 (N_21827,N_17325,N_13314);
and U21828 (N_21828,N_13487,N_16890);
or U21829 (N_21829,N_13372,N_14981);
and U21830 (N_21830,N_15576,N_13330);
and U21831 (N_21831,N_17352,N_15915);
and U21832 (N_21832,N_15284,N_16934);
nand U21833 (N_21833,N_15492,N_17078);
xnor U21834 (N_21834,N_16073,N_13977);
xor U21835 (N_21835,N_16911,N_14032);
nor U21836 (N_21836,N_14249,N_13139);
nand U21837 (N_21837,N_16309,N_14538);
nand U21838 (N_21838,N_15339,N_18351);
nand U21839 (N_21839,N_17627,N_15816);
nor U21840 (N_21840,N_16398,N_15429);
and U21841 (N_21841,N_15645,N_15782);
xor U21842 (N_21842,N_12660,N_15688);
and U21843 (N_21843,N_16531,N_15784);
and U21844 (N_21844,N_17766,N_18664);
or U21845 (N_21845,N_15105,N_15777);
nor U21846 (N_21846,N_14737,N_15295);
xor U21847 (N_21847,N_15841,N_18477);
and U21848 (N_21848,N_18066,N_15555);
or U21849 (N_21849,N_18276,N_14069);
and U21850 (N_21850,N_18132,N_17402);
nand U21851 (N_21851,N_17423,N_15741);
or U21852 (N_21852,N_17848,N_14541);
or U21853 (N_21853,N_17019,N_15385);
or U21854 (N_21854,N_18748,N_14272);
nor U21855 (N_21855,N_17494,N_17032);
and U21856 (N_21856,N_14567,N_15452);
or U21857 (N_21857,N_15871,N_15141);
nand U21858 (N_21858,N_17050,N_14888);
nor U21859 (N_21859,N_12532,N_15157);
xor U21860 (N_21860,N_14439,N_14565);
and U21861 (N_21861,N_16568,N_14589);
and U21862 (N_21862,N_17411,N_15884);
and U21863 (N_21863,N_13136,N_12973);
nor U21864 (N_21864,N_15788,N_18700);
or U21865 (N_21865,N_14826,N_15156);
xor U21866 (N_21866,N_13936,N_17498);
nand U21867 (N_21867,N_15432,N_17726);
nor U21868 (N_21868,N_16396,N_16922);
or U21869 (N_21869,N_13500,N_16233);
or U21870 (N_21870,N_17353,N_16592);
or U21871 (N_21871,N_17832,N_12839);
xor U21872 (N_21872,N_16984,N_15586);
nand U21873 (N_21873,N_13408,N_16018);
nand U21874 (N_21874,N_13527,N_16470);
or U21875 (N_21875,N_16848,N_18153);
and U21876 (N_21876,N_14840,N_17237);
nor U21877 (N_21877,N_14641,N_14682);
or U21878 (N_21878,N_17896,N_15542);
nor U21879 (N_21879,N_15944,N_17655);
or U21880 (N_21880,N_15340,N_17914);
and U21881 (N_21881,N_15904,N_16847);
nor U21882 (N_21882,N_15532,N_15076);
nand U21883 (N_21883,N_17895,N_13774);
and U21884 (N_21884,N_14632,N_17548);
xnor U21885 (N_21885,N_13430,N_17792);
nor U21886 (N_21886,N_13266,N_16447);
or U21887 (N_21887,N_16026,N_13237);
nor U21888 (N_21888,N_17913,N_17493);
nor U21889 (N_21889,N_16644,N_14886);
nand U21890 (N_21890,N_14853,N_14840);
nand U21891 (N_21891,N_13536,N_16710);
or U21892 (N_21892,N_14485,N_17270);
or U21893 (N_21893,N_17693,N_13378);
and U21894 (N_21894,N_14017,N_12681);
or U21895 (N_21895,N_13455,N_17942);
nor U21896 (N_21896,N_18607,N_18113);
and U21897 (N_21897,N_12602,N_15498);
or U21898 (N_21898,N_15878,N_12866);
and U21899 (N_21899,N_13665,N_12568);
xnor U21900 (N_21900,N_15728,N_18000);
xor U21901 (N_21901,N_12594,N_12950);
or U21902 (N_21902,N_16448,N_15429);
nor U21903 (N_21903,N_13692,N_17425);
and U21904 (N_21904,N_15023,N_18220);
nor U21905 (N_21905,N_18256,N_18476);
or U21906 (N_21906,N_16953,N_13844);
and U21907 (N_21907,N_18742,N_13006);
nor U21908 (N_21908,N_15482,N_14291);
xnor U21909 (N_21909,N_16976,N_14241);
nor U21910 (N_21910,N_13814,N_15327);
and U21911 (N_21911,N_14528,N_16262);
or U21912 (N_21912,N_13026,N_14931);
nand U21913 (N_21913,N_15634,N_15726);
or U21914 (N_21914,N_17321,N_17485);
nor U21915 (N_21915,N_17175,N_15925);
or U21916 (N_21916,N_16429,N_17718);
nor U21917 (N_21917,N_17949,N_17259);
and U21918 (N_21918,N_17217,N_16508);
nand U21919 (N_21919,N_14241,N_16959);
xnor U21920 (N_21920,N_15407,N_13430);
nand U21921 (N_21921,N_14475,N_17998);
nand U21922 (N_21922,N_13197,N_14572);
or U21923 (N_21923,N_17344,N_15241);
nor U21924 (N_21924,N_14482,N_13545);
or U21925 (N_21925,N_12602,N_15556);
or U21926 (N_21926,N_15804,N_17265);
nor U21927 (N_21927,N_15352,N_14914);
or U21928 (N_21928,N_12569,N_16956);
and U21929 (N_21929,N_14717,N_17098);
nor U21930 (N_21930,N_15060,N_14551);
and U21931 (N_21931,N_14614,N_14864);
or U21932 (N_21932,N_14188,N_12837);
or U21933 (N_21933,N_17485,N_15914);
nand U21934 (N_21934,N_18027,N_14673);
xor U21935 (N_21935,N_14701,N_17928);
and U21936 (N_21936,N_14936,N_16420);
nand U21937 (N_21937,N_15989,N_13751);
nand U21938 (N_21938,N_18497,N_18537);
nand U21939 (N_21939,N_15929,N_17086);
nand U21940 (N_21940,N_18133,N_14170);
and U21941 (N_21941,N_14983,N_13291);
or U21942 (N_21942,N_16285,N_14161);
nand U21943 (N_21943,N_15360,N_15489);
and U21944 (N_21944,N_14368,N_12770);
nor U21945 (N_21945,N_13426,N_13949);
nand U21946 (N_21946,N_15837,N_18509);
and U21947 (N_21947,N_17048,N_14934);
or U21948 (N_21948,N_13985,N_17203);
and U21949 (N_21949,N_15470,N_14061);
and U21950 (N_21950,N_13958,N_15351);
nand U21951 (N_21951,N_13902,N_12954);
xor U21952 (N_21952,N_13960,N_16957);
and U21953 (N_21953,N_18316,N_17086);
nor U21954 (N_21954,N_14972,N_17628);
and U21955 (N_21955,N_18249,N_13103);
nor U21956 (N_21956,N_15025,N_15741);
and U21957 (N_21957,N_16327,N_15697);
nor U21958 (N_21958,N_18388,N_13849);
nor U21959 (N_21959,N_18197,N_12929);
and U21960 (N_21960,N_18708,N_17382);
or U21961 (N_21961,N_14935,N_17454);
and U21962 (N_21962,N_14486,N_17563);
nand U21963 (N_21963,N_18375,N_17267);
nand U21964 (N_21964,N_16835,N_17512);
or U21965 (N_21965,N_15114,N_15018);
nor U21966 (N_21966,N_14011,N_12697);
and U21967 (N_21967,N_16911,N_14868);
nand U21968 (N_21968,N_15531,N_18206);
nand U21969 (N_21969,N_16751,N_13419);
nand U21970 (N_21970,N_13280,N_16248);
and U21971 (N_21971,N_14122,N_12940);
and U21972 (N_21972,N_15180,N_17944);
and U21973 (N_21973,N_16449,N_13067);
nand U21974 (N_21974,N_14197,N_14433);
nor U21975 (N_21975,N_17940,N_17800);
or U21976 (N_21976,N_18620,N_15622);
or U21977 (N_21977,N_12541,N_15454);
nor U21978 (N_21978,N_13413,N_15177);
nand U21979 (N_21979,N_14076,N_17099);
nand U21980 (N_21980,N_17942,N_15691);
and U21981 (N_21981,N_13504,N_17376);
or U21982 (N_21982,N_15277,N_16758);
nor U21983 (N_21983,N_15070,N_18697);
xor U21984 (N_21984,N_15100,N_17282);
and U21985 (N_21985,N_13461,N_17119);
or U21986 (N_21986,N_13772,N_15448);
nor U21987 (N_21987,N_18592,N_14948);
and U21988 (N_21988,N_17785,N_12873);
nor U21989 (N_21989,N_17029,N_14659);
xnor U21990 (N_21990,N_16365,N_14748);
or U21991 (N_21991,N_16304,N_13222);
nor U21992 (N_21992,N_16157,N_13613);
and U21993 (N_21993,N_17277,N_12732);
or U21994 (N_21994,N_15405,N_15913);
or U21995 (N_21995,N_16707,N_18284);
nor U21996 (N_21996,N_14208,N_12871);
nand U21997 (N_21997,N_17280,N_13507);
nand U21998 (N_21998,N_13688,N_18304);
or U21999 (N_21999,N_18563,N_14111);
or U22000 (N_22000,N_13254,N_15074);
nand U22001 (N_22001,N_15738,N_14024);
nor U22002 (N_22002,N_17257,N_17695);
nand U22003 (N_22003,N_14814,N_16271);
nand U22004 (N_22004,N_17031,N_16089);
and U22005 (N_22005,N_15210,N_17325);
xnor U22006 (N_22006,N_16230,N_18124);
and U22007 (N_22007,N_18643,N_12895);
and U22008 (N_22008,N_16742,N_14401);
or U22009 (N_22009,N_14461,N_16068);
or U22010 (N_22010,N_16980,N_15005);
nand U22011 (N_22011,N_17371,N_15853);
nor U22012 (N_22012,N_18279,N_17714);
and U22013 (N_22013,N_14389,N_16544);
or U22014 (N_22014,N_12964,N_15731);
and U22015 (N_22015,N_13087,N_15276);
or U22016 (N_22016,N_14876,N_16446);
nand U22017 (N_22017,N_13580,N_18459);
nand U22018 (N_22018,N_18112,N_14755);
and U22019 (N_22019,N_15259,N_18347);
nand U22020 (N_22020,N_18073,N_17386);
or U22021 (N_22021,N_17144,N_14131);
nand U22022 (N_22022,N_16948,N_14654);
or U22023 (N_22023,N_14205,N_15997);
nor U22024 (N_22024,N_14918,N_17501);
nor U22025 (N_22025,N_15326,N_15752);
nor U22026 (N_22026,N_12946,N_13056);
nand U22027 (N_22027,N_16944,N_13808);
and U22028 (N_22028,N_18632,N_16955);
and U22029 (N_22029,N_17600,N_14253);
and U22030 (N_22030,N_14171,N_16094);
and U22031 (N_22031,N_14073,N_13025);
nand U22032 (N_22032,N_17114,N_13001);
nor U22033 (N_22033,N_17392,N_18444);
nor U22034 (N_22034,N_17874,N_16504);
nor U22035 (N_22035,N_17517,N_15304);
nand U22036 (N_22036,N_12774,N_12810);
nor U22037 (N_22037,N_17308,N_14274);
and U22038 (N_22038,N_18518,N_14114);
and U22039 (N_22039,N_16568,N_14808);
nor U22040 (N_22040,N_14317,N_18365);
or U22041 (N_22041,N_16202,N_13595);
and U22042 (N_22042,N_16281,N_18743);
or U22043 (N_22043,N_16670,N_14361);
nand U22044 (N_22044,N_15406,N_14260);
or U22045 (N_22045,N_16629,N_12682);
nor U22046 (N_22046,N_14902,N_17847);
nand U22047 (N_22047,N_17694,N_12979);
nand U22048 (N_22048,N_17633,N_15086);
and U22049 (N_22049,N_17562,N_18283);
xnor U22050 (N_22050,N_13664,N_18224);
nor U22051 (N_22051,N_14527,N_16731);
nor U22052 (N_22052,N_16041,N_18719);
xnor U22053 (N_22053,N_15621,N_17291);
and U22054 (N_22054,N_14087,N_14874);
and U22055 (N_22055,N_12911,N_13173);
nor U22056 (N_22056,N_13503,N_13096);
nand U22057 (N_22057,N_12627,N_12559);
nand U22058 (N_22058,N_18241,N_15517);
nor U22059 (N_22059,N_16389,N_17687);
and U22060 (N_22060,N_18560,N_17797);
and U22061 (N_22061,N_16679,N_14137);
and U22062 (N_22062,N_17715,N_13914);
or U22063 (N_22063,N_15319,N_15298);
and U22064 (N_22064,N_16908,N_15972);
nand U22065 (N_22065,N_18254,N_15663);
or U22066 (N_22066,N_14942,N_16047);
nor U22067 (N_22067,N_18288,N_12647);
and U22068 (N_22068,N_13249,N_16007);
nand U22069 (N_22069,N_15659,N_13254);
nor U22070 (N_22070,N_17252,N_17659);
and U22071 (N_22071,N_12787,N_18666);
xor U22072 (N_22072,N_18117,N_14914);
nand U22073 (N_22073,N_15088,N_15893);
or U22074 (N_22074,N_17893,N_14206);
nand U22075 (N_22075,N_14874,N_18450);
nor U22076 (N_22076,N_15548,N_16402);
nand U22077 (N_22077,N_17807,N_12629);
nand U22078 (N_22078,N_13940,N_13143);
or U22079 (N_22079,N_15117,N_17552);
xor U22080 (N_22080,N_17807,N_15409);
nor U22081 (N_22081,N_14312,N_16787);
xnor U22082 (N_22082,N_15651,N_18304);
nor U22083 (N_22083,N_17190,N_15100);
and U22084 (N_22084,N_14895,N_17047);
or U22085 (N_22085,N_14229,N_18489);
and U22086 (N_22086,N_15657,N_14878);
nand U22087 (N_22087,N_13310,N_17936);
nand U22088 (N_22088,N_12774,N_16465);
and U22089 (N_22089,N_15282,N_14307);
and U22090 (N_22090,N_16436,N_15479);
and U22091 (N_22091,N_17520,N_17824);
nand U22092 (N_22092,N_18499,N_13574);
nand U22093 (N_22093,N_18329,N_15393);
nand U22094 (N_22094,N_15336,N_18344);
nor U22095 (N_22095,N_17755,N_13698);
xor U22096 (N_22096,N_13748,N_15633);
and U22097 (N_22097,N_12736,N_13503);
xor U22098 (N_22098,N_13706,N_18532);
or U22099 (N_22099,N_17854,N_15910);
and U22100 (N_22100,N_18717,N_15165);
nor U22101 (N_22101,N_15457,N_14079);
nand U22102 (N_22102,N_16710,N_16403);
nand U22103 (N_22103,N_16371,N_12576);
nand U22104 (N_22104,N_14575,N_15944);
nor U22105 (N_22105,N_16996,N_14089);
nand U22106 (N_22106,N_18435,N_17285);
nor U22107 (N_22107,N_15399,N_13359);
nor U22108 (N_22108,N_14981,N_16366);
and U22109 (N_22109,N_16031,N_12671);
nor U22110 (N_22110,N_12506,N_14144);
nand U22111 (N_22111,N_16543,N_16439);
or U22112 (N_22112,N_18594,N_13368);
xnor U22113 (N_22113,N_13108,N_14709);
nand U22114 (N_22114,N_14674,N_14068);
and U22115 (N_22115,N_16234,N_16300);
xnor U22116 (N_22116,N_16278,N_16810);
or U22117 (N_22117,N_14691,N_16033);
or U22118 (N_22118,N_14047,N_14152);
nor U22119 (N_22119,N_13384,N_18192);
and U22120 (N_22120,N_18366,N_17237);
and U22121 (N_22121,N_15535,N_13558);
and U22122 (N_22122,N_17310,N_18050);
and U22123 (N_22123,N_15501,N_15039);
or U22124 (N_22124,N_14540,N_13314);
nand U22125 (N_22125,N_12676,N_15153);
nor U22126 (N_22126,N_12622,N_14280);
and U22127 (N_22127,N_15059,N_16438);
xor U22128 (N_22128,N_16901,N_14353);
or U22129 (N_22129,N_15207,N_18406);
nand U22130 (N_22130,N_13006,N_18677);
nor U22131 (N_22131,N_17340,N_16589);
nor U22132 (N_22132,N_13767,N_17281);
and U22133 (N_22133,N_16321,N_16873);
or U22134 (N_22134,N_14839,N_18066);
or U22135 (N_22135,N_14160,N_14346);
xor U22136 (N_22136,N_15986,N_14790);
and U22137 (N_22137,N_15045,N_17298);
nor U22138 (N_22138,N_16896,N_13909);
nand U22139 (N_22139,N_14851,N_13194);
and U22140 (N_22140,N_12623,N_18430);
nor U22141 (N_22141,N_13424,N_15819);
nor U22142 (N_22142,N_18644,N_17018);
nand U22143 (N_22143,N_13407,N_16381);
or U22144 (N_22144,N_16986,N_16239);
and U22145 (N_22145,N_14372,N_17446);
and U22146 (N_22146,N_18345,N_13776);
or U22147 (N_22147,N_14303,N_18093);
and U22148 (N_22148,N_18586,N_18334);
nor U22149 (N_22149,N_12962,N_14583);
or U22150 (N_22150,N_16803,N_16245);
and U22151 (N_22151,N_15127,N_18276);
nand U22152 (N_22152,N_15282,N_17470);
nand U22153 (N_22153,N_15247,N_14934);
or U22154 (N_22154,N_17362,N_12517);
nor U22155 (N_22155,N_16727,N_12946);
xnor U22156 (N_22156,N_18385,N_15246);
xnor U22157 (N_22157,N_16944,N_16119);
and U22158 (N_22158,N_15022,N_14799);
xor U22159 (N_22159,N_15869,N_15540);
or U22160 (N_22160,N_16356,N_13003);
and U22161 (N_22161,N_14718,N_14526);
nand U22162 (N_22162,N_17818,N_16384);
nand U22163 (N_22163,N_16009,N_17119);
and U22164 (N_22164,N_13415,N_17949);
nor U22165 (N_22165,N_17773,N_15661);
or U22166 (N_22166,N_14859,N_17766);
nand U22167 (N_22167,N_12534,N_12871);
or U22168 (N_22168,N_15186,N_18738);
and U22169 (N_22169,N_16128,N_17141);
or U22170 (N_22170,N_16496,N_17804);
nand U22171 (N_22171,N_17064,N_16581);
or U22172 (N_22172,N_13131,N_17098);
and U22173 (N_22173,N_18310,N_14995);
nand U22174 (N_22174,N_15113,N_15592);
nor U22175 (N_22175,N_12688,N_13782);
nand U22176 (N_22176,N_13600,N_14651);
nand U22177 (N_22177,N_16730,N_17313);
xor U22178 (N_22178,N_18150,N_17140);
nand U22179 (N_22179,N_13322,N_16865);
nand U22180 (N_22180,N_14997,N_17348);
xnor U22181 (N_22181,N_17750,N_14491);
and U22182 (N_22182,N_15091,N_14617);
or U22183 (N_22183,N_14574,N_17944);
or U22184 (N_22184,N_12804,N_17499);
nor U22185 (N_22185,N_17343,N_13740);
nor U22186 (N_22186,N_18514,N_14365);
nand U22187 (N_22187,N_17828,N_16336);
or U22188 (N_22188,N_12725,N_18026);
or U22189 (N_22189,N_17873,N_17918);
nand U22190 (N_22190,N_16447,N_14708);
and U22191 (N_22191,N_12536,N_15991);
nor U22192 (N_22192,N_17447,N_14664);
nand U22193 (N_22193,N_12744,N_13759);
or U22194 (N_22194,N_17378,N_18748);
nor U22195 (N_22195,N_15489,N_16550);
or U22196 (N_22196,N_16289,N_14423);
or U22197 (N_22197,N_14120,N_18172);
nor U22198 (N_22198,N_13660,N_15794);
nand U22199 (N_22199,N_15721,N_13773);
and U22200 (N_22200,N_17176,N_14299);
nand U22201 (N_22201,N_15894,N_16059);
nor U22202 (N_22202,N_14944,N_14073);
nor U22203 (N_22203,N_17626,N_15370);
and U22204 (N_22204,N_12930,N_18045);
xor U22205 (N_22205,N_13815,N_16598);
or U22206 (N_22206,N_14635,N_14299);
and U22207 (N_22207,N_14955,N_16214);
and U22208 (N_22208,N_16482,N_15826);
nand U22209 (N_22209,N_15533,N_16964);
and U22210 (N_22210,N_14259,N_13885);
nor U22211 (N_22211,N_15903,N_17300);
nand U22212 (N_22212,N_17381,N_14414);
and U22213 (N_22213,N_17351,N_12743);
nand U22214 (N_22214,N_14389,N_14055);
and U22215 (N_22215,N_15021,N_17140);
xor U22216 (N_22216,N_18596,N_17862);
or U22217 (N_22217,N_14029,N_12649);
xor U22218 (N_22218,N_14502,N_13890);
nor U22219 (N_22219,N_14477,N_13278);
xnor U22220 (N_22220,N_15265,N_16417);
or U22221 (N_22221,N_15421,N_17988);
and U22222 (N_22222,N_16264,N_12823);
and U22223 (N_22223,N_16026,N_16073);
or U22224 (N_22224,N_15100,N_15832);
xnor U22225 (N_22225,N_17056,N_16465);
and U22226 (N_22226,N_13803,N_17422);
nor U22227 (N_22227,N_13842,N_18224);
or U22228 (N_22228,N_16387,N_17489);
or U22229 (N_22229,N_16846,N_18382);
nand U22230 (N_22230,N_14913,N_15472);
and U22231 (N_22231,N_12591,N_14273);
nor U22232 (N_22232,N_17026,N_13470);
and U22233 (N_22233,N_14196,N_18037);
or U22234 (N_22234,N_13756,N_14052);
nor U22235 (N_22235,N_14520,N_15559);
or U22236 (N_22236,N_16901,N_15423);
or U22237 (N_22237,N_14765,N_17249);
or U22238 (N_22238,N_13374,N_18380);
and U22239 (N_22239,N_14172,N_14811);
nor U22240 (N_22240,N_18720,N_16044);
nor U22241 (N_22241,N_18007,N_14874);
xnor U22242 (N_22242,N_13911,N_13490);
or U22243 (N_22243,N_16897,N_15779);
nand U22244 (N_22244,N_17871,N_16988);
nor U22245 (N_22245,N_14259,N_13964);
xor U22246 (N_22246,N_16201,N_12542);
and U22247 (N_22247,N_18545,N_17849);
nor U22248 (N_22248,N_17195,N_17776);
nand U22249 (N_22249,N_12757,N_14724);
and U22250 (N_22250,N_14201,N_18433);
xnor U22251 (N_22251,N_17134,N_16800);
nand U22252 (N_22252,N_15043,N_16583);
nor U22253 (N_22253,N_14784,N_16178);
or U22254 (N_22254,N_18401,N_15904);
and U22255 (N_22255,N_12711,N_16117);
nor U22256 (N_22256,N_12670,N_13003);
and U22257 (N_22257,N_13473,N_17096);
nor U22258 (N_22258,N_14967,N_16400);
nor U22259 (N_22259,N_18134,N_15681);
xnor U22260 (N_22260,N_15607,N_17820);
or U22261 (N_22261,N_14058,N_12982);
nor U22262 (N_22262,N_15403,N_12939);
xor U22263 (N_22263,N_13468,N_14741);
and U22264 (N_22264,N_14851,N_15520);
or U22265 (N_22265,N_16528,N_18730);
nor U22266 (N_22266,N_18309,N_12869);
nor U22267 (N_22267,N_13677,N_14373);
or U22268 (N_22268,N_14113,N_14161);
and U22269 (N_22269,N_18425,N_12968);
and U22270 (N_22270,N_18465,N_17751);
and U22271 (N_22271,N_15672,N_15400);
nor U22272 (N_22272,N_18218,N_16515);
and U22273 (N_22273,N_16727,N_15980);
and U22274 (N_22274,N_17126,N_14276);
xor U22275 (N_22275,N_12588,N_18653);
and U22276 (N_22276,N_15254,N_12713);
and U22277 (N_22277,N_16803,N_14320);
xnor U22278 (N_22278,N_14497,N_15262);
and U22279 (N_22279,N_13586,N_17369);
and U22280 (N_22280,N_16636,N_17719);
xnor U22281 (N_22281,N_17658,N_15294);
and U22282 (N_22282,N_15266,N_18362);
and U22283 (N_22283,N_13706,N_12692);
xor U22284 (N_22284,N_14777,N_15960);
and U22285 (N_22285,N_16237,N_18582);
nor U22286 (N_22286,N_16837,N_15128);
nor U22287 (N_22287,N_13955,N_15603);
and U22288 (N_22288,N_17778,N_12792);
and U22289 (N_22289,N_13110,N_18468);
or U22290 (N_22290,N_15882,N_18286);
or U22291 (N_22291,N_16458,N_14181);
nand U22292 (N_22292,N_13038,N_17274);
nor U22293 (N_22293,N_16877,N_14531);
xor U22294 (N_22294,N_14695,N_14388);
or U22295 (N_22295,N_13229,N_14503);
nand U22296 (N_22296,N_16449,N_17113);
and U22297 (N_22297,N_12726,N_15512);
nor U22298 (N_22298,N_18133,N_13545);
or U22299 (N_22299,N_12928,N_14781);
nand U22300 (N_22300,N_17514,N_17810);
nor U22301 (N_22301,N_17327,N_12662);
xnor U22302 (N_22302,N_16810,N_13407);
or U22303 (N_22303,N_12531,N_17103);
nand U22304 (N_22304,N_17091,N_17558);
nor U22305 (N_22305,N_15228,N_12782);
xor U22306 (N_22306,N_13811,N_15806);
nor U22307 (N_22307,N_18384,N_18278);
or U22308 (N_22308,N_17907,N_17190);
and U22309 (N_22309,N_16594,N_17595);
nand U22310 (N_22310,N_13327,N_13207);
nand U22311 (N_22311,N_16677,N_18400);
xor U22312 (N_22312,N_15669,N_18631);
xnor U22313 (N_22313,N_18592,N_16215);
nor U22314 (N_22314,N_15634,N_13959);
or U22315 (N_22315,N_17904,N_17471);
nand U22316 (N_22316,N_15500,N_15878);
xor U22317 (N_22317,N_13758,N_16599);
nor U22318 (N_22318,N_17860,N_13907);
and U22319 (N_22319,N_12724,N_17643);
nor U22320 (N_22320,N_12874,N_15443);
or U22321 (N_22321,N_16657,N_18160);
nand U22322 (N_22322,N_17411,N_14564);
nand U22323 (N_22323,N_16087,N_18464);
and U22324 (N_22324,N_12972,N_16899);
xor U22325 (N_22325,N_14970,N_17401);
or U22326 (N_22326,N_16376,N_17763);
xnor U22327 (N_22327,N_13589,N_17824);
nor U22328 (N_22328,N_16905,N_16042);
and U22329 (N_22329,N_13830,N_15112);
nand U22330 (N_22330,N_16877,N_17146);
or U22331 (N_22331,N_17709,N_16276);
nand U22332 (N_22332,N_12967,N_18095);
and U22333 (N_22333,N_14426,N_16118);
or U22334 (N_22334,N_18628,N_16827);
nor U22335 (N_22335,N_14535,N_13703);
nand U22336 (N_22336,N_13091,N_13431);
nor U22337 (N_22337,N_13377,N_18332);
nor U22338 (N_22338,N_18606,N_13936);
and U22339 (N_22339,N_17527,N_18711);
nand U22340 (N_22340,N_16971,N_17055);
and U22341 (N_22341,N_15631,N_15487);
nor U22342 (N_22342,N_14440,N_17752);
and U22343 (N_22343,N_13796,N_13798);
nand U22344 (N_22344,N_13588,N_14459);
xor U22345 (N_22345,N_12567,N_18674);
xor U22346 (N_22346,N_15520,N_18101);
xnor U22347 (N_22347,N_18380,N_16841);
or U22348 (N_22348,N_17273,N_13552);
nand U22349 (N_22349,N_13488,N_12585);
and U22350 (N_22350,N_18585,N_12696);
or U22351 (N_22351,N_14437,N_16637);
nor U22352 (N_22352,N_12598,N_12642);
nand U22353 (N_22353,N_15565,N_15773);
nor U22354 (N_22354,N_18082,N_16477);
nor U22355 (N_22355,N_16789,N_16982);
and U22356 (N_22356,N_14781,N_12796);
nor U22357 (N_22357,N_16509,N_12677);
nor U22358 (N_22358,N_16641,N_15284);
nand U22359 (N_22359,N_15090,N_14855);
nand U22360 (N_22360,N_14778,N_15715);
or U22361 (N_22361,N_16566,N_16171);
nor U22362 (N_22362,N_17555,N_18216);
nor U22363 (N_22363,N_12866,N_16471);
nor U22364 (N_22364,N_16615,N_14598);
nand U22365 (N_22365,N_17715,N_18594);
nor U22366 (N_22366,N_15994,N_15264);
xnor U22367 (N_22367,N_13770,N_13764);
nand U22368 (N_22368,N_18425,N_13962);
or U22369 (N_22369,N_17427,N_17209);
nor U22370 (N_22370,N_17390,N_17027);
xnor U22371 (N_22371,N_12796,N_16370);
nor U22372 (N_22372,N_14132,N_13457);
and U22373 (N_22373,N_15030,N_18679);
and U22374 (N_22374,N_17144,N_15608);
nor U22375 (N_22375,N_13236,N_16675);
nand U22376 (N_22376,N_12866,N_18689);
or U22377 (N_22377,N_13925,N_13584);
or U22378 (N_22378,N_17849,N_16481);
nand U22379 (N_22379,N_15042,N_13133);
or U22380 (N_22380,N_14570,N_12951);
or U22381 (N_22381,N_14624,N_17133);
xor U22382 (N_22382,N_15996,N_15347);
nor U22383 (N_22383,N_14719,N_14382);
or U22384 (N_22384,N_17225,N_18329);
and U22385 (N_22385,N_13672,N_18021);
or U22386 (N_22386,N_16448,N_16077);
nor U22387 (N_22387,N_15115,N_15644);
or U22388 (N_22388,N_16605,N_15998);
nand U22389 (N_22389,N_14425,N_12662);
nor U22390 (N_22390,N_13323,N_17963);
nand U22391 (N_22391,N_18639,N_15888);
nor U22392 (N_22392,N_14013,N_17809);
nor U22393 (N_22393,N_17361,N_14321);
nand U22394 (N_22394,N_13374,N_16186);
nand U22395 (N_22395,N_18312,N_15873);
nor U22396 (N_22396,N_18126,N_14965);
or U22397 (N_22397,N_13683,N_16102);
nor U22398 (N_22398,N_18332,N_17453);
nand U22399 (N_22399,N_12806,N_16777);
nand U22400 (N_22400,N_13065,N_13569);
nand U22401 (N_22401,N_12999,N_18693);
or U22402 (N_22402,N_16051,N_16745);
and U22403 (N_22403,N_17816,N_13392);
nand U22404 (N_22404,N_14790,N_18201);
and U22405 (N_22405,N_17050,N_13539);
or U22406 (N_22406,N_17345,N_18667);
and U22407 (N_22407,N_17803,N_17335);
or U22408 (N_22408,N_12856,N_12832);
or U22409 (N_22409,N_14741,N_17766);
nand U22410 (N_22410,N_17349,N_15501);
and U22411 (N_22411,N_14146,N_17414);
nand U22412 (N_22412,N_16478,N_15097);
nand U22413 (N_22413,N_17627,N_18653);
nand U22414 (N_22414,N_18519,N_18365);
and U22415 (N_22415,N_12613,N_18114);
or U22416 (N_22416,N_15911,N_14546);
or U22417 (N_22417,N_18525,N_12962);
nand U22418 (N_22418,N_15505,N_13745);
xnor U22419 (N_22419,N_16027,N_15459);
and U22420 (N_22420,N_18193,N_15563);
nand U22421 (N_22421,N_15133,N_15056);
and U22422 (N_22422,N_16818,N_13733);
or U22423 (N_22423,N_16416,N_13021);
or U22424 (N_22424,N_16623,N_16434);
and U22425 (N_22425,N_14737,N_17419);
and U22426 (N_22426,N_16024,N_18353);
nand U22427 (N_22427,N_13919,N_16535);
and U22428 (N_22428,N_13430,N_16778);
nor U22429 (N_22429,N_15193,N_18415);
xor U22430 (N_22430,N_18189,N_14255);
nor U22431 (N_22431,N_15091,N_18204);
nand U22432 (N_22432,N_13026,N_16895);
or U22433 (N_22433,N_12847,N_18519);
or U22434 (N_22434,N_14321,N_17031);
nor U22435 (N_22435,N_18362,N_12781);
nor U22436 (N_22436,N_18280,N_15847);
or U22437 (N_22437,N_17626,N_16698);
or U22438 (N_22438,N_17522,N_12954);
xor U22439 (N_22439,N_18280,N_13066);
and U22440 (N_22440,N_18228,N_15725);
nand U22441 (N_22441,N_18463,N_15084);
nand U22442 (N_22442,N_12964,N_16997);
nor U22443 (N_22443,N_17013,N_17257);
or U22444 (N_22444,N_17248,N_17800);
or U22445 (N_22445,N_15689,N_14537);
nand U22446 (N_22446,N_12785,N_17994);
and U22447 (N_22447,N_18321,N_16024);
nand U22448 (N_22448,N_16224,N_14492);
nor U22449 (N_22449,N_17136,N_17702);
xnor U22450 (N_22450,N_17708,N_17816);
nor U22451 (N_22451,N_13870,N_15655);
and U22452 (N_22452,N_13120,N_16469);
and U22453 (N_22453,N_17275,N_16805);
xnor U22454 (N_22454,N_13394,N_13514);
or U22455 (N_22455,N_15018,N_17065);
nor U22456 (N_22456,N_14935,N_13572);
nand U22457 (N_22457,N_15827,N_18424);
nor U22458 (N_22458,N_12874,N_13964);
and U22459 (N_22459,N_16800,N_13526);
nor U22460 (N_22460,N_17201,N_13168);
or U22461 (N_22461,N_13554,N_13421);
nor U22462 (N_22462,N_18008,N_17583);
or U22463 (N_22463,N_12880,N_14313);
or U22464 (N_22464,N_15606,N_12946);
and U22465 (N_22465,N_16417,N_17581);
xnor U22466 (N_22466,N_18345,N_18141);
and U22467 (N_22467,N_14332,N_15380);
and U22468 (N_22468,N_17315,N_16147);
and U22469 (N_22469,N_18677,N_13495);
or U22470 (N_22470,N_12708,N_14611);
or U22471 (N_22471,N_16178,N_18321);
nor U22472 (N_22472,N_12505,N_13442);
or U22473 (N_22473,N_16102,N_14155);
nor U22474 (N_22474,N_18475,N_13107);
or U22475 (N_22475,N_14235,N_14603);
and U22476 (N_22476,N_16280,N_14335);
nor U22477 (N_22477,N_17204,N_16834);
xor U22478 (N_22478,N_14946,N_14001);
nand U22479 (N_22479,N_18330,N_14820);
and U22480 (N_22480,N_18408,N_15246);
nor U22481 (N_22481,N_18040,N_17001);
and U22482 (N_22482,N_15988,N_14609);
or U22483 (N_22483,N_18717,N_15861);
nand U22484 (N_22484,N_17040,N_17659);
and U22485 (N_22485,N_14926,N_12693);
and U22486 (N_22486,N_18349,N_12989);
and U22487 (N_22487,N_18585,N_14659);
xnor U22488 (N_22488,N_18183,N_15581);
nand U22489 (N_22489,N_16837,N_14341);
or U22490 (N_22490,N_17596,N_17247);
or U22491 (N_22491,N_13664,N_13852);
and U22492 (N_22492,N_18290,N_14428);
or U22493 (N_22493,N_13171,N_14403);
nand U22494 (N_22494,N_14685,N_12853);
or U22495 (N_22495,N_18674,N_15386);
and U22496 (N_22496,N_17016,N_18652);
or U22497 (N_22497,N_15740,N_12525);
nor U22498 (N_22498,N_16040,N_18211);
nor U22499 (N_22499,N_14611,N_18394);
and U22500 (N_22500,N_18372,N_17168);
nand U22501 (N_22501,N_17350,N_14664);
and U22502 (N_22502,N_13643,N_16712);
nand U22503 (N_22503,N_16418,N_12776);
nand U22504 (N_22504,N_15689,N_13859);
and U22505 (N_22505,N_17459,N_13279);
nand U22506 (N_22506,N_15361,N_13959);
and U22507 (N_22507,N_14947,N_12961);
or U22508 (N_22508,N_15639,N_16519);
or U22509 (N_22509,N_13091,N_15449);
nor U22510 (N_22510,N_13232,N_13718);
nand U22511 (N_22511,N_14671,N_13492);
or U22512 (N_22512,N_18046,N_18385);
and U22513 (N_22513,N_12852,N_13903);
and U22514 (N_22514,N_17768,N_16961);
and U22515 (N_22515,N_15375,N_16102);
nand U22516 (N_22516,N_18607,N_15674);
and U22517 (N_22517,N_16088,N_13354);
xnor U22518 (N_22518,N_17514,N_16068);
or U22519 (N_22519,N_16544,N_17714);
nand U22520 (N_22520,N_15728,N_17540);
and U22521 (N_22521,N_15551,N_14534);
nor U22522 (N_22522,N_14092,N_14042);
or U22523 (N_22523,N_14361,N_14174);
nor U22524 (N_22524,N_14479,N_18532);
nand U22525 (N_22525,N_14169,N_15063);
nor U22526 (N_22526,N_12618,N_12779);
or U22527 (N_22527,N_16161,N_16290);
or U22528 (N_22528,N_15864,N_15597);
and U22529 (N_22529,N_13240,N_13531);
nor U22530 (N_22530,N_16006,N_14458);
nand U22531 (N_22531,N_12510,N_16187);
nand U22532 (N_22532,N_16293,N_18412);
nor U22533 (N_22533,N_15624,N_12676);
and U22534 (N_22534,N_18131,N_16835);
nand U22535 (N_22535,N_17803,N_17478);
or U22536 (N_22536,N_14207,N_12789);
or U22537 (N_22537,N_12762,N_14078);
nor U22538 (N_22538,N_13511,N_17539);
xnor U22539 (N_22539,N_16717,N_16368);
or U22540 (N_22540,N_14652,N_13412);
nor U22541 (N_22541,N_17519,N_16861);
nor U22542 (N_22542,N_14886,N_16982);
and U22543 (N_22543,N_15261,N_17687);
or U22544 (N_22544,N_17229,N_18145);
or U22545 (N_22545,N_12979,N_15316);
nand U22546 (N_22546,N_14617,N_13430);
or U22547 (N_22547,N_14961,N_18560);
nor U22548 (N_22548,N_12984,N_13044);
and U22549 (N_22549,N_18312,N_14755);
xor U22550 (N_22550,N_13677,N_16780);
xnor U22551 (N_22551,N_15029,N_17929);
or U22552 (N_22552,N_14467,N_14003);
nand U22553 (N_22553,N_17527,N_13830);
and U22554 (N_22554,N_17703,N_17581);
and U22555 (N_22555,N_16152,N_15421);
or U22556 (N_22556,N_12509,N_14260);
nand U22557 (N_22557,N_15868,N_17799);
and U22558 (N_22558,N_18215,N_15795);
nand U22559 (N_22559,N_12981,N_12563);
nand U22560 (N_22560,N_16888,N_18321);
nor U22561 (N_22561,N_13385,N_13266);
nand U22562 (N_22562,N_15036,N_13881);
nand U22563 (N_22563,N_14478,N_16964);
xnor U22564 (N_22564,N_13175,N_17981);
or U22565 (N_22565,N_17018,N_15020);
nand U22566 (N_22566,N_15291,N_17992);
nor U22567 (N_22567,N_18286,N_17050);
nor U22568 (N_22568,N_12552,N_14652);
nand U22569 (N_22569,N_15466,N_15979);
and U22570 (N_22570,N_12902,N_16713);
nand U22571 (N_22571,N_12610,N_18296);
xnor U22572 (N_22572,N_18389,N_17157);
nor U22573 (N_22573,N_16210,N_17603);
nand U22574 (N_22574,N_17957,N_17858);
xor U22575 (N_22575,N_13440,N_17932);
or U22576 (N_22576,N_16143,N_14685);
or U22577 (N_22577,N_13507,N_18270);
or U22578 (N_22578,N_14627,N_16621);
nor U22579 (N_22579,N_17832,N_13739);
or U22580 (N_22580,N_16201,N_17205);
xnor U22581 (N_22581,N_14045,N_13320);
and U22582 (N_22582,N_16582,N_14262);
and U22583 (N_22583,N_17243,N_13359);
nor U22584 (N_22584,N_13205,N_17596);
nor U22585 (N_22585,N_18672,N_14503);
or U22586 (N_22586,N_15434,N_12644);
and U22587 (N_22587,N_13498,N_13675);
or U22588 (N_22588,N_18498,N_14086);
or U22589 (N_22589,N_17802,N_12839);
or U22590 (N_22590,N_15929,N_18556);
nand U22591 (N_22591,N_14895,N_13193);
or U22592 (N_22592,N_16070,N_16372);
xnor U22593 (N_22593,N_16380,N_18396);
or U22594 (N_22594,N_14914,N_13027);
nand U22595 (N_22595,N_13993,N_18376);
nor U22596 (N_22596,N_14405,N_14554);
nand U22597 (N_22597,N_12892,N_14020);
nand U22598 (N_22598,N_17385,N_17740);
nand U22599 (N_22599,N_16131,N_15847);
and U22600 (N_22600,N_13763,N_16989);
and U22601 (N_22601,N_12538,N_16199);
xnor U22602 (N_22602,N_18230,N_17114);
xor U22603 (N_22603,N_16344,N_14778);
and U22604 (N_22604,N_15827,N_18096);
nor U22605 (N_22605,N_15397,N_13963);
nor U22606 (N_22606,N_17393,N_14764);
nor U22607 (N_22607,N_13429,N_16884);
nor U22608 (N_22608,N_16067,N_14972);
nand U22609 (N_22609,N_14499,N_16594);
nand U22610 (N_22610,N_16183,N_12827);
nand U22611 (N_22611,N_18218,N_14120);
or U22612 (N_22612,N_15374,N_14999);
nor U22613 (N_22613,N_17687,N_14618);
and U22614 (N_22614,N_18677,N_17443);
nand U22615 (N_22615,N_18260,N_14389);
or U22616 (N_22616,N_14729,N_13724);
or U22617 (N_22617,N_17033,N_16739);
nor U22618 (N_22618,N_18165,N_13883);
nand U22619 (N_22619,N_15364,N_13737);
nor U22620 (N_22620,N_13220,N_16333);
or U22621 (N_22621,N_12712,N_13678);
nand U22622 (N_22622,N_15310,N_16095);
or U22623 (N_22623,N_17639,N_13805);
xnor U22624 (N_22624,N_14324,N_13365);
xnor U22625 (N_22625,N_17394,N_17649);
nor U22626 (N_22626,N_14178,N_12580);
and U22627 (N_22627,N_15933,N_14648);
nor U22628 (N_22628,N_14793,N_12614);
nand U22629 (N_22629,N_12696,N_15722);
nor U22630 (N_22630,N_14462,N_18502);
xnor U22631 (N_22631,N_17773,N_14299);
or U22632 (N_22632,N_16730,N_15025);
nor U22633 (N_22633,N_12963,N_13712);
nor U22634 (N_22634,N_18271,N_17377);
or U22635 (N_22635,N_12863,N_15631);
nand U22636 (N_22636,N_16414,N_14922);
or U22637 (N_22637,N_12587,N_13044);
xor U22638 (N_22638,N_15410,N_13848);
and U22639 (N_22639,N_13883,N_17604);
or U22640 (N_22640,N_13348,N_15950);
nor U22641 (N_22641,N_15280,N_13989);
and U22642 (N_22642,N_17574,N_16205);
nor U22643 (N_22643,N_17454,N_16495);
nand U22644 (N_22644,N_16191,N_16074);
nor U22645 (N_22645,N_15029,N_13710);
nand U22646 (N_22646,N_18576,N_14338);
nor U22647 (N_22647,N_18378,N_15528);
xnor U22648 (N_22648,N_16682,N_14792);
or U22649 (N_22649,N_14691,N_16344);
and U22650 (N_22650,N_15039,N_13824);
or U22651 (N_22651,N_18176,N_15309);
and U22652 (N_22652,N_17341,N_14395);
nand U22653 (N_22653,N_16913,N_14297);
or U22654 (N_22654,N_15927,N_14839);
and U22655 (N_22655,N_15483,N_12927);
and U22656 (N_22656,N_14572,N_16603);
and U22657 (N_22657,N_15532,N_17390);
or U22658 (N_22658,N_17402,N_15499);
and U22659 (N_22659,N_16793,N_17406);
nor U22660 (N_22660,N_16942,N_18312);
nor U22661 (N_22661,N_18147,N_16047);
nand U22662 (N_22662,N_12826,N_15738);
and U22663 (N_22663,N_17020,N_14518);
nor U22664 (N_22664,N_15779,N_17369);
nand U22665 (N_22665,N_17821,N_17843);
xor U22666 (N_22666,N_13134,N_15545);
xnor U22667 (N_22667,N_14475,N_12995);
nand U22668 (N_22668,N_17688,N_12610);
nor U22669 (N_22669,N_12827,N_12622);
nor U22670 (N_22670,N_12533,N_18445);
or U22671 (N_22671,N_16618,N_14497);
xnor U22672 (N_22672,N_16161,N_15943);
and U22673 (N_22673,N_18063,N_12806);
xnor U22674 (N_22674,N_16517,N_16454);
nor U22675 (N_22675,N_16663,N_15335);
nor U22676 (N_22676,N_12612,N_15618);
and U22677 (N_22677,N_16616,N_16234);
nand U22678 (N_22678,N_17506,N_18345);
and U22679 (N_22679,N_14957,N_18504);
nor U22680 (N_22680,N_16269,N_13053);
or U22681 (N_22681,N_17094,N_16009);
and U22682 (N_22682,N_16519,N_14956);
and U22683 (N_22683,N_13629,N_17285);
and U22684 (N_22684,N_18747,N_17847);
and U22685 (N_22685,N_17307,N_17433);
nand U22686 (N_22686,N_17116,N_17142);
nand U22687 (N_22687,N_15648,N_17028);
nor U22688 (N_22688,N_17675,N_14566);
nor U22689 (N_22689,N_13973,N_12788);
and U22690 (N_22690,N_14679,N_15954);
or U22691 (N_22691,N_16925,N_13059);
or U22692 (N_22692,N_12665,N_16068);
and U22693 (N_22693,N_12965,N_12654);
nand U22694 (N_22694,N_18464,N_17991);
xnor U22695 (N_22695,N_14723,N_16196);
nand U22696 (N_22696,N_16185,N_18308);
or U22697 (N_22697,N_17377,N_14651);
xor U22698 (N_22698,N_14632,N_16161);
xnor U22699 (N_22699,N_14851,N_15717);
nor U22700 (N_22700,N_18572,N_14234);
and U22701 (N_22701,N_13785,N_17857);
and U22702 (N_22702,N_18643,N_18669);
nand U22703 (N_22703,N_17432,N_13622);
and U22704 (N_22704,N_15895,N_17857);
and U22705 (N_22705,N_18719,N_15793);
and U22706 (N_22706,N_16810,N_16216);
nand U22707 (N_22707,N_17798,N_16617);
xnor U22708 (N_22708,N_14571,N_18522);
nor U22709 (N_22709,N_15226,N_13245);
nand U22710 (N_22710,N_12547,N_15361);
and U22711 (N_22711,N_17405,N_14075);
nand U22712 (N_22712,N_18626,N_13065);
and U22713 (N_22713,N_16278,N_14708);
or U22714 (N_22714,N_14197,N_15850);
and U22715 (N_22715,N_17087,N_14074);
nand U22716 (N_22716,N_13480,N_15812);
and U22717 (N_22717,N_14515,N_17518);
or U22718 (N_22718,N_13928,N_17854);
or U22719 (N_22719,N_13361,N_17477);
nor U22720 (N_22720,N_17645,N_13747);
or U22721 (N_22721,N_17775,N_14202);
nor U22722 (N_22722,N_14215,N_18183);
or U22723 (N_22723,N_18556,N_17747);
nor U22724 (N_22724,N_15447,N_18708);
or U22725 (N_22725,N_18071,N_17094);
or U22726 (N_22726,N_15561,N_13866);
nand U22727 (N_22727,N_14225,N_14825);
and U22728 (N_22728,N_15268,N_16193);
or U22729 (N_22729,N_13349,N_14787);
or U22730 (N_22730,N_14726,N_16300);
or U22731 (N_22731,N_15190,N_12786);
nor U22732 (N_22732,N_16956,N_14693);
nor U22733 (N_22733,N_13798,N_17003);
nor U22734 (N_22734,N_17580,N_14625);
and U22735 (N_22735,N_18367,N_18062);
nand U22736 (N_22736,N_14993,N_12555);
or U22737 (N_22737,N_17646,N_15101);
nor U22738 (N_22738,N_15193,N_15882);
and U22739 (N_22739,N_12727,N_16777);
nand U22740 (N_22740,N_12806,N_17017);
nor U22741 (N_22741,N_14774,N_17640);
nor U22742 (N_22742,N_14724,N_13745);
nor U22743 (N_22743,N_17646,N_17141);
nor U22744 (N_22744,N_18524,N_15725);
xnor U22745 (N_22745,N_14214,N_17305);
or U22746 (N_22746,N_15767,N_16950);
nor U22747 (N_22747,N_17857,N_14551);
or U22748 (N_22748,N_16098,N_15527);
and U22749 (N_22749,N_13045,N_17666);
nand U22750 (N_22750,N_18379,N_12779);
nand U22751 (N_22751,N_15990,N_13646);
and U22752 (N_22752,N_18311,N_17172);
or U22753 (N_22753,N_18699,N_14892);
or U22754 (N_22754,N_15727,N_18001);
nand U22755 (N_22755,N_15613,N_14853);
nor U22756 (N_22756,N_17092,N_15171);
nand U22757 (N_22757,N_18252,N_12520);
nand U22758 (N_22758,N_13974,N_17331);
and U22759 (N_22759,N_17693,N_18105);
and U22760 (N_22760,N_15314,N_14555);
and U22761 (N_22761,N_17202,N_17606);
and U22762 (N_22762,N_15448,N_15429);
nand U22763 (N_22763,N_15193,N_17232);
nor U22764 (N_22764,N_17740,N_17005);
or U22765 (N_22765,N_14448,N_14828);
and U22766 (N_22766,N_15412,N_18153);
or U22767 (N_22767,N_16520,N_15285);
or U22768 (N_22768,N_17678,N_14042);
nor U22769 (N_22769,N_12901,N_16842);
nor U22770 (N_22770,N_16627,N_17250);
xnor U22771 (N_22771,N_14855,N_13000);
and U22772 (N_22772,N_17132,N_13332);
and U22773 (N_22773,N_13433,N_17343);
nand U22774 (N_22774,N_16307,N_18082);
nor U22775 (N_22775,N_14137,N_13405);
or U22776 (N_22776,N_16274,N_18279);
and U22777 (N_22777,N_13524,N_17703);
nand U22778 (N_22778,N_15898,N_17431);
nor U22779 (N_22779,N_16097,N_13415);
or U22780 (N_22780,N_15591,N_16376);
and U22781 (N_22781,N_18298,N_14259);
and U22782 (N_22782,N_16627,N_14729);
nand U22783 (N_22783,N_15201,N_14267);
or U22784 (N_22784,N_13129,N_18174);
nand U22785 (N_22785,N_17284,N_12806);
nand U22786 (N_22786,N_15239,N_16362);
nand U22787 (N_22787,N_18459,N_17829);
and U22788 (N_22788,N_14901,N_13611);
or U22789 (N_22789,N_13233,N_17544);
nor U22790 (N_22790,N_17480,N_15685);
and U22791 (N_22791,N_14993,N_14182);
nor U22792 (N_22792,N_18445,N_15666);
nand U22793 (N_22793,N_18473,N_14089);
and U22794 (N_22794,N_16512,N_18307);
xnor U22795 (N_22795,N_12900,N_18048);
nand U22796 (N_22796,N_14849,N_17693);
or U22797 (N_22797,N_15127,N_17403);
nor U22798 (N_22798,N_15088,N_13572);
and U22799 (N_22799,N_13802,N_17106);
or U22800 (N_22800,N_13103,N_17095);
nand U22801 (N_22801,N_13934,N_17979);
nor U22802 (N_22802,N_13192,N_14943);
xor U22803 (N_22803,N_17824,N_14767);
nor U22804 (N_22804,N_16988,N_15371);
nand U22805 (N_22805,N_17150,N_18042);
nor U22806 (N_22806,N_16031,N_13795);
or U22807 (N_22807,N_16077,N_17465);
xnor U22808 (N_22808,N_16815,N_15668);
nor U22809 (N_22809,N_16550,N_17817);
nor U22810 (N_22810,N_16495,N_17630);
xor U22811 (N_22811,N_13438,N_14714);
and U22812 (N_22812,N_13939,N_14404);
and U22813 (N_22813,N_13342,N_17862);
or U22814 (N_22814,N_18554,N_18180);
and U22815 (N_22815,N_16980,N_15022);
nor U22816 (N_22816,N_17238,N_17326);
xor U22817 (N_22817,N_17371,N_15085);
nor U22818 (N_22818,N_13028,N_15575);
nand U22819 (N_22819,N_15090,N_14984);
nand U22820 (N_22820,N_13047,N_18157);
nand U22821 (N_22821,N_16840,N_16382);
nor U22822 (N_22822,N_12933,N_14186);
xnor U22823 (N_22823,N_13158,N_12939);
and U22824 (N_22824,N_15443,N_14584);
nand U22825 (N_22825,N_13120,N_17590);
nor U22826 (N_22826,N_18265,N_18396);
nand U22827 (N_22827,N_14527,N_17559);
and U22828 (N_22828,N_12978,N_16057);
or U22829 (N_22829,N_15009,N_18177);
and U22830 (N_22830,N_14763,N_17780);
nand U22831 (N_22831,N_12772,N_16491);
and U22832 (N_22832,N_16299,N_13417);
nor U22833 (N_22833,N_15199,N_16019);
nand U22834 (N_22834,N_17947,N_14333);
nor U22835 (N_22835,N_13937,N_13253);
nor U22836 (N_22836,N_18288,N_16360);
and U22837 (N_22837,N_14225,N_16907);
or U22838 (N_22838,N_16699,N_16242);
and U22839 (N_22839,N_16334,N_16733);
xnor U22840 (N_22840,N_16955,N_14431);
nor U22841 (N_22841,N_18504,N_18489);
and U22842 (N_22842,N_17347,N_16368);
nand U22843 (N_22843,N_17650,N_17142);
and U22844 (N_22844,N_18590,N_16540);
and U22845 (N_22845,N_18656,N_14041);
and U22846 (N_22846,N_17259,N_18345);
and U22847 (N_22847,N_18663,N_17748);
nand U22848 (N_22848,N_14835,N_16536);
xor U22849 (N_22849,N_14029,N_13123);
and U22850 (N_22850,N_17836,N_17373);
nand U22851 (N_22851,N_14177,N_12782);
or U22852 (N_22852,N_14231,N_17586);
or U22853 (N_22853,N_14017,N_16274);
nor U22854 (N_22854,N_14859,N_12640);
nand U22855 (N_22855,N_17532,N_15519);
nor U22856 (N_22856,N_15882,N_18372);
and U22857 (N_22857,N_13683,N_15560);
or U22858 (N_22858,N_13696,N_13634);
or U22859 (N_22859,N_18330,N_16411);
xnor U22860 (N_22860,N_14990,N_16967);
nand U22861 (N_22861,N_18617,N_17217);
nor U22862 (N_22862,N_15970,N_17277);
nand U22863 (N_22863,N_15876,N_17823);
nand U22864 (N_22864,N_14438,N_15069);
or U22865 (N_22865,N_15910,N_13772);
nor U22866 (N_22866,N_18331,N_16063);
and U22867 (N_22867,N_17396,N_13478);
and U22868 (N_22868,N_17305,N_13860);
or U22869 (N_22869,N_14836,N_15251);
or U22870 (N_22870,N_17111,N_17952);
xnor U22871 (N_22871,N_15636,N_13521);
nand U22872 (N_22872,N_14534,N_17609);
nor U22873 (N_22873,N_15020,N_17502);
nor U22874 (N_22874,N_13438,N_16404);
and U22875 (N_22875,N_15109,N_14895);
nand U22876 (N_22876,N_14726,N_12742);
nor U22877 (N_22877,N_16416,N_14051);
nand U22878 (N_22878,N_12770,N_18461);
and U22879 (N_22879,N_18566,N_15469);
or U22880 (N_22880,N_17190,N_13010);
and U22881 (N_22881,N_14995,N_15228);
nand U22882 (N_22882,N_15694,N_13514);
nor U22883 (N_22883,N_17509,N_14893);
and U22884 (N_22884,N_15311,N_13172);
and U22885 (N_22885,N_12672,N_17449);
nand U22886 (N_22886,N_16520,N_13502);
or U22887 (N_22887,N_14382,N_16268);
or U22888 (N_22888,N_15138,N_13182);
nand U22889 (N_22889,N_18226,N_13969);
nand U22890 (N_22890,N_14786,N_13319);
nor U22891 (N_22891,N_17331,N_17277);
and U22892 (N_22892,N_14074,N_17753);
nand U22893 (N_22893,N_17467,N_16937);
xnor U22894 (N_22894,N_18661,N_13411);
nand U22895 (N_22895,N_14011,N_14397);
or U22896 (N_22896,N_13980,N_17206);
nor U22897 (N_22897,N_12802,N_14373);
nand U22898 (N_22898,N_15315,N_14169);
or U22899 (N_22899,N_13102,N_16680);
xor U22900 (N_22900,N_17218,N_16105);
and U22901 (N_22901,N_15861,N_14928);
and U22902 (N_22902,N_15904,N_14605);
and U22903 (N_22903,N_15705,N_14574);
nor U22904 (N_22904,N_13827,N_12779);
and U22905 (N_22905,N_17339,N_15388);
xor U22906 (N_22906,N_14423,N_17642);
nand U22907 (N_22907,N_13900,N_14577);
nor U22908 (N_22908,N_17360,N_13194);
nor U22909 (N_22909,N_16367,N_14267);
nand U22910 (N_22910,N_13247,N_12737);
nand U22911 (N_22911,N_14684,N_16607);
nand U22912 (N_22912,N_18255,N_15197);
and U22913 (N_22913,N_15921,N_14196);
and U22914 (N_22914,N_14371,N_16986);
nor U22915 (N_22915,N_14658,N_14396);
xnor U22916 (N_22916,N_14646,N_15419);
or U22917 (N_22917,N_12826,N_15763);
or U22918 (N_22918,N_16068,N_14059);
and U22919 (N_22919,N_13629,N_13392);
or U22920 (N_22920,N_16518,N_16384);
and U22921 (N_22921,N_14917,N_18389);
nor U22922 (N_22922,N_13456,N_18183);
nor U22923 (N_22923,N_13968,N_16804);
nand U22924 (N_22924,N_17717,N_13891);
nor U22925 (N_22925,N_17906,N_15570);
or U22926 (N_22926,N_18217,N_14998);
xnor U22927 (N_22927,N_15472,N_16363);
xnor U22928 (N_22928,N_14625,N_17057);
or U22929 (N_22929,N_13655,N_12822);
and U22930 (N_22930,N_13688,N_13027);
nor U22931 (N_22931,N_13838,N_17937);
or U22932 (N_22932,N_12585,N_12736);
and U22933 (N_22933,N_18643,N_12886);
or U22934 (N_22934,N_12661,N_13998);
nor U22935 (N_22935,N_13847,N_13987);
nand U22936 (N_22936,N_14323,N_13976);
or U22937 (N_22937,N_16256,N_16932);
and U22938 (N_22938,N_15721,N_18409);
or U22939 (N_22939,N_15743,N_18611);
or U22940 (N_22940,N_15538,N_15901);
nor U22941 (N_22941,N_15875,N_14423);
nor U22942 (N_22942,N_17322,N_15523);
and U22943 (N_22943,N_16730,N_13919);
and U22944 (N_22944,N_17571,N_15897);
or U22945 (N_22945,N_16494,N_15546);
xor U22946 (N_22946,N_15395,N_18460);
nor U22947 (N_22947,N_12958,N_16936);
nand U22948 (N_22948,N_12655,N_17856);
nand U22949 (N_22949,N_18252,N_14959);
or U22950 (N_22950,N_16662,N_18246);
or U22951 (N_22951,N_13827,N_15360);
and U22952 (N_22952,N_12741,N_15385);
or U22953 (N_22953,N_15435,N_14672);
nor U22954 (N_22954,N_16913,N_13263);
nand U22955 (N_22955,N_16112,N_15675);
and U22956 (N_22956,N_14311,N_13367);
nor U22957 (N_22957,N_17153,N_14820);
and U22958 (N_22958,N_18317,N_18445);
nand U22959 (N_22959,N_18553,N_13905);
nor U22960 (N_22960,N_17136,N_14188);
or U22961 (N_22961,N_13307,N_15624);
and U22962 (N_22962,N_13482,N_13195);
and U22963 (N_22963,N_16108,N_13297);
and U22964 (N_22964,N_17447,N_16867);
xnor U22965 (N_22965,N_14588,N_15495);
nand U22966 (N_22966,N_12771,N_13170);
nor U22967 (N_22967,N_12564,N_18667);
nor U22968 (N_22968,N_17680,N_16104);
nand U22969 (N_22969,N_14545,N_13804);
and U22970 (N_22970,N_14613,N_16667);
nand U22971 (N_22971,N_16384,N_16050);
nor U22972 (N_22972,N_17628,N_18535);
or U22973 (N_22973,N_12833,N_18693);
and U22974 (N_22974,N_16285,N_13913);
and U22975 (N_22975,N_17176,N_16481);
nand U22976 (N_22976,N_14975,N_16988);
nor U22977 (N_22977,N_13390,N_16746);
nor U22978 (N_22978,N_17579,N_18723);
nor U22979 (N_22979,N_16200,N_16855);
and U22980 (N_22980,N_18028,N_16180);
nand U22981 (N_22981,N_15472,N_14030);
nor U22982 (N_22982,N_14478,N_18576);
or U22983 (N_22983,N_16325,N_17387);
or U22984 (N_22984,N_17334,N_13972);
or U22985 (N_22985,N_18243,N_14680);
and U22986 (N_22986,N_15321,N_13219);
nand U22987 (N_22987,N_17558,N_18269);
or U22988 (N_22988,N_13546,N_16455);
or U22989 (N_22989,N_15970,N_18091);
or U22990 (N_22990,N_15611,N_17959);
xnor U22991 (N_22991,N_18417,N_16077);
nand U22992 (N_22992,N_14679,N_14386);
xnor U22993 (N_22993,N_13567,N_14152);
nand U22994 (N_22994,N_14688,N_13988);
and U22995 (N_22995,N_17833,N_14006);
or U22996 (N_22996,N_18277,N_16381);
and U22997 (N_22997,N_18666,N_13799);
or U22998 (N_22998,N_15692,N_13857);
nand U22999 (N_22999,N_18622,N_18083);
or U23000 (N_23000,N_14662,N_15748);
or U23001 (N_23001,N_18421,N_17752);
or U23002 (N_23002,N_14071,N_17487);
or U23003 (N_23003,N_17321,N_15770);
nand U23004 (N_23004,N_13770,N_17618);
or U23005 (N_23005,N_12586,N_14977);
nor U23006 (N_23006,N_14301,N_12570);
and U23007 (N_23007,N_16033,N_13374);
nor U23008 (N_23008,N_13259,N_18467);
nor U23009 (N_23009,N_18254,N_18398);
or U23010 (N_23010,N_16944,N_15690);
nand U23011 (N_23011,N_17842,N_15129);
nor U23012 (N_23012,N_16444,N_13603);
nor U23013 (N_23013,N_13437,N_17620);
and U23014 (N_23014,N_16153,N_14513);
or U23015 (N_23015,N_16589,N_16695);
nor U23016 (N_23016,N_16014,N_15867);
nand U23017 (N_23017,N_18004,N_14784);
or U23018 (N_23018,N_17897,N_14949);
nor U23019 (N_23019,N_14662,N_15893);
nand U23020 (N_23020,N_13936,N_15817);
nor U23021 (N_23021,N_13669,N_17124);
nor U23022 (N_23022,N_16167,N_16120);
or U23023 (N_23023,N_13838,N_15498);
nand U23024 (N_23024,N_15304,N_15175);
nand U23025 (N_23025,N_18187,N_14296);
xnor U23026 (N_23026,N_14065,N_15193);
nand U23027 (N_23027,N_16823,N_13016);
xnor U23028 (N_23028,N_17543,N_18148);
nor U23029 (N_23029,N_17162,N_14010);
nand U23030 (N_23030,N_13913,N_13140);
or U23031 (N_23031,N_14455,N_15071);
xor U23032 (N_23032,N_18552,N_13024);
nor U23033 (N_23033,N_17916,N_17074);
and U23034 (N_23034,N_14746,N_15297);
xnor U23035 (N_23035,N_15533,N_16426);
and U23036 (N_23036,N_16649,N_14481);
nor U23037 (N_23037,N_14603,N_18285);
nor U23038 (N_23038,N_17367,N_17806);
or U23039 (N_23039,N_18534,N_17729);
nand U23040 (N_23040,N_17514,N_17461);
or U23041 (N_23041,N_14495,N_16387);
or U23042 (N_23042,N_18150,N_15657);
and U23043 (N_23043,N_13252,N_15291);
nor U23044 (N_23044,N_14098,N_18244);
xor U23045 (N_23045,N_17063,N_15169);
xor U23046 (N_23046,N_17515,N_17162);
nand U23047 (N_23047,N_18656,N_18103);
and U23048 (N_23048,N_18014,N_13868);
and U23049 (N_23049,N_16625,N_18022);
and U23050 (N_23050,N_18149,N_12985);
and U23051 (N_23051,N_17850,N_14602);
nor U23052 (N_23052,N_15996,N_17118);
nor U23053 (N_23053,N_16804,N_16525);
nor U23054 (N_23054,N_18373,N_17032);
or U23055 (N_23055,N_15351,N_15997);
nor U23056 (N_23056,N_14666,N_14450);
nor U23057 (N_23057,N_17638,N_17767);
nor U23058 (N_23058,N_18088,N_13084);
nand U23059 (N_23059,N_15651,N_16145);
or U23060 (N_23060,N_17262,N_12623);
nor U23061 (N_23061,N_14819,N_12918);
or U23062 (N_23062,N_13817,N_12786);
nand U23063 (N_23063,N_14287,N_18349);
nand U23064 (N_23064,N_13600,N_17729);
and U23065 (N_23065,N_17419,N_16256);
or U23066 (N_23066,N_15226,N_14271);
or U23067 (N_23067,N_17859,N_14743);
and U23068 (N_23068,N_16592,N_13672);
and U23069 (N_23069,N_13785,N_12614);
nor U23070 (N_23070,N_16147,N_14049);
nand U23071 (N_23071,N_16686,N_15199);
nand U23072 (N_23072,N_15299,N_14448);
nand U23073 (N_23073,N_12752,N_18553);
nand U23074 (N_23074,N_16140,N_16107);
or U23075 (N_23075,N_17765,N_14124);
and U23076 (N_23076,N_18529,N_13819);
or U23077 (N_23077,N_15640,N_15302);
nand U23078 (N_23078,N_14264,N_16122);
nand U23079 (N_23079,N_17056,N_13925);
and U23080 (N_23080,N_16020,N_16880);
nand U23081 (N_23081,N_15809,N_16230);
and U23082 (N_23082,N_16325,N_18530);
nor U23083 (N_23083,N_13009,N_12975);
nor U23084 (N_23084,N_18456,N_14080);
or U23085 (N_23085,N_12986,N_13701);
and U23086 (N_23086,N_18397,N_17726);
nand U23087 (N_23087,N_15999,N_12718);
nand U23088 (N_23088,N_12557,N_18054);
xor U23089 (N_23089,N_14807,N_18634);
and U23090 (N_23090,N_17162,N_12891);
and U23091 (N_23091,N_13848,N_15840);
nor U23092 (N_23092,N_16224,N_12721);
or U23093 (N_23093,N_16014,N_12927);
nand U23094 (N_23094,N_15371,N_15333);
or U23095 (N_23095,N_15403,N_15328);
and U23096 (N_23096,N_15355,N_15079);
xnor U23097 (N_23097,N_13149,N_14319);
nand U23098 (N_23098,N_12658,N_13059);
or U23099 (N_23099,N_17032,N_16122);
xor U23100 (N_23100,N_17488,N_17295);
nor U23101 (N_23101,N_16867,N_17519);
nand U23102 (N_23102,N_16308,N_16552);
and U23103 (N_23103,N_15001,N_17757);
xnor U23104 (N_23104,N_14063,N_15307);
nor U23105 (N_23105,N_12585,N_14120);
and U23106 (N_23106,N_12714,N_17464);
or U23107 (N_23107,N_13333,N_14906);
nand U23108 (N_23108,N_14084,N_13080);
and U23109 (N_23109,N_14881,N_14607);
nor U23110 (N_23110,N_13435,N_13800);
and U23111 (N_23111,N_18239,N_17879);
xor U23112 (N_23112,N_18248,N_18650);
nand U23113 (N_23113,N_15556,N_14938);
and U23114 (N_23114,N_16172,N_17489);
and U23115 (N_23115,N_14215,N_12793);
and U23116 (N_23116,N_15577,N_18446);
and U23117 (N_23117,N_17786,N_16476);
and U23118 (N_23118,N_17880,N_17368);
or U23119 (N_23119,N_16977,N_12933);
xor U23120 (N_23120,N_12717,N_17753);
and U23121 (N_23121,N_12711,N_15188);
and U23122 (N_23122,N_13725,N_15195);
and U23123 (N_23123,N_18024,N_16152);
or U23124 (N_23124,N_13026,N_15857);
and U23125 (N_23125,N_16475,N_16404);
and U23126 (N_23126,N_18092,N_14191);
xor U23127 (N_23127,N_17407,N_14190);
nand U23128 (N_23128,N_16829,N_16307);
or U23129 (N_23129,N_17322,N_13490);
nor U23130 (N_23130,N_16860,N_14167);
xor U23131 (N_23131,N_16858,N_15023);
and U23132 (N_23132,N_13027,N_17517);
and U23133 (N_23133,N_18395,N_15934);
xor U23134 (N_23134,N_13571,N_16812);
nor U23135 (N_23135,N_14214,N_14356);
nand U23136 (N_23136,N_17212,N_18253);
and U23137 (N_23137,N_13387,N_12800);
nor U23138 (N_23138,N_17083,N_17960);
nand U23139 (N_23139,N_17946,N_17964);
and U23140 (N_23140,N_18380,N_15033);
or U23141 (N_23141,N_14248,N_16836);
or U23142 (N_23142,N_16949,N_12984);
or U23143 (N_23143,N_14854,N_12722);
or U23144 (N_23144,N_16911,N_18661);
xnor U23145 (N_23145,N_18392,N_15207);
nand U23146 (N_23146,N_14346,N_15160);
nor U23147 (N_23147,N_14392,N_12758);
nor U23148 (N_23148,N_17981,N_12738);
nand U23149 (N_23149,N_15056,N_12725);
or U23150 (N_23150,N_12590,N_18083);
and U23151 (N_23151,N_17958,N_17055);
and U23152 (N_23152,N_14264,N_17760);
nor U23153 (N_23153,N_17095,N_15383);
nor U23154 (N_23154,N_13390,N_17866);
nand U23155 (N_23155,N_15420,N_17250);
nor U23156 (N_23156,N_12632,N_18616);
nor U23157 (N_23157,N_16403,N_15147);
nand U23158 (N_23158,N_18608,N_16434);
or U23159 (N_23159,N_12726,N_18672);
nor U23160 (N_23160,N_15424,N_12779);
nor U23161 (N_23161,N_15029,N_14290);
nand U23162 (N_23162,N_15346,N_17759);
nand U23163 (N_23163,N_15044,N_17855);
nor U23164 (N_23164,N_16720,N_17954);
nand U23165 (N_23165,N_17102,N_15712);
nand U23166 (N_23166,N_14749,N_15222);
and U23167 (N_23167,N_14010,N_13392);
nor U23168 (N_23168,N_17818,N_14057);
and U23169 (N_23169,N_12564,N_15621);
or U23170 (N_23170,N_13368,N_12523);
or U23171 (N_23171,N_13569,N_15235);
nor U23172 (N_23172,N_13156,N_16869);
and U23173 (N_23173,N_17700,N_13351);
and U23174 (N_23174,N_17525,N_14467);
nor U23175 (N_23175,N_12606,N_15393);
xor U23176 (N_23176,N_15761,N_18638);
nor U23177 (N_23177,N_13987,N_14746);
nor U23178 (N_23178,N_18521,N_15162);
or U23179 (N_23179,N_15003,N_14110);
xor U23180 (N_23180,N_15427,N_13547);
and U23181 (N_23181,N_15127,N_17633);
and U23182 (N_23182,N_17140,N_13815);
nand U23183 (N_23183,N_13222,N_17702);
or U23184 (N_23184,N_18224,N_17357);
or U23185 (N_23185,N_14066,N_12748);
nor U23186 (N_23186,N_13347,N_16013);
nor U23187 (N_23187,N_16237,N_15083);
and U23188 (N_23188,N_13144,N_12769);
nand U23189 (N_23189,N_13378,N_16866);
nor U23190 (N_23190,N_13644,N_14740);
nor U23191 (N_23191,N_18495,N_15843);
and U23192 (N_23192,N_15889,N_15804);
nor U23193 (N_23193,N_15231,N_17560);
nor U23194 (N_23194,N_16426,N_15307);
nor U23195 (N_23195,N_15670,N_13384);
nand U23196 (N_23196,N_17108,N_14984);
nand U23197 (N_23197,N_17703,N_14638);
nand U23198 (N_23198,N_18446,N_15534);
or U23199 (N_23199,N_14525,N_12528);
and U23200 (N_23200,N_13103,N_14124);
xor U23201 (N_23201,N_16881,N_14629);
nand U23202 (N_23202,N_13100,N_17247);
or U23203 (N_23203,N_18413,N_16065);
or U23204 (N_23204,N_15537,N_16837);
and U23205 (N_23205,N_13304,N_16642);
nor U23206 (N_23206,N_17135,N_16197);
or U23207 (N_23207,N_16280,N_18170);
xor U23208 (N_23208,N_13231,N_18441);
or U23209 (N_23209,N_15712,N_15515);
or U23210 (N_23210,N_16165,N_14963);
nor U23211 (N_23211,N_14685,N_14469);
or U23212 (N_23212,N_17995,N_15257);
nand U23213 (N_23213,N_18077,N_16507);
xor U23214 (N_23214,N_14659,N_15598);
and U23215 (N_23215,N_16151,N_15705);
nor U23216 (N_23216,N_15023,N_18681);
nand U23217 (N_23217,N_16076,N_13774);
nand U23218 (N_23218,N_15037,N_16126);
and U23219 (N_23219,N_13784,N_16782);
or U23220 (N_23220,N_17187,N_17609);
and U23221 (N_23221,N_17198,N_17422);
nand U23222 (N_23222,N_18112,N_14480);
or U23223 (N_23223,N_17000,N_17597);
nor U23224 (N_23224,N_14840,N_13043);
or U23225 (N_23225,N_13553,N_16898);
nand U23226 (N_23226,N_14142,N_16587);
and U23227 (N_23227,N_17345,N_17968);
nor U23228 (N_23228,N_12901,N_16055);
nand U23229 (N_23229,N_18724,N_18477);
and U23230 (N_23230,N_17924,N_15832);
or U23231 (N_23231,N_14707,N_12706);
or U23232 (N_23232,N_15997,N_14677);
nor U23233 (N_23233,N_13219,N_14517);
and U23234 (N_23234,N_12681,N_13064);
and U23235 (N_23235,N_14702,N_18684);
nor U23236 (N_23236,N_14782,N_14350);
and U23237 (N_23237,N_16879,N_18183);
nor U23238 (N_23238,N_16377,N_13873);
nor U23239 (N_23239,N_17738,N_17111);
nor U23240 (N_23240,N_13345,N_18154);
xnor U23241 (N_23241,N_12721,N_15187);
or U23242 (N_23242,N_17442,N_15372);
nor U23243 (N_23243,N_15790,N_13467);
nand U23244 (N_23244,N_13560,N_13219);
or U23245 (N_23245,N_12613,N_12543);
nand U23246 (N_23246,N_17520,N_17262);
nand U23247 (N_23247,N_16496,N_17810);
nor U23248 (N_23248,N_15690,N_15139);
nand U23249 (N_23249,N_18375,N_16685);
and U23250 (N_23250,N_15320,N_17500);
and U23251 (N_23251,N_12958,N_14830);
or U23252 (N_23252,N_16767,N_13899);
and U23253 (N_23253,N_17360,N_14225);
or U23254 (N_23254,N_13811,N_17444);
nor U23255 (N_23255,N_12989,N_15890);
nor U23256 (N_23256,N_17150,N_14376);
or U23257 (N_23257,N_14077,N_14037);
or U23258 (N_23258,N_15646,N_12642);
and U23259 (N_23259,N_12806,N_16313);
and U23260 (N_23260,N_14303,N_14548);
or U23261 (N_23261,N_18692,N_13542);
nand U23262 (N_23262,N_13775,N_14141);
or U23263 (N_23263,N_18223,N_16665);
and U23264 (N_23264,N_15557,N_13651);
and U23265 (N_23265,N_15983,N_16042);
or U23266 (N_23266,N_13181,N_16566);
xnor U23267 (N_23267,N_16658,N_13012);
nand U23268 (N_23268,N_17082,N_14661);
and U23269 (N_23269,N_13991,N_14274);
nor U23270 (N_23270,N_14581,N_14393);
or U23271 (N_23271,N_17608,N_17613);
and U23272 (N_23272,N_18486,N_12536);
or U23273 (N_23273,N_17164,N_15963);
nor U23274 (N_23274,N_15066,N_13413);
and U23275 (N_23275,N_14613,N_13920);
nor U23276 (N_23276,N_14501,N_17225);
and U23277 (N_23277,N_12777,N_16422);
or U23278 (N_23278,N_12533,N_15654);
or U23279 (N_23279,N_17318,N_18308);
nor U23280 (N_23280,N_16189,N_13407);
xor U23281 (N_23281,N_15756,N_13706);
nor U23282 (N_23282,N_18086,N_17076);
nor U23283 (N_23283,N_12651,N_16854);
nand U23284 (N_23284,N_16107,N_16186);
nor U23285 (N_23285,N_17223,N_12700);
and U23286 (N_23286,N_12525,N_18241);
nand U23287 (N_23287,N_18076,N_12988);
nor U23288 (N_23288,N_14013,N_16057);
nor U23289 (N_23289,N_17656,N_18628);
xor U23290 (N_23290,N_14782,N_18473);
or U23291 (N_23291,N_13269,N_13886);
nand U23292 (N_23292,N_15628,N_17123);
and U23293 (N_23293,N_17909,N_14752);
nand U23294 (N_23294,N_16170,N_16304);
nor U23295 (N_23295,N_14617,N_14383);
or U23296 (N_23296,N_13468,N_12733);
xor U23297 (N_23297,N_12947,N_15272);
and U23298 (N_23298,N_16571,N_14147);
and U23299 (N_23299,N_16068,N_18108);
and U23300 (N_23300,N_16695,N_17299);
and U23301 (N_23301,N_13977,N_17900);
nand U23302 (N_23302,N_17133,N_16517);
and U23303 (N_23303,N_17025,N_14403);
or U23304 (N_23304,N_14601,N_18613);
nand U23305 (N_23305,N_15568,N_14106);
nand U23306 (N_23306,N_17695,N_15178);
nand U23307 (N_23307,N_16414,N_15596);
or U23308 (N_23308,N_13509,N_15207);
xnor U23309 (N_23309,N_16735,N_17342);
nand U23310 (N_23310,N_17260,N_15484);
xnor U23311 (N_23311,N_13596,N_17409);
and U23312 (N_23312,N_17111,N_13254);
and U23313 (N_23313,N_14088,N_13658);
nand U23314 (N_23314,N_16812,N_13719);
or U23315 (N_23315,N_12990,N_15615);
nor U23316 (N_23316,N_14538,N_14682);
nor U23317 (N_23317,N_17397,N_12676);
nor U23318 (N_23318,N_17054,N_14814);
and U23319 (N_23319,N_15708,N_14971);
or U23320 (N_23320,N_15653,N_16736);
or U23321 (N_23321,N_17093,N_17504);
and U23322 (N_23322,N_14123,N_14920);
and U23323 (N_23323,N_16538,N_17542);
and U23324 (N_23324,N_13403,N_14857);
nand U23325 (N_23325,N_14078,N_12504);
or U23326 (N_23326,N_17501,N_16422);
nand U23327 (N_23327,N_18196,N_12896);
and U23328 (N_23328,N_14528,N_17303);
nand U23329 (N_23329,N_16115,N_16975);
or U23330 (N_23330,N_13553,N_18172);
nor U23331 (N_23331,N_18065,N_17520);
nor U23332 (N_23332,N_17686,N_17781);
nand U23333 (N_23333,N_13572,N_14226);
nor U23334 (N_23334,N_16100,N_13170);
nor U23335 (N_23335,N_16188,N_16473);
and U23336 (N_23336,N_15888,N_13006);
nand U23337 (N_23337,N_14882,N_12698);
nor U23338 (N_23338,N_13591,N_13498);
nand U23339 (N_23339,N_13356,N_13442);
or U23340 (N_23340,N_13248,N_16031);
nor U23341 (N_23341,N_15455,N_12579);
nor U23342 (N_23342,N_13495,N_16792);
xnor U23343 (N_23343,N_12851,N_16663);
and U23344 (N_23344,N_15767,N_14576);
nand U23345 (N_23345,N_14767,N_12556);
xnor U23346 (N_23346,N_12955,N_17580);
xor U23347 (N_23347,N_14718,N_15427);
nand U23348 (N_23348,N_17950,N_15311);
nand U23349 (N_23349,N_17853,N_14930);
nor U23350 (N_23350,N_16223,N_12513);
nand U23351 (N_23351,N_13799,N_17459);
or U23352 (N_23352,N_13460,N_15506);
or U23353 (N_23353,N_17502,N_16889);
xnor U23354 (N_23354,N_13940,N_13585);
nand U23355 (N_23355,N_17892,N_13179);
nand U23356 (N_23356,N_16029,N_17085);
nor U23357 (N_23357,N_13298,N_13183);
and U23358 (N_23358,N_12544,N_15461);
nand U23359 (N_23359,N_13955,N_15295);
or U23360 (N_23360,N_14793,N_12673);
or U23361 (N_23361,N_16887,N_18723);
nand U23362 (N_23362,N_16027,N_13939);
and U23363 (N_23363,N_15675,N_13590);
or U23364 (N_23364,N_13107,N_16678);
nand U23365 (N_23365,N_14918,N_18070);
xnor U23366 (N_23366,N_16525,N_13070);
xnor U23367 (N_23367,N_15037,N_15567);
nand U23368 (N_23368,N_14441,N_15541);
and U23369 (N_23369,N_16766,N_13288);
nand U23370 (N_23370,N_18316,N_18055);
and U23371 (N_23371,N_14541,N_16235);
xor U23372 (N_23372,N_16130,N_17830);
nor U23373 (N_23373,N_13358,N_15573);
and U23374 (N_23374,N_16687,N_13417);
xnor U23375 (N_23375,N_13283,N_14175);
nor U23376 (N_23376,N_18146,N_16437);
nand U23377 (N_23377,N_18133,N_17195);
and U23378 (N_23378,N_17275,N_12735);
or U23379 (N_23379,N_17376,N_16052);
or U23380 (N_23380,N_16685,N_16372);
nor U23381 (N_23381,N_16966,N_17013);
or U23382 (N_23382,N_18736,N_17087);
or U23383 (N_23383,N_14083,N_16690);
or U23384 (N_23384,N_13170,N_18521);
and U23385 (N_23385,N_14217,N_17211);
and U23386 (N_23386,N_18112,N_16884);
nor U23387 (N_23387,N_13850,N_16302);
nand U23388 (N_23388,N_16364,N_15049);
xnor U23389 (N_23389,N_16857,N_13838);
or U23390 (N_23390,N_17723,N_14179);
nor U23391 (N_23391,N_14880,N_12794);
nand U23392 (N_23392,N_17891,N_15485);
and U23393 (N_23393,N_17595,N_18472);
nor U23394 (N_23394,N_18713,N_17997);
nor U23395 (N_23395,N_14758,N_14800);
nor U23396 (N_23396,N_12574,N_14685);
or U23397 (N_23397,N_18243,N_16400);
nand U23398 (N_23398,N_18510,N_17363);
and U23399 (N_23399,N_12725,N_16873);
and U23400 (N_23400,N_18400,N_14754);
nand U23401 (N_23401,N_17722,N_16128);
nor U23402 (N_23402,N_12741,N_15925);
nor U23403 (N_23403,N_17051,N_18707);
and U23404 (N_23404,N_18740,N_18207);
and U23405 (N_23405,N_15313,N_17142);
xor U23406 (N_23406,N_17155,N_14516);
and U23407 (N_23407,N_16970,N_17159);
or U23408 (N_23408,N_15498,N_14752);
or U23409 (N_23409,N_17253,N_15984);
or U23410 (N_23410,N_17463,N_15521);
nor U23411 (N_23411,N_15332,N_18715);
nand U23412 (N_23412,N_12655,N_17777);
and U23413 (N_23413,N_14598,N_17594);
nor U23414 (N_23414,N_13204,N_14742);
or U23415 (N_23415,N_17162,N_12914);
or U23416 (N_23416,N_13421,N_18597);
nor U23417 (N_23417,N_12666,N_15040);
and U23418 (N_23418,N_14614,N_18593);
or U23419 (N_23419,N_17939,N_17528);
nand U23420 (N_23420,N_18612,N_17642);
or U23421 (N_23421,N_18363,N_14150);
and U23422 (N_23422,N_12748,N_14238);
nor U23423 (N_23423,N_13826,N_15391);
or U23424 (N_23424,N_18594,N_13280);
nor U23425 (N_23425,N_13220,N_15032);
nand U23426 (N_23426,N_13084,N_17903);
and U23427 (N_23427,N_16759,N_13002);
nand U23428 (N_23428,N_15660,N_14020);
or U23429 (N_23429,N_14473,N_14666);
nor U23430 (N_23430,N_18280,N_14401);
or U23431 (N_23431,N_17977,N_17726);
nor U23432 (N_23432,N_12732,N_18736);
or U23433 (N_23433,N_17268,N_12796);
or U23434 (N_23434,N_17158,N_15316);
nor U23435 (N_23435,N_18342,N_14999);
xor U23436 (N_23436,N_14315,N_15461);
and U23437 (N_23437,N_15875,N_12938);
xor U23438 (N_23438,N_17308,N_16377);
or U23439 (N_23439,N_14263,N_14430);
and U23440 (N_23440,N_16014,N_14964);
nor U23441 (N_23441,N_13546,N_15695);
and U23442 (N_23442,N_15320,N_14997);
nand U23443 (N_23443,N_16306,N_17312);
nor U23444 (N_23444,N_14106,N_16562);
and U23445 (N_23445,N_14111,N_15881);
nor U23446 (N_23446,N_13901,N_17017);
nor U23447 (N_23447,N_17677,N_13168);
nor U23448 (N_23448,N_18519,N_14781);
nand U23449 (N_23449,N_14865,N_17799);
nand U23450 (N_23450,N_15602,N_16388);
nand U23451 (N_23451,N_18348,N_18044);
nand U23452 (N_23452,N_15780,N_17865);
or U23453 (N_23453,N_13453,N_15644);
nor U23454 (N_23454,N_16002,N_16140);
nand U23455 (N_23455,N_14701,N_12876);
xnor U23456 (N_23456,N_14830,N_14726);
nor U23457 (N_23457,N_12955,N_17880);
xor U23458 (N_23458,N_13061,N_18573);
nor U23459 (N_23459,N_15235,N_15503);
or U23460 (N_23460,N_14737,N_16614);
nor U23461 (N_23461,N_16944,N_16495);
and U23462 (N_23462,N_14792,N_12585);
and U23463 (N_23463,N_13204,N_13006);
nor U23464 (N_23464,N_16262,N_14081);
nand U23465 (N_23465,N_12955,N_17676);
nand U23466 (N_23466,N_15833,N_15670);
nand U23467 (N_23467,N_15320,N_15773);
xnor U23468 (N_23468,N_15503,N_16758);
nor U23469 (N_23469,N_15841,N_12974);
and U23470 (N_23470,N_18547,N_12966);
nor U23471 (N_23471,N_14046,N_14742);
nand U23472 (N_23472,N_18529,N_16922);
or U23473 (N_23473,N_15308,N_14422);
nor U23474 (N_23474,N_12772,N_14481);
nand U23475 (N_23475,N_13212,N_13071);
and U23476 (N_23476,N_12686,N_12813);
and U23477 (N_23477,N_16102,N_14122);
nor U23478 (N_23478,N_16616,N_15390);
or U23479 (N_23479,N_12907,N_18627);
nor U23480 (N_23480,N_16289,N_13853);
or U23481 (N_23481,N_13813,N_17910);
nor U23482 (N_23482,N_15603,N_15669);
nor U23483 (N_23483,N_13777,N_18414);
or U23484 (N_23484,N_12889,N_13464);
nor U23485 (N_23485,N_15047,N_15272);
or U23486 (N_23486,N_12931,N_16292);
nand U23487 (N_23487,N_15653,N_18322);
nand U23488 (N_23488,N_17541,N_15993);
and U23489 (N_23489,N_15046,N_18747);
nor U23490 (N_23490,N_15597,N_12640);
and U23491 (N_23491,N_15632,N_12555);
nand U23492 (N_23492,N_13164,N_13236);
nand U23493 (N_23493,N_16354,N_15185);
and U23494 (N_23494,N_14654,N_14882);
or U23495 (N_23495,N_13138,N_17109);
nand U23496 (N_23496,N_16970,N_17348);
or U23497 (N_23497,N_15194,N_13731);
nand U23498 (N_23498,N_17359,N_16893);
and U23499 (N_23499,N_16777,N_12692);
xnor U23500 (N_23500,N_14441,N_17909);
xor U23501 (N_23501,N_12840,N_14305);
or U23502 (N_23502,N_16936,N_15018);
nor U23503 (N_23503,N_13979,N_16629);
nand U23504 (N_23504,N_18639,N_15474);
nor U23505 (N_23505,N_14509,N_14626);
or U23506 (N_23506,N_17743,N_16085);
nor U23507 (N_23507,N_13677,N_17019);
or U23508 (N_23508,N_16751,N_13407);
and U23509 (N_23509,N_15523,N_18271);
nand U23510 (N_23510,N_16171,N_13982);
nand U23511 (N_23511,N_12646,N_15370);
and U23512 (N_23512,N_16248,N_15269);
nor U23513 (N_23513,N_17985,N_16409);
or U23514 (N_23514,N_18546,N_17178);
nand U23515 (N_23515,N_16728,N_13798);
or U23516 (N_23516,N_12948,N_13256);
and U23517 (N_23517,N_18031,N_15285);
nor U23518 (N_23518,N_18151,N_15231);
and U23519 (N_23519,N_14736,N_18001);
nand U23520 (N_23520,N_13998,N_14213);
and U23521 (N_23521,N_17344,N_16367);
and U23522 (N_23522,N_16775,N_14384);
or U23523 (N_23523,N_13877,N_14521);
nand U23524 (N_23524,N_16003,N_14221);
xor U23525 (N_23525,N_13145,N_13125);
nor U23526 (N_23526,N_13471,N_14319);
nor U23527 (N_23527,N_16729,N_15589);
or U23528 (N_23528,N_16026,N_13853);
or U23529 (N_23529,N_17341,N_14632);
and U23530 (N_23530,N_15676,N_12576);
or U23531 (N_23531,N_17854,N_14297);
nand U23532 (N_23532,N_18443,N_15134);
xnor U23533 (N_23533,N_13594,N_12516);
nor U23534 (N_23534,N_18473,N_15610);
nand U23535 (N_23535,N_13344,N_17861);
or U23536 (N_23536,N_15198,N_16667);
xor U23537 (N_23537,N_16441,N_15031);
nor U23538 (N_23538,N_14340,N_17703);
xor U23539 (N_23539,N_14741,N_15455);
or U23540 (N_23540,N_17001,N_15995);
nand U23541 (N_23541,N_13118,N_15924);
or U23542 (N_23542,N_15106,N_17756);
nor U23543 (N_23543,N_17174,N_18023);
nor U23544 (N_23544,N_17405,N_12845);
nand U23545 (N_23545,N_18447,N_14423);
or U23546 (N_23546,N_13659,N_14337);
and U23547 (N_23547,N_17356,N_13998);
xor U23548 (N_23548,N_13563,N_13296);
and U23549 (N_23549,N_13420,N_12543);
nand U23550 (N_23550,N_17394,N_14135);
and U23551 (N_23551,N_13736,N_16800);
or U23552 (N_23552,N_12983,N_17380);
or U23553 (N_23553,N_14400,N_13312);
nand U23554 (N_23554,N_15051,N_17731);
nor U23555 (N_23555,N_13069,N_15185);
nand U23556 (N_23556,N_15814,N_14647);
nand U23557 (N_23557,N_15758,N_16780);
xor U23558 (N_23558,N_16953,N_16131);
nor U23559 (N_23559,N_16141,N_16160);
nand U23560 (N_23560,N_16793,N_14430);
nand U23561 (N_23561,N_13140,N_13822);
nor U23562 (N_23562,N_15609,N_14699);
nor U23563 (N_23563,N_14850,N_17477);
nand U23564 (N_23564,N_14642,N_13645);
nand U23565 (N_23565,N_18370,N_14477);
and U23566 (N_23566,N_16545,N_14711);
nor U23567 (N_23567,N_15240,N_17582);
or U23568 (N_23568,N_15223,N_15028);
nand U23569 (N_23569,N_15078,N_13276);
xor U23570 (N_23570,N_13585,N_18060);
nor U23571 (N_23571,N_16069,N_16070);
or U23572 (N_23572,N_18364,N_13377);
xnor U23573 (N_23573,N_14066,N_17630);
nand U23574 (N_23574,N_15232,N_16869);
and U23575 (N_23575,N_13917,N_17574);
or U23576 (N_23576,N_13297,N_14351);
and U23577 (N_23577,N_18002,N_15031);
nand U23578 (N_23578,N_17998,N_15161);
or U23579 (N_23579,N_16219,N_17062);
and U23580 (N_23580,N_17736,N_17465);
nor U23581 (N_23581,N_13617,N_16438);
xor U23582 (N_23582,N_16057,N_14506);
or U23583 (N_23583,N_15520,N_13354);
xor U23584 (N_23584,N_17330,N_13159);
and U23585 (N_23585,N_16529,N_15812);
xor U23586 (N_23586,N_13714,N_16280);
or U23587 (N_23587,N_13059,N_12717);
and U23588 (N_23588,N_16086,N_13632);
nand U23589 (N_23589,N_14922,N_13846);
nor U23590 (N_23590,N_17065,N_12772);
and U23591 (N_23591,N_16080,N_18399);
nand U23592 (N_23592,N_14282,N_14451);
nor U23593 (N_23593,N_18444,N_17651);
nor U23594 (N_23594,N_17456,N_13997);
or U23595 (N_23595,N_13371,N_16503);
and U23596 (N_23596,N_12927,N_18111);
xor U23597 (N_23597,N_17873,N_17255);
or U23598 (N_23598,N_15448,N_16106);
or U23599 (N_23599,N_17463,N_12687);
and U23600 (N_23600,N_17657,N_14985);
and U23601 (N_23601,N_12692,N_17585);
or U23602 (N_23602,N_17520,N_14063);
nor U23603 (N_23603,N_17666,N_18592);
nand U23604 (N_23604,N_12786,N_16893);
and U23605 (N_23605,N_15164,N_15256);
or U23606 (N_23606,N_16297,N_18337);
nand U23607 (N_23607,N_15770,N_17803);
nor U23608 (N_23608,N_14986,N_18522);
or U23609 (N_23609,N_15269,N_18415);
nor U23610 (N_23610,N_16186,N_16056);
and U23611 (N_23611,N_17273,N_15150);
nand U23612 (N_23612,N_15051,N_15856);
or U23613 (N_23613,N_14874,N_14345);
nor U23614 (N_23614,N_14755,N_18428);
nor U23615 (N_23615,N_17440,N_15731);
nand U23616 (N_23616,N_17051,N_12953);
nor U23617 (N_23617,N_14116,N_17888);
and U23618 (N_23618,N_15321,N_15895);
and U23619 (N_23619,N_15145,N_18637);
and U23620 (N_23620,N_14902,N_12967);
and U23621 (N_23621,N_16347,N_18280);
nor U23622 (N_23622,N_13669,N_17469);
nand U23623 (N_23623,N_18676,N_14044);
or U23624 (N_23624,N_16686,N_16557);
or U23625 (N_23625,N_18103,N_13967);
xor U23626 (N_23626,N_15243,N_17827);
and U23627 (N_23627,N_13283,N_14000);
and U23628 (N_23628,N_15794,N_17474);
and U23629 (N_23629,N_16360,N_16178);
xor U23630 (N_23630,N_15238,N_14092);
nor U23631 (N_23631,N_12619,N_15613);
and U23632 (N_23632,N_14911,N_17111);
xnor U23633 (N_23633,N_14541,N_15683);
nand U23634 (N_23634,N_14358,N_14367);
nand U23635 (N_23635,N_18634,N_13381);
xnor U23636 (N_23636,N_17110,N_13788);
and U23637 (N_23637,N_12933,N_18348);
nand U23638 (N_23638,N_13097,N_16526);
nand U23639 (N_23639,N_15076,N_14684);
and U23640 (N_23640,N_14310,N_18682);
or U23641 (N_23641,N_12890,N_18399);
nand U23642 (N_23642,N_15943,N_14641);
or U23643 (N_23643,N_16364,N_17217);
and U23644 (N_23644,N_15666,N_16398);
nand U23645 (N_23645,N_12870,N_18673);
or U23646 (N_23646,N_14514,N_17912);
nand U23647 (N_23647,N_17918,N_13213);
and U23648 (N_23648,N_13009,N_13693);
or U23649 (N_23649,N_14978,N_14966);
and U23650 (N_23650,N_12930,N_17340);
nor U23651 (N_23651,N_14234,N_15776);
nand U23652 (N_23652,N_15037,N_15406);
and U23653 (N_23653,N_15125,N_13432);
nand U23654 (N_23654,N_13413,N_15823);
nand U23655 (N_23655,N_13557,N_17026);
or U23656 (N_23656,N_18568,N_18546);
or U23657 (N_23657,N_14907,N_17102);
xor U23658 (N_23658,N_18050,N_13823);
nor U23659 (N_23659,N_16701,N_17489);
or U23660 (N_23660,N_14756,N_12752);
and U23661 (N_23661,N_14254,N_18363);
and U23662 (N_23662,N_14433,N_13143);
nor U23663 (N_23663,N_17055,N_17523);
xor U23664 (N_23664,N_17267,N_12588);
or U23665 (N_23665,N_17179,N_12672);
nand U23666 (N_23666,N_15481,N_18697);
or U23667 (N_23667,N_14475,N_16970);
nand U23668 (N_23668,N_13374,N_18309);
or U23669 (N_23669,N_12648,N_14753);
and U23670 (N_23670,N_13500,N_17931);
nand U23671 (N_23671,N_14398,N_14372);
xor U23672 (N_23672,N_13182,N_16896);
or U23673 (N_23673,N_13327,N_14144);
xnor U23674 (N_23674,N_18241,N_18743);
or U23675 (N_23675,N_15388,N_17513);
nand U23676 (N_23676,N_12542,N_17890);
xor U23677 (N_23677,N_14572,N_14279);
and U23678 (N_23678,N_12910,N_16523);
or U23679 (N_23679,N_15136,N_13644);
or U23680 (N_23680,N_15988,N_14872);
xor U23681 (N_23681,N_18451,N_17051);
or U23682 (N_23682,N_18663,N_14706);
xor U23683 (N_23683,N_18191,N_14102);
or U23684 (N_23684,N_16351,N_16099);
nand U23685 (N_23685,N_13606,N_17294);
nand U23686 (N_23686,N_15751,N_15494);
xnor U23687 (N_23687,N_16801,N_15065);
nand U23688 (N_23688,N_17352,N_18254);
nand U23689 (N_23689,N_16624,N_14151);
or U23690 (N_23690,N_16847,N_14365);
nand U23691 (N_23691,N_17158,N_15886);
nor U23692 (N_23692,N_17829,N_15257);
or U23693 (N_23693,N_18132,N_14628);
or U23694 (N_23694,N_15181,N_14414);
nand U23695 (N_23695,N_12868,N_18674);
and U23696 (N_23696,N_17517,N_12858);
and U23697 (N_23697,N_16396,N_13471);
nor U23698 (N_23698,N_13972,N_15386);
or U23699 (N_23699,N_16006,N_16192);
and U23700 (N_23700,N_16257,N_15255);
and U23701 (N_23701,N_14487,N_13053);
or U23702 (N_23702,N_15364,N_18134);
or U23703 (N_23703,N_14836,N_13014);
nor U23704 (N_23704,N_15846,N_12547);
and U23705 (N_23705,N_12556,N_14063);
or U23706 (N_23706,N_15184,N_13457);
or U23707 (N_23707,N_18577,N_14620);
nand U23708 (N_23708,N_16658,N_18740);
or U23709 (N_23709,N_17938,N_14005);
nand U23710 (N_23710,N_12833,N_12743);
nand U23711 (N_23711,N_15207,N_13185);
nor U23712 (N_23712,N_18077,N_16122);
and U23713 (N_23713,N_16942,N_13637);
and U23714 (N_23714,N_14871,N_13310);
nand U23715 (N_23715,N_18048,N_15066);
nor U23716 (N_23716,N_16973,N_16639);
nand U23717 (N_23717,N_12937,N_16545);
xnor U23718 (N_23718,N_18265,N_18223);
and U23719 (N_23719,N_17016,N_16874);
nand U23720 (N_23720,N_16732,N_16775);
nor U23721 (N_23721,N_14951,N_16591);
xnor U23722 (N_23722,N_13204,N_17572);
or U23723 (N_23723,N_12524,N_16248);
nor U23724 (N_23724,N_15141,N_12608);
and U23725 (N_23725,N_16124,N_16236);
and U23726 (N_23726,N_13002,N_14816);
xor U23727 (N_23727,N_15928,N_18039);
and U23728 (N_23728,N_15440,N_16790);
nand U23729 (N_23729,N_15850,N_13036);
and U23730 (N_23730,N_18636,N_15232);
and U23731 (N_23731,N_13421,N_15766);
nand U23732 (N_23732,N_16987,N_16845);
xor U23733 (N_23733,N_15330,N_15199);
nand U23734 (N_23734,N_14182,N_13123);
nor U23735 (N_23735,N_13425,N_15950);
or U23736 (N_23736,N_13085,N_12921);
xnor U23737 (N_23737,N_18036,N_13255);
and U23738 (N_23738,N_12888,N_16266);
xor U23739 (N_23739,N_13637,N_17741);
nand U23740 (N_23740,N_16848,N_15242);
or U23741 (N_23741,N_17464,N_13091);
or U23742 (N_23742,N_13962,N_18383);
nand U23743 (N_23743,N_16550,N_14671);
nor U23744 (N_23744,N_16883,N_18537);
and U23745 (N_23745,N_14098,N_15301);
nand U23746 (N_23746,N_16572,N_15415);
and U23747 (N_23747,N_18558,N_15699);
or U23748 (N_23748,N_14410,N_15613);
or U23749 (N_23749,N_12963,N_18310);
nand U23750 (N_23750,N_17974,N_13259);
nand U23751 (N_23751,N_12821,N_15713);
nor U23752 (N_23752,N_18353,N_18749);
and U23753 (N_23753,N_14084,N_16086);
and U23754 (N_23754,N_17877,N_17889);
and U23755 (N_23755,N_15049,N_18519);
or U23756 (N_23756,N_18118,N_13679);
or U23757 (N_23757,N_14661,N_18543);
nor U23758 (N_23758,N_16977,N_13092);
or U23759 (N_23759,N_13715,N_15453);
nand U23760 (N_23760,N_15060,N_13039);
nor U23761 (N_23761,N_12794,N_15450);
nand U23762 (N_23762,N_18575,N_13415);
nand U23763 (N_23763,N_14892,N_17816);
xor U23764 (N_23764,N_13322,N_15389);
nor U23765 (N_23765,N_15913,N_15866);
and U23766 (N_23766,N_13685,N_17077);
and U23767 (N_23767,N_16491,N_16812);
nor U23768 (N_23768,N_14523,N_18728);
xnor U23769 (N_23769,N_13507,N_14316);
xnor U23770 (N_23770,N_13470,N_16393);
nor U23771 (N_23771,N_13050,N_17739);
and U23772 (N_23772,N_12922,N_18179);
or U23773 (N_23773,N_13441,N_16281);
or U23774 (N_23774,N_16111,N_15122);
nor U23775 (N_23775,N_18264,N_14735);
nand U23776 (N_23776,N_14196,N_13992);
nor U23777 (N_23777,N_15818,N_12988);
nand U23778 (N_23778,N_12614,N_18497);
xor U23779 (N_23779,N_14669,N_16778);
or U23780 (N_23780,N_13827,N_13321);
and U23781 (N_23781,N_18419,N_18316);
xnor U23782 (N_23782,N_18497,N_17731);
nor U23783 (N_23783,N_17325,N_13470);
and U23784 (N_23784,N_14283,N_12949);
or U23785 (N_23785,N_14881,N_15574);
and U23786 (N_23786,N_18725,N_16707);
or U23787 (N_23787,N_14145,N_12667);
nand U23788 (N_23788,N_17412,N_18644);
and U23789 (N_23789,N_15286,N_13675);
nand U23790 (N_23790,N_18494,N_14549);
or U23791 (N_23791,N_15950,N_16881);
or U23792 (N_23792,N_16363,N_18404);
nand U23793 (N_23793,N_16100,N_14228);
nand U23794 (N_23794,N_17908,N_14665);
or U23795 (N_23795,N_13581,N_13234);
nor U23796 (N_23796,N_17083,N_13475);
or U23797 (N_23797,N_12833,N_12770);
and U23798 (N_23798,N_15062,N_16777);
nand U23799 (N_23799,N_16198,N_12716);
nand U23800 (N_23800,N_14522,N_17724);
nor U23801 (N_23801,N_14547,N_14955);
nor U23802 (N_23802,N_14951,N_15179);
nand U23803 (N_23803,N_15790,N_18027);
or U23804 (N_23804,N_15518,N_12843);
and U23805 (N_23805,N_13142,N_13808);
nand U23806 (N_23806,N_15647,N_18705);
and U23807 (N_23807,N_17049,N_13989);
or U23808 (N_23808,N_14474,N_12990);
nand U23809 (N_23809,N_12599,N_16993);
and U23810 (N_23810,N_17608,N_15464);
and U23811 (N_23811,N_14338,N_13899);
or U23812 (N_23812,N_14165,N_13025);
nand U23813 (N_23813,N_15670,N_14751);
xnor U23814 (N_23814,N_13873,N_17997);
nor U23815 (N_23815,N_16614,N_17033);
nand U23816 (N_23816,N_14852,N_13676);
or U23817 (N_23817,N_13044,N_12849);
nand U23818 (N_23818,N_17719,N_16753);
nor U23819 (N_23819,N_18308,N_16410);
and U23820 (N_23820,N_16462,N_18381);
and U23821 (N_23821,N_16658,N_13291);
nor U23822 (N_23822,N_15854,N_18151);
and U23823 (N_23823,N_16195,N_17763);
xnor U23824 (N_23824,N_13117,N_16792);
xor U23825 (N_23825,N_18164,N_18430);
or U23826 (N_23826,N_14582,N_12955);
nand U23827 (N_23827,N_18665,N_14831);
and U23828 (N_23828,N_17604,N_15567);
nand U23829 (N_23829,N_18154,N_17534);
and U23830 (N_23830,N_17978,N_15843);
nand U23831 (N_23831,N_18648,N_13555);
and U23832 (N_23832,N_16890,N_17865);
xor U23833 (N_23833,N_15929,N_15633);
nor U23834 (N_23834,N_13829,N_17927);
or U23835 (N_23835,N_14676,N_12906);
or U23836 (N_23836,N_14848,N_14677);
or U23837 (N_23837,N_18013,N_13472);
nor U23838 (N_23838,N_12576,N_18085);
nand U23839 (N_23839,N_15483,N_13787);
nor U23840 (N_23840,N_17010,N_16480);
and U23841 (N_23841,N_14681,N_15234);
nand U23842 (N_23842,N_13179,N_14566);
or U23843 (N_23843,N_13189,N_18108);
xor U23844 (N_23844,N_14806,N_15171);
nand U23845 (N_23845,N_15435,N_14162);
and U23846 (N_23846,N_16296,N_13279);
or U23847 (N_23847,N_13929,N_18471);
or U23848 (N_23848,N_16513,N_13371);
and U23849 (N_23849,N_17857,N_16462);
nand U23850 (N_23850,N_15869,N_14687);
xnor U23851 (N_23851,N_18556,N_12754);
nand U23852 (N_23852,N_16611,N_15823);
nand U23853 (N_23853,N_14302,N_13258);
and U23854 (N_23854,N_17511,N_12602);
or U23855 (N_23855,N_16318,N_16361);
nor U23856 (N_23856,N_14701,N_14877);
nand U23857 (N_23857,N_14318,N_13696);
xnor U23858 (N_23858,N_12850,N_15433);
nand U23859 (N_23859,N_13388,N_17211);
or U23860 (N_23860,N_18591,N_17283);
nand U23861 (N_23861,N_16943,N_17248);
and U23862 (N_23862,N_15527,N_17778);
nor U23863 (N_23863,N_17047,N_17846);
or U23864 (N_23864,N_17430,N_12829);
nand U23865 (N_23865,N_17502,N_13388);
or U23866 (N_23866,N_15012,N_17498);
nand U23867 (N_23867,N_16772,N_14399);
or U23868 (N_23868,N_18307,N_16019);
nand U23869 (N_23869,N_14314,N_14974);
nor U23870 (N_23870,N_16241,N_18231);
and U23871 (N_23871,N_13379,N_14399);
nand U23872 (N_23872,N_13796,N_14314);
nor U23873 (N_23873,N_15973,N_13645);
or U23874 (N_23874,N_14387,N_18144);
and U23875 (N_23875,N_15947,N_12672);
and U23876 (N_23876,N_16349,N_15296);
and U23877 (N_23877,N_15758,N_14664);
nor U23878 (N_23878,N_16403,N_14412);
nor U23879 (N_23879,N_13753,N_15567);
nor U23880 (N_23880,N_17234,N_18454);
nand U23881 (N_23881,N_18588,N_15460);
and U23882 (N_23882,N_16978,N_15817);
or U23883 (N_23883,N_16497,N_13071);
nand U23884 (N_23884,N_12954,N_15015);
xnor U23885 (N_23885,N_16604,N_17847);
nor U23886 (N_23886,N_15450,N_15483);
nand U23887 (N_23887,N_18284,N_17083);
or U23888 (N_23888,N_17881,N_13081);
nor U23889 (N_23889,N_14120,N_13778);
nand U23890 (N_23890,N_18646,N_14187);
nor U23891 (N_23891,N_15252,N_13791);
nor U23892 (N_23892,N_14302,N_15042);
and U23893 (N_23893,N_17502,N_14961);
nor U23894 (N_23894,N_16729,N_15507);
nand U23895 (N_23895,N_12631,N_16713);
nor U23896 (N_23896,N_16070,N_14334);
or U23897 (N_23897,N_16614,N_16504);
or U23898 (N_23898,N_13241,N_18023);
nand U23899 (N_23899,N_16708,N_13418);
nand U23900 (N_23900,N_17072,N_14849);
xor U23901 (N_23901,N_15634,N_17320);
nor U23902 (N_23902,N_12820,N_15901);
nor U23903 (N_23903,N_16585,N_17512);
xnor U23904 (N_23904,N_18421,N_15177);
nor U23905 (N_23905,N_18274,N_15165);
or U23906 (N_23906,N_12706,N_14714);
or U23907 (N_23907,N_17533,N_17060);
or U23908 (N_23908,N_13813,N_14432);
nand U23909 (N_23909,N_13742,N_14328);
and U23910 (N_23910,N_12802,N_17923);
nor U23911 (N_23911,N_17467,N_14775);
and U23912 (N_23912,N_14964,N_15519);
xor U23913 (N_23913,N_16288,N_12638);
and U23914 (N_23914,N_18216,N_13180);
nor U23915 (N_23915,N_12890,N_17885);
nand U23916 (N_23916,N_15337,N_14473);
nor U23917 (N_23917,N_15025,N_13307);
and U23918 (N_23918,N_18501,N_17181);
or U23919 (N_23919,N_16821,N_14235);
nor U23920 (N_23920,N_16998,N_13607);
nor U23921 (N_23921,N_14569,N_13802);
nand U23922 (N_23922,N_18050,N_17213);
or U23923 (N_23923,N_16375,N_17206);
nor U23924 (N_23924,N_17777,N_18732);
and U23925 (N_23925,N_13957,N_15152);
nor U23926 (N_23926,N_15207,N_13786);
nor U23927 (N_23927,N_14659,N_15730);
xnor U23928 (N_23928,N_12705,N_13757);
and U23929 (N_23929,N_17100,N_14157);
and U23930 (N_23930,N_14569,N_13502);
nand U23931 (N_23931,N_16299,N_18322);
nor U23932 (N_23932,N_14403,N_13442);
nor U23933 (N_23933,N_14757,N_18732);
or U23934 (N_23934,N_13931,N_17072);
nand U23935 (N_23935,N_18164,N_12764);
or U23936 (N_23936,N_17646,N_17533);
nor U23937 (N_23937,N_16234,N_16728);
or U23938 (N_23938,N_17842,N_14354);
nor U23939 (N_23939,N_18467,N_17883);
nand U23940 (N_23940,N_13370,N_16890);
nand U23941 (N_23941,N_16383,N_13074);
nand U23942 (N_23942,N_17178,N_15697);
nor U23943 (N_23943,N_14183,N_16180);
or U23944 (N_23944,N_12744,N_14249);
and U23945 (N_23945,N_18184,N_14937);
or U23946 (N_23946,N_16767,N_18514);
and U23947 (N_23947,N_16384,N_17328);
nor U23948 (N_23948,N_17213,N_16345);
nor U23949 (N_23949,N_14747,N_16588);
nor U23950 (N_23950,N_18091,N_13975);
nor U23951 (N_23951,N_15740,N_15611);
nand U23952 (N_23952,N_16509,N_12562);
xor U23953 (N_23953,N_15868,N_18051);
nor U23954 (N_23954,N_13687,N_17812);
or U23955 (N_23955,N_16488,N_13661);
nand U23956 (N_23956,N_15608,N_18492);
nor U23957 (N_23957,N_15733,N_15138);
nor U23958 (N_23958,N_14477,N_15699);
and U23959 (N_23959,N_13562,N_12850);
nor U23960 (N_23960,N_16128,N_13660);
nor U23961 (N_23961,N_14751,N_13490);
nor U23962 (N_23962,N_15574,N_14549);
xnor U23963 (N_23963,N_14495,N_18322);
nand U23964 (N_23964,N_17622,N_13943);
or U23965 (N_23965,N_16769,N_13896);
and U23966 (N_23966,N_18716,N_15574);
and U23967 (N_23967,N_13890,N_17988);
nor U23968 (N_23968,N_13403,N_13127);
nand U23969 (N_23969,N_15394,N_17993);
or U23970 (N_23970,N_14539,N_17339);
nor U23971 (N_23971,N_13594,N_14939);
nor U23972 (N_23972,N_14450,N_14299);
nand U23973 (N_23973,N_14112,N_17317);
nor U23974 (N_23974,N_15797,N_16229);
nor U23975 (N_23975,N_14662,N_17757);
xor U23976 (N_23976,N_14875,N_15893);
nand U23977 (N_23977,N_17631,N_17638);
nand U23978 (N_23978,N_14203,N_16188);
xor U23979 (N_23979,N_14059,N_14014);
or U23980 (N_23980,N_17729,N_17066);
nand U23981 (N_23981,N_12642,N_17459);
or U23982 (N_23982,N_15041,N_17782);
nand U23983 (N_23983,N_16273,N_13617);
nor U23984 (N_23984,N_15574,N_13925);
nand U23985 (N_23985,N_18714,N_15781);
or U23986 (N_23986,N_13166,N_13019);
and U23987 (N_23987,N_17448,N_18129);
xnor U23988 (N_23988,N_14746,N_16213);
nor U23989 (N_23989,N_18418,N_15501);
nand U23990 (N_23990,N_13233,N_18315);
nand U23991 (N_23991,N_12675,N_16315);
nor U23992 (N_23992,N_14686,N_17433);
nand U23993 (N_23993,N_15704,N_16172);
and U23994 (N_23994,N_17676,N_15486);
nor U23995 (N_23995,N_16321,N_15292);
nand U23996 (N_23996,N_12725,N_17728);
and U23997 (N_23997,N_15111,N_13479);
nor U23998 (N_23998,N_17878,N_13297);
xor U23999 (N_23999,N_18315,N_17288);
and U24000 (N_24000,N_12511,N_13094);
or U24001 (N_24001,N_14451,N_15590);
or U24002 (N_24002,N_12634,N_15773);
or U24003 (N_24003,N_13339,N_16696);
or U24004 (N_24004,N_15099,N_16906);
nand U24005 (N_24005,N_16028,N_16185);
nor U24006 (N_24006,N_15071,N_17477);
and U24007 (N_24007,N_18418,N_18066);
and U24008 (N_24008,N_16746,N_16554);
xnor U24009 (N_24009,N_14498,N_18345);
or U24010 (N_24010,N_12539,N_14900);
xnor U24011 (N_24011,N_16595,N_13960);
and U24012 (N_24012,N_15794,N_13432);
and U24013 (N_24013,N_13499,N_15305);
nand U24014 (N_24014,N_15251,N_12756);
or U24015 (N_24015,N_16964,N_14626);
and U24016 (N_24016,N_14612,N_14178);
nand U24017 (N_24017,N_15129,N_15703);
or U24018 (N_24018,N_13632,N_18618);
nor U24019 (N_24019,N_18238,N_15598);
nor U24020 (N_24020,N_13441,N_14694);
and U24021 (N_24021,N_14828,N_13688);
nor U24022 (N_24022,N_12664,N_17404);
and U24023 (N_24023,N_16227,N_14732);
and U24024 (N_24024,N_17223,N_17623);
and U24025 (N_24025,N_12667,N_18377);
nor U24026 (N_24026,N_16102,N_15445);
xor U24027 (N_24027,N_17234,N_14738);
and U24028 (N_24028,N_13173,N_16111);
or U24029 (N_24029,N_13870,N_14748);
or U24030 (N_24030,N_18403,N_17055);
nand U24031 (N_24031,N_13303,N_13443);
or U24032 (N_24032,N_14234,N_13994);
or U24033 (N_24033,N_16429,N_14040);
xnor U24034 (N_24034,N_13181,N_13567);
xor U24035 (N_24035,N_15903,N_17943);
nand U24036 (N_24036,N_18140,N_13264);
and U24037 (N_24037,N_15831,N_14737);
and U24038 (N_24038,N_13798,N_16798);
nand U24039 (N_24039,N_16422,N_17596);
and U24040 (N_24040,N_13083,N_13243);
nand U24041 (N_24041,N_12974,N_16877);
or U24042 (N_24042,N_16559,N_18693);
nor U24043 (N_24043,N_17722,N_12972);
nand U24044 (N_24044,N_16550,N_13797);
xnor U24045 (N_24045,N_12789,N_13992);
and U24046 (N_24046,N_13836,N_15640);
and U24047 (N_24047,N_17010,N_16172);
and U24048 (N_24048,N_15908,N_17197);
nor U24049 (N_24049,N_13592,N_14839);
nand U24050 (N_24050,N_14689,N_15119);
and U24051 (N_24051,N_17437,N_15737);
or U24052 (N_24052,N_17878,N_17810);
nand U24053 (N_24053,N_16120,N_17432);
and U24054 (N_24054,N_12973,N_15461);
nor U24055 (N_24055,N_15870,N_13849);
nor U24056 (N_24056,N_18036,N_17640);
nor U24057 (N_24057,N_12852,N_16068);
nand U24058 (N_24058,N_14334,N_16382);
nor U24059 (N_24059,N_15075,N_13405);
and U24060 (N_24060,N_13441,N_16015);
or U24061 (N_24061,N_13360,N_17463);
or U24062 (N_24062,N_13993,N_18211);
nor U24063 (N_24063,N_16400,N_17189);
or U24064 (N_24064,N_14955,N_14380);
nand U24065 (N_24065,N_17752,N_17290);
or U24066 (N_24066,N_15130,N_12557);
nor U24067 (N_24067,N_13383,N_17614);
or U24068 (N_24068,N_16042,N_18666);
or U24069 (N_24069,N_17475,N_15473);
or U24070 (N_24070,N_17759,N_17293);
and U24071 (N_24071,N_13765,N_16655);
or U24072 (N_24072,N_15196,N_15407);
or U24073 (N_24073,N_15023,N_14690);
nand U24074 (N_24074,N_18060,N_15073);
xor U24075 (N_24075,N_17349,N_18328);
or U24076 (N_24076,N_14541,N_16158);
nand U24077 (N_24077,N_13853,N_13994);
nand U24078 (N_24078,N_13160,N_12891);
nand U24079 (N_24079,N_17505,N_17144);
nand U24080 (N_24080,N_16550,N_18309);
and U24081 (N_24081,N_12592,N_14584);
nor U24082 (N_24082,N_17948,N_12819);
xnor U24083 (N_24083,N_16850,N_15865);
or U24084 (N_24084,N_18426,N_17258);
or U24085 (N_24085,N_14521,N_17366);
or U24086 (N_24086,N_16322,N_16635);
or U24087 (N_24087,N_18256,N_16162);
or U24088 (N_24088,N_18261,N_12799);
nor U24089 (N_24089,N_17223,N_15151);
xor U24090 (N_24090,N_13114,N_16293);
nor U24091 (N_24091,N_17737,N_16970);
and U24092 (N_24092,N_15052,N_18199);
and U24093 (N_24093,N_14081,N_18632);
and U24094 (N_24094,N_17733,N_13283);
xnor U24095 (N_24095,N_13440,N_18360);
or U24096 (N_24096,N_14345,N_16218);
nand U24097 (N_24097,N_13491,N_16773);
nor U24098 (N_24098,N_15808,N_14683);
nand U24099 (N_24099,N_17785,N_18147);
nand U24100 (N_24100,N_15603,N_18533);
xor U24101 (N_24101,N_18580,N_12716);
or U24102 (N_24102,N_18712,N_16719);
and U24103 (N_24103,N_13136,N_16435);
nor U24104 (N_24104,N_14861,N_16793);
nand U24105 (N_24105,N_15222,N_17608);
nor U24106 (N_24106,N_17906,N_16524);
or U24107 (N_24107,N_17923,N_18237);
and U24108 (N_24108,N_17187,N_16607);
and U24109 (N_24109,N_14765,N_14437);
nor U24110 (N_24110,N_16453,N_13634);
nand U24111 (N_24111,N_13883,N_12545);
xnor U24112 (N_24112,N_13185,N_16473);
nor U24113 (N_24113,N_15670,N_16237);
nor U24114 (N_24114,N_17814,N_18271);
xor U24115 (N_24115,N_14822,N_15760);
nor U24116 (N_24116,N_14461,N_17245);
and U24117 (N_24117,N_14071,N_14210);
nand U24118 (N_24118,N_17914,N_15098);
nand U24119 (N_24119,N_16022,N_17499);
or U24120 (N_24120,N_14774,N_14579);
and U24121 (N_24121,N_14207,N_15151);
or U24122 (N_24122,N_14668,N_13756);
or U24123 (N_24123,N_17152,N_14354);
nand U24124 (N_24124,N_18219,N_16658);
xnor U24125 (N_24125,N_15459,N_12825);
or U24126 (N_24126,N_14974,N_12850);
or U24127 (N_24127,N_17360,N_15574);
nand U24128 (N_24128,N_15957,N_16543);
nand U24129 (N_24129,N_15202,N_13876);
or U24130 (N_24130,N_13324,N_15546);
or U24131 (N_24131,N_13277,N_13020);
or U24132 (N_24132,N_17983,N_18212);
or U24133 (N_24133,N_16806,N_15737);
and U24134 (N_24134,N_12936,N_13363);
and U24135 (N_24135,N_17367,N_13467);
nor U24136 (N_24136,N_18257,N_12546);
or U24137 (N_24137,N_13072,N_16130);
nand U24138 (N_24138,N_15771,N_18552);
or U24139 (N_24139,N_12844,N_13966);
nand U24140 (N_24140,N_17790,N_13299);
nor U24141 (N_24141,N_12813,N_16227);
nand U24142 (N_24142,N_13943,N_18571);
nor U24143 (N_24143,N_18189,N_17217);
or U24144 (N_24144,N_12813,N_16885);
xor U24145 (N_24145,N_14397,N_14940);
xor U24146 (N_24146,N_12608,N_14561);
and U24147 (N_24147,N_14361,N_15006);
and U24148 (N_24148,N_15450,N_14051);
and U24149 (N_24149,N_16287,N_18230);
or U24150 (N_24150,N_17626,N_14328);
and U24151 (N_24151,N_12507,N_15114);
or U24152 (N_24152,N_16833,N_14284);
or U24153 (N_24153,N_12824,N_13743);
nor U24154 (N_24154,N_17879,N_16951);
and U24155 (N_24155,N_13009,N_16889);
nand U24156 (N_24156,N_14321,N_15783);
or U24157 (N_24157,N_13644,N_16265);
nand U24158 (N_24158,N_18194,N_17663);
xnor U24159 (N_24159,N_12698,N_16181);
or U24160 (N_24160,N_13969,N_18382);
and U24161 (N_24161,N_15122,N_15325);
and U24162 (N_24162,N_17874,N_18182);
nor U24163 (N_24163,N_17940,N_16867);
nor U24164 (N_24164,N_13323,N_17958);
nand U24165 (N_24165,N_14368,N_13276);
nand U24166 (N_24166,N_15551,N_13831);
nor U24167 (N_24167,N_17026,N_13379);
or U24168 (N_24168,N_14887,N_16883);
nand U24169 (N_24169,N_18683,N_15999);
or U24170 (N_24170,N_14437,N_17801);
nor U24171 (N_24171,N_16556,N_17704);
nand U24172 (N_24172,N_17192,N_15763);
nor U24173 (N_24173,N_15045,N_17306);
nor U24174 (N_24174,N_16011,N_17885);
and U24175 (N_24175,N_14713,N_12714);
or U24176 (N_24176,N_14074,N_12805);
nor U24177 (N_24177,N_14877,N_16544);
and U24178 (N_24178,N_15588,N_12596);
nand U24179 (N_24179,N_14831,N_16285);
nand U24180 (N_24180,N_18702,N_14389);
or U24181 (N_24181,N_16806,N_17503);
nand U24182 (N_24182,N_15995,N_16821);
nand U24183 (N_24183,N_16200,N_12607);
nand U24184 (N_24184,N_17554,N_17689);
or U24185 (N_24185,N_12670,N_13146);
nor U24186 (N_24186,N_15284,N_16930);
nand U24187 (N_24187,N_15480,N_14871);
or U24188 (N_24188,N_18026,N_15368);
nand U24189 (N_24189,N_12638,N_17045);
nand U24190 (N_24190,N_17736,N_16535);
xnor U24191 (N_24191,N_13877,N_15337);
and U24192 (N_24192,N_13757,N_14917);
nor U24193 (N_24193,N_18077,N_17299);
nand U24194 (N_24194,N_17921,N_17408);
and U24195 (N_24195,N_15719,N_14791);
or U24196 (N_24196,N_13894,N_15636);
nand U24197 (N_24197,N_13164,N_14298);
or U24198 (N_24198,N_16605,N_16248);
nor U24199 (N_24199,N_14102,N_18344);
or U24200 (N_24200,N_17895,N_17357);
nor U24201 (N_24201,N_16201,N_15512);
or U24202 (N_24202,N_18468,N_16377);
nand U24203 (N_24203,N_14045,N_14423);
or U24204 (N_24204,N_13439,N_13149);
and U24205 (N_24205,N_13312,N_18028);
nand U24206 (N_24206,N_13857,N_18051);
nand U24207 (N_24207,N_18280,N_15570);
or U24208 (N_24208,N_14795,N_17947);
and U24209 (N_24209,N_16363,N_17131);
and U24210 (N_24210,N_17929,N_13965);
nand U24211 (N_24211,N_14963,N_17358);
nor U24212 (N_24212,N_14540,N_14560);
and U24213 (N_24213,N_17613,N_17477);
nor U24214 (N_24214,N_13776,N_15916);
or U24215 (N_24215,N_12573,N_13184);
and U24216 (N_24216,N_16242,N_18522);
and U24217 (N_24217,N_17399,N_16567);
and U24218 (N_24218,N_14311,N_17518);
nor U24219 (N_24219,N_18193,N_14347);
nand U24220 (N_24220,N_15240,N_17537);
and U24221 (N_24221,N_14819,N_12903);
or U24222 (N_24222,N_17352,N_15690);
and U24223 (N_24223,N_12692,N_15831);
or U24224 (N_24224,N_15037,N_15472);
and U24225 (N_24225,N_15764,N_13578);
xor U24226 (N_24226,N_18421,N_16106);
nand U24227 (N_24227,N_16276,N_17149);
nand U24228 (N_24228,N_14310,N_13342);
nand U24229 (N_24229,N_14411,N_13465);
or U24230 (N_24230,N_14006,N_16659);
or U24231 (N_24231,N_15596,N_16765);
nor U24232 (N_24232,N_13930,N_14085);
nor U24233 (N_24233,N_16713,N_18360);
or U24234 (N_24234,N_16994,N_18368);
or U24235 (N_24235,N_14945,N_16043);
or U24236 (N_24236,N_14526,N_13689);
or U24237 (N_24237,N_13665,N_15360);
xor U24238 (N_24238,N_13568,N_14311);
and U24239 (N_24239,N_16638,N_14017);
or U24240 (N_24240,N_16164,N_15629);
or U24241 (N_24241,N_16857,N_18432);
or U24242 (N_24242,N_14814,N_15414);
and U24243 (N_24243,N_17429,N_16132);
nand U24244 (N_24244,N_17125,N_17507);
and U24245 (N_24245,N_15481,N_15769);
nand U24246 (N_24246,N_16690,N_17521);
nand U24247 (N_24247,N_15882,N_13697);
and U24248 (N_24248,N_17313,N_16634);
or U24249 (N_24249,N_13179,N_14418);
and U24250 (N_24250,N_13100,N_13449);
nand U24251 (N_24251,N_17714,N_15812);
nor U24252 (N_24252,N_16848,N_13936);
or U24253 (N_24253,N_16119,N_14976);
nor U24254 (N_24254,N_13399,N_13984);
nor U24255 (N_24255,N_18423,N_17482);
and U24256 (N_24256,N_15287,N_12501);
or U24257 (N_24257,N_18266,N_16777);
nor U24258 (N_24258,N_17850,N_17643);
nor U24259 (N_24259,N_15552,N_15811);
and U24260 (N_24260,N_13697,N_16786);
and U24261 (N_24261,N_17702,N_12618);
nor U24262 (N_24262,N_15691,N_17336);
or U24263 (N_24263,N_12863,N_15390);
or U24264 (N_24264,N_16530,N_17821);
nor U24265 (N_24265,N_14168,N_16789);
and U24266 (N_24266,N_12593,N_12910);
and U24267 (N_24267,N_13959,N_15112);
or U24268 (N_24268,N_14766,N_18010);
nand U24269 (N_24269,N_15836,N_17258);
nand U24270 (N_24270,N_15873,N_17999);
nor U24271 (N_24271,N_12650,N_18549);
or U24272 (N_24272,N_17479,N_16573);
nor U24273 (N_24273,N_17871,N_17450);
nor U24274 (N_24274,N_13654,N_15161);
xor U24275 (N_24275,N_15166,N_15984);
nand U24276 (N_24276,N_17258,N_18429);
and U24277 (N_24277,N_14220,N_13906);
xor U24278 (N_24278,N_13547,N_18260);
nor U24279 (N_24279,N_17603,N_14475);
xnor U24280 (N_24280,N_18203,N_15215);
nor U24281 (N_24281,N_18674,N_17138);
nor U24282 (N_24282,N_14593,N_16332);
or U24283 (N_24283,N_16479,N_14506);
nor U24284 (N_24284,N_15785,N_13065);
nor U24285 (N_24285,N_12991,N_13175);
and U24286 (N_24286,N_15883,N_13060);
and U24287 (N_24287,N_18376,N_16284);
nor U24288 (N_24288,N_18172,N_17598);
nor U24289 (N_24289,N_12600,N_15798);
nand U24290 (N_24290,N_15663,N_14501);
or U24291 (N_24291,N_18400,N_12769);
nand U24292 (N_24292,N_15569,N_18132);
xnor U24293 (N_24293,N_17831,N_17627);
nor U24294 (N_24294,N_18139,N_13742);
nor U24295 (N_24295,N_13636,N_14975);
nor U24296 (N_24296,N_17241,N_13161);
xnor U24297 (N_24297,N_18281,N_14549);
nor U24298 (N_24298,N_14083,N_17933);
nand U24299 (N_24299,N_13895,N_17519);
and U24300 (N_24300,N_17920,N_18668);
xor U24301 (N_24301,N_16201,N_17449);
nor U24302 (N_24302,N_15276,N_16641);
nand U24303 (N_24303,N_15889,N_15229);
nor U24304 (N_24304,N_18210,N_18074);
or U24305 (N_24305,N_15546,N_15082);
nor U24306 (N_24306,N_18410,N_14913);
and U24307 (N_24307,N_16456,N_18264);
or U24308 (N_24308,N_13378,N_13794);
and U24309 (N_24309,N_12893,N_16566);
nand U24310 (N_24310,N_16562,N_17296);
or U24311 (N_24311,N_14461,N_13738);
nor U24312 (N_24312,N_16170,N_13179);
nand U24313 (N_24313,N_15190,N_12575);
and U24314 (N_24314,N_15031,N_16434);
nor U24315 (N_24315,N_13850,N_17596);
or U24316 (N_24316,N_13559,N_15604);
or U24317 (N_24317,N_17976,N_12525);
and U24318 (N_24318,N_14515,N_17102);
or U24319 (N_24319,N_13297,N_18048);
and U24320 (N_24320,N_13710,N_18197);
or U24321 (N_24321,N_16978,N_16853);
nand U24322 (N_24322,N_17364,N_14545);
nor U24323 (N_24323,N_14804,N_18229);
nor U24324 (N_24324,N_16650,N_15565);
nand U24325 (N_24325,N_16359,N_16641);
or U24326 (N_24326,N_13909,N_17058);
or U24327 (N_24327,N_12578,N_13997);
or U24328 (N_24328,N_13256,N_14117);
nand U24329 (N_24329,N_14310,N_15800);
and U24330 (N_24330,N_18104,N_17220);
nand U24331 (N_24331,N_16882,N_13704);
and U24332 (N_24332,N_13983,N_18115);
and U24333 (N_24333,N_14305,N_15016);
xnor U24334 (N_24334,N_15763,N_13802);
nor U24335 (N_24335,N_16274,N_18523);
nand U24336 (N_24336,N_16241,N_16803);
or U24337 (N_24337,N_15429,N_17389);
xor U24338 (N_24338,N_18092,N_17545);
xor U24339 (N_24339,N_17420,N_15424);
nor U24340 (N_24340,N_17822,N_18246);
and U24341 (N_24341,N_14781,N_12613);
xnor U24342 (N_24342,N_16010,N_16888);
nand U24343 (N_24343,N_12986,N_18359);
nand U24344 (N_24344,N_17574,N_16736);
nand U24345 (N_24345,N_15237,N_14936);
nor U24346 (N_24346,N_12651,N_17120);
nor U24347 (N_24347,N_13554,N_17723);
or U24348 (N_24348,N_15376,N_15084);
nand U24349 (N_24349,N_13507,N_13057);
and U24350 (N_24350,N_17162,N_13084);
xnor U24351 (N_24351,N_15511,N_14878);
and U24352 (N_24352,N_16765,N_12653);
or U24353 (N_24353,N_17567,N_18061);
and U24354 (N_24354,N_15704,N_16324);
or U24355 (N_24355,N_16170,N_13995);
nand U24356 (N_24356,N_15972,N_17176);
xor U24357 (N_24357,N_14558,N_16761);
and U24358 (N_24358,N_14175,N_15696);
or U24359 (N_24359,N_18209,N_14866);
nand U24360 (N_24360,N_13505,N_14090);
or U24361 (N_24361,N_18208,N_14890);
nor U24362 (N_24362,N_12992,N_13508);
nor U24363 (N_24363,N_15499,N_18200);
or U24364 (N_24364,N_15449,N_16909);
xnor U24365 (N_24365,N_17544,N_16608);
and U24366 (N_24366,N_13301,N_18414);
nand U24367 (N_24367,N_16752,N_15068);
xnor U24368 (N_24368,N_16682,N_16408);
nor U24369 (N_24369,N_18127,N_18617);
nand U24370 (N_24370,N_15553,N_18505);
nand U24371 (N_24371,N_14932,N_12665);
nor U24372 (N_24372,N_18273,N_13818);
nor U24373 (N_24373,N_13619,N_18302);
nor U24374 (N_24374,N_16189,N_15029);
nor U24375 (N_24375,N_16724,N_18646);
nor U24376 (N_24376,N_18087,N_13762);
xor U24377 (N_24377,N_15526,N_16974);
and U24378 (N_24378,N_17134,N_16298);
nand U24379 (N_24379,N_17768,N_14558);
and U24380 (N_24380,N_17114,N_18256);
or U24381 (N_24381,N_17083,N_18106);
and U24382 (N_24382,N_16621,N_17597);
nor U24383 (N_24383,N_18000,N_13812);
nand U24384 (N_24384,N_13870,N_12902);
nand U24385 (N_24385,N_12798,N_15884);
or U24386 (N_24386,N_15062,N_12904);
and U24387 (N_24387,N_17186,N_15301);
nand U24388 (N_24388,N_17444,N_15797);
or U24389 (N_24389,N_13163,N_16855);
and U24390 (N_24390,N_17539,N_13618);
or U24391 (N_24391,N_14944,N_13830);
nand U24392 (N_24392,N_14172,N_17685);
nor U24393 (N_24393,N_13425,N_14636);
nand U24394 (N_24394,N_16803,N_14966);
nand U24395 (N_24395,N_14988,N_14226);
and U24396 (N_24396,N_16360,N_16727);
nand U24397 (N_24397,N_14570,N_15002);
and U24398 (N_24398,N_13044,N_16490);
nor U24399 (N_24399,N_15952,N_14768);
nor U24400 (N_24400,N_14497,N_13400);
nand U24401 (N_24401,N_13183,N_18149);
nand U24402 (N_24402,N_15183,N_16909);
and U24403 (N_24403,N_18224,N_17230);
nand U24404 (N_24404,N_13917,N_15562);
and U24405 (N_24405,N_16416,N_17730);
or U24406 (N_24406,N_13497,N_15068);
nand U24407 (N_24407,N_17835,N_16929);
and U24408 (N_24408,N_17721,N_14258);
nand U24409 (N_24409,N_17539,N_18473);
or U24410 (N_24410,N_18362,N_18295);
or U24411 (N_24411,N_18243,N_13997);
or U24412 (N_24412,N_16219,N_16114);
or U24413 (N_24413,N_12610,N_17501);
xnor U24414 (N_24414,N_14621,N_15322);
nor U24415 (N_24415,N_15063,N_17874);
nor U24416 (N_24416,N_17121,N_13743);
and U24417 (N_24417,N_18204,N_18293);
or U24418 (N_24418,N_14991,N_16799);
and U24419 (N_24419,N_14548,N_18013);
and U24420 (N_24420,N_14058,N_12764);
nand U24421 (N_24421,N_14724,N_15778);
xor U24422 (N_24422,N_16534,N_17578);
and U24423 (N_24423,N_15589,N_16983);
nand U24424 (N_24424,N_15006,N_13566);
or U24425 (N_24425,N_15648,N_16392);
xnor U24426 (N_24426,N_18404,N_18734);
or U24427 (N_24427,N_16131,N_12692);
xor U24428 (N_24428,N_15683,N_14869);
nor U24429 (N_24429,N_18393,N_16555);
xor U24430 (N_24430,N_17593,N_14810);
xnor U24431 (N_24431,N_15233,N_18530);
nand U24432 (N_24432,N_17850,N_13071);
or U24433 (N_24433,N_13450,N_12569);
nor U24434 (N_24434,N_14152,N_18247);
or U24435 (N_24435,N_15620,N_13971);
nand U24436 (N_24436,N_17033,N_18660);
and U24437 (N_24437,N_12781,N_14980);
and U24438 (N_24438,N_12827,N_16513);
nor U24439 (N_24439,N_14179,N_17443);
nand U24440 (N_24440,N_17127,N_14477);
or U24441 (N_24441,N_14479,N_15809);
or U24442 (N_24442,N_16619,N_15767);
nand U24443 (N_24443,N_13856,N_15403);
or U24444 (N_24444,N_16332,N_15200);
or U24445 (N_24445,N_15561,N_17601);
nor U24446 (N_24446,N_12954,N_16631);
nor U24447 (N_24447,N_14896,N_17816);
nand U24448 (N_24448,N_16146,N_14136);
nand U24449 (N_24449,N_17226,N_16995);
nand U24450 (N_24450,N_15258,N_16236);
xor U24451 (N_24451,N_13067,N_14763);
nand U24452 (N_24452,N_16486,N_16475);
or U24453 (N_24453,N_14003,N_14862);
nor U24454 (N_24454,N_17761,N_17816);
or U24455 (N_24455,N_13539,N_17948);
or U24456 (N_24456,N_16385,N_13215);
nand U24457 (N_24457,N_16125,N_14991);
nor U24458 (N_24458,N_14088,N_12544);
or U24459 (N_24459,N_18234,N_17347);
nand U24460 (N_24460,N_13239,N_13119);
and U24461 (N_24461,N_17811,N_13099);
nor U24462 (N_24462,N_12812,N_15818);
and U24463 (N_24463,N_13684,N_12676);
and U24464 (N_24464,N_16523,N_17252);
or U24465 (N_24465,N_17955,N_18078);
nor U24466 (N_24466,N_12907,N_12700);
or U24467 (N_24467,N_17023,N_17904);
and U24468 (N_24468,N_18452,N_14924);
nor U24469 (N_24469,N_13076,N_12907);
nor U24470 (N_24470,N_16155,N_17964);
or U24471 (N_24471,N_16600,N_17300);
or U24472 (N_24472,N_17507,N_15011);
xnor U24473 (N_24473,N_14999,N_12756);
nor U24474 (N_24474,N_17899,N_15081);
nand U24475 (N_24475,N_18686,N_13727);
or U24476 (N_24476,N_14630,N_14590);
xor U24477 (N_24477,N_18369,N_15419);
and U24478 (N_24478,N_17431,N_14106);
or U24479 (N_24479,N_15457,N_13884);
nor U24480 (N_24480,N_15297,N_13698);
or U24481 (N_24481,N_14481,N_13052);
or U24482 (N_24482,N_18558,N_17441);
or U24483 (N_24483,N_13890,N_15308);
nor U24484 (N_24484,N_12818,N_13389);
xor U24485 (N_24485,N_18681,N_14003);
and U24486 (N_24486,N_13318,N_15802);
xnor U24487 (N_24487,N_13057,N_14565);
nand U24488 (N_24488,N_12768,N_16636);
xnor U24489 (N_24489,N_18219,N_12884);
or U24490 (N_24490,N_17244,N_14046);
nand U24491 (N_24491,N_16456,N_16766);
and U24492 (N_24492,N_13804,N_16700);
or U24493 (N_24493,N_16005,N_14154);
nor U24494 (N_24494,N_16366,N_14927);
xor U24495 (N_24495,N_18054,N_14854);
and U24496 (N_24496,N_15635,N_17508);
xnor U24497 (N_24497,N_18377,N_17488);
and U24498 (N_24498,N_17364,N_16284);
and U24499 (N_24499,N_14009,N_13698);
or U24500 (N_24500,N_14505,N_16535);
and U24501 (N_24501,N_13293,N_16224);
nand U24502 (N_24502,N_13887,N_18107);
nand U24503 (N_24503,N_15058,N_15015);
nand U24504 (N_24504,N_14283,N_12721);
and U24505 (N_24505,N_16136,N_17166);
or U24506 (N_24506,N_15233,N_14748);
nand U24507 (N_24507,N_14806,N_12846);
nand U24508 (N_24508,N_13776,N_14573);
nor U24509 (N_24509,N_14111,N_16311);
or U24510 (N_24510,N_15919,N_17576);
and U24511 (N_24511,N_15760,N_15703);
or U24512 (N_24512,N_18446,N_17617);
or U24513 (N_24513,N_13664,N_13749);
nor U24514 (N_24514,N_14051,N_13796);
nand U24515 (N_24515,N_12876,N_14475);
nand U24516 (N_24516,N_18296,N_17659);
or U24517 (N_24517,N_16845,N_14110);
and U24518 (N_24518,N_17162,N_13940);
or U24519 (N_24519,N_15836,N_13364);
nand U24520 (N_24520,N_17083,N_13002);
xnor U24521 (N_24521,N_15551,N_15550);
or U24522 (N_24522,N_16574,N_15048);
nand U24523 (N_24523,N_13789,N_16864);
nand U24524 (N_24524,N_15057,N_16618);
and U24525 (N_24525,N_14433,N_14026);
or U24526 (N_24526,N_13828,N_13189);
and U24527 (N_24527,N_16014,N_15615);
and U24528 (N_24528,N_17391,N_14921);
nor U24529 (N_24529,N_15539,N_13457);
or U24530 (N_24530,N_14435,N_16959);
nor U24531 (N_24531,N_14451,N_16979);
nor U24532 (N_24532,N_14195,N_13597);
and U24533 (N_24533,N_13029,N_13325);
nand U24534 (N_24534,N_15387,N_14152);
or U24535 (N_24535,N_16144,N_15977);
and U24536 (N_24536,N_17263,N_14306);
nor U24537 (N_24537,N_15836,N_12994);
or U24538 (N_24538,N_17214,N_18323);
or U24539 (N_24539,N_16767,N_16475);
nand U24540 (N_24540,N_18735,N_18671);
or U24541 (N_24541,N_14896,N_13286);
or U24542 (N_24542,N_15544,N_13390);
and U24543 (N_24543,N_17824,N_15685);
or U24544 (N_24544,N_13384,N_15813);
xor U24545 (N_24545,N_18535,N_13655);
nand U24546 (N_24546,N_13454,N_16571);
or U24547 (N_24547,N_18544,N_16685);
or U24548 (N_24548,N_13277,N_13640);
and U24549 (N_24549,N_16792,N_12671);
nand U24550 (N_24550,N_15624,N_14028);
and U24551 (N_24551,N_17181,N_15322);
or U24552 (N_24552,N_12632,N_13635);
or U24553 (N_24553,N_15439,N_12766);
nor U24554 (N_24554,N_18068,N_14873);
nand U24555 (N_24555,N_17706,N_17105);
nand U24556 (N_24556,N_17780,N_17651);
or U24557 (N_24557,N_17882,N_12911);
and U24558 (N_24558,N_12978,N_16570);
or U24559 (N_24559,N_14043,N_13539);
nand U24560 (N_24560,N_15301,N_16314);
nor U24561 (N_24561,N_13566,N_16660);
nor U24562 (N_24562,N_14895,N_17214);
and U24563 (N_24563,N_12554,N_12903);
or U24564 (N_24564,N_14618,N_12716);
nand U24565 (N_24565,N_13393,N_13427);
nand U24566 (N_24566,N_13255,N_14020);
or U24567 (N_24567,N_14484,N_15183);
or U24568 (N_24568,N_13932,N_13278);
and U24569 (N_24569,N_13957,N_15869);
or U24570 (N_24570,N_18431,N_12995);
nor U24571 (N_24571,N_18031,N_16797);
nand U24572 (N_24572,N_13067,N_15963);
and U24573 (N_24573,N_17990,N_13208);
or U24574 (N_24574,N_18066,N_16935);
and U24575 (N_24575,N_16262,N_15885);
nor U24576 (N_24576,N_13342,N_15843);
nor U24577 (N_24577,N_14221,N_14794);
and U24578 (N_24578,N_17577,N_16303);
and U24579 (N_24579,N_18195,N_13135);
nor U24580 (N_24580,N_17665,N_17514);
nor U24581 (N_24581,N_13255,N_14783);
or U24582 (N_24582,N_12685,N_16992);
and U24583 (N_24583,N_16029,N_17696);
nor U24584 (N_24584,N_13364,N_15989);
or U24585 (N_24585,N_13995,N_13556);
or U24586 (N_24586,N_13655,N_13940);
nand U24587 (N_24587,N_16121,N_15824);
and U24588 (N_24588,N_14457,N_18686);
or U24589 (N_24589,N_17930,N_18182);
nand U24590 (N_24590,N_14504,N_16986);
nand U24591 (N_24591,N_15291,N_13177);
and U24592 (N_24592,N_14335,N_17869);
and U24593 (N_24593,N_16899,N_18265);
or U24594 (N_24594,N_16636,N_17456);
nor U24595 (N_24595,N_17183,N_17893);
and U24596 (N_24596,N_17748,N_17833);
and U24597 (N_24597,N_15661,N_17318);
nand U24598 (N_24598,N_17390,N_17163);
or U24599 (N_24599,N_13881,N_17078);
nor U24600 (N_24600,N_16716,N_16197);
nand U24601 (N_24601,N_15165,N_18332);
nor U24602 (N_24602,N_15704,N_12668);
or U24603 (N_24603,N_13921,N_14766);
xor U24604 (N_24604,N_15426,N_14063);
nor U24605 (N_24605,N_17059,N_14807);
and U24606 (N_24606,N_17637,N_13657);
nand U24607 (N_24607,N_15736,N_16099);
nand U24608 (N_24608,N_16119,N_17782);
and U24609 (N_24609,N_16807,N_12546);
nand U24610 (N_24610,N_16242,N_12633);
or U24611 (N_24611,N_12710,N_17591);
nand U24612 (N_24612,N_15105,N_18156);
xnor U24613 (N_24613,N_16439,N_17466);
xnor U24614 (N_24614,N_14837,N_17141);
and U24615 (N_24615,N_13551,N_18124);
nand U24616 (N_24616,N_15104,N_12706);
nand U24617 (N_24617,N_16799,N_14238);
nand U24618 (N_24618,N_14790,N_14247);
xnor U24619 (N_24619,N_17516,N_18653);
and U24620 (N_24620,N_17817,N_15775);
xor U24621 (N_24621,N_17676,N_15420);
and U24622 (N_24622,N_16378,N_15497);
nand U24623 (N_24623,N_15487,N_18517);
nor U24624 (N_24624,N_17385,N_15081);
nand U24625 (N_24625,N_13639,N_18403);
nor U24626 (N_24626,N_16495,N_16223);
or U24627 (N_24627,N_15675,N_13049);
nor U24628 (N_24628,N_17425,N_16700);
or U24629 (N_24629,N_15440,N_12913);
nand U24630 (N_24630,N_18393,N_15877);
nand U24631 (N_24631,N_15096,N_13938);
or U24632 (N_24632,N_12817,N_17509);
nand U24633 (N_24633,N_17141,N_14758);
or U24634 (N_24634,N_14248,N_12877);
or U24635 (N_24635,N_14152,N_17172);
and U24636 (N_24636,N_14156,N_16191);
and U24637 (N_24637,N_16303,N_13713);
or U24638 (N_24638,N_15289,N_16683);
nor U24639 (N_24639,N_16286,N_18104);
or U24640 (N_24640,N_15059,N_16129);
nand U24641 (N_24641,N_12840,N_14795);
nand U24642 (N_24642,N_12938,N_14763);
and U24643 (N_24643,N_14653,N_14069);
nand U24644 (N_24644,N_15773,N_14513);
nand U24645 (N_24645,N_18230,N_18653);
and U24646 (N_24646,N_15534,N_17179);
nand U24647 (N_24647,N_16878,N_15335);
nor U24648 (N_24648,N_18677,N_16366);
nor U24649 (N_24649,N_15120,N_13672);
nor U24650 (N_24650,N_15490,N_14792);
and U24651 (N_24651,N_18134,N_14267);
or U24652 (N_24652,N_15591,N_15403);
nor U24653 (N_24653,N_16349,N_15882);
and U24654 (N_24654,N_13246,N_14782);
and U24655 (N_24655,N_12706,N_18163);
nand U24656 (N_24656,N_17422,N_16595);
nand U24657 (N_24657,N_16380,N_18684);
nand U24658 (N_24658,N_14828,N_14743);
xor U24659 (N_24659,N_13949,N_18212);
nand U24660 (N_24660,N_15636,N_16854);
or U24661 (N_24661,N_15666,N_14620);
or U24662 (N_24662,N_17587,N_16902);
nand U24663 (N_24663,N_13860,N_17216);
nand U24664 (N_24664,N_13255,N_13031);
nor U24665 (N_24665,N_16277,N_17053);
nand U24666 (N_24666,N_17917,N_13162);
or U24667 (N_24667,N_13776,N_16987);
nor U24668 (N_24668,N_12783,N_16606);
xor U24669 (N_24669,N_15831,N_15263);
nor U24670 (N_24670,N_12836,N_15703);
and U24671 (N_24671,N_16613,N_17025);
nor U24672 (N_24672,N_17351,N_13411);
nor U24673 (N_24673,N_17349,N_15106);
nor U24674 (N_24674,N_17608,N_17885);
nand U24675 (N_24675,N_18710,N_13467);
xor U24676 (N_24676,N_18224,N_13215);
and U24677 (N_24677,N_18025,N_15518);
and U24678 (N_24678,N_14777,N_16422);
or U24679 (N_24679,N_15081,N_18281);
xor U24680 (N_24680,N_14766,N_16047);
or U24681 (N_24681,N_18132,N_17165);
and U24682 (N_24682,N_14674,N_16082);
nand U24683 (N_24683,N_12593,N_14969);
nand U24684 (N_24684,N_18071,N_13602);
nor U24685 (N_24685,N_15559,N_13003);
or U24686 (N_24686,N_13164,N_18628);
and U24687 (N_24687,N_16849,N_16084);
or U24688 (N_24688,N_12526,N_18391);
nand U24689 (N_24689,N_17846,N_12714);
nand U24690 (N_24690,N_15126,N_17676);
nor U24691 (N_24691,N_16793,N_17729);
nor U24692 (N_24692,N_13554,N_14196);
nand U24693 (N_24693,N_15977,N_13484);
nand U24694 (N_24694,N_16854,N_16679);
nand U24695 (N_24695,N_15547,N_16950);
and U24696 (N_24696,N_18747,N_17749);
nand U24697 (N_24697,N_14655,N_15820);
nand U24698 (N_24698,N_17198,N_13434);
xor U24699 (N_24699,N_17555,N_15957);
nor U24700 (N_24700,N_18289,N_15927);
and U24701 (N_24701,N_15369,N_18241);
or U24702 (N_24702,N_17946,N_15450);
nor U24703 (N_24703,N_13279,N_18438);
xor U24704 (N_24704,N_17928,N_13462);
nand U24705 (N_24705,N_12987,N_14829);
or U24706 (N_24706,N_14960,N_13888);
or U24707 (N_24707,N_17917,N_17511);
nand U24708 (N_24708,N_13646,N_14219);
nor U24709 (N_24709,N_15418,N_18302);
nand U24710 (N_24710,N_14879,N_13773);
and U24711 (N_24711,N_13847,N_18130);
nand U24712 (N_24712,N_16028,N_13646);
or U24713 (N_24713,N_18472,N_14021);
and U24714 (N_24714,N_12715,N_18626);
and U24715 (N_24715,N_14913,N_13220);
and U24716 (N_24716,N_12720,N_14368);
and U24717 (N_24717,N_14982,N_15424);
or U24718 (N_24718,N_16376,N_14610);
xor U24719 (N_24719,N_15539,N_16917);
or U24720 (N_24720,N_14913,N_16422);
or U24721 (N_24721,N_15236,N_18725);
or U24722 (N_24722,N_13671,N_14542);
nand U24723 (N_24723,N_15943,N_18637);
nor U24724 (N_24724,N_16957,N_12516);
or U24725 (N_24725,N_14990,N_13217);
and U24726 (N_24726,N_13804,N_12886);
xor U24727 (N_24727,N_12993,N_16005);
or U24728 (N_24728,N_13021,N_14125);
nand U24729 (N_24729,N_14552,N_14419);
and U24730 (N_24730,N_12625,N_16724);
nor U24731 (N_24731,N_18641,N_17716);
or U24732 (N_24732,N_13433,N_14807);
and U24733 (N_24733,N_12756,N_15605);
nor U24734 (N_24734,N_15078,N_15510);
nand U24735 (N_24735,N_18316,N_13199);
nand U24736 (N_24736,N_14545,N_16270);
nand U24737 (N_24737,N_15622,N_18098);
or U24738 (N_24738,N_13013,N_14861);
or U24739 (N_24739,N_15517,N_18460);
or U24740 (N_24740,N_14978,N_18560);
nand U24741 (N_24741,N_14504,N_15978);
and U24742 (N_24742,N_17099,N_17683);
nand U24743 (N_24743,N_18608,N_17292);
and U24744 (N_24744,N_15451,N_14585);
or U24745 (N_24745,N_18720,N_16603);
nor U24746 (N_24746,N_18207,N_17074);
or U24747 (N_24747,N_13563,N_15588);
xor U24748 (N_24748,N_14236,N_13553);
nor U24749 (N_24749,N_14963,N_15997);
or U24750 (N_24750,N_13050,N_14710);
and U24751 (N_24751,N_18707,N_14157);
nor U24752 (N_24752,N_13422,N_16847);
nand U24753 (N_24753,N_15965,N_17447);
xnor U24754 (N_24754,N_15966,N_18704);
nor U24755 (N_24755,N_16289,N_18315);
or U24756 (N_24756,N_14931,N_18151);
nand U24757 (N_24757,N_16781,N_13238);
and U24758 (N_24758,N_14833,N_18680);
or U24759 (N_24759,N_12829,N_14079);
nor U24760 (N_24760,N_12679,N_16948);
xnor U24761 (N_24761,N_15801,N_13537);
nand U24762 (N_24762,N_14306,N_18411);
nand U24763 (N_24763,N_13589,N_13361);
and U24764 (N_24764,N_16901,N_17299);
and U24765 (N_24765,N_18236,N_15785);
or U24766 (N_24766,N_15283,N_15366);
nand U24767 (N_24767,N_13335,N_16528);
or U24768 (N_24768,N_13167,N_13262);
or U24769 (N_24769,N_12964,N_15680);
nor U24770 (N_24770,N_14635,N_14734);
and U24771 (N_24771,N_14682,N_13727);
or U24772 (N_24772,N_12964,N_14433);
nand U24773 (N_24773,N_17946,N_14047);
or U24774 (N_24774,N_14302,N_15872);
nand U24775 (N_24775,N_18229,N_12919);
nand U24776 (N_24776,N_13802,N_15346);
xor U24777 (N_24777,N_14748,N_14145);
or U24778 (N_24778,N_15596,N_15604);
nor U24779 (N_24779,N_16583,N_16258);
or U24780 (N_24780,N_16543,N_15244);
xnor U24781 (N_24781,N_16558,N_18374);
and U24782 (N_24782,N_13203,N_13747);
nor U24783 (N_24783,N_17300,N_15785);
nor U24784 (N_24784,N_12746,N_14549);
nor U24785 (N_24785,N_18427,N_12708);
nand U24786 (N_24786,N_15641,N_12658);
or U24787 (N_24787,N_16095,N_18625);
nand U24788 (N_24788,N_17697,N_12938);
nor U24789 (N_24789,N_16967,N_16780);
or U24790 (N_24790,N_18670,N_13471);
nor U24791 (N_24791,N_15372,N_15541);
nand U24792 (N_24792,N_15924,N_14612);
and U24793 (N_24793,N_13387,N_17463);
or U24794 (N_24794,N_15270,N_16318);
nand U24795 (N_24795,N_14894,N_17479);
and U24796 (N_24796,N_14231,N_14379);
nand U24797 (N_24797,N_18517,N_14650);
or U24798 (N_24798,N_14676,N_13407);
xnor U24799 (N_24799,N_16975,N_13503);
or U24800 (N_24800,N_14560,N_13535);
nand U24801 (N_24801,N_15460,N_12520);
or U24802 (N_24802,N_18000,N_12690);
nor U24803 (N_24803,N_17159,N_16112);
xnor U24804 (N_24804,N_18335,N_18521);
nor U24805 (N_24805,N_15476,N_14597);
and U24806 (N_24806,N_13642,N_13338);
or U24807 (N_24807,N_17357,N_15528);
nor U24808 (N_24808,N_15314,N_13036);
xnor U24809 (N_24809,N_15326,N_12602);
and U24810 (N_24810,N_18279,N_12877);
xnor U24811 (N_24811,N_14067,N_13187);
xnor U24812 (N_24812,N_12741,N_16194);
xor U24813 (N_24813,N_15747,N_17507);
nand U24814 (N_24814,N_13161,N_13525);
or U24815 (N_24815,N_13149,N_17461);
or U24816 (N_24816,N_13394,N_15481);
or U24817 (N_24817,N_13694,N_14626);
and U24818 (N_24818,N_13139,N_15774);
nor U24819 (N_24819,N_14095,N_13741);
or U24820 (N_24820,N_18488,N_12793);
nand U24821 (N_24821,N_16484,N_16267);
nand U24822 (N_24822,N_16974,N_14326);
and U24823 (N_24823,N_18662,N_16016);
or U24824 (N_24824,N_16507,N_13366);
and U24825 (N_24825,N_14242,N_14569);
nor U24826 (N_24826,N_14377,N_16147);
and U24827 (N_24827,N_12757,N_17583);
or U24828 (N_24828,N_13618,N_17525);
nand U24829 (N_24829,N_14038,N_14433);
xnor U24830 (N_24830,N_17648,N_16184);
and U24831 (N_24831,N_17887,N_16661);
nor U24832 (N_24832,N_15604,N_13051);
xor U24833 (N_24833,N_16471,N_17652);
and U24834 (N_24834,N_12878,N_17467);
and U24835 (N_24835,N_15714,N_12790);
xnor U24836 (N_24836,N_17736,N_18711);
xnor U24837 (N_24837,N_17390,N_14248);
xnor U24838 (N_24838,N_17530,N_14394);
and U24839 (N_24839,N_13529,N_13754);
or U24840 (N_24840,N_15948,N_13385);
and U24841 (N_24841,N_17490,N_14604);
and U24842 (N_24842,N_13563,N_14388);
nand U24843 (N_24843,N_13085,N_15467);
and U24844 (N_24844,N_17881,N_13503);
nand U24845 (N_24845,N_13197,N_17574);
nand U24846 (N_24846,N_12881,N_14611);
nor U24847 (N_24847,N_17612,N_14288);
or U24848 (N_24848,N_16884,N_15250);
or U24849 (N_24849,N_14338,N_15684);
nor U24850 (N_24850,N_17232,N_13303);
nand U24851 (N_24851,N_15050,N_18459);
nor U24852 (N_24852,N_15302,N_15229);
nor U24853 (N_24853,N_12944,N_17611);
nand U24854 (N_24854,N_13696,N_15843);
or U24855 (N_24855,N_15145,N_13364);
nand U24856 (N_24856,N_17029,N_17372);
or U24857 (N_24857,N_17651,N_14447);
nor U24858 (N_24858,N_18405,N_17374);
and U24859 (N_24859,N_14026,N_13061);
and U24860 (N_24860,N_13039,N_18266);
or U24861 (N_24861,N_17660,N_18700);
xnor U24862 (N_24862,N_13413,N_15220);
nand U24863 (N_24863,N_18540,N_14505);
and U24864 (N_24864,N_15268,N_12880);
nor U24865 (N_24865,N_12680,N_14387);
and U24866 (N_24866,N_15737,N_13360);
nor U24867 (N_24867,N_15699,N_16873);
nand U24868 (N_24868,N_13751,N_15126);
and U24869 (N_24869,N_18407,N_13845);
nand U24870 (N_24870,N_16092,N_12833);
nand U24871 (N_24871,N_14333,N_15073);
nor U24872 (N_24872,N_13926,N_16108);
and U24873 (N_24873,N_12942,N_14370);
nand U24874 (N_24874,N_16036,N_17395);
nand U24875 (N_24875,N_12522,N_15103);
nand U24876 (N_24876,N_18319,N_18262);
nand U24877 (N_24877,N_18704,N_18039);
nand U24878 (N_24878,N_13650,N_15950);
and U24879 (N_24879,N_14129,N_16973);
and U24880 (N_24880,N_13754,N_17993);
xnor U24881 (N_24881,N_16092,N_17751);
nor U24882 (N_24882,N_14138,N_13860);
and U24883 (N_24883,N_12911,N_15318);
nand U24884 (N_24884,N_18356,N_18408);
and U24885 (N_24885,N_17578,N_15407);
or U24886 (N_24886,N_15143,N_15652);
nor U24887 (N_24887,N_16838,N_15103);
nand U24888 (N_24888,N_16087,N_18469);
or U24889 (N_24889,N_17288,N_16017);
or U24890 (N_24890,N_12551,N_13746);
nand U24891 (N_24891,N_17746,N_14912);
or U24892 (N_24892,N_14026,N_18749);
nor U24893 (N_24893,N_14121,N_13494);
or U24894 (N_24894,N_13611,N_13741);
xor U24895 (N_24895,N_16634,N_17435);
xnor U24896 (N_24896,N_15007,N_18017);
or U24897 (N_24897,N_14066,N_13623);
nand U24898 (N_24898,N_12871,N_12746);
xnor U24899 (N_24899,N_17133,N_14133);
or U24900 (N_24900,N_16299,N_16664);
and U24901 (N_24901,N_16523,N_14824);
nor U24902 (N_24902,N_18497,N_17999);
and U24903 (N_24903,N_14812,N_14832);
xnor U24904 (N_24904,N_18048,N_16942);
nand U24905 (N_24905,N_14979,N_16346);
nand U24906 (N_24906,N_17846,N_17892);
nand U24907 (N_24907,N_14983,N_17910);
nor U24908 (N_24908,N_17785,N_13766);
nand U24909 (N_24909,N_13504,N_15215);
or U24910 (N_24910,N_18281,N_17359);
nand U24911 (N_24911,N_17905,N_12589);
or U24912 (N_24912,N_14575,N_12523);
nand U24913 (N_24913,N_16349,N_14956);
or U24914 (N_24914,N_17539,N_17803);
and U24915 (N_24915,N_14113,N_16042);
and U24916 (N_24916,N_15103,N_15004);
xnor U24917 (N_24917,N_16693,N_16217);
or U24918 (N_24918,N_14986,N_14292);
xor U24919 (N_24919,N_15354,N_18052);
or U24920 (N_24920,N_12532,N_12509);
nand U24921 (N_24921,N_13892,N_15596);
or U24922 (N_24922,N_17422,N_13757);
and U24923 (N_24923,N_18598,N_14572);
nand U24924 (N_24924,N_15705,N_16290);
nand U24925 (N_24925,N_16866,N_12895);
or U24926 (N_24926,N_17579,N_16611);
or U24927 (N_24927,N_17548,N_15888);
or U24928 (N_24928,N_15533,N_18053);
nand U24929 (N_24929,N_18112,N_17337);
and U24930 (N_24930,N_15390,N_15747);
or U24931 (N_24931,N_13715,N_12727);
or U24932 (N_24932,N_17619,N_16641);
nor U24933 (N_24933,N_17428,N_18733);
nor U24934 (N_24934,N_16344,N_18574);
nor U24935 (N_24935,N_12591,N_15837);
nand U24936 (N_24936,N_16632,N_14923);
nor U24937 (N_24937,N_18398,N_14943);
nand U24938 (N_24938,N_18365,N_18282);
nand U24939 (N_24939,N_16721,N_15887);
or U24940 (N_24940,N_16946,N_17964);
or U24941 (N_24941,N_17198,N_18732);
or U24942 (N_24942,N_16347,N_13865);
nor U24943 (N_24943,N_15870,N_18405);
nand U24944 (N_24944,N_15142,N_16590);
nor U24945 (N_24945,N_15818,N_16358);
or U24946 (N_24946,N_18157,N_18047);
nor U24947 (N_24947,N_16137,N_18353);
or U24948 (N_24948,N_12916,N_14499);
nand U24949 (N_24949,N_13731,N_16344);
and U24950 (N_24950,N_12900,N_14306);
or U24951 (N_24951,N_18293,N_17471);
nand U24952 (N_24952,N_18515,N_12951);
and U24953 (N_24953,N_17486,N_15658);
nand U24954 (N_24954,N_16105,N_13326);
nor U24955 (N_24955,N_17708,N_15590);
and U24956 (N_24956,N_12513,N_17952);
xnor U24957 (N_24957,N_17947,N_14626);
and U24958 (N_24958,N_13298,N_16092);
or U24959 (N_24959,N_17228,N_17983);
or U24960 (N_24960,N_14192,N_17819);
nand U24961 (N_24961,N_15982,N_18624);
xnor U24962 (N_24962,N_12700,N_17891);
nor U24963 (N_24963,N_12646,N_17725);
nand U24964 (N_24964,N_16842,N_13100);
nand U24965 (N_24965,N_13423,N_14941);
or U24966 (N_24966,N_16001,N_16130);
nor U24967 (N_24967,N_13990,N_14321);
nor U24968 (N_24968,N_16390,N_14091);
or U24969 (N_24969,N_12724,N_17198);
xnor U24970 (N_24970,N_17901,N_15646);
and U24971 (N_24971,N_12749,N_14268);
nand U24972 (N_24972,N_13772,N_14614);
or U24973 (N_24973,N_12526,N_12929);
nor U24974 (N_24974,N_15608,N_12971);
nor U24975 (N_24975,N_15597,N_15344);
nor U24976 (N_24976,N_15358,N_16538);
or U24977 (N_24977,N_15504,N_16221);
nor U24978 (N_24978,N_15581,N_12852);
or U24979 (N_24979,N_18481,N_13571);
nand U24980 (N_24980,N_18126,N_15850);
nand U24981 (N_24981,N_18225,N_13395);
nor U24982 (N_24982,N_18190,N_16458);
or U24983 (N_24983,N_14603,N_17119);
and U24984 (N_24984,N_17384,N_18261);
nor U24985 (N_24985,N_13825,N_15786);
xor U24986 (N_24986,N_16221,N_13859);
and U24987 (N_24987,N_17638,N_18313);
nor U24988 (N_24988,N_15758,N_15638);
or U24989 (N_24989,N_16592,N_15206);
nand U24990 (N_24990,N_13201,N_14425);
nand U24991 (N_24991,N_15752,N_17749);
or U24992 (N_24992,N_15459,N_13446);
or U24993 (N_24993,N_13315,N_18197);
nand U24994 (N_24994,N_14705,N_15203);
xor U24995 (N_24995,N_15953,N_15518);
and U24996 (N_24996,N_13727,N_17834);
or U24997 (N_24997,N_13412,N_14323);
and U24998 (N_24998,N_16706,N_12698);
or U24999 (N_24999,N_17880,N_16109);
xor UO_0 (O_0,N_19290,N_22677);
nor UO_1 (O_1,N_19748,N_21952);
and UO_2 (O_2,N_24075,N_19547);
nor UO_3 (O_3,N_20712,N_24867);
or UO_4 (O_4,N_24301,N_21393);
nand UO_5 (O_5,N_24297,N_22413);
and UO_6 (O_6,N_24674,N_19638);
or UO_7 (O_7,N_21764,N_20109);
nor UO_8 (O_8,N_22308,N_18788);
nor UO_9 (O_9,N_22017,N_23041);
and UO_10 (O_10,N_22469,N_21846);
nand UO_11 (O_11,N_21179,N_24058);
nand UO_12 (O_12,N_22109,N_20007);
and UO_13 (O_13,N_20591,N_22801);
nand UO_14 (O_14,N_18997,N_20063);
or UO_15 (O_15,N_20596,N_23886);
xor UO_16 (O_16,N_23232,N_24994);
nand UO_17 (O_17,N_19084,N_22221);
and UO_18 (O_18,N_18758,N_22035);
xor UO_19 (O_19,N_24062,N_21932);
and UO_20 (O_20,N_20643,N_19966);
nor UO_21 (O_21,N_22423,N_19999);
nand UO_22 (O_22,N_22593,N_24208);
nor UO_23 (O_23,N_21675,N_20048);
and UO_24 (O_24,N_23540,N_24496);
nand UO_25 (O_25,N_20309,N_19258);
nand UO_26 (O_26,N_19913,N_21849);
or UO_27 (O_27,N_23358,N_24389);
nor UO_28 (O_28,N_22831,N_24683);
or UO_29 (O_29,N_18797,N_18925);
nand UO_30 (O_30,N_24762,N_19579);
or UO_31 (O_31,N_23266,N_22482);
nor UO_32 (O_32,N_24272,N_23103);
or UO_33 (O_33,N_24395,N_20069);
nor UO_34 (O_34,N_20363,N_24376);
or UO_35 (O_35,N_18852,N_24702);
and UO_36 (O_36,N_19811,N_21446);
or UO_37 (O_37,N_19301,N_21954);
or UO_38 (O_38,N_21170,N_24767);
xor UO_39 (O_39,N_20411,N_23624);
xnor UO_40 (O_40,N_24436,N_21200);
nor UO_41 (O_41,N_22274,N_21279);
nand UO_42 (O_42,N_19670,N_22425);
and UO_43 (O_43,N_22373,N_22323);
nor UO_44 (O_44,N_21079,N_18943);
nand UO_45 (O_45,N_19956,N_19327);
nor UO_46 (O_46,N_24919,N_19259);
nor UO_47 (O_47,N_22954,N_19420);
and UO_48 (O_48,N_22754,N_23872);
or UO_49 (O_49,N_21149,N_24267);
and UO_50 (O_50,N_20100,N_21231);
and UO_51 (O_51,N_22152,N_18848);
xnor UO_52 (O_52,N_20305,N_23117);
and UO_53 (O_53,N_24235,N_24789);
nand UO_54 (O_54,N_21616,N_24617);
nor UO_55 (O_55,N_24644,N_19789);
xnor UO_56 (O_56,N_22865,N_19433);
nor UO_57 (O_57,N_18813,N_24010);
and UO_58 (O_58,N_23815,N_19366);
and UO_59 (O_59,N_21361,N_20548);
nor UO_60 (O_60,N_21196,N_22355);
or UO_61 (O_61,N_22263,N_21374);
and UO_62 (O_62,N_20814,N_21907);
nor UO_63 (O_63,N_21888,N_21914);
nand UO_64 (O_64,N_22184,N_22023);
nor UO_65 (O_65,N_19632,N_23602);
nor UO_66 (O_66,N_22526,N_23067);
xnor UO_67 (O_67,N_22050,N_24055);
and UO_68 (O_68,N_19168,N_23464);
and UO_69 (O_69,N_20447,N_20239);
nand UO_70 (O_70,N_19263,N_23944);
and UO_71 (O_71,N_19198,N_23833);
xor UO_72 (O_72,N_20269,N_24465);
and UO_73 (O_73,N_24050,N_21514);
nor UO_74 (O_74,N_22694,N_21582);
or UO_75 (O_75,N_21229,N_24845);
nor UO_76 (O_76,N_22494,N_20810);
nand UO_77 (O_77,N_21745,N_21937);
nor UO_78 (O_78,N_24836,N_20292);
nor UO_79 (O_79,N_20738,N_20113);
nor UO_80 (O_80,N_18857,N_20682);
nand UO_81 (O_81,N_19431,N_19372);
nand UO_82 (O_82,N_20718,N_23056);
nand UO_83 (O_83,N_21873,N_24345);
and UO_84 (O_84,N_24823,N_22385);
xor UO_85 (O_85,N_23854,N_19663);
nor UO_86 (O_86,N_21776,N_20703);
xor UO_87 (O_87,N_19466,N_19523);
nand UO_88 (O_88,N_24794,N_24647);
or UO_89 (O_89,N_19088,N_21870);
or UO_90 (O_90,N_20646,N_18985);
and UO_91 (O_91,N_20138,N_20502);
nand UO_92 (O_92,N_24183,N_21795);
nand UO_93 (O_93,N_22443,N_21469);
nor UO_94 (O_94,N_22257,N_23859);
nand UO_95 (O_95,N_20369,N_20689);
xor UO_96 (O_96,N_21126,N_24390);
or UO_97 (O_97,N_23921,N_23714);
or UO_98 (O_98,N_19147,N_19878);
or UO_99 (O_99,N_24385,N_21023);
nand UO_100 (O_100,N_24689,N_22405);
or UO_101 (O_101,N_19584,N_20012);
or UO_102 (O_102,N_22293,N_19337);
nand UO_103 (O_103,N_18884,N_19480);
nor UO_104 (O_104,N_24853,N_21920);
or UO_105 (O_105,N_22275,N_20389);
nand UO_106 (O_106,N_22234,N_22852);
and UO_107 (O_107,N_23260,N_24810);
xor UO_108 (O_108,N_20800,N_19273);
or UO_109 (O_109,N_23591,N_23218);
nor UO_110 (O_110,N_19759,N_21842);
or UO_111 (O_111,N_23834,N_22468);
nand UO_112 (O_112,N_20938,N_21329);
and UO_113 (O_113,N_22097,N_21695);
nand UO_114 (O_114,N_20350,N_23814);
nor UO_115 (O_115,N_21669,N_22487);
xor UO_116 (O_116,N_22799,N_19234);
and UO_117 (O_117,N_19041,N_20412);
nand UO_118 (O_118,N_20526,N_20356);
nand UO_119 (O_119,N_19116,N_20788);
xor UO_120 (O_120,N_20910,N_22091);
nor UO_121 (O_121,N_22421,N_23380);
nor UO_122 (O_122,N_21479,N_20038);
or UO_123 (O_123,N_21533,N_21017);
or UO_124 (O_124,N_22939,N_19176);
nand UO_125 (O_125,N_24935,N_21255);
nor UO_126 (O_126,N_21995,N_20155);
nor UO_127 (O_127,N_20805,N_23630);
and UO_128 (O_128,N_21663,N_20264);
or UO_129 (O_129,N_24007,N_23954);
and UO_130 (O_130,N_22563,N_20937);
or UO_131 (O_131,N_23556,N_23076);
or UO_132 (O_132,N_21302,N_23100);
or UO_133 (O_133,N_23793,N_24338);
nor UO_134 (O_134,N_23632,N_23610);
xor UO_135 (O_135,N_19896,N_19861);
and UO_136 (O_136,N_23025,N_21878);
or UO_137 (O_137,N_23010,N_23482);
nand UO_138 (O_138,N_21004,N_19608);
nor UO_139 (O_139,N_20653,N_19774);
and UO_140 (O_140,N_20501,N_22656);
xor UO_141 (O_141,N_21890,N_19743);
nand UO_142 (O_142,N_19997,N_19024);
and UO_143 (O_143,N_23766,N_22816);
and UO_144 (O_144,N_23702,N_20694);
or UO_145 (O_145,N_23561,N_22684);
nor UO_146 (O_146,N_18869,N_19838);
nand UO_147 (O_147,N_23410,N_22905);
or UO_148 (O_148,N_18860,N_19413);
nor UO_149 (O_149,N_19143,N_20260);
nor UO_150 (O_150,N_23916,N_20115);
nor UO_151 (O_151,N_22340,N_21169);
nor UO_152 (O_152,N_21847,N_23284);
or UO_153 (O_153,N_20507,N_22796);
xor UO_154 (O_154,N_20234,N_21500);
nand UO_155 (O_155,N_20301,N_20806);
nor UO_156 (O_156,N_20439,N_22245);
nor UO_157 (O_157,N_22332,N_23652);
or UO_158 (O_158,N_22155,N_22927);
nand UO_159 (O_159,N_24956,N_18835);
nand UO_160 (O_160,N_24841,N_23760);
nand UO_161 (O_161,N_21307,N_21268);
or UO_162 (O_162,N_19639,N_21592);
or UO_163 (O_163,N_18954,N_21265);
and UO_164 (O_164,N_21584,N_23492);
or UO_165 (O_165,N_24808,N_23170);
or UO_166 (O_166,N_22216,N_20931);
and UO_167 (O_167,N_19318,N_22897);
and UO_168 (O_168,N_20750,N_21159);
nand UO_169 (O_169,N_23520,N_19531);
or UO_170 (O_170,N_21357,N_22010);
or UO_171 (O_171,N_24393,N_20908);
nor UO_172 (O_172,N_23106,N_24472);
nand UO_173 (O_173,N_24622,N_20986);
nand UO_174 (O_174,N_23631,N_19219);
nand UO_175 (O_175,N_21190,N_23345);
and UO_176 (O_176,N_22698,N_21397);
nor UO_177 (O_177,N_21778,N_19596);
nand UO_178 (O_178,N_24106,N_18955);
xor UO_179 (O_179,N_24260,N_21820);
nor UO_180 (O_180,N_20499,N_22807);
nand UO_181 (O_181,N_23213,N_24157);
nand UO_182 (O_182,N_20097,N_21175);
or UO_183 (O_183,N_23017,N_23767);
nor UO_184 (O_184,N_19817,N_23215);
or UO_185 (O_185,N_22864,N_23565);
or UO_186 (O_186,N_19892,N_24586);
or UO_187 (O_187,N_19158,N_22045);
xor UO_188 (O_188,N_24285,N_24462);
or UO_189 (O_189,N_18847,N_20261);
nor UO_190 (O_190,N_19825,N_24030);
nor UO_191 (O_191,N_24599,N_23034);
or UO_192 (O_192,N_20817,N_19625);
nand UO_193 (O_193,N_18762,N_21986);
or UO_194 (O_194,N_24502,N_21997);
nand UO_195 (O_195,N_23033,N_24961);
and UO_196 (O_196,N_23341,N_24950);
and UO_197 (O_197,N_22687,N_24121);
and UO_198 (O_198,N_23276,N_22933);
nor UO_199 (O_199,N_23882,N_24219);
or UO_200 (O_200,N_22614,N_21595);
and UO_201 (O_201,N_19524,N_22131);
or UO_202 (O_202,N_23523,N_24607);
and UO_203 (O_203,N_21762,N_23808);
nand UO_204 (O_204,N_24513,N_22146);
nor UO_205 (O_205,N_20206,N_23969);
and UO_206 (O_206,N_22895,N_23467);
or UO_207 (O_207,N_22439,N_18876);
nand UO_208 (O_208,N_20864,N_21390);
xnor UO_209 (O_209,N_23753,N_20397);
nand UO_210 (O_210,N_22298,N_20714);
nand UO_211 (O_211,N_23933,N_23537);
nand UO_212 (O_212,N_21713,N_21781);
or UO_213 (O_213,N_23008,N_19173);
nor UO_214 (O_214,N_23762,N_22959);
or UO_215 (O_215,N_23328,N_19631);
nand UO_216 (O_216,N_19474,N_24084);
and UO_217 (O_217,N_24669,N_24336);
nand UO_218 (O_218,N_18969,N_18894);
and UO_219 (O_219,N_23927,N_24437);
and UO_220 (O_220,N_21975,N_22832);
nor UO_221 (O_221,N_22726,N_22122);
nor UO_222 (O_222,N_19800,N_20642);
nor UO_223 (O_223,N_23583,N_24339);
nor UO_224 (O_224,N_22744,N_18948);
or UO_225 (O_225,N_23279,N_20154);
xor UO_226 (O_226,N_20713,N_19796);
or UO_227 (O_227,N_23183,N_23309);
xnor UO_228 (O_228,N_21074,N_24865);
nand UO_229 (O_229,N_18770,N_19945);
nor UO_230 (O_230,N_20594,N_22690);
nand UO_231 (O_231,N_18939,N_18972);
xnor UO_232 (O_232,N_22775,N_22032);
nand UO_233 (O_233,N_21771,N_21022);
and UO_234 (O_234,N_21142,N_20025);
and UO_235 (O_235,N_24282,N_24474);
nand UO_236 (O_236,N_21788,N_19814);
or UO_237 (O_237,N_24952,N_19768);
or UO_238 (O_238,N_24929,N_23127);
xor UO_239 (O_239,N_24250,N_24658);
nor UO_240 (O_240,N_23671,N_19356);
or UO_241 (O_241,N_23349,N_24141);
or UO_242 (O_242,N_19949,N_19029);
nor UO_243 (O_243,N_20583,N_23490);
nand UO_244 (O_244,N_21354,N_23163);
nand UO_245 (O_245,N_19298,N_19442);
or UO_246 (O_246,N_19752,N_24125);
or UO_247 (O_247,N_22403,N_23507);
nand UO_248 (O_248,N_23030,N_19943);
or UO_249 (O_249,N_22474,N_21092);
and UO_250 (O_250,N_24655,N_19499);
or UO_251 (O_251,N_19963,N_21915);
nand UO_252 (O_252,N_19912,N_21038);
nor UO_253 (O_253,N_21706,N_24374);
nor UO_254 (O_254,N_23242,N_19113);
xor UO_255 (O_255,N_22202,N_22024);
nand UO_256 (O_256,N_20423,N_19472);
nand UO_257 (O_257,N_23498,N_20276);
and UO_258 (O_258,N_19870,N_24163);
and UO_259 (O_259,N_19281,N_23454);
nor UO_260 (O_260,N_22608,N_23607);
or UO_261 (O_261,N_23891,N_21630);
xor UO_262 (O_262,N_19174,N_21666);
nor UO_263 (O_263,N_18755,N_21962);
and UO_264 (O_264,N_20459,N_24998);
nand UO_265 (O_265,N_23511,N_24812);
or UO_266 (O_266,N_21109,N_19765);
or UO_267 (O_267,N_21739,N_23670);
or UO_268 (O_268,N_21087,N_24680);
or UO_269 (O_269,N_23070,N_21144);
nor UO_270 (O_270,N_24917,N_21116);
or UO_271 (O_271,N_21330,N_22845);
or UO_272 (O_272,N_24608,N_22359);
or UO_273 (O_273,N_24850,N_18789);
nand UO_274 (O_274,N_19646,N_19773);
nand UO_275 (O_275,N_21931,N_20984);
and UO_276 (O_276,N_24298,N_21451);
or UO_277 (O_277,N_20228,N_19107);
nor UO_278 (O_278,N_20925,N_20809);
nor UO_279 (O_279,N_24415,N_22956);
nand UO_280 (O_280,N_24792,N_19206);
xnor UO_281 (O_281,N_23184,N_22064);
nor UO_282 (O_282,N_18964,N_21194);
nand UO_283 (O_283,N_21634,N_24127);
nand UO_284 (O_284,N_24790,N_20739);
and UO_285 (O_285,N_22696,N_24862);
nand UO_286 (O_286,N_20869,N_22885);
nor UO_287 (O_287,N_23364,N_20059);
or UO_288 (O_288,N_21902,N_20359);
or UO_289 (O_289,N_20517,N_23759);
or UO_290 (O_290,N_21122,N_20651);
nor UO_291 (O_291,N_20859,N_19192);
nor UO_292 (O_292,N_22736,N_22358);
nor UO_293 (O_293,N_21216,N_24601);
xnor UO_294 (O_294,N_22418,N_23210);
nand UO_295 (O_295,N_18844,N_20953);
nand UO_296 (O_296,N_19929,N_20119);
or UO_297 (O_297,N_21204,N_21345);
nand UO_298 (O_298,N_24198,N_20926);
nand UO_299 (O_299,N_21935,N_21039);
and UO_300 (O_300,N_23515,N_22366);
nor UO_301 (O_301,N_24284,N_19255);
and UO_302 (O_302,N_20999,N_24604);
or UO_303 (O_303,N_20802,N_19724);
or UO_304 (O_304,N_22853,N_24726);
or UO_305 (O_305,N_23443,N_21948);
and UO_306 (O_306,N_19660,N_24426);
nand UO_307 (O_307,N_20153,N_20328);
nand UO_308 (O_308,N_22001,N_23627);
or UO_309 (O_309,N_21515,N_22942);
or UO_310 (O_310,N_23155,N_22923);
and UO_311 (O_311,N_23636,N_24510);
nor UO_312 (O_312,N_22868,N_19766);
nand UO_313 (O_313,N_23227,N_19621);
or UO_314 (O_314,N_23771,N_24087);
nand UO_315 (O_315,N_22795,N_23222);
and UO_316 (O_316,N_24673,N_21277);
nand UO_317 (O_317,N_19441,N_24334);
or UO_318 (O_318,N_20665,N_22028);
xnor UO_319 (O_319,N_23468,N_21972);
or UO_320 (O_320,N_18864,N_23057);
and UO_321 (O_321,N_22518,N_20799);
nand UO_322 (O_322,N_22241,N_20491);
and UO_323 (O_323,N_20798,N_24944);
nor UO_324 (O_324,N_24581,N_19676);
xor UO_325 (O_325,N_21601,N_19790);
nor UO_326 (O_326,N_22349,N_21893);
nor UO_327 (O_327,N_23174,N_23091);
nand UO_328 (O_328,N_22603,N_22396);
nor UO_329 (O_329,N_19244,N_19548);
nand UO_330 (O_330,N_22128,N_24572);
xnor UO_331 (O_331,N_19037,N_21976);
or UO_332 (O_332,N_21084,N_22722);
and UO_333 (O_333,N_21650,N_22640);
nor UO_334 (O_334,N_23480,N_23974);
or UO_335 (O_335,N_24748,N_23699);
nor UO_336 (O_336,N_23893,N_21368);
nor UO_337 (O_337,N_24066,N_18937);
nor UO_338 (O_338,N_21969,N_20108);
and UO_339 (O_339,N_22090,N_22305);
nor UO_340 (O_340,N_18913,N_24981);
and UO_341 (O_341,N_21955,N_22512);
nand UO_342 (O_342,N_21383,N_20701);
nor UO_343 (O_343,N_18968,N_19783);
and UO_344 (O_344,N_22579,N_23271);
nand UO_345 (O_345,N_19277,N_22306);
or UO_346 (O_346,N_20024,N_23423);
or UO_347 (O_347,N_18980,N_20962);
and UO_348 (O_348,N_22107,N_23798);
and UO_349 (O_349,N_20963,N_24053);
nand UO_350 (O_350,N_20341,N_23653);
nor UO_351 (O_351,N_19716,N_22337);
or UO_352 (O_352,N_24276,N_19730);
or UO_353 (O_353,N_24940,N_24730);
nand UO_354 (O_354,N_22963,N_19726);
xor UO_355 (O_355,N_19391,N_22438);
or UO_356 (O_356,N_21574,N_19935);
nand UO_357 (O_357,N_23246,N_22536);
or UO_358 (O_358,N_23367,N_24154);
and UO_359 (O_359,N_23340,N_24686);
and UO_360 (O_360,N_24356,N_23288);
and UO_361 (O_361,N_20277,N_20014);
nand UO_362 (O_362,N_18772,N_19846);
or UO_363 (O_363,N_20275,N_24980);
nand UO_364 (O_364,N_22891,N_20466);
or UO_365 (O_365,N_24490,N_20374);
nand UO_366 (O_366,N_23665,N_23118);
xnor UO_367 (O_367,N_21271,N_24086);
xnor UO_368 (O_368,N_22573,N_19236);
and UO_369 (O_369,N_21562,N_22909);
nand UO_370 (O_370,N_20479,N_24482);
xnor UO_371 (O_371,N_22917,N_18883);
nand UO_372 (O_372,N_23822,N_22078);
nand UO_373 (O_373,N_24147,N_22772);
and UO_374 (O_374,N_20855,N_21363);
or UO_375 (O_375,N_20598,N_24216);
nor UO_376 (O_376,N_24924,N_24223);
or UO_377 (O_377,N_22653,N_18927);
or UO_378 (O_378,N_22611,N_20998);
nor UO_379 (O_379,N_21798,N_22598);
or UO_380 (O_380,N_20890,N_24857);
nor UO_381 (O_381,N_21911,N_20948);
or UO_382 (O_382,N_23153,N_19426);
and UO_383 (O_383,N_22618,N_23721);
or UO_384 (O_384,N_19493,N_19640);
and UO_385 (O_385,N_24238,N_24570);
or UO_386 (O_386,N_22871,N_21703);
or UO_387 (O_387,N_24380,N_21880);
and UO_388 (O_388,N_20238,N_22681);
and UO_389 (O_389,N_21026,N_21884);
and UO_390 (O_390,N_21230,N_24975);
and UO_391 (O_391,N_23790,N_23357);
nor UO_392 (O_392,N_21989,N_20819);
and UO_393 (O_393,N_19951,N_21490);
and UO_394 (O_394,N_23749,N_22743);
and UO_395 (O_395,N_24469,N_19847);
nor UO_396 (O_396,N_22977,N_20784);
nand UO_397 (O_397,N_21202,N_20876);
or UO_398 (O_398,N_21530,N_21389);
and UO_399 (O_399,N_19105,N_21001);
and UO_400 (O_400,N_23533,N_21481);
nand UO_401 (O_401,N_22084,N_24544);
nor UO_402 (O_402,N_19863,N_19598);
nor UO_403 (O_403,N_23092,N_23737);
or UO_404 (O_404,N_24384,N_22367);
xor UO_405 (O_405,N_22372,N_21544);
xor UO_406 (O_406,N_23880,N_20372);
xor UO_407 (O_407,N_20270,N_22935);
and UO_408 (O_408,N_22544,N_20595);
or UO_409 (O_409,N_19957,N_19611);
nor UO_410 (O_410,N_20314,N_22451);
nand UO_411 (O_411,N_19042,N_19060);
nor UO_412 (O_412,N_23786,N_20046);
nor UO_413 (O_413,N_19486,N_23298);
and UO_414 (O_414,N_24365,N_22582);
nor UO_415 (O_415,N_21964,N_19934);
nand UO_416 (O_416,N_18756,N_23383);
nor UO_417 (O_417,N_22502,N_23449);
nand UO_418 (O_418,N_24441,N_21783);
nor UO_419 (O_419,N_20271,N_20451);
nor UO_420 (O_420,N_21661,N_21339);
xnor UO_421 (O_421,N_24577,N_22719);
or UO_422 (O_422,N_23292,N_21898);
or UO_423 (O_423,N_23501,N_19291);
and UO_424 (O_424,N_20352,N_19497);
nand UO_425 (O_425,N_22409,N_24180);
nand UO_426 (O_426,N_24871,N_21266);
or UO_427 (O_427,N_23861,N_20061);
nand UO_428 (O_428,N_20253,N_24910);
or UO_429 (O_429,N_20203,N_21258);
or UO_430 (O_430,N_19534,N_21919);
nand UO_431 (O_431,N_20959,N_23144);
nor UO_432 (O_432,N_19001,N_20807);
nand UO_433 (O_433,N_19705,N_18872);
or UO_434 (O_434,N_23447,N_23804);
nand UO_435 (O_435,N_20149,N_19858);
nand UO_436 (O_436,N_23018,N_22918);
nand UO_437 (O_437,N_22191,N_23796);
and UO_438 (O_438,N_21747,N_22183);
xor UO_439 (O_439,N_22075,N_24511);
or UO_440 (O_440,N_24971,N_24880);
and UO_441 (O_441,N_19996,N_20398);
and UO_442 (O_442,N_21212,N_23505);
and UO_443 (O_443,N_19224,N_20143);
or UO_444 (O_444,N_24671,N_24034);
and UO_445 (O_445,N_24012,N_21575);
nand UO_446 (O_446,N_19344,N_23356);
and UO_447 (O_447,N_19848,N_24771);
or UO_448 (O_448,N_19262,N_24909);
and UO_449 (O_449,N_21934,N_22448);
nand UO_450 (O_450,N_22988,N_20354);
or UO_451 (O_451,N_24040,N_23128);
nand UO_452 (O_452,N_21335,N_21647);
nor UO_453 (O_453,N_21016,N_23419);
or UO_454 (O_454,N_24552,N_22609);
xor UO_455 (O_455,N_19837,N_22440);
xnor UO_456 (O_456,N_21447,N_22125);
xor UO_457 (O_457,N_20462,N_24884);
and UO_458 (O_458,N_24005,N_23952);
nand UO_459 (O_459,N_21894,N_21572);
and UO_460 (O_460,N_20762,N_24768);
or UO_461 (O_461,N_24592,N_22251);
xor UO_462 (O_462,N_21014,N_21106);
or UO_463 (O_463,N_23970,N_19215);
or UO_464 (O_464,N_21596,N_19756);
nor UO_465 (O_465,N_24931,N_24772);
nand UO_466 (O_466,N_24269,N_21567);
nor UO_467 (O_467,N_21879,N_23840);
nand UO_468 (O_468,N_24100,N_23313);
or UO_469 (O_469,N_20569,N_20322);
nor UO_470 (O_470,N_23172,N_21114);
nor UO_471 (O_471,N_19542,N_21631);
xnor UO_472 (O_472,N_21951,N_24951);
xor UO_473 (O_473,N_21498,N_23105);
nand UO_474 (O_474,N_23810,N_23877);
or UO_475 (O_475,N_20641,N_18784);
or UO_476 (O_476,N_21484,N_19960);
nand UO_477 (O_477,N_23794,N_22670);
nand UO_478 (O_478,N_21509,N_24933);
and UO_479 (O_479,N_23735,N_22560);
or UO_480 (O_480,N_21396,N_22546);
nor UO_481 (O_481,N_23677,N_20834);
or UO_482 (O_482,N_21233,N_19958);
and UO_483 (O_483,N_22974,N_23757);
nand UO_484 (O_484,N_23578,N_23945);
nor UO_485 (O_485,N_22397,N_21243);
and UO_486 (O_486,N_20934,N_22786);
nor UO_487 (O_487,N_19217,N_24964);
nor UO_488 (O_488,N_23712,N_21709);
nor UO_489 (O_489,N_24700,N_22718);
nand UO_490 (O_490,N_21378,N_21725);
xor UO_491 (O_491,N_19894,N_24203);
nand UO_492 (O_492,N_19127,N_24143);
or UO_493 (O_493,N_19229,N_22822);
xnor UO_494 (O_494,N_23307,N_24028);
or UO_495 (O_495,N_19475,N_19136);
and UO_496 (O_496,N_22995,N_24535);
or UO_497 (O_497,N_24049,N_21164);
and UO_498 (O_498,N_24728,N_20041);
and UO_499 (O_499,N_19564,N_20773);
nor UO_500 (O_500,N_20733,N_19799);
nand UO_501 (O_501,N_19414,N_19066);
and UO_502 (O_502,N_19877,N_20376);
nor UO_503 (O_503,N_24512,N_22713);
or UO_504 (O_504,N_23637,N_20939);
nor UO_505 (O_505,N_19794,N_23590);
nand UO_506 (O_506,N_21585,N_19137);
or UO_507 (O_507,N_20645,N_18839);
and UO_508 (O_508,N_19227,N_22230);
or UO_509 (O_509,N_24863,N_20637);
nor UO_510 (O_510,N_23216,N_20630);
or UO_511 (O_511,N_21576,N_24116);
nor UO_512 (O_512,N_21333,N_24675);
or UO_513 (O_513,N_24286,N_21323);
or UO_514 (O_514,N_21154,N_21994);
nand UO_515 (O_515,N_24230,N_23154);
nor UO_516 (O_516,N_23598,N_20988);
nor UO_517 (O_517,N_23680,N_22641);
nand UO_518 (O_518,N_19321,N_24126);
nand UO_519 (O_519,N_21464,N_22334);
or UO_520 (O_520,N_21786,N_24188);
or UO_521 (O_521,N_19040,N_19944);
nor UO_522 (O_522,N_21423,N_20961);
or UO_523 (O_523,N_21441,N_24885);
nand UO_524 (O_524,N_21598,N_24400);
nor UO_525 (O_525,N_18929,N_24947);
or UO_526 (O_526,N_22163,N_21727);
and UO_527 (O_527,N_22051,N_22511);
or UO_528 (O_528,N_20302,N_21228);
or UO_529 (O_529,N_19099,N_22347);
and UO_530 (O_530,N_21403,N_24283);
and UO_531 (O_531,N_20408,N_19252);
nand UO_532 (O_532,N_23263,N_19855);
or UO_533 (O_533,N_20922,N_24263);
or UO_534 (O_534,N_21968,N_22769);
and UO_535 (O_535,N_22287,N_20036);
nand UO_536 (O_536,N_22011,N_24195);
nor UO_537 (O_537,N_24322,N_19354);
or UO_538 (O_538,N_24859,N_21273);
nand UO_539 (O_539,N_24588,N_19429);
nor UO_540 (O_540,N_19339,N_21413);
or UO_541 (O_541,N_22826,N_21220);
nand UO_542 (O_542,N_21181,N_20344);
or UO_543 (O_543,N_23539,N_24806);
and UO_544 (O_544,N_22790,N_24002);
and UO_545 (O_545,N_20405,N_19423);
and UO_546 (O_546,N_22140,N_22843);
nor UO_547 (O_547,N_23428,N_24388);
nor UO_548 (O_548,N_23059,N_24044);
or UO_549 (O_549,N_22180,N_21431);
and UO_550 (O_550,N_21215,N_23685);
or UO_551 (O_551,N_19378,N_23301);
and UO_552 (O_552,N_21205,N_24838);
or UO_553 (O_553,N_19562,N_24559);
nand UO_554 (O_554,N_20393,N_23426);
or UO_555 (O_555,N_22061,N_22406);
and UO_556 (O_556,N_19507,N_21434);
and UO_557 (O_557,N_24457,N_19775);
nand UO_558 (O_558,N_22415,N_20870);
and UO_559 (O_559,N_23729,N_21201);
or UO_560 (O_560,N_23711,N_22950);
and UO_561 (O_561,N_24009,N_21387);
nor UO_562 (O_562,N_22254,N_21254);
nand UO_563 (O_563,N_24015,N_22492);
and UO_564 (O_564,N_22490,N_23188);
nor UO_565 (O_565,N_19854,N_22758);
or UO_566 (O_566,N_20213,N_19888);
nor UO_567 (O_567,N_21055,N_23165);
and UO_568 (O_568,N_19388,N_18766);
nor UO_569 (O_569,N_19182,N_19427);
or UO_570 (O_570,N_20446,N_20603);
nand UO_571 (O_571,N_19435,N_19605);
nor UO_572 (O_572,N_23087,N_20457);
and UO_573 (O_573,N_24209,N_20697);
or UO_574 (O_574,N_24366,N_22198);
xnor UO_575 (O_575,N_24755,N_21163);
or UO_576 (O_576,N_20445,N_18888);
nor UO_577 (O_577,N_22206,N_21622);
xor UO_578 (O_578,N_19241,N_19525);
nor UO_579 (O_579,N_22411,N_21086);
or UO_580 (O_580,N_24618,N_23414);
and UO_581 (O_581,N_22712,N_20853);
nand UO_582 (O_582,N_23881,N_20066);
or UO_583 (O_583,N_22734,N_24882);
xor UO_584 (O_584,N_21527,N_23803);
and UO_585 (O_585,N_20165,N_22803);
and UO_586 (O_586,N_18991,N_21837);
or UO_587 (O_587,N_24632,N_20118);
xnor UO_588 (O_588,N_23534,N_24459);
or UO_589 (O_589,N_24417,N_20312);
nor UO_590 (O_590,N_24732,N_22095);
nor UO_591 (O_591,N_19094,N_24184);
nor UO_592 (O_592,N_19589,N_24760);
nand UO_593 (O_593,N_22931,N_23335);
and UO_594 (O_594,N_23255,N_22297);
or UO_595 (O_595,N_20485,N_23248);
or UO_596 (O_596,N_18841,N_20333);
nor UO_597 (O_597,N_20081,N_24358);
nor UO_598 (O_598,N_20087,N_20174);
or UO_599 (O_599,N_23205,N_22009);
and UO_600 (O_600,N_20690,N_24346);
and UO_601 (O_601,N_24699,N_19309);
and UO_602 (O_602,N_20137,N_19090);
nor UO_603 (O_603,N_18780,N_20324);
and UO_604 (O_604,N_21473,N_22624);
and UO_605 (O_605,N_23466,N_24977);
and UO_606 (O_606,N_19307,N_23422);
and UO_607 (O_607,N_22928,N_23199);
or UO_608 (O_608,N_24778,N_20198);
or UO_609 (O_609,N_19463,N_24450);
nand UO_610 (O_610,N_19221,N_20547);
nor UO_611 (O_611,N_23016,N_19314);
nand UO_612 (O_612,N_19563,N_20387);
nand UO_613 (O_613,N_22747,N_21037);
nor UO_614 (O_614,N_19939,N_23618);
and UO_615 (O_615,N_24557,N_22232);
or UO_616 (O_616,N_23640,N_19648);
nor UO_617 (O_617,N_24996,N_20818);
and UO_618 (O_618,N_22629,N_23698);
and UO_619 (O_619,N_23541,N_19494);
nand UO_620 (O_620,N_21612,N_20424);
nand UO_621 (O_621,N_19897,N_24239);
nor UO_622 (O_622,N_18854,N_20555);
and UO_623 (O_623,N_21063,N_21684);
nor UO_624 (O_624,N_24307,N_19628);
nand UO_625 (O_625,N_19816,N_21863);
and UO_626 (O_626,N_20563,N_21714);
nand UO_627 (O_627,N_20418,N_19249);
nor UO_628 (O_628,N_21723,N_18771);
nor UO_629 (O_629,N_22112,N_21824);
xnor UO_630 (O_630,N_22063,N_21104);
or UO_631 (O_631,N_19432,N_23772);
or UO_632 (O_632,N_19578,N_23312);
nor UO_633 (O_633,N_24386,N_22505);
nor UO_634 (O_634,N_23024,N_23542);
and UO_635 (O_635,N_19689,N_18875);
and UO_636 (O_636,N_18936,N_23936);
or UO_637 (O_637,N_20022,N_24063);
and UO_638 (O_638,N_24793,N_24887);
or UO_639 (O_639,N_19380,N_20873);
and UO_640 (O_640,N_18805,N_22621);
and UO_641 (O_641,N_19447,N_24036);
or UO_642 (O_642,N_19211,N_19017);
and UO_643 (O_643,N_22904,N_21272);
nor UO_644 (O_644,N_21281,N_22806);
and UO_645 (O_645,N_20947,N_18816);
and UO_646 (O_646,N_18910,N_23930);
nand UO_647 (O_647,N_21152,N_21791);
xor UO_648 (O_648,N_24955,N_23378);
nor UO_649 (O_649,N_24396,N_18833);
nor UO_650 (O_650,N_24442,N_24361);
and UO_651 (O_651,N_21280,N_20592);
or UO_652 (O_652,N_21736,N_23156);
nor UO_653 (O_653,N_20654,N_23268);
or UO_654 (O_654,N_23826,N_19925);
or UO_655 (O_655,N_21301,N_19142);
or UO_656 (O_656,N_24061,N_20375);
or UO_657 (O_657,N_24247,N_21415);
or UO_658 (O_658,N_21865,N_20029);
nand UO_659 (O_659,N_20565,N_20862);
and UO_660 (O_660,N_23362,N_18983);
nor UO_661 (O_661,N_22794,N_18790);
nor UO_662 (O_662,N_21029,N_20628);
and UO_663 (O_663,N_18862,N_23332);
or UO_664 (O_664,N_21529,N_20146);
nand UO_665 (O_665,N_21691,N_20020);
or UO_666 (O_666,N_21685,N_19723);
nor UO_667 (O_667,N_22196,N_21465);
or UO_668 (O_668,N_21318,N_22833);
xor UO_669 (O_669,N_24712,N_20659);
or UO_670 (O_670,N_19819,N_20205);
or UO_671 (O_671,N_19591,N_19362);
nand UO_672 (O_672,N_24350,N_19446);
nor UO_673 (O_673,N_19843,N_23845);
or UO_674 (O_674,N_21250,N_24019);
nor UO_675 (O_675,N_20559,N_22631);
or UO_676 (O_676,N_24470,N_22315);
nor UO_677 (O_677,N_21147,N_20527);
xnor UO_678 (O_678,N_22761,N_20704);
or UO_679 (O_679,N_24029,N_21681);
xnor UO_680 (O_680,N_18815,N_22626);
or UO_681 (O_681,N_23713,N_24295);
or UO_682 (O_682,N_23303,N_19928);
xnor UO_683 (O_683,N_19376,N_20413);
xnor UO_684 (O_684,N_19351,N_24288);
and UO_685 (O_685,N_22062,N_23251);
or UO_686 (O_686,N_19469,N_24418);
nand UO_687 (O_687,N_24636,N_24439);
nor UO_688 (O_688,N_21047,N_24508);
or UO_689 (O_689,N_23250,N_19069);
nor UO_690 (O_690,N_22160,N_23506);
xnor UO_691 (O_691,N_18942,N_19379);
xor UO_692 (O_692,N_22660,N_24266);
and UO_693 (O_693,N_19609,N_23141);
or UO_694 (O_694,N_21297,N_19641);
or UO_695 (O_695,N_20223,N_21445);
nand UO_696 (O_696,N_24659,N_18990);
or UO_697 (O_697,N_20500,N_20161);
nand UO_698 (O_698,N_23875,N_21508);
and UO_699 (O_699,N_20506,N_22244);
or UO_700 (O_700,N_24970,N_19149);
xnor UO_701 (O_701,N_22764,N_22079);
nor UO_702 (O_702,N_24896,N_20151);
nand UO_703 (O_703,N_24852,N_20018);
or UO_704 (O_704,N_20972,N_23249);
and UO_705 (O_705,N_21236,N_19830);
nor UO_706 (O_706,N_19851,N_18909);
and UO_707 (O_707,N_22893,N_22217);
or UO_708 (O_708,N_24670,N_21000);
and UO_709 (O_709,N_22089,N_21343);
or UO_710 (O_710,N_23582,N_21662);
nand UO_711 (O_711,N_23950,N_19313);
nor UO_712 (O_712,N_23646,N_22975);
and UO_713 (O_713,N_24079,N_21558);
nand UO_714 (O_714,N_22086,N_23190);
or UO_715 (O_715,N_23589,N_22985);
xor UO_716 (O_716,N_23728,N_22788);
and UO_717 (O_717,N_19947,N_22226);
or UO_718 (O_718,N_22111,N_19141);
or UO_719 (O_719,N_21551,N_23734);
and UO_720 (O_720,N_22185,N_22302);
nor UO_721 (O_721,N_19653,N_21751);
and UO_722 (O_722,N_24801,N_24523);
and UO_723 (O_723,N_20743,N_22798);
nand UO_724 (O_724,N_20943,N_22255);
and UO_725 (O_725,N_21299,N_19271);
nor UO_726 (O_726,N_23320,N_23740);
and UO_727 (O_727,N_21814,N_19043);
and UO_728 (O_728,N_21524,N_21720);
xnor UO_729 (O_729,N_24703,N_21070);
nand UO_730 (O_730,N_23855,N_23717);
xor UO_731 (O_731,N_18973,N_19642);
nand UO_732 (O_732,N_24256,N_23557);
nand UO_733 (O_733,N_21131,N_22265);
and UO_734 (O_734,N_18928,N_18995);
nor UO_735 (O_735,N_22386,N_19284);
and UO_736 (O_736,N_21525,N_19189);
or UO_737 (O_737,N_22678,N_22797);
nor UO_738 (O_738,N_21502,N_21646);
nand UO_739 (O_739,N_21545,N_20175);
or UO_740 (O_740,N_23075,N_23524);
nand UO_741 (O_741,N_20804,N_20226);
or UO_742 (O_742,N_22751,N_24681);
nand UO_743 (O_743,N_19842,N_18779);
nor UO_744 (O_744,N_22981,N_21629);
or UO_745 (O_745,N_20104,N_21119);
xor UO_746 (O_746,N_19436,N_19006);
or UO_747 (O_747,N_22834,N_24739);
nand UO_748 (O_748,N_24411,N_23832);
and UO_749 (O_749,N_20460,N_23236);
and UO_750 (O_750,N_21077,N_24488);
or UO_751 (O_751,N_22471,N_22344);
or UO_752 (O_752,N_23563,N_19719);
nand UO_753 (O_753,N_20034,N_24661);
nand UO_754 (O_754,N_19686,N_21436);
xor UO_755 (O_755,N_21471,N_22116);
nand UO_756 (O_756,N_21938,N_22307);
nor UO_757 (O_757,N_22984,N_21260);
or UO_758 (O_758,N_22676,N_20378);
nand UO_759 (O_759,N_24353,N_22514);
nor UO_760 (O_760,N_23956,N_22683);
xor UO_761 (O_761,N_24568,N_18782);
or UO_762 (O_762,N_22994,N_20147);
nor UO_763 (O_763,N_22416,N_21577);
and UO_764 (O_764,N_21184,N_24567);
xnor UO_765 (O_765,N_20842,N_22219);
or UO_766 (O_766,N_22291,N_22919);
or UO_767 (O_767,N_23837,N_22783);
or UO_768 (O_768,N_20588,N_21493);
or UO_769 (O_769,N_23823,N_24109);
nand UO_770 (O_770,N_19728,N_24046);
nor UO_771 (O_771,N_21304,N_20032);
and UO_772 (O_772,N_23682,N_19681);
xor UO_773 (O_773,N_20557,N_22130);
or UO_774 (O_774,N_21328,N_23894);
and UO_775 (O_775,N_23391,N_18777);
and UO_776 (O_776,N_21953,N_22674);
nor UO_777 (O_777,N_19590,N_21827);
nand UO_778 (O_778,N_19355,N_22320);
nand UO_779 (O_779,N_20662,N_23816);
and UO_780 (O_780,N_23197,N_21283);
or UO_781 (O_781,N_22153,N_24821);
or UO_782 (O_782,N_20663,N_21806);
and UO_783 (O_783,N_20043,N_24554);
and UO_784 (O_784,N_19096,N_22628);
or UO_785 (O_785,N_19079,N_19390);
nor UO_786 (O_786,N_23139,N_23159);
nor UO_787 (O_787,N_19108,N_24162);
or UO_788 (O_788,N_22938,N_22577);
nand UO_789 (O_789,N_22780,N_20370);
and UO_790 (O_790,N_24813,N_24185);
and UO_791 (O_791,N_19574,N_23453);
or UO_792 (O_792,N_19100,N_19991);
xor UO_793 (O_793,N_19083,N_19288);
nor UO_794 (O_794,N_23939,N_20306);
nand UO_795 (O_795,N_21552,N_21606);
nor UO_796 (O_796,N_23966,N_23874);
nor UO_797 (O_797,N_22414,N_22019);
or UO_798 (O_798,N_23107,N_19214);
xor UO_799 (O_799,N_23243,N_20649);
and UO_800 (O_800,N_20236,N_21282);
or UO_801 (O_801,N_20135,N_19613);
nor UO_802 (O_802,N_22508,N_20878);
or UO_803 (O_803,N_20207,N_20741);
nor UO_804 (O_804,N_22335,N_20783);
nand UO_805 (O_805,N_20140,N_24501);
or UO_806 (O_806,N_18868,N_22071);
and UO_807 (O_807,N_20158,N_23194);
and UO_808 (O_808,N_20550,N_23596);
nand UO_809 (O_809,N_20317,N_22958);
nand UO_810 (O_810,N_19157,N_20102);
nand UO_811 (O_811,N_20872,N_22708);
nor UO_812 (O_812,N_23503,N_20184);
nand UO_813 (O_813,N_20077,N_21470);
and UO_814 (O_814,N_24693,N_22154);
nor UO_815 (O_815,N_19286,N_20556);
and UO_816 (O_816,N_24811,N_19328);
or UO_817 (O_817,N_21660,N_22225);
and UO_818 (O_818,N_23623,N_22352);
and UO_819 (O_819,N_21729,N_21550);
and UO_820 (O_820,N_23252,N_22319);
or UO_821 (O_821,N_23280,N_22968);
or UO_822 (O_822,N_21866,N_19246);
and UO_823 (O_823,N_24805,N_21665);
or UO_824 (O_824,N_19687,N_21350);
and UO_825 (O_825,N_23707,N_22652);
or UO_826 (O_826,N_20830,N_23071);
and UO_827 (O_827,N_18897,N_21054);
and UO_828 (O_828,N_19014,N_19635);
and UO_829 (O_829,N_20579,N_21043);
nor UO_830 (O_830,N_23972,N_19603);
nor UO_831 (O_831,N_22632,N_18793);
nand UO_832 (O_832,N_21936,N_19265);
and UO_833 (O_833,N_20431,N_19065);
nor UO_834 (O_834,N_23658,N_23850);
and UO_835 (O_835,N_20037,N_20503);
nand UO_836 (O_836,N_19509,N_23876);
and UO_837 (O_837,N_19057,N_18920);
and UO_838 (O_838,N_21442,N_20148);
and UO_839 (O_839,N_24171,N_24540);
nand UO_840 (O_840,N_23078,N_19489);
and UO_841 (O_841,N_22143,N_21796);
xnor UO_842 (O_842,N_24445,N_22951);
nor UO_843 (O_843,N_23634,N_24685);
nor UO_844 (O_844,N_22589,N_23704);
nor UO_845 (O_845,N_19154,N_24915);
or UO_846 (O_846,N_19845,N_20789);
or UO_847 (O_847,N_23379,N_19829);
nand UO_848 (O_848,N_19932,N_22325);
nand UO_849 (O_849,N_20060,N_23705);
nand UO_850 (O_850,N_24521,N_20044);
nand UO_851 (O_851,N_23581,N_19502);
nor UO_852 (O_852,N_19936,N_23369);
nor UO_853 (O_853,N_22498,N_21672);
or UO_854 (O_854,N_24816,N_22311);
and UO_855 (O_855,N_22817,N_23095);
nor UO_856 (O_856,N_23111,N_22213);
nor UO_857 (O_857,N_24132,N_19086);
and UO_858 (O_858,N_19655,N_23011);
or UO_859 (O_859,N_20257,N_20636);
and UO_860 (O_860,N_19471,N_21908);
nor UO_861 (O_861,N_19541,N_24562);
nor UO_862 (O_862,N_19012,N_22663);
and UO_863 (O_863,N_22752,N_24927);
nor UO_864 (O_864,N_20026,N_21240);
nor UO_865 (O_865,N_20086,N_20991);
xnor UO_866 (O_866,N_22164,N_23764);
nor UO_867 (O_867,N_22874,N_24763);
nor UO_868 (O_868,N_22215,N_19727);
and UO_869 (O_869,N_19092,N_19401);
nand UO_870 (O_870,N_21700,N_19979);
nor UO_871 (O_871,N_24543,N_21810);
nor UO_872 (O_872,N_22496,N_21214);
nor UO_873 (O_873,N_19806,N_24281);
or UO_874 (O_874,N_20284,N_23483);
and UO_875 (O_875,N_20828,N_24024);
or UO_876 (O_876,N_22489,N_22570);
or UO_877 (O_877,N_23878,N_21366);
nor UO_878 (O_878,N_18787,N_22515);
nand UO_879 (O_879,N_22310,N_24820);
nor UO_880 (O_880,N_21083,N_21158);
and UO_881 (O_881,N_23809,N_24299);
or UO_882 (O_882,N_21988,N_19439);
nand UO_883 (O_883,N_20520,N_23259);
and UO_884 (O_884,N_20366,N_21787);
and UO_885 (O_885,N_19114,N_21373);
nand UO_886 (O_886,N_24134,N_21716);
and UO_887 (O_887,N_20785,N_23026);
and UO_888 (O_888,N_18981,N_24017);
nor UO_889 (O_889,N_21850,N_22279);
and UO_890 (O_890,N_23436,N_22840);
or UO_891 (O_891,N_23645,N_22920);
or UO_892 (O_892,N_22277,N_24207);
or UO_893 (O_893,N_19400,N_23747);
nand UO_894 (O_894,N_20776,N_23385);
nand UO_895 (O_895,N_21604,N_19782);
nor UO_896 (O_896,N_23696,N_23151);
and UO_897 (O_897,N_24735,N_21717);
and UO_898 (O_898,N_23072,N_19821);
nor UO_899 (O_899,N_19778,N_20316);
or UO_900 (O_900,N_23985,N_24795);
and UO_901 (O_901,N_18824,N_24443);
nand UO_902 (O_902,N_21557,N_23684);
nand UO_903 (O_903,N_20202,N_23412);
or UO_904 (O_904,N_20541,N_19988);
and UO_905 (O_905,N_23007,N_18908);
nand UO_906 (O_906,N_20681,N_23406);
nand UO_907 (O_907,N_21680,N_20896);
nand UO_908 (O_908,N_23867,N_20062);
and UO_909 (O_909,N_21334,N_19891);
xnor UO_910 (O_910,N_22564,N_22706);
and UO_911 (O_911,N_21696,N_21005);
xnor UO_912 (O_912,N_20346,N_22092);
or UO_913 (O_913,N_20181,N_23355);
or UO_914 (O_914,N_21391,N_19011);
nor UO_915 (O_915,N_23600,N_24452);
nor UO_916 (O_916,N_19018,N_23976);
and UO_917 (O_917,N_20224,N_23293);
or UO_918 (O_918,N_20906,N_20683);
xor UO_919 (O_919,N_24637,N_21803);
and UO_920 (O_920,N_20467,N_19005);
nor UO_921 (O_921,N_18881,N_21025);
and UO_922 (O_922,N_21353,N_19212);
nor UO_923 (O_923,N_21439,N_19438);
nor UO_924 (O_924,N_18893,N_20120);
nand UO_925 (O_925,N_20587,N_22638);
and UO_926 (O_926,N_24268,N_23439);
and UO_927 (O_927,N_19931,N_20954);
and UO_928 (O_928,N_19552,N_22401);
nand UO_929 (O_929,N_22088,N_22188);
xnor UO_930 (O_930,N_20377,N_23217);
nand UO_931 (O_931,N_20340,N_20955);
nor UO_932 (O_932,N_19968,N_20008);
xor UO_933 (O_933,N_22800,N_24477);
nor UO_934 (O_934,N_20742,N_21293);
nor UO_935 (O_935,N_19964,N_19076);
xor UO_936 (O_936,N_21499,N_20676);
or UO_937 (O_937,N_22742,N_23318);
and UO_938 (O_938,N_24217,N_21452);
nor UO_939 (O_939,N_22876,N_23228);
xnor UO_940 (O_940,N_21712,N_20249);
or UO_941 (O_941,N_22646,N_24253);
or UO_942 (O_942,N_22280,N_24144);
nand UO_943 (O_943,N_22375,N_20671);
and UO_944 (O_944,N_21495,N_24547);
xor UO_945 (O_945,N_22149,N_20106);
nor UO_946 (O_946,N_23452,N_21587);
nor UO_947 (O_947,N_22535,N_21658);
and UO_948 (O_948,N_24566,N_18941);
and UO_949 (O_949,N_19772,N_20514);
nor UO_950 (O_950,N_19371,N_20821);
nor UO_951 (O_951,N_22760,N_19887);
nor UO_952 (O_952,N_22911,N_24803);
nand UO_953 (O_953,N_23065,N_21395);
xor UO_954 (O_954,N_22271,N_23647);
nor UO_955 (O_955,N_19731,N_22026);
and UO_956 (O_956,N_19349,N_19540);
or UO_957 (O_957,N_23130,N_21782);
or UO_958 (O_958,N_20856,N_24289);
nor UO_959 (O_959,N_19034,N_21088);
and UO_960 (O_960,N_23296,N_24556);
nor UO_961 (O_961,N_22617,N_22456);
nand UO_962 (O_962,N_18778,N_20495);
nand UO_963 (O_963,N_23115,N_21674);
nand UO_964 (O_964,N_24324,N_23046);
nor UO_965 (O_965,N_20054,N_20924);
nand UO_966 (O_966,N_23143,N_24925);
nand UO_967 (O_967,N_20848,N_22491);
nor UO_968 (O_968,N_20907,N_24111);
or UO_969 (O_969,N_22877,N_21564);
nand UO_970 (O_970,N_20777,N_18863);
nand UO_971 (O_971,N_24291,N_21538);
nor UO_972 (O_972,N_22724,N_22695);
xnor UO_973 (O_973,N_21437,N_24791);
nor UO_974 (O_974,N_24842,N_22539);
nand UO_975 (O_975,N_21044,N_19419);
and UO_976 (O_976,N_23836,N_23176);
nor UO_977 (O_977,N_23664,N_20311);
or UO_978 (O_978,N_19074,N_21108);
nand UO_979 (O_979,N_19952,N_19410);
and UO_980 (O_980,N_20390,N_19862);
and UO_981 (O_981,N_21448,N_20734);
nor UO_982 (O_982,N_24378,N_22837);
xnor UO_983 (O_983,N_19144,N_20538);
or UO_984 (O_984,N_22701,N_21942);
and UO_985 (O_985,N_21056,N_22604);
or UO_986 (O_986,N_24624,N_22828);
and UO_987 (O_987,N_22662,N_22937);
or UO_988 (O_988,N_19882,N_21311);
nand UO_989 (O_989,N_19477,N_18829);
xor UO_990 (O_990,N_24107,N_20707);
nor UO_991 (O_991,N_24047,N_19735);
and UO_992 (O_992,N_22043,N_23961);
nand UO_993 (O_993,N_19059,N_23181);
nor UO_994 (O_994,N_19230,N_18919);
nand UO_995 (O_995,N_23997,N_22846);
nor UO_996 (O_996,N_20000,N_20875);
nand UO_997 (O_997,N_20127,N_22437);
and UO_998 (O_998,N_21140,N_22273);
or UO_999 (O_999,N_23278,N_22506);
nand UO_1000 (O_1000,N_20607,N_23710);
or UO_1001 (O_1001,N_24904,N_24877);
nand UO_1002 (O_1002,N_19506,N_23088);
or UO_1003 (O_1003,N_23424,N_22336);
or UO_1004 (O_1004,N_22784,N_19884);
xor UO_1005 (O_1005,N_22878,N_19254);
or UO_1006 (O_1006,N_24486,N_19197);
nand UO_1007 (O_1007,N_19225,N_23529);
nand UO_1008 (O_1008,N_19444,N_20942);
or UO_1009 (O_1009,N_23890,N_21113);
or UO_1010 (O_1010,N_19734,N_19278);
or UO_1011 (O_1011,N_21453,N_19513);
nand UO_1012 (O_1012,N_20825,N_20216);
and UO_1013 (O_1013,N_21694,N_24213);
nor UO_1014 (O_1014,N_22791,N_20103);
and UO_1015 (O_1015,N_24911,N_19656);
nand UO_1016 (O_1016,N_24362,N_18821);
xnor UO_1017 (O_1017,N_19527,N_19063);
and UO_1018 (O_1018,N_21565,N_21459);
or UO_1019 (O_1019,N_21325,N_19970);
and UO_1020 (O_1020,N_19375,N_23904);
nand UO_1021 (O_1021,N_19440,N_23865);
xor UO_1022 (O_1022,N_22351,N_22052);
nor UO_1023 (O_1023,N_24600,N_19311);
nand UO_1024 (O_1024,N_24869,N_24310);
and UO_1025 (O_1025,N_22326,N_22667);
and UO_1026 (O_1026,N_20909,N_22969);
and UO_1027 (O_1027,N_20617,N_21697);
nand UO_1028 (O_1028,N_21422,N_19844);
nor UO_1029 (O_1029,N_21900,N_19898);
xnor UO_1030 (O_1030,N_19580,N_23585);
nand UO_1031 (O_1031,N_22887,N_20182);
and UO_1032 (O_1032,N_23686,N_22745);
or UO_1033 (O_1033,N_21965,N_23193);
nor UO_1034 (O_1034,N_22284,N_23125);
nand UO_1035 (O_1035,N_19261,N_20291);
nor UO_1036 (O_1036,N_23456,N_19550);
nand UO_1037 (O_1037,N_24953,N_19750);
nor UO_1038 (O_1038,N_24633,N_21809);
and UO_1039 (O_1039,N_24710,N_18752);
xor UO_1040 (O_1040,N_23869,N_24348);
nor UO_1041 (O_1041,N_20212,N_22133);
or UO_1042 (O_1042,N_19633,N_22331);
and UO_1043 (O_1043,N_24891,N_21275);
nand UO_1044 (O_1044,N_24137,N_20779);
and UO_1045 (O_1045,N_18904,N_20417);
or UO_1046 (O_1046,N_21327,N_20983);
xnor UO_1047 (O_1047,N_23943,N_20836);
nor UO_1048 (O_1048,N_23400,N_19365);
or UO_1049 (O_1049,N_20797,N_22317);
nand UO_1050 (O_1050,N_24123,N_19117);
nand UO_1051 (O_1051,N_23363,N_24844);
nand UO_1052 (O_1052,N_20774,N_22399);
and UO_1053 (O_1053,N_21420,N_21375);
or UO_1054 (O_1054,N_23545,N_23421);
nand UO_1055 (O_1055,N_20710,N_23182);
or UO_1056 (O_1056,N_19268,N_20240);
and UO_1057 (O_1057,N_24479,N_24672);
nand UO_1058 (O_1058,N_24518,N_22256);
and UO_1059 (O_1059,N_23397,N_22766);
xnor UO_1060 (O_1060,N_23178,N_20917);
and UO_1061 (O_1061,N_22258,N_22072);
or UO_1062 (O_1062,N_18911,N_24236);
or UO_1063 (O_1063,N_22395,N_20726);
nor UO_1064 (O_1064,N_19155,N_19383);
nand UO_1065 (O_1065,N_24202,N_21193);
nand UO_1066 (O_1066,N_24425,N_22303);
or UO_1067 (O_1067,N_19699,N_18808);
or UO_1068 (O_1068,N_23543,N_21749);
nor UO_1069 (O_1069,N_20492,N_21057);
nor UO_1070 (O_1070,N_22278,N_21733);
or UO_1071 (O_1071,N_20162,N_21042);
or UO_1072 (O_1072,N_19455,N_23042);
nand UO_1073 (O_1073,N_20973,N_24173);
nor UO_1074 (O_1074,N_21349,N_21813);
nand UO_1075 (O_1075,N_20157,N_21766);
nand UO_1076 (O_1076,N_24555,N_23413);
or UO_1077 (O_1077,N_20326,N_23396);
nor UO_1078 (O_1078,N_18794,N_19058);
nor UO_1079 (O_1079,N_22821,N_24349);
or UO_1080 (O_1080,N_21555,N_23964);
nor UO_1081 (O_1081,N_24609,N_20968);
nor UO_1082 (O_1082,N_24225,N_24456);
nand UO_1083 (O_1083,N_22247,N_23359);
nand UO_1084 (O_1084,N_19742,N_22457);
nor UO_1085 (O_1085,N_21921,N_23258);
nand UO_1086 (O_1086,N_21639,N_20286);
nor UO_1087 (O_1087,N_24902,N_22460);
and UO_1088 (O_1088,N_20122,N_19201);
and UO_1089 (O_1089,N_22316,N_20754);
or UO_1090 (O_1090,N_23599,N_19749);
or UO_1091 (O_1091,N_20770,N_18917);
nor UO_1092 (O_1092,N_22812,N_20262);
nand UO_1093 (O_1093,N_20456,N_24519);
xor UO_1094 (O_1094,N_23668,N_19163);
and UO_1095 (O_1095,N_22523,N_20214);
nor UO_1096 (O_1096,N_19959,N_23286);
nor UO_1097 (O_1097,N_24611,N_22600);
xor UO_1098 (O_1098,N_19595,N_18807);
xor UO_1099 (O_1099,N_24705,N_18764);
nand UO_1100 (O_1100,N_18947,N_22150);
nor UO_1101 (O_1101,N_20247,N_21300);
nor UO_1102 (O_1102,N_23931,N_22720);
nand UO_1103 (O_1103,N_21513,N_19153);
nand UO_1104 (O_1104,N_19586,N_24115);
or UO_1105 (O_1105,N_23992,N_19020);
nor UO_1106 (O_1106,N_22455,N_23019);
nor UO_1107 (O_1107,N_21750,N_24138);
and UO_1108 (O_1108,N_19164,N_19736);
or UO_1109 (O_1109,N_24153,N_23868);
or UO_1110 (O_1110,N_19710,N_23895);
nor UO_1111 (O_1111,N_24011,N_20794);
nor UO_1112 (O_1112,N_23848,N_21917);
and UO_1113 (O_1113,N_22999,N_22630);
nand UO_1114 (O_1114,N_23846,N_22220);
nand UO_1115 (O_1115,N_23361,N_19673);
nor UO_1116 (O_1116,N_21069,N_24851);
and UO_1117 (O_1117,N_24421,N_24916);
or UO_1118 (O_1118,N_23940,N_22572);
and UO_1119 (O_1119,N_23327,N_19050);
and UO_1120 (O_1120,N_19161,N_22556);
or UO_1121 (O_1121,N_19899,N_22042);
nand UO_1122 (O_1122,N_19002,N_19559);
and UO_1123 (O_1123,N_22104,N_22613);
nand UO_1124 (O_1124,N_24140,N_23902);
nand UO_1125 (O_1125,N_23678,N_19630);
and UO_1126 (O_1126,N_22172,N_23373);
xor UO_1127 (O_1127,N_23192,N_24759);
nor UO_1128 (O_1128,N_20132,N_23167);
and UO_1129 (O_1129,N_22655,N_19233);
and UO_1130 (O_1130,N_24595,N_24514);
and UO_1131 (O_1131,N_21270,N_20688);
xor UO_1132 (O_1132,N_24071,N_22645);
or UO_1133 (O_1133,N_23457,N_20263);
and UO_1134 (O_1134,N_19701,N_24776);
nor UO_1135 (O_1135,N_23888,N_23828);
and UO_1136 (O_1136,N_21506,N_19245);
nor UO_1137 (O_1137,N_19624,N_21306);
nor UO_1138 (O_1138,N_23152,N_21794);
or UO_1139 (O_1139,N_24471,N_24494);
and UO_1140 (O_1140,N_21162,N_18801);
nand UO_1141 (O_1141,N_18961,N_21021);
and UO_1142 (O_1142,N_24876,N_24177);
and UO_1143 (O_1143,N_22212,N_22264);
nand UO_1144 (O_1144,N_22036,N_24234);
and UO_1145 (O_1145,N_21209,N_19831);
and UO_1146 (O_1146,N_21637,N_23745);
nand UO_1147 (O_1147,N_24539,N_20528);
nand UO_1148 (O_1148,N_20861,N_18999);
and UO_1149 (O_1149,N_22996,N_24835);
nand UO_1150 (O_1150,N_19055,N_23508);
or UO_1151 (O_1151,N_23430,N_19303);
nand UO_1152 (O_1152,N_23960,N_22785);
nor UO_1153 (O_1153,N_20248,N_24242);
nor UO_1154 (O_1154,N_22825,N_24325);
nor UO_1155 (O_1155,N_22567,N_20904);
nor UO_1156 (O_1156,N_21136,N_19428);
and UO_1157 (O_1157,N_19572,N_19826);
nand UO_1158 (O_1158,N_24398,N_18832);
or UO_1159 (O_1159,N_23014,N_20589);
or UO_1160 (O_1160,N_22531,N_24634);
nor UO_1161 (O_1161,N_20839,N_19715);
nand UO_1162 (O_1162,N_22941,N_22952);
nor UO_1163 (O_1163,N_18922,N_18775);
xnor UO_1164 (O_1164,N_23132,N_20505);
and UO_1165 (O_1165,N_21833,N_21759);
nand UO_1166 (O_1166,N_24706,N_20428);
or UO_1167 (O_1167,N_22458,N_22186);
or UO_1168 (O_1168,N_22209,N_19300);
nor UO_1169 (O_1169,N_21659,N_23674);
or UO_1170 (O_1170,N_23765,N_19009);
nand UO_1171 (O_1171,N_22353,N_19190);
nor UO_1172 (O_1172,N_20051,N_23986);
xor UO_1173 (O_1173,N_21839,N_22157);
or UO_1174 (O_1174,N_22228,N_19602);
nand UO_1175 (O_1175,N_19023,N_19537);
or UO_1176 (O_1176,N_23587,N_23681);
nor UO_1177 (O_1177,N_22607,N_21728);
or UO_1178 (O_1178,N_19160,N_20835);
nor UO_1179 (O_1179,N_22269,N_24355);
nand UO_1180 (O_1180,N_23499,N_22081);
or UO_1181 (O_1181,N_21417,N_20070);
and UO_1182 (O_1182,N_22364,N_20693);
and UO_1183 (O_1183,N_20897,N_19343);
and UO_1184 (O_1184,N_21933,N_22098);
or UO_1185 (O_1185,N_24651,N_19620);
or UO_1186 (O_1186,N_24766,N_22997);
nand UO_1187 (O_1187,N_23864,N_19296);
xor UO_1188 (O_1188,N_24293,N_19503);
nor UO_1189 (O_1189,N_24945,N_22945);
or UO_1190 (O_1190,N_23336,N_19294);
and UO_1191 (O_1191,N_24383,N_22553);
and UO_1192 (O_1192,N_19798,N_23171);
and UO_1193 (O_1193,N_21899,N_21034);
xnor UO_1194 (O_1194,N_24178,N_21421);
or UO_1195 (O_1195,N_21505,N_18898);
or UO_1196 (O_1196,N_20191,N_22016);
nor UO_1197 (O_1197,N_23724,N_22236);
and UO_1198 (O_1198,N_20126,N_23993);
nand UO_1199 (O_1199,N_23863,N_19569);
and UO_1200 (O_1200,N_24992,N_21462);
and UO_1201 (O_1201,N_20480,N_24797);
nand UO_1202 (O_1202,N_24447,N_21085);
or UO_1203 (O_1203,N_19047,N_24332);
or UO_1204 (O_1204,N_20033,N_19459);
nor UO_1205 (O_1205,N_24150,N_22121);
and UO_1206 (O_1206,N_22200,N_22113);
nand UO_1207 (O_1207,N_23434,N_21408);
and UO_1208 (O_1208,N_20373,N_24340);
or UO_1209 (O_1209,N_19490,N_22644);
nand UO_1210 (O_1210,N_22866,N_21075);
or UO_1211 (O_1211,N_20031,N_20123);
xor UO_1212 (O_1212,N_23831,N_20442);
nand UO_1213 (O_1213,N_22569,N_24312);
nand UO_1214 (O_1214,N_20449,N_19993);
nand UO_1215 (O_1215,N_21218,N_20650);
xnor UO_1216 (O_1216,N_24831,N_22242);
and UO_1217 (O_1217,N_20235,N_22485);
nor UO_1218 (O_1218,N_22055,N_19360);
and UO_1219 (O_1219,N_21805,N_22540);
nand UO_1220 (O_1220,N_19470,N_24782);
or UO_1221 (O_1221,N_20440,N_19709);
or UO_1222 (O_1222,N_22123,N_22165);
and UO_1223 (O_1223,N_24736,N_20857);
nand UO_1224 (O_1224,N_24151,N_24654);
nand UO_1225 (O_1225,N_24573,N_23273);
or UO_1226 (O_1226,N_24991,N_23900);
and UO_1227 (O_1227,N_21645,N_24731);
nor UO_1228 (O_1228,N_22327,N_19138);
nor UO_1229 (O_1229,N_20837,N_23564);
and UO_1230 (O_1230,N_20432,N_24666);
and UO_1231 (O_1231,N_20325,N_22103);
nor UO_1232 (O_1232,N_23547,N_23060);
nor UO_1233 (O_1233,N_24641,N_24799);
nand UO_1234 (O_1234,N_21793,N_21491);
and UO_1235 (O_1235,N_19199,N_20357);
and UO_1236 (O_1236,N_21138,N_21435);
or UO_1237 (O_1237,N_21111,N_19077);
and UO_1238 (O_1238,N_20652,N_24073);
nand UO_1239 (O_1239,N_20673,N_19703);
nor UO_1240 (O_1240,N_24856,N_23473);
nor UO_1241 (O_1241,N_20772,N_23350);
or UO_1242 (O_1242,N_21399,N_22224);
xor UO_1243 (O_1243,N_18804,N_19647);
or UO_1244 (O_1244,N_22137,N_22654);
or UO_1245 (O_1245,N_18820,N_24215);
nor UO_1246 (O_1246,N_23862,N_22749);
or UO_1247 (O_1247,N_24170,N_23020);
nor UO_1248 (O_1248,N_22899,N_21523);
nand UO_1249 (O_1249,N_21239,N_20611);
or UO_1250 (O_1250,N_19053,N_20769);
nor UO_1251 (O_1251,N_24051,N_24176);
xor UO_1252 (O_1252,N_22827,N_21732);
nor UO_1253 (O_1253,N_19185,N_22557);
nand UO_1254 (O_1254,N_22387,N_19967);
or UO_1255 (O_1255,N_19095,N_22830);
or UO_1256 (O_1256,N_22973,N_19179);
nor UO_1257 (O_1257,N_18962,N_24967);
or UO_1258 (O_1258,N_21123,N_19202);
nand UO_1259 (O_1259,N_22432,N_21924);
nor UO_1260 (O_1260,N_22333,N_24006);
and UO_1261 (O_1261,N_24545,N_21704);
or UO_1262 (O_1262,N_21690,N_21825);
nor UO_1263 (O_1263,N_22768,N_24826);
xor UO_1264 (O_1264,N_22168,N_24394);
and UO_1265 (O_1265,N_22249,N_21688);
or UO_1266 (O_1266,N_24621,N_21740);
and UO_1267 (O_1267,N_20171,N_23330);
nor UO_1268 (O_1268,N_23517,N_20496);
nand UO_1269 (O_1269,N_19467,N_18783);
or UO_1270 (O_1270,N_23064,N_23584);
nor UO_1271 (O_1271,N_21362,N_20658);
nor UO_1272 (O_1272,N_24985,N_23733);
and UO_1273 (O_1273,N_21386,N_20966);
nand UO_1274 (O_1274,N_23386,N_20065);
or UO_1275 (O_1275,N_19517,N_20230);
nor UO_1276 (O_1276,N_22725,N_23755);
nand UO_1277 (O_1277,N_20124,N_21377);
nor UO_1278 (O_1278,N_22029,N_24847);
or UO_1279 (O_1279,N_21568,N_24343);
nand UO_1280 (O_1280,N_18926,N_20186);
and UO_1281 (O_1281,N_24294,N_23580);
nand UO_1282 (O_1282,N_23980,N_23390);
nor UO_1283 (O_1283,N_20315,N_24561);
nand UO_1284 (O_1284,N_24427,N_22727);
or UO_1285 (O_1285,N_24434,N_21430);
nand UO_1286 (O_1286,N_22509,N_23270);
and UO_1287 (O_1287,N_20522,N_21456);
or UO_1288 (O_1288,N_19533,N_22120);
and UO_1289 (O_1289,N_18965,N_20078);
or UO_1290 (O_1290,N_24499,N_21168);
or UO_1291 (O_1291,N_22507,N_21178);
nor UO_1292 (O_1292,N_23977,N_23066);
and UO_1293 (O_1293,N_19657,N_21488);
and UO_1294 (O_1294,N_19683,N_21549);
or UO_1295 (O_1295,N_18812,N_21428);
and UO_1296 (O_1296,N_19228,N_19106);
and UO_1297 (O_1297,N_22187,N_23516);
nor UO_1298 (O_1298,N_23643,N_20723);
xnor UO_1299 (O_1299,N_21040,N_19359);
and UO_1300 (O_1300,N_23257,N_19933);
and UO_1301 (O_1301,N_22881,N_20932);
and UO_1302 (O_1302,N_23560,N_21157);
xnor UO_1303 (O_1303,N_23932,N_20180);
nand UO_1304 (O_1304,N_23311,N_20684);
or UO_1305 (O_1305,N_20791,N_20512);
nor UO_1306 (O_1306,N_19942,N_19181);
nand UO_1307 (O_1307,N_22966,N_21007);
nor UO_1308 (O_1308,N_24807,N_22517);
and UO_1309 (O_1309,N_20096,N_23898);
nand UO_1310 (O_1310,N_21980,N_23114);
xor UO_1311 (O_1311,N_19780,N_19704);
nor UO_1312 (O_1312,N_21651,N_19649);
and UO_1313 (O_1313,N_22077,N_22859);
nand UO_1314 (O_1314,N_21388,N_19482);
or UO_1315 (O_1315,N_24405,N_21068);
or UO_1316 (O_1316,N_23471,N_22033);
or UO_1317 (O_1317,N_24515,N_23947);
or UO_1318 (O_1318,N_22993,N_23469);
and UO_1319 (O_1319,N_19304,N_20655);
nand UO_1320 (O_1320,N_23185,N_19393);
or UO_1321 (O_1321,N_24280,N_22668);
or UO_1322 (O_1322,N_21653,N_24788);
nand UO_1323 (O_1323,N_20172,N_22503);
nand UO_1324 (O_1324,N_20766,N_21414);
nor UO_1325 (O_1325,N_19914,N_21765);
and UO_1326 (O_1326,N_24889,N_24972);
or UO_1327 (O_1327,N_19054,N_20893);
nand UO_1328 (O_1328,N_24698,N_24906);
or UO_1329 (O_1329,N_22869,N_24773);
nand UO_1330 (O_1330,N_22268,N_24098);
nor UO_1331 (O_1331,N_23666,N_23294);
nand UO_1332 (O_1332,N_21559,N_24720);
nand UO_1333 (O_1333,N_21982,N_19906);
or UO_1334 (O_1334,N_23281,N_20930);
nor UO_1335 (O_1335,N_24076,N_23609);
nand UO_1336 (O_1336,N_21748,N_18803);
and UO_1337 (O_1337,N_23342,N_21261);
and UO_1338 (O_1338,N_24912,N_19865);
nor UO_1339 (O_1339,N_18989,N_20433);
or UO_1340 (O_1340,N_18825,N_21187);
nor UO_1341 (O_1341,N_23393,N_19529);
nand UO_1342 (O_1342,N_19087,N_23438);
and UO_1343 (O_1343,N_19022,N_20453);
nand UO_1344 (O_1344,N_19788,N_24190);
nor UO_1345 (O_1345,N_23701,N_22648);
nor UO_1346 (O_1346,N_20211,N_19815);
or UO_1347 (O_1347,N_22936,N_24495);
xor UO_1348 (O_1348,N_21182,N_21718);
and UO_1349 (O_1349,N_23604,N_19272);
nor UO_1350 (O_1350,N_18800,N_19382);
nor UO_1351 (O_1351,N_23510,N_24690);
and UO_1352 (O_1352,N_19374,N_24467);
or UO_1353 (O_1353,N_23179,N_23437);
nor UO_1354 (O_1354,N_21224,N_21098);
or UO_1355 (O_1355,N_23168,N_21365);
nand UO_1356 (O_1356,N_20016,N_22127);
xor UO_1357 (O_1357,N_20170,N_21715);
nand UO_1358 (O_1358,N_22452,N_22661);
or UO_1359 (O_1359,N_23425,N_24870);
nand UO_1360 (O_1360,N_19405,N_23722);
xor UO_1361 (O_1361,N_19082,N_21489);
or UO_1362 (O_1362,N_20225,N_21843);
nand UO_1363 (O_1363,N_24715,N_24750);
and UO_1364 (O_1364,N_20166,N_21267);
xor UO_1365 (O_1365,N_23459,N_22948);
nand UO_1366 (O_1366,N_23813,N_23673);
or UO_1367 (O_1367,N_19324,N_23858);
or UO_1368 (O_1368,N_19978,N_20912);
nand UO_1369 (O_1369,N_21141,N_21012);
or UO_1370 (O_1370,N_23230,N_19104);
or UO_1371 (O_1371,N_20509,N_22204);
nand UO_1372 (O_1372,N_20345,N_21352);
and UO_1373 (O_1373,N_21425,N_20551);
nand UO_1374 (O_1374,N_20581,N_21051);
nand UO_1375 (O_1375,N_24643,N_23189);
nand UO_1376 (O_1376,N_20437,N_24161);
or UO_1377 (O_1377,N_21779,N_22166);
nand UO_1378 (O_1378,N_24220,N_19357);
xnor UO_1379 (O_1379,N_24254,N_23922);
nand UO_1380 (O_1380,N_22015,N_21133);
and UO_1381 (O_1381,N_23054,N_21812);
and UO_1382 (O_1382,N_18899,N_24431);
nor UO_1383 (O_1383,N_20992,N_19747);
nand UO_1384 (O_1384,N_24905,N_21983);
and UO_1385 (O_1385,N_24549,N_20699);
nand UO_1386 (O_1386,N_23244,N_23769);
and UO_1387 (O_1387,N_19348,N_23959);
or UO_1388 (O_1388,N_22616,N_23427);
or UO_1389 (O_1389,N_22637,N_19737);
or UO_1390 (O_1390,N_19634,N_24387);
nand UO_1391 (O_1391,N_22142,N_21197);
or UO_1392 (O_1392,N_19449,N_21614);
nor UO_1393 (O_1393,N_22101,N_19700);
nor UO_1394 (O_1394,N_22639,N_21648);
and UO_1395 (O_1395,N_22642,N_22376);
and UO_1396 (O_1396,N_23180,N_20525);
nor UO_1397 (O_1397,N_19538,N_22446);
or UO_1398 (O_1398,N_24316,N_22756);
nand UO_1399 (O_1399,N_20244,N_19131);
and UO_1400 (O_1400,N_23919,N_24895);
and UO_1401 (O_1401,N_19662,N_20474);
nor UO_1402 (O_1402,N_20822,N_21677);
or UO_1403 (O_1403,N_22447,N_19751);
and UO_1404 (O_1404,N_24729,N_22208);
nand UO_1405 (O_1405,N_22965,N_21476);
and UO_1406 (O_1406,N_23145,N_20533);
nand UO_1407 (O_1407,N_24119,N_23013);
xor UO_1408 (O_1408,N_23500,N_24652);
or UO_1409 (O_1409,N_24149,N_23491);
or UO_1410 (O_1410,N_21132,N_22093);
nor UO_1411 (O_1411,N_22470,N_20490);
nand UO_1412 (O_1412,N_23021,N_21830);
nor UO_1413 (O_1413,N_20816,N_22703);
nor UO_1414 (O_1414,N_21981,N_23824);
xor UO_1415 (O_1415,N_18998,N_19992);
nand UO_1416 (O_1416,N_22066,N_21380);
nor UO_1417 (O_1417,N_21922,N_24890);
or UO_1418 (O_1418,N_18767,N_19422);
xor UO_1419 (O_1419,N_20458,N_24428);
nor UO_1420 (O_1420,N_24635,N_22998);
or UO_1421 (O_1421,N_20604,N_19575);
nand UO_1422 (O_1422,N_23329,N_23137);
nor UO_1423 (O_1423,N_23663,N_23138);
nand UO_1424 (O_1424,N_19123,N_23234);
and UO_1425 (O_1425,N_22233,N_21419);
and UO_1426 (O_1426,N_23723,N_21235);
or UO_1427 (O_1427,N_24965,N_22357);
nand UO_1428 (O_1428,N_23116,N_18916);
nor UO_1429 (O_1429,N_22804,N_22906);
nor UO_1430 (O_1430,N_20183,N_24754);
nand UO_1431 (O_1431,N_18791,N_22329);
and UO_1432 (O_1432,N_20843,N_20755);
nor UO_1433 (O_1433,N_19787,N_19684);
nand UO_1434 (O_1434,N_21532,N_23461);
xnor UO_1435 (O_1435,N_24966,N_21859);
and UO_1436 (O_1436,N_22171,N_23497);
nand UO_1437 (O_1437,N_20716,N_19027);
xnor UO_1438 (O_1438,N_19505,N_22907);
nand UO_1439 (O_1439,N_21944,N_20392);
xor UO_1440 (O_1440,N_24781,N_22341);
and UO_1441 (O_1441,N_19010,N_21885);
or UO_1442 (O_1442,N_22848,N_23283);
or UO_1443 (O_1443,N_20027,N_20796);
nor UO_1444 (O_1444,N_22148,N_19813);
and UO_1445 (O_1445,N_21192,N_21234);
nand UO_1446 (O_1446,N_20648,N_19145);
nor UO_1447 (O_1447,N_19597,N_24938);
nor UO_1448 (O_1448,N_22243,N_21742);
and UO_1449 (O_1449,N_20781,N_24888);
or UO_1450 (O_1450,N_23572,N_22704);
nor UO_1451 (O_1451,N_18880,N_24783);
xnor UO_1452 (O_1452,N_23206,N_20993);
xnor UO_1453 (O_1453,N_23324,N_22218);
or UO_1454 (O_1454,N_24612,N_19514);
nand UO_1455 (O_1455,N_20450,N_23642);
or UO_1456 (O_1456,N_24210,N_21101);
or UO_1457 (O_1457,N_19972,N_22659);
and UO_1458 (O_1458,N_24200,N_19073);
nor UO_1459 (O_1459,N_19607,N_20736);
nand UO_1460 (O_1460,N_21548,N_23208);
nor UO_1461 (O_1461,N_24245,N_23789);
or UO_1462 (O_1462,N_22538,N_20534);
and UO_1463 (O_1463,N_23039,N_21895);
and UO_1464 (O_1464,N_21036,N_22561);
xnor UO_1465 (O_1465,N_20711,N_18851);
and UO_1466 (O_1466,N_21360,N_20542);
xor UO_1467 (O_1467,N_20337,N_22199);
and UO_1468 (O_1468,N_22117,N_22379);
and UO_1469 (O_1469,N_24679,N_20178);
nor UO_1470 (O_1470,N_23200,N_24099);
and UO_1471 (O_1471,N_23983,N_19864);
nand UO_1472 (O_1472,N_21486,N_24900);
nor UO_1473 (O_1473,N_23405,N_24565);
xor UO_1474 (O_1474,N_21058,N_24642);
nor UO_1475 (O_1475,N_19920,N_23038);
and UO_1476 (O_1476,N_21726,N_23687);
nor UO_1477 (O_1477,N_19240,N_20748);
and UO_1478 (O_1478,N_23962,N_19193);
nor UO_1479 (O_1479,N_18993,N_19685);
nand UO_1480 (O_1480,N_19146,N_21511);
and UO_1481 (O_1481,N_23558,N_18866);
nor UO_1482 (O_1482,N_23245,N_21167);
and UO_1483 (O_1483,N_21990,N_19694);
and UO_1484 (O_1484,N_19969,N_22856);
or UO_1485 (O_1485,N_19953,N_23669);
nand UO_1486 (O_1486,N_22813,N_20624);
and UO_1487 (O_1487,N_19995,N_22096);
or UO_1488 (O_1488,N_19839,N_24290);
nor UO_1489 (O_1489,N_24373,N_20811);
and UO_1490 (O_1490,N_20778,N_20443);
and UO_1491 (O_1491,N_21537,N_21857);
or UO_1492 (O_1492,N_20144,N_20215);
or UO_1493 (O_1493,N_20274,N_22392);
xnor UO_1494 (O_1494,N_24112,N_20028);
and UO_1495 (O_1495,N_21957,N_22880);
nor UO_1496 (O_1496,N_24224,N_24949);
or UO_1497 (O_1497,N_19828,N_22953);
and UO_1498 (O_1498,N_23203,N_23136);
nand UO_1499 (O_1499,N_19172,N_19124);
nor UO_1500 (O_1500,N_23371,N_20902);
or UO_1501 (O_1501,N_19820,N_24973);
nand UO_1502 (O_1502,N_18867,N_24694);
and UO_1503 (O_1503,N_20220,N_22282);
xor UO_1504 (O_1504,N_20768,N_21457);
or UO_1505 (O_1505,N_19045,N_22145);
or UO_1506 (O_1506,N_19251,N_24741);
and UO_1507 (O_1507,N_23844,N_22252);
nor UO_1508 (O_1508,N_23027,N_21785);
nand UO_1509 (O_1509,N_23022,N_22771);
and UO_1510 (O_1510,N_21053,N_19336);
and UO_1511 (O_1511,N_24583,N_24901);
nor UO_1512 (O_1512,N_23310,N_23999);
nor UO_1513 (O_1513,N_18785,N_21251);
nor UO_1514 (O_1514,N_24538,N_24662);
nand UO_1515 (O_1515,N_20444,N_21010);
nor UO_1516 (O_1516,N_24743,N_23763);
and UO_1517 (O_1517,N_20858,N_21657);
and UO_1518 (O_1518,N_21227,N_23908);
nand UO_1519 (O_1519,N_21171,N_20279);
and UO_1520 (O_1520,N_23768,N_22177);
nor UO_1521 (O_1521,N_21737,N_19126);
nor UO_1522 (O_1522,N_24201,N_19353);
nand UO_1523 (O_1523,N_18765,N_23308);
and UO_1524 (O_1524,N_19386,N_21923);
and UO_1525 (O_1525,N_21553,N_21816);
nor UO_1526 (O_1526,N_22750,N_23884);
and UO_1527 (O_1527,N_23475,N_22591);
nand UO_1528 (O_1528,N_24579,N_20747);
or UO_1529 (O_1529,N_22543,N_22330);
nand UO_1530 (O_1530,N_20976,N_19392);
xnor UO_1531 (O_1531,N_20913,N_20058);
xnor UO_1532 (O_1532,N_23402,N_21099);
or UO_1533 (O_1533,N_24453,N_21191);
and UO_1534 (O_1534,N_19841,N_20477);
or UO_1535 (O_1535,N_21367,N_22549);
xor UO_1536 (O_1536,N_23693,N_21103);
nor UO_1537 (O_1537,N_21512,N_23968);
xor UO_1538 (O_1538,N_24483,N_23648);
and UO_1539 (O_1539,N_23544,N_19501);
or UO_1540 (O_1540,N_19218,N_22658);
or UO_1541 (O_1541,N_22739,N_22926);
nor UO_1542 (O_1542,N_19576,N_19672);
xnor UO_1543 (O_1543,N_20210,N_22170);
or UO_1544 (O_1544,N_20952,N_21569);
nand UO_1545 (O_1545,N_18792,N_22466);
nor UO_1546 (O_1546,N_19808,N_23053);
or UO_1547 (O_1547,N_20429,N_19758);
xor UO_1548 (O_1548,N_24541,N_19036);
nor UO_1549 (O_1549,N_22510,N_23988);
or UO_1550 (O_1550,N_24894,N_19675);
xnor UO_1551 (O_1551,N_23924,N_19911);
xor UO_1552 (O_1552,N_22021,N_21211);
nor UO_1553 (O_1553,N_19545,N_22354);
and UO_1554 (O_1554,N_19725,N_22240);
nand UO_1555 (O_1555,N_24113,N_18781);
or UO_1556 (O_1556,N_20945,N_23870);
or UO_1557 (O_1557,N_23852,N_22384);
xor UO_1558 (O_1558,N_19326,N_24623);
and UO_1559 (O_1559,N_20233,N_21583);
and UO_1560 (O_1560,N_22820,N_19797);
nand UO_1561 (O_1561,N_21248,N_22342);
nor UO_1562 (O_1562,N_22227,N_19051);
and UO_1563 (O_1563,N_22855,N_19902);
nand UO_1564 (O_1564,N_19156,N_21589);
and UO_1565 (O_1565,N_24438,N_22006);
nand UO_1566 (O_1566,N_22664,N_20074);
xor UO_1567 (O_1567,N_21232,N_20093);
or UO_1568 (O_1568,N_23552,N_19395);
or UO_1569 (O_1569,N_24603,N_23787);
nor UO_1570 (O_1570,N_20098,N_20021);
xnor UO_1571 (O_1571,N_20382,N_21289);
nand UO_1572 (O_1572,N_22106,N_19492);
or UO_1573 (O_1573,N_19900,N_24023);
nand UO_1574 (O_1574,N_24718,N_19102);
nand UO_1575 (O_1575,N_19549,N_21636);
xnor UO_1576 (O_1576,N_22584,N_20960);
or UO_1577 (O_1577,N_21358,N_21840);
nor UO_1578 (O_1578,N_23987,N_23633);
nand UO_1579 (O_1579,N_21066,N_22309);
nand UO_1580 (O_1580,N_22693,N_22657);
and UO_1581 (O_1581,N_24211,N_20951);
or UO_1582 (O_1582,N_20616,N_22861);
nand UO_1583 (O_1583,N_23559,N_20252);
nand UO_1584 (O_1584,N_22700,N_19269);
nor UO_1585 (O_1585,N_24252,N_21752);
or UO_1586 (O_1586,N_21970,N_19986);
and UO_1587 (O_1587,N_19612,N_24108);
and UO_1588 (O_1588,N_18934,N_19556);
nand UO_1589 (O_1589,N_21356,N_20486);
or UO_1590 (O_1590,N_23812,N_21253);
or UO_1591 (O_1591,N_22361,N_23853);
nand UO_1592 (O_1592,N_19184,N_20971);
or UO_1593 (O_1593,N_22067,N_20112);
nor UO_1594 (O_1594,N_22961,N_22134);
and UO_1595 (O_1595,N_23157,N_22070);
xor UO_1596 (O_1596,N_19744,N_20970);
or UO_1597 (O_1597,N_24168,N_23546);
xnor UO_1598 (O_1598,N_18900,N_20156);
xor UO_1599 (O_1599,N_20290,N_21418);
nand UO_1600 (O_1600,N_19981,N_18992);
nand UO_1601 (O_1601,N_18761,N_23638);
or UO_1602 (O_1602,N_20883,N_22838);
xor UO_1603 (O_1603,N_21174,N_21370);
and UO_1604 (O_1604,N_23866,N_21656);
or UO_1605 (O_1605,N_23819,N_18861);
or UO_1606 (O_1606,N_19453,N_19622);
nor UO_1607 (O_1607,N_21032,N_21432);
and UO_1608 (O_1608,N_22231,N_20482);
and UO_1609 (O_1609,N_21337,N_24758);
or UO_1610 (O_1610,N_20729,N_20177);
and UO_1611 (O_1611,N_23202,N_23055);
and UO_1612 (O_1612,N_21655,N_19216);
xor UO_1613 (O_1613,N_21472,N_19406);
and UO_1614 (O_1614,N_18849,N_22338);
and UO_1615 (O_1615,N_21819,N_22565);
and UO_1616 (O_1616,N_24187,N_24517);
or UO_1617 (O_1617,N_22815,N_20511);
xnor UO_1618 (O_1618,N_21507,N_24233);
and UO_1619 (O_1619,N_24692,N_23857);
nand UO_1620 (O_1620,N_20730,N_21081);
nor UO_1621 (O_1621,N_23967,N_22903);
or UO_1622 (O_1622,N_20001,N_23370);
or UO_1623 (O_1623,N_19785,N_24574);
nor UO_1624 (O_1624,N_24409,N_23800);
nand UO_1625 (O_1625,N_20803,N_20323);
nand UO_1626 (O_1626,N_24770,N_23446);
nand UO_1627 (O_1627,N_19237,N_24159);
nor UO_1628 (O_1628,N_20343,N_23700);
nand UO_1629 (O_1629,N_24410,N_23162);
nor UO_1630 (O_1630,N_24932,N_20293);
or UO_1631 (O_1631,N_24648,N_19930);
xor UO_1632 (O_1632,N_19478,N_19610);
and UO_1633 (O_1633,N_24296,N_23240);
xor UO_1634 (O_1634,N_19515,N_19200);
nor UO_1635 (O_1635,N_21219,N_19881);
nand UO_1636 (O_1636,N_24408,N_24323);
nor UO_1637 (O_1637,N_21223,N_21909);
or UO_1638 (O_1638,N_24018,N_24923);
nor UO_1639 (O_1639,N_22283,N_20887);
and UO_1640 (O_1640,N_21406,N_22738);
nor UO_1641 (O_1641,N_20055,N_20780);
nor UO_1642 (O_1642,N_22262,N_20879);
xor UO_1643 (O_1643,N_20076,N_20605);
nor UO_1644 (O_1644,N_20827,N_20702);
or UO_1645 (O_1645,N_19132,N_18951);
nand UO_1646 (O_1646,N_23937,N_19120);
xnor UO_1647 (O_1647,N_19111,N_21460);
nand UO_1648 (O_1648,N_21906,N_21930);
or UO_1649 (O_1649,N_23161,N_22901);
or UO_1650 (O_1650,N_21410,N_19582);
and UO_1651 (O_1651,N_21643,N_24986);
or UO_1652 (O_1652,N_22588,N_20911);
and UO_1653 (O_1653,N_20965,N_19760);
nand UO_1654 (O_1654,N_24327,N_21943);
or UO_1655 (O_1655,N_19162,N_23195);
or UO_1656 (O_1656,N_22944,N_23028);
or UO_1657 (O_1657,N_24533,N_24979);
or UO_1658 (O_1658,N_24368,N_23514);
and UO_1659 (O_1659,N_23339,N_24003);
nor UO_1660 (O_1660,N_24148,N_18810);
nor UO_1661 (O_1661,N_22481,N_23343);
nor UO_1662 (O_1662,N_22777,N_20173);
and UO_1663 (O_1663,N_20964,N_23975);
xor UO_1664 (O_1664,N_24667,N_19905);
nor UO_1665 (O_1665,N_23984,N_23392);
nand UO_1666 (O_1666,N_23043,N_22007);
and UO_1667 (O_1667,N_22201,N_21775);
nor UO_1668 (O_1668,N_19713,N_19812);
or UO_1669 (O_1669,N_24874,N_18855);
nand UO_1670 (O_1670,N_21013,N_18774);
nand UO_1671 (O_1671,N_21979,N_24090);
or UO_1672 (O_1672,N_24616,N_23134);
or UO_1673 (O_1673,N_20273,N_20661);
nand UO_1674 (O_1674,N_24749,N_21165);
and UO_1675 (O_1675,N_22461,N_24043);
and UO_1676 (O_1676,N_19767,N_20187);
nand UO_1677 (O_1677,N_21247,N_24682);
nand UO_1678 (O_1678,N_19456,N_21615);
and UO_1679 (O_1679,N_20621,N_19822);
nor UO_1680 (O_1680,N_21117,N_22762);
nor UO_1681 (O_1681,N_21881,N_20691);
nand UO_1682 (O_1682,N_23169,N_23005);
or UO_1683 (O_1683,N_21172,N_24412);
and UO_1684 (O_1684,N_24309,N_23879);
nand UO_1685 (O_1685,N_24987,N_24839);
and UO_1686 (O_1686,N_19654,N_18958);
or UO_1687 (O_1687,N_20685,N_21701);
or UO_1688 (O_1688,N_23791,N_19093);
nand UO_1689 (O_1689,N_23429,N_20243);
xor UO_1690 (O_1690,N_22612,N_23448);
nor UO_1691 (O_1691,N_19717,N_20082);
or UO_1692 (O_1692,N_20265,N_21242);
nand UO_1693 (O_1693,N_19247,N_21454);
xnor UO_1694 (O_1694,N_22916,N_21482);
nor UO_1695 (O_1695,N_24424,N_23377);
and UO_1696 (O_1696,N_19140,N_20088);
nand UO_1697 (O_1697,N_22522,N_24668);
or UO_1698 (O_1698,N_24227,N_24742);
and UO_1699 (O_1699,N_18887,N_19889);
nor UO_1700 (O_1700,N_19411,N_22454);
and UO_1701 (O_1701,N_24167,N_24056);
nand UO_1702 (O_1702,N_20150,N_24130);
nor UO_1703 (O_1703,N_24837,N_19973);
or UO_1704 (O_1704,N_20242,N_24520);
and UO_1705 (O_1705,N_23905,N_21405);
nor UO_1706 (O_1706,N_20410,N_24819);
nand UO_1707 (O_1707,N_20981,N_21346);
or UO_1708 (O_1708,N_22467,N_22368);
or UO_1709 (O_1709,N_20130,N_20310);
or UO_1710 (O_1710,N_23750,N_24721);
or UO_1711 (O_1711,N_24704,N_20901);
and UO_1712 (O_1712,N_20900,N_18921);
or UO_1713 (O_1713,N_20863,N_24397);
nor UO_1714 (O_1714,N_19373,N_19008);
nor UO_1715 (O_1715,N_18978,N_19682);
nor UO_1716 (O_1716,N_19793,N_19971);
nor UO_1717 (O_1717,N_20091,N_24526);
nor UO_1718 (O_1718,N_19479,N_21315);
xor UO_1719 (O_1719,N_20094,N_23594);
or UO_1720 (O_1720,N_20582,N_19239);
nor UO_1721 (O_1721,N_24243,N_19904);
or UO_1722 (O_1722,N_21379,N_23608);
nor UO_1723 (O_1723,N_22842,N_23829);
and UO_1724 (O_1724,N_21262,N_23742);
or UO_1725 (O_1725,N_24593,N_23901);
nand UO_1726 (O_1726,N_18957,N_21959);
nor UO_1727 (O_1727,N_24946,N_19496);
or UO_1728 (O_1728,N_18932,N_20833);
nor UO_1729 (O_1729,N_20321,N_24274);
nor UO_1730 (O_1730,N_20430,N_23732);
and UO_1731 (O_1731,N_24300,N_22537);
and UO_1732 (O_1732,N_20297,N_20997);
nor UO_1733 (O_1733,N_21398,N_19128);
nand UO_1734 (O_1734,N_23126,N_23238);
or UO_1735 (O_1735,N_19052,N_20222);
and UO_1736 (O_1736,N_24978,N_21112);
nand UO_1737 (O_1737,N_21627,N_24531);
or UO_1738 (O_1738,N_18773,N_20753);
nor UO_1739 (O_1739,N_18828,N_21588);
or UO_1740 (O_1740,N_21153,N_24101);
and UO_1741 (O_1741,N_24315,N_19316);
or UO_1742 (O_1742,N_19927,N_20396);
and UO_1743 (O_1743,N_23445,N_19771);
nor UO_1744 (O_1744,N_23526,N_23382);
nand UO_1745 (O_1745,N_23909,N_20197);
nor UO_1746 (O_1746,N_24033,N_22054);
or UO_1747 (O_1747,N_21188,N_21698);
and UO_1748 (O_1748,N_22504,N_19722);
xor UO_1749 (O_1749,N_22300,N_21520);
nor UO_1750 (O_1750,N_22139,N_24337);
and UO_1751 (O_1751,N_23331,N_18830);
xnor UO_1752 (O_1752,N_21291,N_20590);
nand UO_1753 (O_1753,N_24725,N_19409);
xor UO_1754 (O_1754,N_19895,N_24451);
xor UO_1755 (O_1755,N_19922,N_22711);
or UO_1756 (O_1756,N_21185,N_22890);
nor UO_1757 (O_1757,N_24096,N_24591);
or UO_1758 (O_1758,N_19910,N_21541);
and UO_1759 (O_1759,N_24246,N_22495);
and UO_1760 (O_1760,N_18753,N_22141);
nor UO_1761 (O_1761,N_21466,N_22472);
xor UO_1762 (O_1762,N_24466,N_21161);
nand UO_1763 (O_1763,N_21264,N_24752);
xor UO_1764 (O_1764,N_22394,N_23518);
nand UO_1765 (O_1765,N_21176,N_23649);
nand UO_1766 (O_1766,N_20391,N_19256);
and UO_1767 (O_1767,N_23509,N_19030);
and UO_1768 (O_1768,N_24402,N_22689);
or UO_1769 (O_1769,N_21605,N_23697);
and UO_1770 (O_1770,N_21483,N_22987);
or UO_1771 (O_1771,N_22147,N_20289);
xnor UO_1772 (O_1772,N_21625,N_19282);
and UO_1773 (O_1773,N_21166,N_19702);
nor UO_1774 (O_1774,N_22046,N_23709);
nor UO_1775 (O_1775,N_24193,N_20744);
nand UO_1776 (O_1776,N_24360,N_20510);
nand UO_1777 (O_1777,N_22449,N_19458);
nand UO_1778 (O_1778,N_21811,N_21617);
nand UO_1779 (O_1779,N_21708,N_23792);
and UO_1780 (O_1780,N_22721,N_20488);
and UO_1781 (O_1781,N_23287,N_19740);
or UO_1782 (O_1782,N_20672,N_22883);
nand UO_1783 (O_1783,N_19857,N_19260);
xnor UO_1784 (O_1784,N_21160,N_22889);
nor UO_1785 (O_1785,N_22759,N_19924);
and UO_1786 (O_1786,N_22430,N_22925);
or UO_1787 (O_1787,N_20969,N_24475);
xnor UO_1788 (O_1788,N_20570,N_22419);
nor UO_1789 (O_1789,N_22435,N_22595);
or UO_1790 (O_1790,N_20871,N_23404);
and UO_1791 (O_1791,N_19650,N_23458);
or UO_1792 (O_1792,N_22044,N_23003);
and UO_1793 (O_1793,N_22542,N_20812);
or UO_1794 (O_1794,N_22476,N_22596);
nor UO_1795 (O_1795,N_24563,N_24406);
nor UO_1796 (O_1796,N_21082,N_23775);
nor UO_1797 (O_1797,N_21731,N_22532);
nor UO_1798 (O_1798,N_21797,N_21348);
xnor UO_1799 (O_1799,N_22529,N_23304);
nor UO_1800 (O_1800,N_19974,N_24716);
and UO_1801 (O_1801,N_18819,N_19033);
nand UO_1802 (O_1802,N_24008,N_21619);
nor UO_1803 (O_1803,N_23979,N_19039);
xnor UO_1804 (O_1804,N_23982,N_19711);
nor UO_1805 (O_1805,N_20571,N_21769);
nand UO_1806 (O_1806,N_23752,N_20136);
or UO_1807 (O_1807,N_24777,N_24212);
and UO_1808 (O_1808,N_22731,N_24473);
or UO_1809 (O_1809,N_24873,N_21679);
and UO_1810 (O_1810,N_24414,N_24166);
nor UO_1811 (O_1811,N_18940,N_20201);
nor UO_1812 (O_1812,N_23615,N_19080);
nand UO_1813 (O_1813,N_23571,N_21973);
xnor UO_1814 (O_1814,N_19338,N_20409);
xor UO_1815 (O_1815,N_23465,N_22634);
and UO_1816 (O_1816,N_24585,N_19404);
nor UO_1817 (O_1817,N_24897,N_23289);
nand UO_1818 (O_1818,N_24989,N_19130);
and UO_1819 (O_1819,N_21401,N_24892);
or UO_1820 (O_1820,N_19462,N_20472);
xnor UO_1821 (O_1821,N_24186,N_23639);
or UO_1822 (O_1822,N_23366,N_20380);
or UO_1823 (O_1823,N_24815,N_19048);
and UO_1824 (O_1824,N_21433,N_21078);
nand UO_1825 (O_1825,N_24722,N_19926);
nand UO_1826 (O_1826,N_22321,N_24392);
and UO_1827 (O_1827,N_24020,N_24001);
nor UO_1828 (O_1828,N_20854,N_19757);
xnor UO_1829 (O_1829,N_19473,N_21821);
nor UO_1830 (O_1830,N_24432,N_24677);
and UO_1831 (O_1831,N_23781,N_21828);
nor UO_1832 (O_1832,N_23958,N_24962);
and UO_1833 (O_1833,N_21654,N_21027);
nand UO_1834 (O_1834,N_20218,N_19112);
nor UO_1835 (O_1835,N_22716,N_21424);
or UO_1836 (O_1836,N_24321,N_24372);
and UO_1837 (O_1837,N_22970,N_22590);
nand UO_1838 (O_1838,N_22735,N_24920);
nor UO_1839 (O_1839,N_24128,N_19890);
nand UO_1840 (O_1840,N_22159,N_24613);
and UO_1841 (O_1841,N_21993,N_23567);
nor UO_1842 (O_1842,N_18811,N_24941);
nor UO_1843 (O_1843,N_22562,N_21867);
nand UO_1844 (O_1844,N_19629,N_22566);
and UO_1845 (O_1845,N_21724,N_21912);
or UO_1846 (O_1846,N_21312,N_19786);
and UO_1847 (O_1847,N_20404,N_22991);
and UO_1848 (O_1848,N_21777,N_22578);
and UO_1849 (O_1849,N_23254,N_22463);
and UO_1850 (O_1850,N_19614,N_23521);
nor UO_1851 (O_1851,N_23679,N_22099);
nand UO_1852 (O_1852,N_24206,N_24551);
nand UO_1853 (O_1853,N_23784,N_21340);
or UO_1854 (O_1854,N_24596,N_23323);
xnor UO_1855 (O_1855,N_19871,N_24614);
nor UO_1856 (O_1856,N_23955,N_22697);
nor UO_1857 (O_1857,N_19280,N_18865);
or UO_1858 (O_1858,N_23549,N_23597);
or UO_1859 (O_1859,N_24449,N_19207);
and UO_1860 (O_1860,N_21186,N_19056);
nor UO_1861 (O_1861,N_20052,N_24578);
or UO_1862 (O_1862,N_23032,N_23883);
or UO_1863 (O_1863,N_20967,N_21754);
nand UO_1864 (O_1864,N_24691,N_22276);
nor UO_1865 (O_1865,N_24619,N_19975);
nand UO_1866 (O_1866,N_24701,N_22672);
or UO_1867 (O_1867,N_20192,N_24199);
or UO_1868 (O_1868,N_23738,N_24866);
or UO_1869 (O_1869,N_22377,N_21744);
and UO_1870 (O_1870,N_18798,N_23644);
nand UO_1871 (O_1871,N_20047,N_23849);
xor UO_1872 (O_1872,N_24078,N_23641);
xnor UO_1873 (O_1873,N_24542,N_19368);
nor UO_1874 (O_1874,N_24229,N_18768);
nor UO_1875 (O_1875,N_20294,N_20307);
and UO_1876 (O_1876,N_20985,N_23347);
and UO_1877 (O_1877,N_23776,N_18885);
nand UO_1878 (O_1878,N_20267,N_20979);
and UO_1879 (O_1879,N_23474,N_20193);
nor UO_1880 (O_1880,N_24999,N_21916);
and UO_1881 (O_1881,N_23433,N_20826);
and UO_1882 (O_1882,N_24516,N_24110);
xnor UO_1883 (O_1883,N_24571,N_23920);
and UO_1884 (O_1884,N_19266,N_24164);
and UO_1885 (O_1885,N_21222,N_24205);
and UO_1886 (O_1886,N_21080,N_23000);
xnor UO_1887 (O_1887,N_21676,N_24784);
nor UO_1888 (O_1888,N_24179,N_20686);
or UO_1889 (O_1889,N_21856,N_22900);
and UO_1890 (O_1890,N_20395,N_20308);
and UO_1891 (O_1891,N_19333,N_21642);
or UO_1892 (O_1892,N_23416,N_23211);
or UO_1893 (O_1893,N_24182,N_21381);
nor UO_1894 (O_1894,N_22675,N_19955);
nor UO_1895 (O_1895,N_19818,N_23119);
or UO_1896 (O_1896,N_24403,N_23522);
or UO_1897 (O_1897,N_21705,N_24779);
nand UO_1898 (O_1898,N_21135,N_23949);
or UO_1899 (O_1899,N_20846,N_21946);
nor UO_1900 (O_1900,N_20815,N_18896);
nor UO_1901 (O_1901,N_24025,N_19297);
nor UO_1902 (O_1902,N_23121,N_23741);
nor UO_1903 (O_1903,N_23531,N_23006);
nand UO_1904 (O_1904,N_20231,N_19250);
or UO_1905 (O_1905,N_20455,N_21369);
nor UO_1906 (O_1906,N_23998,N_20095);
and UO_1907 (O_1907,N_22501,N_21570);
or UO_1908 (O_1908,N_23365,N_22060);
nand UO_1909 (O_1909,N_24342,N_18994);
nand UO_1910 (O_1910,N_20468,N_24610);
or UO_1911 (O_1911,N_23532,N_18823);
nand UO_1912 (O_1912,N_21876,N_19139);
or UO_1913 (O_1913,N_21741,N_22398);
or UO_1914 (O_1914,N_21033,N_18971);
or UO_1915 (O_1915,N_19827,N_20217);
and UO_1916 (O_1916,N_20420,N_23479);
and UO_1917 (O_1917,N_24505,N_21404);
or UO_1918 (O_1918,N_22964,N_22318);
nand UO_1919 (O_1919,N_19334,N_19907);
nand UO_1920 (O_1920,N_22374,N_22094);
or UO_1921 (O_1921,N_23375,N_21139);
or UO_1922 (O_1922,N_21664,N_22685);
nor UO_1923 (O_1923,N_20987,N_18870);
or UO_1924 (O_1924,N_20989,N_24939);
and UO_1925 (O_1925,N_19483,N_22434);
nand UO_1926 (O_1926,N_21148,N_18842);
and UO_1927 (O_1927,N_22705,N_23175);
nor UO_1928 (O_1928,N_20845,N_21611);
nor UO_1929 (O_1929,N_20882,N_22671);
nand UO_1930 (O_1930,N_22636,N_19781);
nand UO_1931 (O_1931,N_21536,N_24881);
or UO_1932 (O_1932,N_20889,N_24500);
or UO_1933 (O_1933,N_23129,N_23080);
and UO_1934 (O_1934,N_24504,N_19856);
or UO_1935 (O_1935,N_19840,N_20524);
nor UO_1936 (O_1936,N_22151,N_20471);
and UO_1937 (O_1937,N_18918,N_23112);
xor UO_1938 (O_1938,N_21517,N_19984);
nor UO_1939 (O_1939,N_20367,N_23149);
nand UO_1940 (O_1940,N_21028,N_22580);
nand UO_1941 (O_1941,N_20838,N_20268);
or UO_1942 (O_1942,N_21320,N_24429);
nor UO_1943 (O_1943,N_18889,N_19285);
or UO_1944 (O_1944,N_24413,N_23574);
and UO_1945 (O_1945,N_22393,N_23158);
or UO_1946 (O_1946,N_18984,N_23381);
nand UO_1947 (O_1947,N_19016,N_24684);
nor UO_1948 (O_1948,N_20670,N_21985);
or UO_1949 (O_1949,N_20072,N_19583);
or UO_1950 (O_1950,N_20608,N_24407);
nand UO_1951 (O_1951,N_19666,N_23399);
nand UO_1952 (O_1952,N_23264,N_23272);
and UO_1953 (O_1953,N_20532,N_24481);
nor UO_1954 (O_1954,N_20068,N_18966);
nand UO_1955 (O_1955,N_24713,N_24615);
or UO_1956 (O_1956,N_23611,N_23376);
or UO_1957 (O_1957,N_22714,N_22875);
nor UO_1958 (O_1958,N_20824,N_24582);
and UO_1959 (O_1959,N_20283,N_20384);
or UO_1960 (O_1960,N_21516,N_24039);
nor UO_1961 (O_1961,N_24089,N_19498);
nor UO_1962 (O_1962,N_19824,N_20336);
and UO_1963 (O_1963,N_21784,N_24248);
nor UO_1964 (O_1964,N_20045,N_18915);
or UO_1965 (O_1965,N_24860,N_24303);
and UO_1966 (O_1966,N_22085,N_24082);
or UO_1967 (O_1967,N_20586,N_20898);
or UO_1968 (O_1968,N_23035,N_21292);
nand UO_1969 (O_1969,N_20383,N_20452);
nand UO_1970 (O_1970,N_20674,N_19733);
nand UO_1971 (O_1971,N_19223,N_24678);
and UO_1972 (O_1972,N_20756,N_21581);
or UO_1973 (O_1973,N_20549,N_19937);
and UO_1974 (O_1974,N_18996,N_23455);
and UO_1975 (O_1975,N_19437,N_23290);
and UO_1976 (O_1976,N_23588,N_22682);
nor UO_1977 (O_1977,N_20229,N_22619);
or UO_1978 (O_1978,N_19363,N_23910);
and UO_1979 (O_1979,N_20895,N_18975);
nor UO_1980 (O_1980,N_23486,N_23603);
xnor UO_1981 (O_1981,N_23779,N_22008);
or UO_1982 (O_1982,N_23460,N_21949);
or UO_1983 (O_1983,N_23906,N_23135);
and UO_1984 (O_1984,N_19807,N_19412);
nand UO_1985 (O_1985,N_21858,N_22732);
nand UO_1986 (O_1986,N_20475,N_23527);
xor UO_1987 (O_1987,N_23360,N_23851);
xor UO_1988 (O_1988,N_24222,N_24454);
nor UO_1989 (O_1989,N_21638,N_20629);
nor UO_1990 (O_1990,N_21838,N_24367);
xnor UO_1991 (O_1991,N_20792,N_21067);
nor UO_1992 (O_1992,N_18967,N_19551);
nor UO_1993 (O_1993,N_21978,N_23788);
and UO_1994 (O_1994,N_24165,N_23241);
xor UO_1995 (O_1995,N_20338,N_21800);
nand UO_1996 (O_1996,N_19319,N_22692);
or UO_1997 (O_1997,N_18838,N_23946);
nor UO_1998 (O_1998,N_22286,N_19310);
nor UO_1999 (O_1999,N_20327,N_19159);
and UO_2000 (O_2000,N_22894,N_23487);
nand UO_2001 (O_2001,N_22793,N_24379);
nor UO_2002 (O_2002,N_19532,N_22371);
nand UO_2003 (O_2003,N_22135,N_21276);
or UO_2004 (O_2004,N_23325,N_24104);
or UO_2005 (O_2005,N_18871,N_20706);
xor UO_2006 (O_2006,N_20368,N_21443);
and UO_2007 (O_2007,N_20254,N_20905);
and UO_2008 (O_2008,N_22839,N_20497);
nand UO_2009 (O_2009,N_24333,N_22679);
or UO_2010 (O_2010,N_19394,N_23566);
nand UO_2011 (O_2011,N_21889,N_24194);
nand UO_2012 (O_2012,N_22860,N_18799);
nand UO_2013 (O_2013,N_22774,N_24489);
or UO_2014 (O_2014,N_22388,N_22048);
and UO_2015 (O_2015,N_20841,N_22129);
or UO_2016 (O_2016,N_23302,N_23148);
nand UO_2017 (O_2017,N_21579,N_22723);
nand UO_2018 (O_2018,N_24311,N_20564);
nor UO_2019 (O_2019,N_23683,N_19853);
nor UO_2020 (O_2020,N_20421,N_20530);
nand UO_2021 (O_2021,N_19893,N_24258);
nand UO_2022 (O_2022,N_24605,N_21534);
nor UO_2023 (O_2023,N_21743,N_19119);
and UO_2024 (O_2024,N_23198,N_21008);
nor UO_2025 (O_2025,N_19194,N_21560);
or UO_2026 (O_2026,N_19279,N_18986);
nor UO_2027 (O_2027,N_23660,N_18859);
xor UO_2028 (O_2028,N_21540,N_22189);
and UO_2029 (O_2029,N_22850,N_20438);
nand UO_2030 (O_2030,N_21246,N_20956);
or UO_2031 (O_2031,N_21928,N_19399);
and UO_2032 (O_2032,N_21773,N_24984);
nor UO_2033 (O_2033,N_20419,N_23716);
and UO_2034 (O_2034,N_20232,N_19961);
nor UO_2035 (O_2035,N_20256,N_20537);
and UO_2036 (O_2036,N_19708,N_21826);
nor UO_2037 (O_2037,N_23703,N_22169);
and UO_2038 (O_2038,N_23606,N_23801);
and UO_2039 (O_2039,N_24804,N_23626);
and UO_2040 (O_2040,N_21284,N_18873);
and UO_2041 (O_2041,N_20085,N_21143);
or UO_2042 (O_2042,N_20454,N_19019);
nor UO_2043 (O_2043,N_19518,N_23204);
nor UO_2044 (O_2044,N_21640,N_18938);
nor UO_2045 (O_2045,N_20731,N_21504);
xnor UO_2046 (O_2046,N_19049,N_20478);
or UO_2047 (O_2047,N_23131,N_24976);
or UO_2048 (O_2048,N_19367,N_22741);
nand UO_2049 (O_2049,N_24709,N_21412);
or UO_2050 (O_2050,N_23123,N_24734);
nor UO_2051 (O_2051,N_22030,N_22441);
xnor UO_2052 (O_2052,N_22192,N_22746);
nor UO_2053 (O_2053,N_19553,N_22365);
or UO_2054 (O_2054,N_20928,N_19183);
nor UO_2055 (O_2055,N_21409,N_23297);
and UO_2056 (O_2056,N_22027,N_19320);
and UO_2057 (O_2057,N_23675,N_24422);
xor UO_2058 (O_2058,N_19350,N_23147);
or UO_2059 (O_2059,N_24160,N_23948);
nand UO_2060 (O_2060,N_21321,N_21673);
and UO_2061 (O_2061,N_19407,N_18754);
nor UO_2062 (O_2062,N_23915,N_23795);
or UO_2063 (O_2063,N_19623,N_19600);
or UO_2064 (O_2064,N_22829,N_21667);
nand UO_2065 (O_2065,N_24074,N_22990);
nand UO_2066 (O_2066,N_19915,N_19712);
nand UO_2067 (O_2067,N_23689,N_23860);
nor UO_2068 (O_2068,N_22962,N_20760);
nor UO_2069 (O_2069,N_23830,N_24695);
and UO_2070 (O_2070,N_20470,N_21760);
nand UO_2071 (O_2071,N_19565,N_24000);
nand UO_2072 (O_2072,N_19626,N_19810);
and UO_2073 (O_2073,N_23481,N_19038);
nand UO_2074 (O_2074,N_21091,N_19484);
or UO_2075 (O_2075,N_21217,N_20865);
and UO_2076 (O_2076,N_19652,N_24287);
and UO_2077 (O_2077,N_22493,N_22080);
and UO_2078 (O_2078,N_19434,N_22888);
nor UO_2079 (O_2079,N_20278,N_23463);
nand UO_2080 (O_2080,N_18935,N_24240);
xor UO_2081 (O_2081,N_20042,N_23261);
nor UO_2082 (O_2082,N_20245,N_18987);
or UO_2083 (O_2083,N_21632,N_24769);
nor UO_2084 (O_2084,N_22862,N_21607);
or UO_2085 (O_2085,N_21269,N_22389);
nor UO_2086 (O_2086,N_19690,N_23061);
xor UO_2087 (O_2087,N_24898,N_19276);
nand UO_2088 (O_2088,N_20508,N_23450);
nand UO_2089 (O_2089,N_19323,N_18924);
nor UO_2090 (O_2090,N_20083,N_19295);
and UO_2091 (O_2091,N_22802,N_18795);
nor UO_2092 (O_2092,N_22488,N_19522);
nand UO_2093 (O_2093,N_24118,N_24598);
or UO_2094 (O_2094,N_19248,N_19921);
nor UO_2095 (O_2095,N_20365,N_20521);
or UO_2096 (O_2096,N_20881,N_21521);
nor UO_2097 (O_2097,N_21468,N_22587);
and UO_2098 (O_2098,N_24052,N_20049);
and UO_2099 (O_2099,N_24628,N_23887);
nor UO_2100 (O_2100,N_21180,N_23104);
nor UO_2101 (O_2101,N_22730,N_22910);
nor UO_2102 (O_2102,N_19577,N_21173);
nand UO_2103 (O_2103,N_20994,N_19035);
and UO_2104 (O_2104,N_20918,N_20980);
and UO_2105 (O_2105,N_20272,N_22898);
nor UO_2106 (O_2106,N_24156,N_23818);
or UO_2107 (O_2107,N_24846,N_24665);
or UO_2108 (O_2108,N_22605,N_21853);
or UO_2109 (O_2109,N_24463,N_22003);
or UO_2110 (O_2110,N_18956,N_20866);
and UO_2111 (O_2111,N_24524,N_24145);
and UO_2112 (O_2112,N_24983,N_24244);
and UO_2113 (O_2113,N_24458,N_21467);
nand UO_2114 (O_2114,N_24241,N_24657);
or UO_2115 (O_2115,N_24371,N_18856);
nand UO_2116 (O_2116,N_23995,N_18750);
nand UO_2117 (O_2117,N_23282,N_21693);
xnor UO_2118 (O_2118,N_19536,N_19315);
nand UO_2119 (O_2119,N_18763,N_23233);
nor UO_2120 (O_2120,N_21719,N_20361);
and UO_2121 (O_2121,N_24934,N_23573);
or UO_2122 (O_2122,N_23951,N_20709);
or UO_2123 (O_2123,N_19195,N_20935);
nor UO_2124 (O_2124,N_24840,N_21939);
xnor UO_2125 (O_2125,N_23577,N_19121);
or UO_2126 (O_2126,N_20923,N_20402);
and UO_2127 (O_2127,N_22552,N_20899);
nor UO_2128 (O_2128,N_19909,N_19539);
nand UO_2129 (O_2129,N_19879,N_19880);
nor UO_2130 (O_2130,N_24829,N_21129);
and UO_2131 (O_2131,N_23150,N_20696);
nand UO_2132 (O_2132,N_23398,N_24264);
or UO_2133 (O_2133,N_20619,N_20190);
nand UO_2134 (O_2134,N_23321,N_23777);
nor UO_2135 (O_2135,N_19264,N_24065);
and UO_2136 (O_2136,N_23133,N_21444);
and UO_2137 (O_2137,N_21542,N_21882);
nand UO_2138 (O_2138,N_24560,N_21384);
or UO_2139 (O_2139,N_21613,N_19520);
nor UO_2140 (O_2140,N_18912,N_20599);
nand UO_2141 (O_2141,N_23009,N_19669);
and UO_2142 (O_2142,N_19292,N_21620);
or UO_2143 (O_2143,N_21772,N_20318);
and UO_2144 (O_2144,N_19883,N_22294);
and UO_2145 (O_2145,N_24645,N_24214);
and UO_2146 (O_2146,N_19270,N_24974);
nor UO_2147 (O_2147,N_23841,N_22002);
nor UO_2148 (O_2148,N_20131,N_18963);
and UO_2149 (O_2149,N_24774,N_22450);
nor UO_2150 (O_2150,N_19643,N_19396);
nor UO_2151 (O_2151,N_19739,N_23512);
and UO_2152 (O_2152,N_22857,N_23417);
nor UO_2153 (O_2153,N_20660,N_24584);
nor UO_2154 (O_2154,N_22978,N_19990);
nor UO_2155 (O_2155,N_22787,N_23551);
nand UO_2156 (O_2156,N_21372,N_22382);
and UO_2157 (O_2157,N_23525,N_22378);
nor UO_2158 (O_2158,N_22940,N_24329);
nor UO_2159 (O_2159,N_19109,N_19637);
nor UO_2160 (O_2160,N_23911,N_24037);
xnor UO_2161 (O_2161,N_24054,N_24308);
xnor UO_2162 (O_2162,N_21073,N_19485);
xor UO_2163 (O_2163,N_24597,N_20381);
or UO_2164 (O_2164,N_22132,N_20886);
or UO_2165 (O_2165,N_23269,N_22239);
xor UO_2166 (O_2166,N_19196,N_19658);
nor UO_2167 (O_2167,N_20577,N_19135);
nor UO_2168 (O_2168,N_19062,N_19923);
nor UO_2169 (O_2169,N_19693,N_23160);
or UO_2170 (O_2170,N_19521,N_22292);
or UO_2171 (O_2171,N_24273,N_19103);
nor UO_2172 (O_2172,N_20019,N_21539);
nor UO_2173 (O_2173,N_21480,N_20056);
and UO_2174 (O_2174,N_19555,N_20880);
and UO_2175 (O_2175,N_20585,N_23774);
nand UO_2176 (O_2176,N_19289,N_20728);
and UO_2177 (O_2177,N_20330,N_21128);
nor UO_2178 (O_2178,N_18817,N_23629);
nor UO_2179 (O_2179,N_23140,N_24751);
or UO_2180 (O_2180,N_19762,N_24959);
or UO_2181 (O_2181,N_20364,N_19665);
nor UO_2182 (O_2182,N_22343,N_22459);
and UO_2183 (O_2183,N_23802,N_20282);
and UO_2184 (O_2184,N_19186,N_20195);
and UO_2185 (O_2185,N_19075,N_23613);
and UO_2186 (O_2186,N_19977,N_20758);
nand UO_2187 (O_2187,N_24228,N_19691);
or UO_2188 (O_2188,N_19804,N_18840);
nor UO_2189 (O_2189,N_20099,N_21305);
and UO_2190 (O_2190,N_22555,N_22420);
nand UO_2191 (O_2191,N_19491,N_23113);
nand UO_2192 (O_2192,N_19115,N_21860);
nor UO_2193 (O_2193,N_23621,N_23746);
or UO_2194 (O_2194,N_24796,N_19213);
or UO_2195 (O_2195,N_20515,N_18953);
and UO_2196 (O_2196,N_19696,N_19561);
and UO_2197 (O_2197,N_23274,N_22680);
or UO_2198 (O_2198,N_23622,N_21336);
and UO_2199 (O_2199,N_23957,N_20737);
or UO_2200 (O_2200,N_19508,N_22381);
and UO_2201 (O_2201,N_23351,N_22053);
nand UO_2202 (O_2202,N_23352,N_23267);
and UO_2203 (O_2203,N_23012,N_19618);
and UO_2204 (O_2204,N_24843,N_22483);
or UO_2205 (O_2205,N_19511,N_21355);
or UO_2206 (O_2206,N_19476,N_21072);
nor UO_2207 (O_2207,N_22550,N_24464);
nand UO_2208 (O_2208,N_21426,N_22782);
or UO_2209 (O_2209,N_22983,N_23441);
nand UO_2210 (O_2210,N_24697,N_21125);
nor UO_2211 (O_2211,N_19777,N_24440);
nor UO_2212 (O_2212,N_22422,N_20978);
xnor UO_2213 (O_2213,N_19461,N_19741);
and UO_2214 (O_2214,N_24359,N_21599);
xor UO_2215 (O_2215,N_20355,N_22223);
nor UO_2216 (O_2216,N_23548,N_21402);
nor UO_2217 (O_2217,N_19659,N_19335);
or UO_2218 (O_2218,N_19588,N_20176);
xor UO_2219 (O_2219,N_21999,N_20209);
and UO_2220 (O_2220,N_22486,N_19081);
nand UO_2221 (O_2221,N_19177,N_24232);
nand UO_2222 (O_2222,N_23989,N_22615);
xor UO_2223 (O_2223,N_21510,N_24328);
xnor UO_2224 (O_2224,N_22020,N_23462);
nand UO_2225 (O_2225,N_24155,N_20349);
and UO_2226 (O_2226,N_23004,N_20407);
nand UO_2227 (O_2227,N_21407,N_24530);
or UO_2228 (O_2228,N_20761,N_24014);
and UO_2229 (O_2229,N_19210,N_22559);
xnor UO_2230 (O_2230,N_20885,N_19331);
nand UO_2231 (O_2231,N_22214,N_22879);
nand UO_2232 (O_2232,N_19692,N_19645);
or UO_2233 (O_2233,N_22558,N_20035);
nand UO_2234 (O_2234,N_19674,N_23235);
nand UO_2235 (O_2235,N_23981,N_21901);
nor UO_2236 (O_2236,N_20949,N_20584);
and UO_2237 (O_2237,N_22124,N_21207);
nor UO_2238 (O_2238,N_23695,N_21960);
nand UO_2239 (O_2239,N_24629,N_23847);
nand UO_2240 (O_2240,N_21623,N_18850);
nor UO_2241 (O_2241,N_21591,N_20110);
or UO_2242 (O_2242,N_23692,N_19604);
or UO_2243 (O_2243,N_21966,N_20561);
nor UO_2244 (O_2244,N_20255,N_20558);
nor UO_2245 (O_2245,N_24351,N_24487);
nand UO_2246 (O_2246,N_20675,N_21961);
nor UO_2247 (O_2247,N_23476,N_21861);
nor UO_2248 (O_2248,N_24590,N_20767);
and UO_2249 (O_2249,N_19171,N_21487);
and UO_2250 (O_2250,N_21792,N_20568);
nor UO_2251 (O_2251,N_23659,N_18988);
or UO_2252 (O_2252,N_22290,N_24377);
nor UO_2253 (O_2253,N_20957,N_20593);
and UO_2254 (O_2254,N_20727,N_24747);
or UO_2255 (O_2255,N_22844,N_23897);
nand UO_2256 (O_2256,N_20057,N_23797);
and UO_2257 (O_2257,N_22126,N_24849);
nor UO_2258 (O_2258,N_21347,N_21633);
or UO_2259 (O_2259,N_20982,N_21146);
nor UO_2260 (O_2260,N_22643,N_22238);
and UO_2261 (O_2261,N_22267,N_21392);
nor UO_2262 (O_2262,N_20360,N_19465);
nand UO_2263 (O_2263,N_18877,N_19460);
and UO_2264 (O_2264,N_18826,N_20719);
nand UO_2265 (O_2265,N_19445,N_21244);
or UO_2266 (O_2266,N_22776,N_19385);
and UO_2267 (O_2267,N_24537,N_19636);
nor UO_2268 (O_2268,N_24958,N_24558);
nor UO_2269 (O_2269,N_19678,N_21554);
or UO_2270 (O_2270,N_21061,N_22571);
xor UO_2271 (O_2271,N_24497,N_23838);
and UO_2272 (O_2272,N_20529,N_19755);
nor UO_2273 (O_2273,N_20610,N_19695);
nand UO_2274 (O_2274,N_20936,N_21958);
and UO_2275 (O_2275,N_24676,N_22989);
and UO_2276 (O_2276,N_23601,N_24175);
xnor UO_2277 (O_2277,N_23484,N_19015);
or UO_2278 (O_2278,N_23440,N_22849);
and UO_2279 (O_2279,N_24326,N_19802);
and UO_2280 (O_2280,N_23277,N_23991);
or UO_2281 (O_2281,N_19504,N_21566);
nor UO_2282 (O_2282,N_19448,N_18836);
nor UO_2283 (O_2283,N_19089,N_23990);
and UO_2284 (O_2284,N_21699,N_21974);
and UO_2285 (O_2285,N_24663,N_24013);
nand UO_2286 (O_2286,N_18751,N_19908);
or UO_2287 (O_2287,N_19257,N_22547);
or UO_2288 (O_2288,N_21344,N_21458);
xor UO_2289 (O_2289,N_19332,N_23411);
nor UO_2290 (O_2290,N_20071,N_22957);
nand UO_2291 (O_2291,N_21702,N_23096);
and UO_2292 (O_2292,N_23739,N_22686);
nand UO_2293 (O_2293,N_21252,N_23146);
or UO_2294 (O_2294,N_24854,N_19122);
nor UO_2295 (O_2295,N_21107,N_22851);
nor UO_2296 (O_2296,N_20929,N_19680);
nor UO_2297 (O_2297,N_24344,N_22568);
xor UO_2298 (O_2298,N_20647,N_20687);
nor UO_2299 (O_2299,N_23569,N_23782);
and UO_2300 (O_2300,N_24550,N_20801);
nand UO_2301 (O_2301,N_20618,N_24818);
nand UO_2302 (O_2302,N_22541,N_21789);
or UO_2303 (O_2303,N_20089,N_21597);
nand UO_2304 (O_2304,N_22748,N_24181);
xnor UO_2305 (O_2305,N_22715,N_23971);
nor UO_2306 (O_2306,N_20639,N_20793);
and UO_2307 (O_2307,N_19770,N_20251);
and UO_2308 (O_2308,N_22102,N_19754);
xor UO_2309 (O_2309,N_22979,N_22250);
and UO_2310 (O_2310,N_24982,N_23842);
and UO_2311 (O_2311,N_24872,N_23098);
and UO_2312 (O_2312,N_21730,N_23052);
nor UO_2313 (O_2313,N_21929,N_22108);
nor UO_2314 (O_2314,N_21608,N_21903);
nor UO_2315 (O_2315,N_24740,N_23743);
nor UO_2316 (O_2316,N_19028,N_22858);
and UO_2317 (O_2317,N_24085,N_21062);
or UO_2318 (O_2318,N_19317,N_23827);
and UO_2319 (O_2319,N_19558,N_23472);
or UO_2320 (O_2320,N_23625,N_21644);
nor UO_2321 (O_2321,N_20576,N_24594);
or UO_2322 (O_2322,N_24930,N_22972);
or UO_2323 (O_2323,N_21137,N_21155);
and UO_2324 (O_2324,N_24960,N_23348);
nor UO_2325 (O_2325,N_24802,N_24786);
and UO_2326 (O_2326,N_20121,N_21474);
nor UO_2327 (O_2327,N_20840,N_22810);
or UO_2328 (O_2328,N_19495,N_22433);
and UO_2329 (O_2329,N_21124,N_19481);
nand UO_2330 (O_2330,N_20075,N_24430);
nand UO_2331 (O_2331,N_22976,N_21203);
nor UO_2332 (O_2332,N_19072,N_24068);
nor UO_2333 (O_2333,N_22625,N_20487);
and UO_2334 (O_2334,N_19235,N_23451);
or UO_2335 (O_2335,N_21150,N_19850);
nand UO_2336 (O_2336,N_24589,N_18901);
nand UO_2337 (O_2337,N_21274,N_20422);
and UO_2338 (O_2338,N_24764,N_22346);
nand UO_2339 (O_2339,N_23237,N_24848);
or UO_2340 (O_2340,N_20483,N_21382);
or UO_2341 (O_2341,N_19593,N_21237);
or UO_2342 (O_2342,N_22499,N_23820);
nand UO_2343 (O_2343,N_20179,N_19868);
or UO_2344 (O_2344,N_20543,N_24401);
or UO_2345 (O_2345,N_23124,N_23029);
xnor UO_2346 (O_2346,N_19487,N_20221);
nor UO_2347 (O_2347,N_22947,N_20298);
or UO_2348 (O_2348,N_21177,N_23186);
nor UO_2349 (O_2349,N_21519,N_21910);
nor UO_2350 (O_2350,N_21603,N_21710);
nand UO_2351 (O_2351,N_24265,N_20117);
nor UO_2352 (O_2352,N_24382,N_22161);
and UO_2353 (O_2353,N_19982,N_19209);
or UO_2354 (O_2354,N_23593,N_22709);
xnor UO_2355 (O_2355,N_23953,N_23655);
nor UO_2356 (O_2356,N_20241,N_23002);
nand UO_2357 (O_2357,N_20560,N_21019);
and UO_2358 (O_2358,N_20415,N_19361);
and UO_2359 (O_2359,N_20847,N_20128);
nor UO_2360 (O_2360,N_21818,N_18944);
nand UO_2361 (O_2361,N_19450,N_23925);
and UO_2362 (O_2362,N_23595,N_21429);
nand UO_2363 (O_2363,N_20358,N_23806);
or UO_2364 (O_2364,N_19962,N_24226);
nor UO_2365 (O_2365,N_21492,N_23672);
and UO_2366 (O_2366,N_19500,N_18796);
and UO_2367 (O_2367,N_23300,N_24169);
nor UO_2368 (O_2368,N_20638,N_24825);
nand UO_2369 (O_2369,N_19044,N_19557);
nor UO_2370 (O_2370,N_23562,N_21610);
nor UO_2371 (O_2371,N_24419,N_20940);
or UO_2372 (O_2372,N_22484,N_21738);
nor UO_2373 (O_2373,N_19917,N_19601);
nor UO_2374 (O_2374,N_18982,N_24081);
nor UO_2375 (O_2375,N_19061,N_22100);
nor UO_2376 (O_2376,N_21734,N_20362);
nor UO_2377 (O_2377,N_20640,N_20258);
and UO_2378 (O_2378,N_24649,N_24370);
and UO_2379 (O_2379,N_20142,N_22992);
and UO_2380 (O_2380,N_22519,N_23478);
nand UO_2381 (O_2381,N_23214,N_21626);
or UO_2382 (O_2382,N_24314,N_23914);
xnor UO_2383 (O_2383,N_22270,N_21198);
xnor UO_2384 (O_2384,N_23403,N_20237);
or UO_2385 (O_2385,N_19938,N_22551);
nor UO_2386 (O_2386,N_22424,N_21461);
nand UO_2387 (O_2387,N_19150,N_23570);
nand UO_2388 (O_2388,N_19954,N_22699);
nor UO_2389 (O_2389,N_19792,N_20246);
and UO_2390 (O_2390,N_20339,N_21009);
or UO_2391 (O_2391,N_23785,N_24278);
or UO_2392 (O_2392,N_22836,N_21130);
and UO_2393 (O_2393,N_23656,N_20009);
nand UO_2394 (O_2394,N_19987,N_24004);
or UO_2395 (O_2395,N_21195,N_22156);
and UO_2396 (O_2396,N_22534,N_23754);
nand UO_2397 (O_2397,N_21326,N_24306);
nand UO_2398 (O_2398,N_19571,N_20399);
nor UO_2399 (O_2399,N_21682,N_22462);
or UO_2400 (O_2400,N_20469,N_23262);
or UO_2401 (O_2401,N_20764,N_23073);
or UO_2402 (O_2402,N_21689,N_23305);
nor UO_2403 (O_2403,N_18769,N_22602);
or UO_2404 (O_2404,N_24136,N_24903);
and UO_2405 (O_2405,N_22313,N_24320);
nor UO_2406 (O_2406,N_18814,N_20296);
nand UO_2407 (O_2407,N_24798,N_19823);
and UO_2408 (O_2408,N_19275,N_24830);
nand UO_2409 (O_2409,N_24640,N_24653);
or UO_2410 (O_2410,N_22412,N_19745);
or UO_2411 (O_2411,N_24021,N_22391);
or UO_2412 (O_2412,N_20519,N_19078);
nor UO_2413 (O_2413,N_23196,N_21692);
or UO_2414 (O_2414,N_21064,N_23528);
nand UO_2415 (O_2415,N_24319,N_24733);
nand UO_2416 (O_2416,N_22237,N_24485);
xor UO_2417 (O_2417,N_18759,N_20334);
nor UO_2418 (O_2418,N_24969,N_20535);
or UO_2419 (O_2419,N_21256,N_19226);
xnor UO_2420 (O_2420,N_23550,N_23050);
or UO_2421 (O_2421,N_20163,N_22193);
nor UO_2422 (O_2422,N_20950,N_19852);
and UO_2423 (O_2423,N_22592,N_21485);
xor UO_2424 (O_2424,N_22304,N_21799);
nor UO_2425 (O_2425,N_21780,N_19231);
nand UO_2426 (O_2426,N_23994,N_20860);
and UO_2427 (O_2427,N_23191,N_22548);
nor UO_2428 (O_2428,N_24886,N_19425);
nor UO_2429 (O_2429,N_20635,N_21586);
and UO_2430 (O_2430,N_20406,N_22314);
and UO_2431 (O_2431,N_21031,N_22312);
nor UO_2432 (O_2432,N_20371,N_19795);
or UO_2433 (O_2433,N_22478,N_19000);
nand UO_2434 (O_2434,N_21319,N_20903);
nor UO_2435 (O_2435,N_21670,N_18933);
nor UO_2436 (O_2436,N_19544,N_21494);
or UO_2437 (O_2437,N_19134,N_23023);
xnor UO_2438 (O_2438,N_23758,N_21015);
nor UO_2439 (O_2439,N_20562,N_22934);
nor UO_2440 (O_2440,N_19833,N_20759);
or UO_2441 (O_2441,N_22610,N_24922);
nand UO_2442 (O_2442,N_23727,N_20546);
or UO_2443 (O_2443,N_18834,N_20092);
xor UO_2444 (O_2444,N_19627,N_22781);
or UO_2445 (O_2445,N_23873,N_21303);
or UO_2446 (O_2446,N_24122,N_24364);
nor UO_2447 (O_2447,N_24800,N_20313);
or UO_2448 (O_2448,N_20820,N_21308);
and UO_2449 (O_2449,N_22428,N_23015);
nand UO_2450 (O_2450,N_22442,N_20494);
nor UO_2451 (O_2451,N_20722,N_22811);
and UO_2452 (O_2452,N_21624,N_20602);
xor UO_2453 (O_2453,N_23346,N_22586);
nand UO_2454 (O_2454,N_21338,N_20720);
nor UO_2455 (O_2455,N_20079,N_18907);
and UO_2456 (O_2456,N_19387,N_21561);
nand UO_2457 (O_2457,N_21006,N_20067);
or UO_2458 (O_2458,N_22554,N_19302);
nor UO_2459 (O_2459,N_18818,N_23489);
nand UO_2460 (O_2460,N_24907,N_21097);
or UO_2461 (O_2461,N_19980,N_22574);
nand UO_2462 (O_2462,N_23001,N_21768);
nand UO_2463 (O_2463,N_18923,N_23554);
and UO_2464 (O_2464,N_23108,N_21287);
nor UO_2465 (O_2465,N_23231,N_22083);
nor UO_2466 (O_2466,N_23575,N_23928);
nor UO_2467 (O_2467,N_22808,N_22207);
or UO_2468 (O_2468,N_22049,N_24943);
or UO_2469 (O_2469,N_24908,N_21259);
nor UO_2470 (O_2470,N_24318,N_19688);
and UO_2471 (O_2471,N_23885,N_18809);
and UO_2472 (O_2472,N_23122,N_20133);
or UO_2473 (O_2473,N_22175,N_23817);
xnor UO_2474 (O_2474,N_20580,N_23899);
or UO_2475 (O_2475,N_22362,N_18914);
nand UO_2476 (O_2476,N_23616,N_19384);
nor UO_2477 (O_2477,N_21817,N_23963);
or UO_2478 (O_2478,N_21971,N_18970);
or UO_2479 (O_2479,N_24724,N_24335);
and UO_2480 (O_2480,N_22870,N_24259);
and UO_2481 (O_2481,N_21102,N_20353);
xor UO_2482 (O_2482,N_21121,N_23223);
or UO_2483 (O_2483,N_20877,N_22407);
and UO_2484 (O_2484,N_19021,N_20516);
and UO_2485 (O_2485,N_22037,N_24478);
nor UO_2486 (O_2486,N_20347,N_21501);
nor UO_2487 (O_2487,N_24509,N_18977);
nand UO_2488 (O_2488,N_19941,N_22047);
and UO_2489 (O_2489,N_23907,N_22717);
or UO_2490 (O_2490,N_20250,N_23576);
nor UO_2491 (O_2491,N_23212,N_20613);
nand UO_2492 (O_2492,N_24461,N_19732);
nand UO_2493 (O_2493,N_24817,N_24688);
nor UO_2494 (O_2494,N_21668,N_22194);
xor UO_2495 (O_2495,N_22465,N_20708);
nand UO_2496 (O_2496,N_22295,N_21341);
or UO_2497 (O_2497,N_21059,N_23839);
and UO_2498 (O_2498,N_19720,N_22932);
or UO_2499 (O_2499,N_20567,N_23493);
xnor UO_2500 (O_2500,N_24707,N_21210);
or UO_2501 (O_2501,N_19424,N_23291);
and UO_2502 (O_2502,N_22982,N_19148);
or UO_2503 (O_2503,N_22162,N_19764);
nor UO_2504 (O_2504,N_24341,N_24491);
nor UO_2505 (O_2505,N_21977,N_22882);
nand UO_2506 (O_2506,N_21987,N_22824);
nand UO_2507 (O_2507,N_21313,N_21110);
or UO_2508 (O_2508,N_21298,N_23097);
or UO_2509 (O_2509,N_19873,N_24357);
nand UO_2510 (O_2510,N_19118,N_24381);
or UO_2511 (O_2511,N_19512,N_22410);
or UO_2512 (O_2512,N_22195,N_20116);
or UO_2513 (O_2513,N_19753,N_19064);
xor UO_2514 (O_2514,N_21836,N_19567);
xor UO_2515 (O_2515,N_19166,N_19007);
and UO_2516 (O_2516,N_24404,N_19125);
nor UO_2517 (O_2517,N_21089,N_19950);
or UO_2518 (O_2518,N_19651,N_20107);
nor UO_2519 (O_2519,N_20073,N_22105);
xnor UO_2520 (O_2520,N_24744,N_22943);
and UO_2521 (O_2521,N_21808,N_23337);
nand UO_2522 (O_2522,N_22606,N_18760);
and UO_2523 (O_2523,N_18846,N_21872);
or UO_2524 (O_2524,N_24433,N_23085);
and UO_2525 (O_2525,N_18976,N_19671);
and UO_2526 (O_2526,N_24095,N_19287);
nand UO_2527 (O_2527,N_22755,N_22601);
and UO_2528 (O_2528,N_24883,N_22533);
and UO_2529 (O_2529,N_23923,N_20320);
and UO_2530 (O_2530,N_21652,N_22058);
or UO_2531 (O_2531,N_24638,N_23485);
nor UO_2532 (O_2532,N_21950,N_23488);
and UO_2533 (O_2533,N_23334,N_22040);
nor UO_2534 (O_2534,N_22863,N_24057);
nor UO_2535 (O_2535,N_22651,N_24625);
or UO_2536 (O_2536,N_24745,N_19698);
and UO_2537 (O_2537,N_21578,N_21628);
and UO_2538 (O_2538,N_23926,N_24492);
xor UO_2539 (O_2539,N_21208,N_21918);
or UO_2540 (O_2540,N_22322,N_19220);
and UO_2541 (O_2541,N_20677,N_24757);
or UO_2542 (O_2542,N_20808,N_20342);
or UO_2543 (O_2543,N_20606,N_20493);
nand UO_2544 (O_2544,N_21045,N_21571);
xnor UO_2545 (O_2545,N_20504,N_21011);
xor UO_2546 (O_2546,N_21024,N_24313);
nand UO_2547 (O_2547,N_22041,N_24347);
nor UO_2548 (O_2548,N_21945,N_19151);
and UO_2549 (O_2549,N_20813,N_20884);
and UO_2550 (O_2550,N_19389,N_19175);
or UO_2551 (O_2551,N_20394,N_22847);
nor UO_2552 (O_2552,N_21286,N_23628);
nor UO_2553 (O_2553,N_24968,N_21851);
and UO_2554 (O_2554,N_19329,N_20403);
nand UO_2555 (O_2555,N_20735,N_21416);
nand UO_2556 (O_2556,N_22669,N_19644);
xor UO_2557 (O_2557,N_20626,N_22620);
or UO_2558 (O_2558,N_23408,N_19989);
xor UO_2559 (O_2559,N_24527,N_24031);
or UO_2560 (O_2560,N_22778,N_20189);
or UO_2561 (O_2561,N_21317,N_21035);
and UO_2562 (O_2562,N_21475,N_19325);
or UO_2563 (O_2563,N_21844,N_19615);
nand UO_2564 (O_2564,N_20331,N_21049);
and UO_2565 (O_2565,N_24536,N_21774);
nor UO_2566 (O_2566,N_22513,N_22924);
nor UO_2567 (O_2567,N_20680,N_24575);
or UO_2568 (O_2568,N_24822,N_19454);
and UO_2569 (O_2569,N_20473,N_20129);
nand UO_2570 (O_2570,N_20259,N_20679);
nor UO_2571 (O_2571,N_20849,N_20933);
nor UO_2572 (O_2572,N_20280,N_21580);
nand UO_2573 (O_2573,N_19592,N_22288);
nand UO_2574 (O_2574,N_20427,N_21756);
nor UO_2575 (O_2575,N_24914,N_22479);
and UO_2576 (O_2576,N_23918,N_20627);
nor UO_2577 (O_2577,N_24620,N_19528);
and UO_2578 (O_2578,N_24833,N_22922);
nand UO_2579 (O_2579,N_23718,N_22520);
and UO_2580 (O_2580,N_24277,N_23394);
nor UO_2581 (O_2581,N_21290,N_21963);
nor UO_2582 (O_2582,N_22211,N_20752);
nor UO_2583 (O_2583,N_20295,N_23586);
nor UO_2584 (O_2584,N_21600,N_22174);
nand UO_2585 (O_2585,N_22930,N_24484);
nand UO_2586 (O_2586,N_18882,N_21096);
or UO_2587 (O_2587,N_19661,N_22740);
nand UO_2588 (O_2588,N_20601,N_20288);
nand UO_2589 (O_2589,N_21815,N_19306);
nor UO_2590 (O_2590,N_24317,N_20111);
or UO_2591 (O_2591,N_19834,N_23047);
or UO_2592 (O_2592,N_24687,N_23720);
nor UO_2593 (O_2593,N_23086,N_20436);
nor UO_2594 (O_2594,N_22076,N_22647);
or UO_2595 (O_2595,N_19738,N_24292);
and UO_2596 (O_2596,N_21342,N_23821);
nand UO_2597 (O_2597,N_22665,N_23799);
and UO_2598 (O_2598,N_22205,N_23295);
or UO_2599 (O_2599,N_23093,N_21875);
nor UO_2600 (O_2600,N_19097,N_24775);
or UO_2601 (O_2601,N_19170,N_24022);
nor UO_2602 (O_2602,N_21896,N_23081);
and UO_2603 (O_2603,N_22814,N_19232);
or UO_2604 (O_2604,N_20208,N_21547);
nor UO_2605 (O_2605,N_24420,N_19849);
nor UO_2606 (O_2606,N_19187,N_24091);
nor UO_2607 (O_2607,N_19946,N_20448);
or UO_2608 (O_2608,N_23314,N_21991);
or UO_2609 (O_2609,N_20574,N_22763);
nor UO_2610 (O_2610,N_21887,N_22819);
and UO_2611 (O_2611,N_24937,N_22246);
and UO_2612 (O_2612,N_23326,N_23166);
nor UO_2613 (O_2613,N_23536,N_21449);
xnor UO_2614 (O_2614,N_24097,N_20975);
and UO_2615 (O_2615,N_19835,N_24828);
and UO_2616 (O_2616,N_21127,N_20832);
and UO_2617 (O_2617,N_24753,N_21649);
and UO_2618 (O_2618,N_21967,N_21926);
and UO_2619 (O_2619,N_21503,N_19994);
and UO_2620 (O_2620,N_21052,N_23177);
and UO_2621 (O_2621,N_21249,N_23690);
or UO_2622 (O_2622,N_20168,N_20287);
or UO_2623 (O_2623,N_19761,N_19606);
nor UO_2624 (O_2624,N_20385,N_24196);
xor UO_2625 (O_2625,N_20498,N_22261);
xnor UO_2626 (O_2626,N_21257,N_23495);
xor UO_2627 (O_2627,N_24780,N_20721);
nand UO_2628 (O_2628,N_22034,N_18895);
nand UO_2629 (O_2629,N_24761,N_24787);
xor UO_2630 (O_2630,N_24275,N_23502);
nand UO_2631 (O_2631,N_21095,N_23069);
or UO_2632 (O_2632,N_21046,N_23435);
xnor UO_2633 (O_2633,N_24893,N_22069);
or UO_2634 (O_2634,N_19381,N_22235);
or UO_2635 (O_2635,N_19110,N_19274);
and UO_2636 (O_2636,N_19364,N_23074);
xor UO_2637 (O_2637,N_21245,N_20101);
and UO_2638 (O_2638,N_18879,N_22022);
or UO_2639 (O_2639,N_22955,N_24878);
nor UO_2640 (O_2640,N_23592,N_23306);
and UO_2641 (O_2641,N_20414,N_24069);
or UO_2642 (O_2642,N_22530,N_22527);
and UO_2643 (O_2643,N_21526,N_22182);
and UO_2644 (O_2644,N_22210,N_19976);
nand UO_2645 (O_2645,N_21886,N_20435);
or UO_2646 (O_2646,N_24448,N_24059);
or UO_2647 (O_2647,N_24602,N_18786);
or UO_2648 (O_2648,N_24756,N_21823);
xor UO_2649 (O_2649,N_23555,N_22707);
or UO_2650 (O_2650,N_23442,N_22818);
nor UO_2651 (O_2651,N_20484,N_23811);
nor UO_2652 (O_2652,N_23694,N_19573);
or UO_2653 (O_2653,N_24261,N_23825);
or UO_2654 (O_2654,N_21241,N_23110);
nand UO_2655 (O_2655,N_20715,N_19025);
or UO_2656 (O_2656,N_23676,N_22012);
nor UO_2657 (O_2657,N_21707,N_18930);
and UO_2658 (O_2658,N_21156,N_22383);
and UO_2659 (O_2659,N_22757,N_21621);
nor UO_2660 (O_2660,N_21770,N_23996);
nand UO_2661 (O_2661,N_20152,N_22835);
or UO_2662 (O_2662,N_22272,N_21427);
nand UO_2663 (O_2663,N_24656,N_22260);
nand UO_2664 (O_2664,N_21411,N_20622);
xor UO_2665 (O_2665,N_22429,N_18949);
and UO_2666 (O_2666,N_22005,N_20030);
nand UO_2667 (O_2667,N_23420,N_20927);
xor UO_2668 (O_2668,N_22480,N_19312);
nor UO_2669 (O_2669,N_22789,N_19451);
and UO_2670 (O_2670,N_24174,N_20481);
nor UO_2671 (O_2671,N_24221,N_19464);
nor UO_2672 (O_2672,N_23726,N_21120);
and UO_2673 (O_2673,N_18853,N_22575);
nand UO_2674 (O_2674,N_19784,N_19874);
and UO_2675 (O_2675,N_24375,N_23219);
or UO_2676 (O_2676,N_20765,N_22118);
or UO_2677 (O_2677,N_21807,N_19721);
or UO_2678 (O_2678,N_20612,N_23082);
or UO_2679 (O_2679,N_24785,N_24926);
and UO_2680 (O_2680,N_20668,N_18902);
nor UO_2681 (O_2681,N_23553,N_19776);
and UO_2682 (O_2682,N_24035,N_19801);
or UO_2683 (O_2683,N_24626,N_18878);
or UO_2684 (O_2684,N_20620,N_24391);
nor UO_2685 (O_2685,N_19267,N_21927);
nand UO_2686 (O_2686,N_20787,N_23089);
xnor UO_2687 (O_2687,N_23770,N_19983);
and UO_2688 (O_2688,N_24105,N_19418);
nor UO_2689 (O_2689,N_22792,N_19031);
nor UO_2690 (O_2690,N_19809,N_19535);
nor UO_2691 (O_2691,N_20003,N_24083);
nor UO_2692 (O_2692,N_20544,N_22767);
nand UO_2693 (O_2693,N_21871,N_24172);
and UO_2694 (O_2694,N_19358,N_21998);
nor UO_2695 (O_2695,N_22597,N_22178);
nand UO_2696 (O_2696,N_20623,N_20348);
nand UO_2697 (O_2697,N_23903,N_23444);
nand UO_2698 (O_2698,N_19859,N_20010);
and UO_2699 (O_2699,N_20921,N_19510);
or UO_2700 (O_2700,N_21206,N_23120);
nand UO_2701 (O_2701,N_24117,N_19398);
nand UO_2702 (O_2702,N_19985,N_21892);
nor UO_2703 (O_2703,N_21763,N_22068);
or UO_2704 (O_2704,N_23973,N_21310);
nand UO_2705 (O_2705,N_22728,N_22809);
or UO_2706 (O_2706,N_19568,N_22753);
nand UO_2707 (O_2707,N_19867,N_23719);
nor UO_2708 (O_2708,N_19345,N_22854);
or UO_2709 (O_2709,N_20160,N_22475);
and UO_2710 (O_2710,N_21947,N_19347);
nand UO_2711 (O_2711,N_23568,N_20002);
nand UO_2712 (O_2712,N_21018,N_21048);
nand UO_2713 (O_2713,N_22408,N_21002);
nand UO_2714 (O_2714,N_18845,N_24627);
or UO_2715 (O_2715,N_24218,N_23389);
and UO_2716 (O_2716,N_20531,N_24993);
nand UO_2717 (O_2717,N_22203,N_21134);
or UO_2718 (O_2718,N_20644,N_24723);
or UO_2719 (O_2719,N_24204,N_21686);
or UO_2720 (O_2720,N_20786,N_21518);
or UO_2721 (O_2721,N_22627,N_21897);
or UO_2722 (O_2722,N_22886,N_21263);
nor UO_2723 (O_2723,N_20164,N_20666);
or UO_2724 (O_2724,N_18960,N_21225);
xnor UO_2725 (O_2725,N_21556,N_24995);
and UO_2726 (O_2726,N_24304,N_21868);
xnor UO_2727 (O_2727,N_20852,N_23099);
nor UO_2728 (O_2728,N_22473,N_20185);
nor UO_2729 (O_2729,N_24528,N_20888);
nand UO_2730 (O_2730,N_24197,N_19457);
nor UO_2731 (O_2731,N_24861,N_22400);
nor UO_2732 (O_2732,N_20426,N_24468);
and UO_2733 (O_2733,N_23338,N_19468);
or UO_2734 (O_2734,N_20829,N_23256);
nor UO_2735 (O_2735,N_19352,N_22059);
nor UO_2736 (O_2736,N_24152,N_19222);
or UO_2737 (O_2737,N_24879,N_20084);
xor UO_2738 (O_2738,N_21531,N_19526);
nand UO_2739 (O_2739,N_21213,N_19617);
and UO_2740 (O_2740,N_18806,N_22324);
nand UO_2741 (O_2741,N_23094,N_21758);
nor UO_2742 (O_2742,N_19581,N_23079);
nor UO_2743 (O_2743,N_23942,N_22158);
nand UO_2744 (O_2744,N_21678,N_20634);
nor UO_2745 (O_2745,N_21450,N_19430);
nand UO_2746 (O_2746,N_22057,N_22167);
and UO_2747 (O_2747,N_23780,N_22222);
nor UO_2748 (O_2748,N_19004,N_23031);
and UO_2749 (O_2749,N_20705,N_24525);
nand UO_2750 (O_2750,N_24855,N_22014);
or UO_2751 (O_2751,N_21288,N_21855);
and UO_2752 (O_2752,N_22986,N_21440);
nand UO_2753 (O_2753,N_23432,N_20064);
nor UO_2754 (O_2754,N_24948,N_24330);
nand UO_2755 (O_2755,N_20732,N_24270);
nor UO_2756 (O_2756,N_23938,N_21845);
xor UO_2757 (O_2757,N_22248,N_20227);
or UO_2758 (O_2758,N_21802,N_24503);
or UO_2759 (O_2759,N_18831,N_23929);
and UO_2760 (O_2760,N_21364,N_19746);
nand UO_2761 (O_2761,N_20125,N_24548);
and UO_2762 (O_2762,N_20894,N_19718);
nand UO_2763 (O_2763,N_24630,N_21050);
nor UO_2764 (O_2764,N_19679,N_20388);
and UO_2765 (O_2765,N_23316,N_19668);
or UO_2766 (O_2766,N_20335,N_20914);
or UO_2767 (O_2767,N_22524,N_23494);
or UO_2768 (O_2768,N_24824,N_23614);
and UO_2769 (O_2769,N_19169,N_24135);
nand UO_2770 (O_2770,N_19208,N_24042);
nand UO_2771 (O_2771,N_21573,N_21687);
and UO_2772 (O_2772,N_20425,N_23756);
xnor UO_2773 (O_2773,N_20194,N_20566);
or UO_2774 (O_2774,N_23871,N_22380);
nor UO_2775 (O_2775,N_24660,N_20597);
xor UO_2776 (O_2776,N_24918,N_18757);
nand UO_2777 (O_2777,N_19293,N_22114);
nand UO_2778 (O_2778,N_21602,N_24363);
or UO_2779 (O_2779,N_23504,N_20751);
and UO_2780 (O_2780,N_19697,N_18802);
nor UO_2781 (O_2781,N_24631,N_22929);
nor UO_2782 (O_2782,N_19940,N_24048);
or UO_2783 (O_2783,N_22867,N_24990);
nor UO_2784 (O_2784,N_21463,N_22039);
nand UO_2785 (O_2785,N_19305,N_22453);
or UO_2786 (O_2786,N_21376,N_23209);
xnor UO_2787 (O_2787,N_22581,N_20013);
and UO_2788 (O_2788,N_24279,N_18843);
and UO_2789 (O_2789,N_20090,N_20219);
nand UO_2790 (O_2790,N_21076,N_24129);
or UO_2791 (O_2791,N_22181,N_19667);
nor UO_2792 (O_2792,N_22285,N_22599);
or UO_2793 (O_2793,N_21757,N_23662);
xor UO_2794 (O_2794,N_23207,N_21455);
or UO_2795 (O_2795,N_23333,N_23706);
nor UO_2796 (O_2796,N_21767,N_22773);
nor UO_2797 (O_2797,N_23084,N_18931);
or UO_2798 (O_2798,N_21848,N_22253);
nor UO_2799 (O_2799,N_20023,N_19003);
nand UO_2800 (O_2800,N_19330,N_18822);
nor UO_2801 (O_2801,N_21030,N_22908);
and UO_2802 (O_2802,N_20915,N_21905);
or UO_2803 (O_2803,N_24954,N_24103);
and UO_2804 (O_2804,N_23058,N_24460);
or UO_2805 (O_2805,N_22281,N_21618);
or UO_2806 (O_2806,N_24957,N_19152);
nand UO_2807 (O_2807,N_23221,N_22635);
nand UO_2808 (O_2808,N_19070,N_19178);
or UO_2809 (O_2809,N_19543,N_22545);
and UO_2810 (O_2810,N_21940,N_20464);
or UO_2811 (O_2811,N_22427,N_20299);
nor UO_2812 (O_2812,N_22967,N_22516);
or UO_2813 (O_2813,N_20545,N_22500);
nand UO_2814 (O_2814,N_21309,N_19203);
nand UO_2815 (O_2815,N_21060,N_20657);
or UO_2816 (O_2816,N_21528,N_22356);
nor UO_2817 (O_2817,N_24529,N_22737);
nor UO_2818 (O_2818,N_20319,N_21285);
or UO_2819 (O_2819,N_20995,N_22136);
nand UO_2820 (O_2820,N_23285,N_19707);
nand UO_2821 (O_2821,N_20851,N_19903);
nor UO_2822 (O_2822,N_22299,N_23605);
or UO_2823 (O_2823,N_23496,N_24522);
nor UO_2824 (O_2824,N_22289,N_19416);
nand UO_2825 (O_2825,N_21322,N_19616);
or UO_2826 (O_2826,N_20518,N_19530);
or UO_2827 (O_2827,N_20204,N_19101);
nand UO_2828 (O_2828,N_20523,N_24963);
or UO_2829 (O_2829,N_23247,N_19046);
nand UO_2830 (O_2830,N_23040,N_20831);
or UO_2831 (O_2831,N_21496,N_23395);
nand UO_2832 (O_2832,N_20552,N_22915);
or UO_2833 (O_2833,N_23513,N_20578);
or UO_2834 (O_2834,N_20782,N_24060);
nand UO_2835 (O_2835,N_20867,N_19068);
or UO_2836 (O_2836,N_21761,N_24158);
nand UO_2837 (O_2837,N_23708,N_22144);
nand UO_2838 (O_2838,N_23535,N_23299);
xor UO_2839 (O_2839,N_22073,N_23519);
and UO_2840 (O_2840,N_23037,N_20039);
nor UO_2841 (O_2841,N_20188,N_23062);
and UO_2842 (O_2842,N_23835,N_22013);
or UO_2843 (O_2843,N_21804,N_18906);
nor UO_2844 (O_2844,N_22348,N_23773);
and UO_2845 (O_2845,N_22431,N_21294);
and UO_2846 (O_2846,N_24921,N_24067);
nand UO_2847 (O_2847,N_18905,N_23783);
nor UO_2848 (O_2848,N_24480,N_19560);
xnor UO_2849 (O_2849,N_24737,N_20489);
nand UO_2850 (O_2850,N_23935,N_24045);
nand UO_2851 (O_2851,N_18874,N_24255);
nor UO_2852 (O_2852,N_23275,N_20990);
and UO_2853 (O_2853,N_24146,N_20040);
and UO_2854 (O_2854,N_19283,N_23650);
or UO_2855 (O_2855,N_22902,N_20379);
nand UO_2856 (O_2856,N_20745,N_24038);
nor UO_2857 (O_2857,N_23225,N_21593);
nand UO_2858 (O_2858,N_23101,N_24251);
or UO_2859 (O_2859,N_22770,N_23142);
nor UO_2860 (O_2860,N_22946,N_19763);
nor UO_2861 (O_2861,N_24088,N_24809);
nand UO_2862 (O_2862,N_21822,N_24708);
or UO_2863 (O_2863,N_21925,N_24639);
and UO_2864 (O_2864,N_22688,N_20823);
nand UO_2865 (O_2865,N_18892,N_22138);
nor UO_2866 (O_2866,N_21996,N_21296);
or UO_2867 (O_2867,N_20891,N_22031);
nor UO_2868 (O_2868,N_21877,N_21477);
nor UO_2869 (O_2869,N_21497,N_22087);
nand UO_2870 (O_2870,N_24094,N_21753);
or UO_2871 (O_2871,N_21722,N_21238);
nor UO_2872 (O_2872,N_24070,N_20695);
nor UO_2873 (O_2873,N_22525,N_21065);
nor UO_2874 (O_2874,N_21594,N_23388);
nor UO_2875 (O_2875,N_21100,N_19791);
nand UO_2876 (O_2876,N_22477,N_19377);
and UO_2877 (O_2877,N_22082,N_19322);
or UO_2878 (O_2878,N_23387,N_22190);
nand UO_2879 (O_2879,N_19516,N_23044);
or UO_2880 (O_2880,N_24814,N_20139);
or UO_2881 (O_2881,N_19253,N_23102);
nand UO_2882 (O_2882,N_20199,N_21854);
and UO_2883 (O_2883,N_19965,N_20625);
nor UO_2884 (O_2884,N_22025,N_18979);
xor UO_2885 (O_2885,N_20790,N_19729);
xor UO_2886 (O_2886,N_21874,N_23715);
nor UO_2887 (O_2887,N_22649,N_23431);
nand UO_2888 (O_2888,N_21295,N_21790);
nor UO_2889 (O_2889,N_19402,N_21118);
and UO_2890 (O_2890,N_23913,N_21984);
and UO_2891 (O_2891,N_23651,N_21385);
or UO_2892 (O_2892,N_19619,N_20134);
and UO_2893 (O_2893,N_24120,N_20763);
xnor UO_2894 (O_2894,N_21226,N_23090);
or UO_2895 (O_2895,N_19129,N_21199);
and UO_2896 (O_2896,N_19071,N_23220);
xor UO_2897 (O_2897,N_20717,N_20080);
nand UO_2898 (O_2898,N_23354,N_19919);
and UO_2899 (O_2899,N_19026,N_24498);
nor UO_2900 (O_2900,N_23317,N_20941);
xnor UO_2901 (O_2901,N_22673,N_23265);
nor UO_2902 (O_2902,N_21841,N_23843);
nor UO_2903 (O_2903,N_23635,N_24696);
and UO_2904 (O_2904,N_21478,N_19706);
nor UO_2905 (O_2905,N_22339,N_19417);
nor UO_2906 (O_2906,N_20977,N_23049);
nand UO_2907 (O_2907,N_22733,N_20167);
and UO_2908 (O_2908,N_20304,N_19885);
nand UO_2909 (O_2909,N_21671,N_23173);
and UO_2910 (O_2910,N_20633,N_19519);
or UO_2911 (O_2911,N_24080,N_23736);
nand UO_2912 (O_2912,N_24305,N_20145);
and UO_2913 (O_2913,N_23965,N_24131);
nand UO_2914 (O_2914,N_22402,N_20434);
or UO_2915 (O_2915,N_20698,N_23934);
nor UO_2916 (O_2916,N_22622,N_24834);
and UO_2917 (O_2917,N_24237,N_22521);
nand UO_2918 (O_2918,N_20771,N_20285);
and UO_2919 (O_2919,N_20795,N_24650);
or UO_2920 (O_2920,N_20844,N_19242);
or UO_2921 (O_2921,N_24714,N_22896);
nor UO_2922 (O_2922,N_24899,N_18837);
and UO_2923 (O_2923,N_19369,N_24257);
and UO_2924 (O_2924,N_20017,N_19188);
nand UO_2925 (O_2925,N_24455,N_20200);
and UO_2926 (O_2926,N_22960,N_20575);
nand UO_2927 (O_2927,N_20678,N_20332);
nand UO_2928 (O_2928,N_20573,N_24717);
nand UO_2929 (O_2929,N_19546,N_21331);
nand UO_2930 (O_2930,N_19916,N_23407);
nand UO_2931 (O_2931,N_23731,N_20958);
and UO_2932 (O_2932,N_22363,N_19403);
or UO_2933 (O_2933,N_22873,N_20554);
or UO_2934 (O_2934,N_23657,N_19243);
nor UO_2935 (O_2935,N_20400,N_24858);
or UO_2936 (O_2936,N_21904,N_22369);
and UO_2937 (O_2937,N_22259,N_24646);
and UO_2938 (O_2938,N_19443,N_24331);
nor UO_2939 (O_2939,N_22360,N_18827);
or UO_2940 (O_2940,N_20004,N_22691);
or UO_2941 (O_2941,N_22115,N_21093);
xnor UO_2942 (O_2942,N_20281,N_20011);
or UO_2943 (O_2943,N_22585,N_20465);
or UO_2944 (O_2944,N_21543,N_20600);
nand UO_2945 (O_2945,N_22980,N_20874);
and UO_2946 (O_2946,N_23415,N_24302);
xor UO_2947 (O_2947,N_23051,N_21151);
and UO_2948 (O_2948,N_22018,N_18946);
or UO_2949 (O_2949,N_22038,N_19587);
nor UO_2950 (O_2950,N_20303,N_19397);
or UO_2951 (O_2951,N_22328,N_22004);
and UO_2952 (O_2952,N_24936,N_18886);
nor UO_2953 (O_2953,N_22065,N_22445);
or UO_2954 (O_2954,N_21332,N_20775);
xor UO_2955 (O_2955,N_23917,N_22913);
nand UO_2956 (O_2956,N_22779,N_21869);
or UO_2957 (O_2957,N_24133,N_23892);
or UO_2958 (O_2958,N_21145,N_24369);
and UO_2959 (O_2959,N_24416,N_24576);
nand UO_2960 (O_2960,N_24435,N_22179);
nand UO_2961 (O_2961,N_22765,N_18945);
and UO_2962 (O_2962,N_24875,N_23856);
and UO_2963 (O_2963,N_23470,N_21324);
xor UO_2964 (O_2964,N_23661,N_22702);
or UO_2965 (O_2965,N_22623,N_22404);
and UO_2966 (O_2966,N_21755,N_23730);
nand UO_2967 (O_2967,N_24142,N_23224);
or UO_2968 (O_2968,N_24249,N_20536);
or UO_2969 (O_2969,N_24027,N_21003);
and UO_2970 (O_2970,N_21183,N_24832);
nand UO_2971 (O_2971,N_19714,N_24041);
nand UO_2972 (O_2972,N_19918,N_23063);
nand UO_2973 (O_2973,N_24506,N_20386);
nand UO_2974 (O_2974,N_23620,N_22176);
xnor UO_2975 (O_2975,N_22805,N_23353);
or UO_2976 (O_2976,N_23401,N_22301);
and UO_2977 (O_2977,N_19238,N_19948);
nand UO_2978 (O_2978,N_20105,N_20401);
nand UO_2979 (O_2979,N_24546,N_21711);
and UO_2980 (O_2980,N_23912,N_24493);
nand UO_2981 (O_2981,N_21635,N_21394);
nor UO_2982 (O_2982,N_21105,N_18974);
nor UO_2983 (O_2983,N_19875,N_22119);
nand UO_2984 (O_2984,N_22823,N_24606);
xnor UO_2985 (O_2985,N_24352,N_20539);
nand UO_2986 (O_2986,N_20513,N_24114);
nor UO_2987 (O_2987,N_19832,N_19308);
or UO_2988 (O_2988,N_19452,N_21891);
or UO_2989 (O_2989,N_18950,N_19599);
nor UO_2990 (O_2990,N_23374,N_22650);
nor UO_2991 (O_2991,N_22173,N_21522);
nand UO_2992 (O_2992,N_20916,N_23226);
nand UO_2993 (O_2993,N_20664,N_24354);
and UO_2994 (O_2994,N_24746,N_20946);
nand UO_2995 (O_2995,N_21563,N_23748);
xor UO_2996 (O_2996,N_24738,N_19872);
xor UO_2997 (O_2997,N_23319,N_24064);
nand UO_2998 (O_2998,N_19204,N_24092);
nand UO_2999 (O_2999,N_20351,N_22912);
endmodule