module basic_2500_25000_3000_125_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_406,In_367);
and U1 (N_1,In_2037,In_1595);
and U2 (N_2,In_1908,In_1689);
xor U3 (N_3,In_1928,In_1020);
nand U4 (N_4,In_568,In_1023);
xnor U5 (N_5,In_602,In_2093);
xor U6 (N_6,In_2395,In_2276);
xnor U7 (N_7,In_975,In_1057);
or U8 (N_8,In_1321,In_1053);
nand U9 (N_9,In_1825,In_299);
xor U10 (N_10,In_424,In_1490);
nand U11 (N_11,In_692,In_623);
or U12 (N_12,In_1289,In_1594);
nand U13 (N_13,In_805,In_1921);
and U14 (N_14,In_1076,In_415);
nor U15 (N_15,In_2024,In_183);
and U16 (N_16,In_1345,In_227);
or U17 (N_17,In_455,In_1543);
or U18 (N_18,In_2006,In_437);
xor U19 (N_19,In_2417,In_386);
and U20 (N_20,In_308,In_1501);
xor U21 (N_21,In_1841,In_265);
xnor U22 (N_22,In_201,In_991);
or U23 (N_23,In_1522,In_1961);
and U24 (N_24,In_1215,In_440);
nand U25 (N_25,In_1523,In_2200);
or U26 (N_26,In_941,In_1044);
nor U27 (N_27,In_448,In_1453);
or U28 (N_28,In_1232,In_1794);
and U29 (N_29,In_1141,In_951);
or U30 (N_30,In_1480,In_510);
xor U31 (N_31,In_1484,In_376);
xor U32 (N_32,In_1727,In_1989);
or U33 (N_33,In_1335,In_1265);
nand U34 (N_34,In_798,In_835);
or U35 (N_35,In_1920,In_1884);
and U36 (N_36,In_2092,In_952);
xor U37 (N_37,In_253,In_1801);
or U38 (N_38,In_1770,In_400);
xnor U39 (N_39,In_1082,In_1974);
and U40 (N_40,In_163,In_1912);
or U41 (N_41,In_2321,In_1202);
xnor U42 (N_42,In_2369,In_1676);
xor U43 (N_43,In_1304,In_8);
nand U44 (N_44,In_1336,In_272);
xor U45 (N_45,In_1608,In_1041);
nand U46 (N_46,In_1814,In_1326);
and U47 (N_47,In_2077,In_1476);
xor U48 (N_48,In_2271,In_2224);
xor U49 (N_49,In_1133,In_298);
and U50 (N_50,In_467,In_2013);
nor U51 (N_51,In_138,In_1264);
xor U52 (N_52,In_2349,In_329);
nor U53 (N_53,In_210,In_1173);
or U54 (N_54,In_1433,In_1253);
or U55 (N_55,In_2203,In_615);
xor U56 (N_56,In_1504,In_2394);
or U57 (N_57,In_2236,In_1271);
nand U58 (N_58,In_2097,In_1220);
or U59 (N_59,In_1903,In_1547);
nand U60 (N_60,In_1427,In_1391);
or U61 (N_61,In_870,In_93);
xnor U62 (N_62,In_1243,In_2357);
nor U63 (N_63,In_208,In_1168);
nand U64 (N_64,In_2217,In_2142);
or U65 (N_65,In_2251,In_1347);
nand U66 (N_66,In_238,In_1670);
nand U67 (N_67,In_747,In_620);
and U68 (N_68,In_355,In_101);
nor U69 (N_69,In_1724,In_1333);
xor U70 (N_70,In_674,In_1744);
xnor U71 (N_71,In_2385,In_2477);
xor U72 (N_72,In_1373,In_645);
nand U73 (N_73,In_1281,In_800);
nor U74 (N_74,In_31,In_1119);
nor U75 (N_75,In_689,In_2173);
and U76 (N_76,In_1174,In_2331);
and U77 (N_77,In_2207,In_590);
xor U78 (N_78,In_1367,In_342);
nor U79 (N_79,In_671,In_2310);
or U80 (N_80,In_1455,In_1148);
and U81 (N_81,In_855,In_338);
or U82 (N_82,In_892,In_1306);
nand U83 (N_83,In_1312,In_2322);
nor U84 (N_84,In_2040,In_2038);
or U85 (N_85,In_1792,In_324);
or U86 (N_86,In_1610,In_1596);
nand U87 (N_87,In_2350,In_742);
and U88 (N_88,In_213,In_2463);
or U89 (N_89,In_408,In_488);
xnor U90 (N_90,In_1995,In_769);
nand U91 (N_91,In_1823,In_2247);
or U92 (N_92,In_1551,In_2253);
or U93 (N_93,In_2447,In_1240);
nand U94 (N_94,In_2201,In_2407);
nand U95 (N_95,In_612,In_1688);
and U96 (N_96,In_362,In_548);
nand U97 (N_97,In_1812,In_200);
nand U98 (N_98,In_2191,In_1877);
or U99 (N_99,In_118,In_115);
or U100 (N_100,In_429,In_2289);
and U101 (N_101,In_1886,In_1049);
xor U102 (N_102,In_417,In_1357);
xnor U103 (N_103,In_1355,In_2343);
nor U104 (N_104,In_1157,In_1497);
nor U105 (N_105,In_2177,In_579);
nor U106 (N_106,In_767,In_1130);
xnor U107 (N_107,In_2287,In_1579);
nand U108 (N_108,In_1129,In_533);
xor U109 (N_109,In_1552,In_746);
and U110 (N_110,In_1692,In_149);
nor U111 (N_111,In_750,In_2220);
nand U112 (N_112,In_1668,In_1019);
nor U113 (N_113,In_2157,In_947);
and U114 (N_114,In_1601,In_2258);
or U115 (N_115,In_789,In_2244);
and U116 (N_116,In_913,In_2401);
xor U117 (N_117,In_249,In_148);
or U118 (N_118,In_1245,In_294);
or U119 (N_119,In_1517,In_1590);
nand U120 (N_120,In_2223,In_157);
xor U121 (N_121,In_136,In_1636);
xor U122 (N_122,In_1534,In_682);
nor U123 (N_123,In_1258,In_1774);
or U124 (N_124,In_825,In_923);
nor U125 (N_125,In_1027,In_259);
or U126 (N_126,In_496,In_1796);
or U127 (N_127,In_1766,In_1259);
nor U128 (N_128,In_1307,In_1840);
nor U129 (N_129,In_1645,In_2004);
nand U130 (N_130,In_2269,In_1585);
or U131 (N_131,In_445,In_116);
nor U132 (N_132,In_303,In_2458);
or U133 (N_133,In_2105,In_1519);
or U134 (N_134,In_1156,In_1845);
and U135 (N_135,In_292,In_2160);
xnor U136 (N_136,In_1277,In_999);
xor U137 (N_137,In_1984,In_860);
nor U138 (N_138,In_1923,In_59);
and U139 (N_139,In_1772,In_1211);
or U140 (N_140,In_1820,In_2116);
and U141 (N_141,In_402,In_473);
or U142 (N_142,In_844,In_168);
and U143 (N_143,In_2131,In_304);
nand U144 (N_144,In_756,In_1092);
xnor U145 (N_145,In_460,In_2170);
xnor U146 (N_146,In_1212,In_608);
or U147 (N_147,In_1883,In_1328);
nor U148 (N_148,In_1134,In_2490);
nand U149 (N_149,In_1997,In_2029);
nand U150 (N_150,In_160,In_247);
nand U151 (N_151,In_1379,In_628);
and U152 (N_152,In_2189,In_2378);
xor U153 (N_153,In_1646,In_926);
and U154 (N_154,In_1748,In_1278);
xor U155 (N_155,In_2007,In_1482);
or U156 (N_156,In_2423,In_1809);
xnor U157 (N_157,In_314,In_2424);
and U158 (N_158,In_1496,In_783);
nand U159 (N_159,In_1658,In_1566);
and U160 (N_160,In_214,In_942);
and U161 (N_161,In_1214,In_959);
or U162 (N_162,In_372,In_2121);
xor U163 (N_163,In_1233,In_691);
nor U164 (N_164,In_1806,In_2185);
and U165 (N_165,In_757,In_1745);
xnor U166 (N_166,In_2263,In_262);
xnor U167 (N_167,In_1275,In_147);
and U168 (N_168,In_3,In_956);
nand U169 (N_169,In_1998,In_2483);
and U170 (N_170,In_1127,In_1628);
nor U171 (N_171,In_2133,In_1350);
nand U172 (N_172,In_23,In_1016);
nand U173 (N_173,In_483,In_536);
and U174 (N_174,In_2195,In_1085);
nor U175 (N_175,In_1045,In_494);
nand U176 (N_176,In_466,In_1691);
and U177 (N_177,In_2125,In_1565);
or U178 (N_178,In_954,In_2068);
nand U179 (N_179,In_2485,In_2081);
or U180 (N_180,In_1250,In_1337);
nand U181 (N_181,In_1602,In_1634);
nand U182 (N_182,In_618,In_2104);
xnor U183 (N_183,In_2154,In_935);
xor U184 (N_184,In_105,In_1943);
nor U185 (N_185,In_1858,In_532);
nor U186 (N_186,In_420,In_1381);
and U187 (N_187,In_2044,In_2347);
and U188 (N_188,In_2233,In_1666);
xnor U189 (N_189,In_1423,In_98);
nand U190 (N_190,In_733,In_209);
and U191 (N_191,In_199,In_1224);
nand U192 (N_192,In_2080,In_7);
nand U193 (N_193,In_1471,In_477);
xor U194 (N_194,In_1371,In_1680);
nand U195 (N_195,In_1713,In_1581);
nor U196 (N_196,In_1203,In_847);
nor U197 (N_197,In_1752,In_1349);
nand U198 (N_198,In_457,In_1743);
nor U199 (N_199,In_1818,In_1441);
or U200 (N_200,In_573,In_1408);
or U201 (N_201,In_96,In_1936);
xor U202 (N_202,In_228,N_106);
nor U203 (N_203,In_2179,In_2245);
nor U204 (N_204,N_102,In_1401);
and U205 (N_205,In_1873,In_1159);
xnor U206 (N_206,N_34,N_61);
xor U207 (N_207,In_1370,In_1848);
nand U208 (N_208,In_785,In_1467);
xor U209 (N_209,In_1429,In_1880);
or U210 (N_210,In_1425,In_1817);
and U211 (N_211,In_1536,In_864);
nand U212 (N_212,In_965,In_1922);
and U213 (N_213,In_1574,In_1394);
nor U214 (N_214,In_2323,In_560);
or U215 (N_215,In_2032,In_137);
and U216 (N_216,In_597,In_2293);
nand U217 (N_217,N_124,In_604);
and U218 (N_218,In_1040,In_64);
nand U219 (N_219,In_2309,In_1061);
nor U220 (N_220,In_1520,In_1135);
and U221 (N_221,In_2259,In_831);
or U222 (N_222,In_1623,In_1115);
and U223 (N_223,In_1090,In_899);
nand U224 (N_224,In_1538,In_2384);
and U225 (N_225,N_46,In_1126);
or U226 (N_226,In_1696,In_2240);
or U227 (N_227,In_500,In_180);
and U228 (N_228,N_20,N_183);
nand U229 (N_229,In_1446,In_365);
or U230 (N_230,In_47,In_544);
xnor U231 (N_231,In_851,In_1660);
nor U232 (N_232,In_1607,In_1450);
xor U233 (N_233,In_2396,In_866);
xor U234 (N_234,In_2484,In_1799);
xnor U235 (N_235,N_159,In_1144);
nand U236 (N_236,In_2148,In_2085);
or U237 (N_237,In_2438,In_6);
nor U238 (N_238,In_1638,In_1618);
nor U239 (N_239,In_2302,In_1905);
nor U240 (N_240,In_531,In_2413);
nand U241 (N_241,N_131,In_914);
nor U242 (N_242,In_2460,In_1975);
and U243 (N_243,In_1026,In_1614);
or U244 (N_244,In_145,In_2027);
nand U245 (N_245,In_2100,In_121);
and U246 (N_246,In_268,In_79);
or U247 (N_247,In_1364,In_1470);
and U248 (N_248,In_878,In_87);
or U249 (N_249,In_1681,In_1421);
xnor U250 (N_250,In_822,N_83);
nor U251 (N_251,N_25,In_656);
and U252 (N_252,In_1376,In_468);
and U253 (N_253,In_2445,N_139);
nand U254 (N_254,In_2468,In_749);
nand U255 (N_255,In_1031,In_911);
xor U256 (N_256,In_396,In_2156);
or U257 (N_257,In_279,In_1153);
xnor U258 (N_258,In_1560,In_586);
nand U259 (N_259,In_650,In_2014);
nor U260 (N_260,In_1444,In_267);
nor U261 (N_261,In_619,In_252);
xor U262 (N_262,In_1161,In_2313);
nor U263 (N_263,In_2212,In_699);
nor U264 (N_264,N_24,In_1901);
and U265 (N_265,In_728,In_343);
or U266 (N_266,In_2046,In_1591);
nand U267 (N_267,In_1842,In_1879);
nor U268 (N_268,In_1385,In_921);
nand U269 (N_269,In_436,In_196);
or U270 (N_270,In_1828,In_2346);
or U271 (N_271,In_658,In_546);
nor U272 (N_272,In_2147,In_1657);
and U273 (N_273,In_469,In_1514);
nor U274 (N_274,In_673,In_1548);
nand U275 (N_275,In_1358,In_1051);
nor U276 (N_276,In_1247,In_2480);
or U277 (N_277,In_1545,In_1354);
nor U278 (N_278,In_2172,In_1248);
nor U279 (N_279,In_861,In_2344);
xor U280 (N_280,In_2058,In_1164);
nor U281 (N_281,In_1081,In_647);
or U282 (N_282,In_1736,In_944);
xor U283 (N_283,In_1193,In_1919);
xnor U284 (N_284,In_1485,In_1725);
nor U285 (N_285,In_2214,In_817);
nor U286 (N_286,In_2098,In_1804);
xnor U287 (N_287,In_380,In_690);
xnor U288 (N_288,In_1341,N_191);
nor U289 (N_289,In_1251,In_694);
nand U290 (N_290,In_2108,In_2138);
nor U291 (N_291,In_1437,N_88);
xnor U292 (N_292,In_837,In_1682);
or U293 (N_293,In_111,In_1178);
and U294 (N_294,In_1481,In_434);
xnor U295 (N_295,In_2272,In_1937);
xor U296 (N_296,In_1434,In_462);
nand U297 (N_297,In_2486,In_1968);
nand U298 (N_298,In_334,N_123);
or U299 (N_299,In_1299,In_1656);
nand U300 (N_300,In_2327,N_122);
nand U301 (N_301,In_754,In_2150);
nand U302 (N_302,In_748,In_2473);
nand U303 (N_303,In_519,In_610);
and U304 (N_304,In_676,In_2248);
or U305 (N_305,In_670,In_1900);
nand U306 (N_306,In_727,In_2487);
nor U307 (N_307,In_2096,In_2197);
nand U308 (N_308,In_2283,In_2443);
nand U309 (N_309,In_522,In_29);
xor U310 (N_310,In_2059,In_637);
xor U311 (N_311,N_172,In_2194);
or U312 (N_312,In_912,In_1847);
nand U313 (N_313,In_1719,In_2119);
nor U314 (N_314,In_1555,In_1965);
nor U315 (N_315,In_1196,In_1489);
and U316 (N_316,In_1037,In_2074);
xnor U317 (N_317,In_1521,In_212);
nand U318 (N_318,In_2159,In_592);
or U319 (N_319,In_1301,In_2270);
and U320 (N_320,In_2433,In_1);
or U321 (N_321,In_146,In_2362);
nand U322 (N_322,In_1783,In_1462);
nand U323 (N_323,In_1582,In_2392);
and U324 (N_324,N_115,In_1535);
nor U325 (N_325,In_113,In_1073);
or U326 (N_326,In_1673,In_1571);
and U327 (N_327,In_398,In_1208);
or U328 (N_328,N_150,In_900);
and U329 (N_329,In_17,In_174);
or U330 (N_330,In_2405,N_22);
nor U331 (N_331,In_505,In_194);
nand U332 (N_332,In_281,N_2);
or U333 (N_333,In_1065,In_1241);
or U334 (N_334,In_349,N_44);
xor U335 (N_335,In_1351,In_1558);
or U336 (N_336,In_1518,In_517);
nand U337 (N_337,In_154,In_1916);
and U338 (N_338,In_1276,In_2135);
xor U339 (N_339,In_1762,In_166);
nand U340 (N_340,In_968,In_1765);
xnor U341 (N_341,In_84,In_839);
or U342 (N_342,In_2400,In_405);
xnor U343 (N_343,N_182,In_1641);
xor U344 (N_344,In_840,In_401);
nor U345 (N_345,In_2499,In_2232);
xnor U346 (N_346,In_295,In_1853);
and U347 (N_347,In_1225,In_1851);
nor U348 (N_348,N_3,In_1332);
and U349 (N_349,In_609,In_1894);
xor U350 (N_350,In_1620,In_1459);
and U351 (N_351,In_1457,In_565);
nor U352 (N_352,In_2446,In_1181);
nand U353 (N_353,In_1859,In_915);
xnor U354 (N_354,In_274,In_239);
or U355 (N_355,In_2123,In_882);
and U356 (N_356,In_305,In_129);
or U357 (N_357,In_431,In_1392);
nand U358 (N_358,In_2419,In_1661);
nor U359 (N_359,N_187,In_2469);
nand U360 (N_360,In_234,In_972);
nand U361 (N_361,In_1343,In_744);
nor U362 (N_362,In_929,In_1701);
and U363 (N_363,In_648,In_739);
xnor U364 (N_364,In_566,In_563);
or U365 (N_365,In_2261,In_2102);
nor U366 (N_366,In_495,In_235);
nand U367 (N_367,In_1864,In_2192);
or U368 (N_368,In_2190,N_52);
nand U369 (N_369,In_731,In_677);
nor U370 (N_370,In_503,N_110);
and U371 (N_371,N_32,In_617);
and U372 (N_372,In_1107,In_82);
nor U373 (N_373,In_1896,In_2282);
xor U374 (N_374,In_306,In_2143);
nor U375 (N_375,In_382,In_1800);
or U376 (N_376,In_179,In_1010);
nand U377 (N_377,In_2360,In_634);
and U378 (N_378,In_766,In_762);
and U379 (N_379,In_30,In_649);
xor U380 (N_380,In_1169,In_1707);
nor U381 (N_381,In_28,In_1039);
or U382 (N_382,In_99,In_557);
nand U383 (N_383,In_1263,In_778);
nor U384 (N_384,In_1469,In_1669);
and U385 (N_385,In_1430,In_397);
xnor U386 (N_386,In_1929,In_358);
xor U387 (N_387,In_2218,In_203);
nor U388 (N_388,In_1223,In_893);
nand U389 (N_389,In_1749,In_479);
nand U390 (N_390,In_1603,In_1091);
and U391 (N_391,In_1907,In_311);
or U392 (N_392,In_1147,N_79);
or U393 (N_393,In_1780,In_143);
and U394 (N_394,N_177,In_264);
or U395 (N_395,In_662,In_471);
nand U396 (N_396,In_94,In_2471);
and U397 (N_397,In_384,In_763);
xor U398 (N_398,In_871,In_1317);
xnor U399 (N_399,In_13,In_1340);
nand U400 (N_400,In_1007,In_1992);
or U401 (N_401,N_223,In_1528);
and U402 (N_402,In_188,In_796);
nor U403 (N_403,In_895,In_632);
nor U404 (N_404,In_625,In_297);
and U405 (N_405,N_290,In_1781);
xnor U406 (N_406,In_2110,In_1994);
nor U407 (N_407,N_75,In_344);
nor U408 (N_408,In_127,In_2015);
nand U409 (N_409,In_2091,In_758);
and U410 (N_410,In_95,N_313);
and U411 (N_411,In_791,In_1311);
xnor U412 (N_412,In_2083,In_1750);
and U413 (N_413,N_286,In_2380);
nand U414 (N_414,In_856,In_2453);
nand U415 (N_415,In_1515,In_883);
xor U416 (N_416,In_370,In_884);
xnor U417 (N_417,In_1218,In_1319);
or U418 (N_418,In_640,In_26);
xor U419 (N_419,In_572,In_1687);
or U420 (N_420,N_351,In_1431);
xnor U421 (N_421,In_1128,In_2146);
nand U422 (N_422,N_189,In_1925);
nand U423 (N_423,In_356,In_11);
xnor U424 (N_424,In_540,In_1786);
or U425 (N_425,In_515,In_1881);
or U426 (N_426,In_482,In_506);
xor U427 (N_427,In_687,N_15);
or U428 (N_428,In_225,In_1527);
and U429 (N_429,In_554,In_2178);
nand U430 (N_430,In_360,N_12);
xnor U431 (N_431,In_348,In_939);
nand U432 (N_432,In_641,In_804);
nor U433 (N_433,In_1006,In_881);
or U434 (N_434,In_359,In_24);
nand U435 (N_435,In_435,In_1499);
nand U436 (N_436,In_106,In_1948);
xnor U437 (N_437,In_953,In_1834);
nor U438 (N_438,In_997,N_277);
xor U439 (N_439,In_669,In_2155);
and U440 (N_440,In_2489,In_2051);
nor U441 (N_441,In_1438,In_1717);
nor U442 (N_442,In_1142,In_1298);
nand U443 (N_443,In_1755,In_323);
and U444 (N_444,In_1475,N_30);
nor U445 (N_445,In_221,In_2418);
nand U446 (N_446,In_1541,In_220);
nor U447 (N_447,In_1398,In_1187);
or U448 (N_448,In_896,In_254);
or U449 (N_449,In_924,In_1146);
xnor U450 (N_450,In_1911,In_100);
nor U451 (N_451,In_1509,N_54);
nor U452 (N_452,In_2226,In_78);
xnor U453 (N_453,N_43,In_1000);
xor U454 (N_454,In_869,In_1025);
or U455 (N_455,In_1505,In_131);
xnor U456 (N_456,In_2328,In_374);
and U457 (N_457,In_34,In_2333);
xnor U458 (N_458,In_1200,In_2237);
and U459 (N_459,In_978,In_1860);
and U460 (N_460,In_1447,In_452);
or U461 (N_461,In_1097,In_229);
and U462 (N_462,In_1028,N_84);
and U463 (N_463,In_1891,In_846);
or U464 (N_464,In_389,N_236);
xnor U465 (N_465,N_100,In_917);
nand U466 (N_466,In_1926,In_1604);
and U467 (N_467,N_168,In_1863);
nor U468 (N_468,In_222,N_314);
and U469 (N_469,In_2129,In_409);
and U470 (N_470,N_388,In_2491);
or U471 (N_471,In_1316,In_1758);
or U472 (N_472,In_523,In_10);
and U473 (N_473,N_254,In_1454);
or U474 (N_474,In_40,In_2087);
nand U475 (N_475,In_2334,In_1913);
xor U476 (N_476,In_2295,N_85);
nand U477 (N_477,N_310,In_508);
or U478 (N_478,In_824,In_2026);
and U479 (N_479,In_2340,In_339);
xor U480 (N_480,In_1979,In_1064);
nand U481 (N_481,In_1383,In_2338);
nor U482 (N_482,In_2117,In_1290);
nor U483 (N_483,In_1314,In_1906);
xnor U484 (N_484,In_2383,In_829);
nand U485 (N_485,In_446,In_2285);
and U486 (N_486,In_575,In_1616);
nand U487 (N_487,In_567,In_2249);
or U488 (N_488,In_1393,In_1372);
xnor U489 (N_489,In_948,In_2025);
nand U490 (N_490,N_72,In_1177);
or U491 (N_491,In_696,In_1567);
xor U492 (N_492,In_1932,In_1325);
xnor U493 (N_493,In_1180,In_1753);
nand U494 (N_494,In_1568,In_335);
nand U495 (N_495,In_528,N_339);
xnor U496 (N_496,In_794,In_995);
nand U497 (N_497,N_170,In_2366);
xnor U498 (N_498,In_2075,N_318);
nor U499 (N_499,N_69,In_1071);
xnor U500 (N_500,In_1172,In_458);
xnor U501 (N_501,In_2149,N_142);
and U502 (N_502,In_1990,In_1983);
and U503 (N_503,N_128,In_53);
nand U504 (N_504,In_2071,In_734);
or U505 (N_505,In_2066,In_81);
or U506 (N_506,In_286,In_256);
or U507 (N_507,In_898,In_1261);
nor U508 (N_508,In_1030,In_2294);
nor U509 (N_509,In_2188,In_18);
or U510 (N_510,In_2472,N_157);
xor U511 (N_511,N_173,In_833);
and U512 (N_512,In_2127,In_1001);
or U513 (N_513,In_1985,In_1272);
or U514 (N_514,In_293,In_1056);
xnor U515 (N_515,In_2470,In_2054);
nor U516 (N_516,In_1043,In_961);
xnor U517 (N_517,In_112,In_1139);
xor U518 (N_518,In_1068,In_49);
xnor U519 (N_519,In_2364,N_376);
xnor U520 (N_520,In_940,In_1422);
nor U521 (N_521,In_653,In_1213);
nand U522 (N_522,In_184,In_189);
or U523 (N_523,In_1106,In_375);
xnor U524 (N_524,In_582,N_112);
xnor U525 (N_525,In_2230,In_529);
and U526 (N_526,In_1771,In_2239);
nor U527 (N_527,In_322,In_863);
or U528 (N_528,N_140,In_2427);
nor U529 (N_529,In_1870,In_1318);
nor U530 (N_530,N_126,In_476);
and U531 (N_531,In_2120,N_95);
xor U532 (N_532,In_161,N_203);
xnor U533 (N_533,In_2440,In_2482);
nor U534 (N_534,In_535,N_185);
nor U535 (N_535,In_2167,In_1805);
or U536 (N_536,In_897,In_1739);
or U537 (N_537,In_2332,In_1715);
nor U538 (N_538,In_1024,In_257);
and U539 (N_539,In_2280,In_712);
nor U540 (N_540,In_426,In_449);
and U541 (N_541,In_242,In_858);
nand U542 (N_542,In_444,In_1009);
nor U543 (N_543,In_2016,In_725);
and U544 (N_544,N_328,In_73);
xor U545 (N_545,N_18,In_1274);
nor U546 (N_546,In_478,In_1052);
nand U547 (N_547,N_393,In_1957);
nor U548 (N_548,In_1787,In_2144);
and U549 (N_549,In_1330,In_520);
nand U550 (N_550,N_307,In_1839);
or U551 (N_551,N_210,In_2023);
and U552 (N_552,In_379,In_605);
and U553 (N_553,In_2497,In_243);
nand U554 (N_554,In_58,In_2165);
nor U555 (N_555,In_2166,In_1120);
and U556 (N_556,In_2426,In_2137);
nor U557 (N_557,N_333,In_215);
nand U558 (N_558,In_1930,N_303);
or U559 (N_559,In_1838,In_1827);
and U560 (N_560,In_2474,In_1188);
xor U561 (N_561,N_358,In_20);
xor U562 (N_562,In_2216,In_760);
and U563 (N_563,In_328,In_14);
nor U564 (N_564,N_230,In_1359);
xor U565 (N_565,In_441,In_1524);
or U566 (N_566,N_385,In_2448);
or U567 (N_567,In_1448,In_787);
or U568 (N_568,In_416,In_68);
xnor U569 (N_569,In_1764,In_1899);
xor U570 (N_570,In_1855,In_1526);
and U571 (N_571,N_217,In_117);
xnor U572 (N_572,N_199,In_1953);
or U573 (N_573,In_967,N_389);
xnor U574 (N_574,In_2266,In_1642);
and U575 (N_575,N_28,In_103);
or U576 (N_576,In_868,N_179);
or U577 (N_577,In_1406,In_1201);
and U578 (N_578,In_1400,In_2021);
and U579 (N_579,In_1735,N_96);
and U580 (N_580,In_809,In_321);
nand U581 (N_581,In_422,In_1111);
or U582 (N_582,In_2461,N_227);
xor U583 (N_583,N_276,N_369);
or U584 (N_584,In_1268,In_1122);
nor U585 (N_585,In_1308,In_631);
nor U586 (N_586,In_1693,In_1378);
or U587 (N_587,N_262,In_2094);
nor U588 (N_588,In_2318,N_343);
or U589 (N_589,N_53,In_353);
or U590 (N_590,In_2052,In_1344);
xor U591 (N_591,In_80,N_38);
nand U592 (N_592,In_588,N_163);
and U593 (N_593,N_200,In_1287);
nor U594 (N_594,In_432,In_963);
xnor U595 (N_595,In_427,In_530);
or U596 (N_596,In_48,In_1757);
nand U597 (N_597,In_211,In_1158);
or U598 (N_598,In_1295,In_1163);
nor U599 (N_599,In_318,In_1366);
xnor U600 (N_600,In_1698,In_1305);
nand U601 (N_601,In_345,N_401);
or U602 (N_602,N_536,In_1665);
xor U603 (N_603,In_1632,In_2213);
xnor U604 (N_604,In_1617,In_1492);
or U605 (N_605,In_1915,N_50);
and U606 (N_606,In_1530,In_2030);
or U607 (N_607,In_1409,In_526);
nand U608 (N_608,In_1708,N_573);
and U609 (N_609,N_279,N_475);
nand U610 (N_610,In_1946,In_1293);
or U611 (N_611,In_507,In_594);
nor U612 (N_612,In_433,N_338);
nor U613 (N_613,In_2288,In_1050);
xor U614 (N_614,In_2444,In_616);
nand U615 (N_615,In_2361,N_370);
nor U616 (N_616,N_585,N_147);
or U617 (N_617,In_1138,N_80);
and U618 (N_618,N_575,In_1835);
and U619 (N_619,In_810,In_1532);
nand U620 (N_620,In_1952,N_478);
or U621 (N_621,In_1626,N_444);
nor U622 (N_622,In_2317,In_170);
and U623 (N_623,In_202,In_819);
xor U624 (N_624,In_1960,In_1410);
xnor U625 (N_625,N_582,N_253);
or U626 (N_626,In_702,In_2454);
or U627 (N_627,In_667,In_186);
xor U628 (N_628,N_348,In_801);
nor U629 (N_629,N_289,In_552);
and U630 (N_630,In_418,In_1746);
nor U631 (N_631,N_509,N_48);
xor U632 (N_632,N_425,In_1513);
xnor U633 (N_633,In_2363,N_13);
or U634 (N_634,In_1546,N_90);
or U635 (N_635,N_579,In_1012);
or U636 (N_636,In_2163,In_976);
and U637 (N_637,In_1950,In_1679);
nand U638 (N_638,N_375,In_395);
or U639 (N_639,In_428,In_2275);
nand U640 (N_640,In_1389,In_493);
xnor U641 (N_641,In_1861,N_341);
or U642 (N_642,N_114,N_249);
or U643 (N_643,In_1569,In_1069);
nor U644 (N_644,In_990,In_1468);
xnor U645 (N_645,In_1964,In_803);
xnor U646 (N_646,N_0,N_564);
xor U647 (N_647,In_1959,In_1931);
nand U648 (N_648,N_429,In_1554);
xor U649 (N_649,In_2033,In_1418);
or U650 (N_650,In_2339,In_1365);
xnor U651 (N_651,N_524,N_474);
nand U652 (N_652,In_1353,In_36);
nand U653 (N_653,N_120,N_515);
or U654 (N_654,N_244,N_404);
or U655 (N_655,In_1487,N_438);
or U656 (N_656,In_175,N_505);
nand U657 (N_657,N_574,In_217);
or U658 (N_658,In_695,In_880);
or U659 (N_659,In_1933,In_2134);
nor U660 (N_660,In_2274,In_1987);
and U661 (N_661,In_2073,In_2151);
and U662 (N_662,In_1769,N_458);
nand U663 (N_663,In_1703,In_1356);
nand U664 (N_664,In_1498,In_1777);
xor U665 (N_665,In_430,In_159);
nor U666 (N_666,In_2377,N_299);
or U667 (N_667,N_591,N_511);
xnor U668 (N_668,In_1865,In_414);
and U669 (N_669,In_755,N_459);
and U670 (N_670,N_415,In_683);
xnor U671 (N_671,In_849,In_2001);
nand U672 (N_672,In_464,In_2231);
nand U673 (N_673,In_621,In_622);
xor U674 (N_674,N_340,In_1390);
xor U675 (N_675,In_688,In_1598);
nand U676 (N_676,In_1015,N_516);
nand U677 (N_677,In_603,In_1678);
and U678 (N_678,In_816,N_426);
or U679 (N_679,In_425,In_1486);
nor U680 (N_680,In_65,In_979);
nor U681 (N_681,In_102,In_1910);
nor U682 (N_682,In_1600,In_957);
nor U683 (N_683,In_1267,In_1150);
and U684 (N_684,In_1352,N_308);
xor U685 (N_685,In_1580,In_1677);
nand U686 (N_686,In_1149,N_327);
xnor U687 (N_687,In_164,In_123);
or U688 (N_688,In_1412,In_1714);
nand U689 (N_689,In_331,In_1256);
xnor U690 (N_690,In_2273,In_1399);
and U691 (N_691,In_2397,In_955);
or U692 (N_692,N_98,N_436);
nand U693 (N_693,In_980,In_974);
nor U694 (N_694,In_1198,In_1951);
and U695 (N_695,N_197,In_659);
and U696 (N_696,In_1226,N_87);
or U697 (N_697,In_1776,In_1732);
nand U698 (N_698,In_1118,In_1072);
or U699 (N_699,N_479,N_285);
nand U700 (N_700,N_402,N_473);
nand U701 (N_701,N_551,In_710);
and U702 (N_702,In_390,In_729);
xor U703 (N_703,In_1194,In_54);
or U704 (N_704,N_468,In_1479);
nor U705 (N_705,In_1374,N_502);
xnor U706 (N_706,In_1592,In_2140);
nor U707 (N_707,In_237,N_467);
nor U708 (N_708,In_9,In_1875);
nor U709 (N_709,In_753,In_2371);
nor U710 (N_710,In_1221,In_2246);
nor U711 (N_711,In_626,In_781);
nand U712 (N_712,N_219,In_52);
and U713 (N_713,In_453,In_2303);
nand U714 (N_714,In_1563,In_2183);
or U715 (N_715,N_165,In_1235);
nand U716 (N_716,In_2415,In_107);
xor U717 (N_717,In_4,N_541);
or U718 (N_718,N_543,N_378);
xor U719 (N_719,In_341,In_2031);
nor U720 (N_720,In_693,In_679);
nor U721 (N_721,In_1712,In_1578);
xnor U722 (N_722,In_1934,In_1671);
nand U723 (N_723,In_521,N_86);
nor U724 (N_724,N_325,In_537);
or U725 (N_725,In_438,N_7);
nor U726 (N_726,In_1627,In_2388);
nand U727 (N_727,In_797,In_2070);
and U728 (N_728,In_1048,N_250);
or U729 (N_729,N_550,In_1420);
and U730 (N_730,In_1464,N_162);
nor U731 (N_731,In_2475,In_413);
and U732 (N_732,N_221,In_182);
and U733 (N_733,N_107,In_1967);
or U734 (N_734,In_2341,N_492);
nand U735 (N_735,N_529,In_1363);
xnor U736 (N_736,In_399,In_1404);
nand U737 (N_737,In_336,In_1597);
nand U738 (N_738,N_55,In_598);
xnor U739 (N_739,N_350,N_160);
nor U740 (N_740,In_288,In_705);
xor U741 (N_741,In_1866,In_2130);
or U742 (N_742,In_141,In_1204);
or U743 (N_743,N_158,In_1407);
xor U744 (N_744,In_836,In_1167);
nand U745 (N_745,In_1767,In_169);
xnor U746 (N_746,In_1763,N_130);
xnor U747 (N_747,In_369,N_368);
xor U748 (N_748,N_70,In_1011);
or U749 (N_749,In_561,In_1508);
nor U750 (N_750,In_1080,In_151);
nor U751 (N_751,N_268,N_334);
or U752 (N_752,In_1183,In_1885);
nor U753 (N_753,In_1525,In_661);
xor U754 (N_754,N_584,In_1005);
xnor U755 (N_755,In_1971,N_228);
nand U756 (N_756,In_827,In_128);
and U757 (N_757,In_300,N_209);
nand U758 (N_758,In_289,In_1195);
or U759 (N_759,In_1871,In_2291);
nand U760 (N_760,N_5,In_1331);
xnor U761 (N_761,In_949,N_534);
or U762 (N_762,In_2022,In_549);
nor U763 (N_763,In_1324,In_1639);
or U764 (N_764,In_366,N_154);
and U765 (N_765,N_11,In_1237);
nand U766 (N_766,N_305,In_119);
nor U767 (N_767,In_463,In_1273);
nor U768 (N_768,In_1876,N_403);
nand U769 (N_769,N_36,In_63);
nor U770 (N_770,In_578,N_384);
nand U771 (N_771,N_141,In_1402);
xor U772 (N_772,In_664,In_2286);
or U773 (N_773,In_2000,N_105);
or U774 (N_774,In_346,N_151);
nor U775 (N_775,In_192,In_1694);
or U776 (N_776,In_2202,In_720);
xor U777 (N_777,N_281,In_732);
xnor U778 (N_778,In_2372,In_2430);
or U779 (N_779,In_1442,N_49);
nor U780 (N_780,In_771,In_2162);
or U781 (N_781,In_984,In_1589);
nor U782 (N_782,N_78,In_392);
or U783 (N_783,In_1192,In_412);
nor U784 (N_784,In_1488,In_1611);
nor U785 (N_785,N_477,N_125);
and U786 (N_786,N_176,In_1386);
and U787 (N_787,In_1491,In_450);
xor U788 (N_788,In_2041,In_1612);
nor U789 (N_789,In_1063,N_344);
nand U790 (N_790,In_2153,N_414);
nand U791 (N_791,N_113,In_1461);
or U792 (N_792,In_2356,In_122);
xor U793 (N_793,In_2076,N_568);
nor U794 (N_794,N_267,In_1436);
nand U795 (N_795,In_2043,In_1996);
nand U796 (N_796,In_2086,In_2242);
or U797 (N_797,In_1836,In_489);
nor U798 (N_798,In_988,In_1593);
and U799 (N_799,In_1108,In_2158);
and U800 (N_800,N_471,In_1785);
and U801 (N_801,In_491,In_1074);
and U802 (N_802,N_243,N_722);
xnor U803 (N_803,N_256,In_652);
or U804 (N_804,N_699,In_75);
xnor U805 (N_805,In_518,In_905);
or U806 (N_806,N_514,In_246);
nor U807 (N_807,In_162,In_90);
and U808 (N_808,In_2399,In_908);
xor U809 (N_809,In_901,In_1613);
xor U810 (N_810,In_2297,In_2432);
and U811 (N_811,N_542,N_647);
xnor U812 (N_812,In_187,N_785);
and U813 (N_813,In_852,In_1229);
nor U814 (N_814,In_994,In_2047);
nor U815 (N_815,In_1889,In_1944);
and U816 (N_816,In_638,N_781);
nand U817 (N_817,In_2008,In_2221);
nor U818 (N_818,In_707,In_263);
nand U819 (N_819,N_657,In_60);
xnor U820 (N_820,N_576,In_42);
and U821 (N_821,N_319,In_171);
nand U822 (N_822,N_238,In_1529);
nand U823 (N_823,N_391,In_660);
nand U824 (N_824,In_1465,In_1182);
or U825 (N_825,In_1186,N_506);
nand U826 (N_826,In_16,N_23);
or U827 (N_827,In_2020,N_605);
nor U828 (N_828,In_812,In_987);
xor U829 (N_829,In_511,N_145);
xnor U830 (N_830,In_1917,In_697);
nand U831 (N_831,In_1104,In_2255);
and U832 (N_832,In_1615,In_1342);
xor U833 (N_833,In_173,In_1854);
xor U834 (N_834,In_574,In_589);
nor U835 (N_835,In_153,N_347);
and U836 (N_836,In_2099,N_651);
and U837 (N_837,In_651,N_192);
nor U838 (N_838,N_604,In_543);
nand U839 (N_839,In_2113,In_633);
nand U840 (N_840,N_193,In_1209);
and U841 (N_841,In_1811,In_2456);
and U842 (N_842,In_1405,N_696);
and U843 (N_843,In_1084,In_251);
or U844 (N_844,N_616,N_792);
and U845 (N_845,N_733,N_118);
nor U846 (N_846,N_717,In_718);
nand U847 (N_847,In_717,N_771);
and U848 (N_848,N_271,N_440);
nand U849 (N_849,N_627,In_916);
xnor U850 (N_850,In_1700,In_2126);
nand U851 (N_851,N_510,N_798);
or U852 (N_852,N_19,N_398);
xnor U853 (N_853,In_872,N_357);
xor U854 (N_854,In_2072,In_2495);
or U855 (N_855,N_712,In_2264);
nor U856 (N_856,N_101,In_873);
or U857 (N_857,In_313,N_739);
xor U858 (N_858,N_407,In_1564);
xnor U859 (N_859,N_462,In_351);
nor U860 (N_860,In_1942,N_730);
nor U861 (N_861,In_1510,In_216);
or U862 (N_862,In_2198,In_2082);
or U863 (N_863,In_197,N_546);
nor U864 (N_864,N_490,In_2193);
nor U865 (N_865,N_214,In_828);
nor U866 (N_866,In_403,N_639);
xor U867 (N_867,N_6,N_213);
nor U868 (N_868,N_337,In_423);
and U869 (N_869,In_361,N_504);
nor U870 (N_870,In_1742,N_732);
xor U871 (N_871,In_2481,In_719);
and U872 (N_872,In_224,N_320);
xor U873 (N_873,In_818,In_741);
and U874 (N_874,In_2330,In_1002);
or U875 (N_875,In_1779,In_1981);
xnor U876 (N_876,N_483,In_2436);
or U877 (N_877,N_295,N_606);
or U878 (N_878,N_570,In_657);
and U879 (N_879,N_322,N_485);
xnor U880 (N_880,In_2171,In_2225);
or U881 (N_881,In_1067,In_642);
nand U882 (N_882,N_232,N_494);
nor U883 (N_883,In_2300,In_607);
or U884 (N_884,In_2314,N_169);
or U885 (N_885,N_278,In_2036);
nand U886 (N_886,In_1747,In_1413);
or U887 (N_887,In_1869,In_1892);
nor U888 (N_888,In_83,In_2325);
nor U889 (N_889,N_521,N_215);
nand U890 (N_890,In_1338,N_736);
nand U891 (N_891,In_191,N_745);
and U892 (N_892,In_930,In_2139);
nand U893 (N_893,In_1643,In_1702);
nor U894 (N_894,In_2088,N_371);
nor U895 (N_895,N_270,In_492);
nand U896 (N_896,In_108,N_265);
xor U897 (N_897,N_760,N_646);
xnor U898 (N_898,N_91,N_455);
xnor U899 (N_899,In_1114,In_1047);
and U900 (N_900,In_497,N_715);
nand U901 (N_901,N_618,N_282);
nand U902 (N_902,In_404,In_1868);
and U903 (N_903,N_288,In_889);
or U904 (N_904,In_2496,N_752);
and U905 (N_905,In_591,N_791);
nor U906 (N_906,In_377,In_19);
nand U907 (N_907,N_749,N_316);
nand U908 (N_908,In_1397,In_1544);
nor U909 (N_909,In_774,In_700);
nor U910 (N_910,In_352,In_1285);
nand U911 (N_911,In_1956,N_526);
xor U912 (N_912,In_1587,In_502);
nand U913 (N_913,N_662,In_1690);
xor U914 (N_914,N_164,In_876);
and U915 (N_915,In_1706,In_811);
and U916 (N_916,In_2459,In_2048);
nor U917 (N_917,In_385,In_1055);
nand U918 (N_918,In_1086,N_190);
xor U919 (N_919,In_2359,N_503);
xnor U920 (N_920,In_928,N_640);
xor U921 (N_921,In_629,In_302);
or U922 (N_922,In_716,N_258);
nand U923 (N_923,N_658,In_1935);
or U924 (N_924,In_853,In_1718);
nand U925 (N_925,N_395,In_2181);
nand U926 (N_926,In_2208,In_442);
xor U927 (N_927,N_463,N_196);
xor U928 (N_928,In_1170,In_583);
xor U929 (N_929,In_1112,N_143);
and U930 (N_930,N_608,N_409);
xor U931 (N_931,In_2306,In_1539);
or U932 (N_932,In_782,In_2260);
xnor U933 (N_933,N_596,In_1269);
nand U934 (N_934,N_148,In_1166);
nor U935 (N_935,In_1103,In_1856);
and U936 (N_936,N_291,N_654);
and U937 (N_937,In_986,In_2011);
xnor U938 (N_938,N_421,N_127);
nor U939 (N_939,In_1414,N_587);
xnor U940 (N_940,N_508,N_566);
and U941 (N_941,In_970,In_1843);
and U942 (N_942,N_610,N_321);
nand U943 (N_943,In_177,N_133);
nor U944 (N_944,In_1542,In_1778);
or U945 (N_945,In_903,N_247);
xnor U946 (N_946,In_1205,In_39);
nand U947 (N_947,In_703,In_715);
nand U948 (N_948,N_547,In_1924);
and U949 (N_949,N_108,In_958);
nor U950 (N_950,N_428,N_734);
and U951 (N_951,In_655,In_486);
nor U952 (N_952,In_2109,In_387);
nand U953 (N_953,N_413,In_936);
and U954 (N_954,N_42,In_1280);
xnor U955 (N_955,In_663,N_423);
xnor U956 (N_956,In_1377,N_450);
xnor U957 (N_957,N_597,N_583);
and U958 (N_958,In_2374,In_2365);
nor U959 (N_959,In_1042,In_854);
and U960 (N_960,In_1099,N_174);
and U961 (N_961,In_559,In_2254);
nor U962 (N_962,In_1941,In_261);
and U963 (N_963,In_1003,In_282);
nand U964 (N_964,In_1575,In_850);
and U965 (N_965,In_1096,N_687);
and U966 (N_966,N_225,In_1980);
xnor U967 (N_967,In_1197,In_1257);
xnor U968 (N_968,In_1236,N_694);
and U969 (N_969,In_245,N_275);
and U970 (N_970,N_392,N_73);
nor U971 (N_971,In_1720,In_1302);
nand U972 (N_972,In_539,In_1014);
nand U973 (N_973,In_542,N_558);
nor U974 (N_974,In_1021,In_354);
nor U975 (N_975,In_5,N_155);
or U976 (N_976,In_639,In_2012);
xor U977 (N_977,In_2421,In_1829);
and U978 (N_978,In_1819,In_1644);
and U979 (N_979,In_630,In_2161);
and U980 (N_980,N_703,N_708);
and U981 (N_981,N_445,In_44);
nand U982 (N_982,In_1075,In_231);
or U983 (N_983,In_2403,N_761);
or U984 (N_984,In_2467,In_319);
nor U985 (N_985,In_223,N_469);
and U986 (N_986,In_91,N_601);
and U987 (N_987,In_330,In_611);
nor U988 (N_988,In_368,In_2064);
xnor U989 (N_989,In_776,In_2290);
or U990 (N_990,In_885,In_1029);
or U991 (N_991,In_421,In_874);
or U992 (N_992,In_2324,In_2368);
and U993 (N_993,In_2267,In_1954);
nand U994 (N_994,In_470,In_1382);
or U995 (N_995,In_2009,In_1705);
and U996 (N_996,In_1136,In_1477);
or U997 (N_997,In_2387,N_527);
nand U998 (N_998,In_768,In_730);
or U999 (N_999,N_650,N_218);
and U1000 (N_1000,In_547,In_1348);
xnor U1001 (N_1001,In_1723,In_1789);
or U1002 (N_1002,N_111,In_185);
nor U1003 (N_1003,N_686,In_1759);
nand U1004 (N_1004,In_983,In_1473);
nor U1005 (N_1005,In_193,N_612);
and U1006 (N_1006,In_89,N_747);
nor U1007 (N_1007,N_367,In_2019);
xor U1008 (N_1008,N_571,N_999);
nor U1009 (N_1009,In_1791,In_1038);
nor U1010 (N_1010,In_1088,In_198);
and U1011 (N_1011,N_935,In_1939);
nor U1012 (N_1012,N_971,N_998);
xor U1013 (N_1013,In_1993,In_1058);
and U1014 (N_1014,In_1098,In_2118);
and U1015 (N_1015,N_632,In_1586);
nand U1016 (N_1016,In_996,N_598);
nand U1017 (N_1017,In_743,In_283);
or U1018 (N_1018,In_636,N_801);
and U1019 (N_1019,In_1151,In_1219);
and U1020 (N_1020,N_713,In_1231);
nand U1021 (N_1021,In_920,N_4);
and U1022 (N_1022,N_969,In_2479);
xor U1023 (N_1023,N_836,In_678);
nand U1024 (N_1024,N_963,N_702);
xor U1025 (N_1025,In_1315,In_275);
or U1026 (N_1026,In_2391,N_652);
xnor U1027 (N_1027,N_774,In_562);
nor U1028 (N_1028,N_868,N_711);
nor U1029 (N_1029,N_272,In_888);
and U1030 (N_1030,N_822,N_623);
nor U1031 (N_1031,In_1904,N_29);
xor U1032 (N_1032,N_301,In_1140);
xnor U1033 (N_1033,N_957,In_1572);
nand U1034 (N_1034,In_1621,In_277);
nor U1035 (N_1035,In_971,N_565);
and U1036 (N_1036,In_1165,In_1795);
xnor U1037 (N_1037,In_514,N_507);
or U1038 (N_1038,In_474,In_1557);
nor U1039 (N_1039,N_809,In_1428);
xor U1040 (N_1040,In_1588,In_1432);
nand U1041 (N_1041,In_1443,In_1384);
nor U1042 (N_1042,In_241,N_396);
nand U1043 (N_1043,N_743,In_1449);
or U1044 (N_1044,In_867,In_992);
and U1045 (N_1045,In_2342,In_1451);
nand U1046 (N_1046,In_1184,In_736);
nand U1047 (N_1047,N_500,In_485);
nand U1048 (N_1048,N_673,N_670);
and U1049 (N_1049,N_498,N_729);
and U1050 (N_1050,In_1664,In_934);
xnor U1051 (N_1051,In_981,In_270);
nor U1052 (N_1052,N_355,N_493);
and U1053 (N_1053,In_675,In_859);
nand U1054 (N_1054,In_2406,N_922);
and U1055 (N_1055,N_312,N_679);
xnor U1056 (N_1056,In_973,In_1649);
and U1057 (N_1057,In_2174,In_1988);
xor U1058 (N_1058,In_1210,In_2435);
and U1059 (N_1059,N_408,N_707);
nand U1060 (N_1060,N_261,In_1123);
nor U1061 (N_1061,N_917,In_1503);
and U1062 (N_1062,N_846,In_1857);
nor U1063 (N_1063,In_1495,In_2152);
xnor U1064 (N_1064,N_302,In_1709);
and U1065 (N_1065,N_856,In_919);
nand U1066 (N_1066,In_784,N_780);
nand U1067 (N_1067,N_577,In_2281);
and U1068 (N_1068,In_1362,In_269);
and U1069 (N_1069,In_480,In_1445);
nand U1070 (N_1070,In_2257,N_300);
or U1071 (N_1071,In_795,In_1686);
or U1072 (N_1072,In_672,N_981);
or U1073 (N_1073,N_851,In_1368);
nand U1074 (N_1074,N_251,In_857);
and U1075 (N_1075,In_792,N_136);
or U1076 (N_1076,N_562,In_1977);
nor U1077 (N_1077,N_834,In_722);
nor U1078 (N_1078,N_242,N_390);
nor U1079 (N_1079,In_490,In_2398);
nand U1080 (N_1080,In_1117,N_180);
xnor U1081 (N_1081,In_977,N_926);
or U1082 (N_1082,In_1175,N_452);
nand U1083 (N_1083,In_333,N_789);
and U1084 (N_1084,N_915,In_1733);
or U1085 (N_1085,In_2326,N_976);
nand U1086 (N_1086,In_86,N_21);
xnor U1087 (N_1087,In_2206,N_663);
nand U1088 (N_1088,In_596,N_859);
xor U1089 (N_1089,N_240,N_664);
nand U1090 (N_1090,N_908,In_1113);
or U1091 (N_1091,In_2078,In_685);
xor U1092 (N_1092,In_764,In_1507);
and U1093 (N_1093,N_539,In_2101);
nor U1094 (N_1094,N_235,In_1426);
nand U1095 (N_1095,In_2451,N_464);
or U1096 (N_1096,N_776,In_2355);
and U1097 (N_1097,N_63,In_1387);
nand U1098 (N_1098,In_807,In_1629);
and U1099 (N_1099,N_751,In_1249);
or U1100 (N_1100,In_2379,In_2437);
or U1101 (N_1101,In_894,N_93);
nand U1102 (N_1102,In_1022,N_941);
nor U1103 (N_1103,In_775,In_2053);
or U1104 (N_1104,N_556,N_879);
and U1105 (N_1105,N_76,In_862);
nand U1106 (N_1106,In_907,In_2045);
nand U1107 (N_1107,N_132,In_2441);
or U1108 (N_1108,In_447,N_273);
nor U1109 (N_1109,N_795,N_292);
nor U1110 (N_1110,In_1550,N_67);
or U1111 (N_1111,N_399,In_998);
nor U1112 (N_1112,N_559,In_721);
xor U1113 (N_1113,In_1622,N_635);
nand U1114 (N_1114,In_1808,N_721);
xor U1115 (N_1115,N_97,In_2335);
or U1116 (N_1116,In_841,N_208);
or U1117 (N_1117,In_2412,N_374);
and U1118 (N_1118,In_1802,In_1872);
or U1119 (N_1119,In_1768,In_1017);
and U1120 (N_1120,N_379,In_534);
or U1121 (N_1121,In_1125,In_654);
nand U1122 (N_1122,N_973,In_1822);
or U1123 (N_1123,N_660,N_31);
nor U1124 (N_1124,In_701,N_548);
nor U1125 (N_1125,N_363,In_624);
and U1126 (N_1126,In_1234,In_751);
and U1127 (N_1127,In_266,In_1761);
xor U1128 (N_1128,N_315,In_2268);
and U1129 (N_1129,In_2095,N_719);
and U1130 (N_1130,In_1684,N_910);
nor U1131 (N_1131,N_704,In_2209);
or U1132 (N_1132,In_1292,N_864);
or U1133 (N_1133,N_476,In_1741);
and U1134 (N_1134,N_896,In_584);
xor U1135 (N_1135,In_2010,N_666);
or U1136 (N_1136,In_1375,In_545);
nand U1137 (N_1137,In_309,N_480);
xor U1138 (N_1138,In_1145,N_782);
and U1139 (N_1139,N_754,In_1191);
xor U1140 (N_1140,In_1734,In_2079);
and U1141 (N_1141,In_2002,N_676);
xnor U1142 (N_1142,In_761,In_85);
or U1143 (N_1143,N_178,N_759);
xnor U1144 (N_1144,In_513,N_930);
nor U1145 (N_1145,N_992,N_914);
and U1146 (N_1146,In_126,N_977);
nand U1147 (N_1147,N_644,In_821);
and U1148 (N_1148,In_2003,In_130);
xnor U1149 (N_1149,N_818,N_674);
nor U1150 (N_1150,N_944,In_1849);
xor U1151 (N_1151,In_969,N_51);
or U1152 (N_1152,In_772,N_366);
or U1153 (N_1153,In_271,In_1576);
and U1154 (N_1154,In_790,In_33);
xnor U1155 (N_1155,In_410,In_1246);
nor U1156 (N_1156,In_62,In_1609);
xnor U1157 (N_1157,N_362,In_2204);
or U1158 (N_1158,In_2219,N_773);
and U1159 (N_1159,In_2416,In_291);
and U1160 (N_1160,N_447,N_726);
nand U1161 (N_1161,N_807,In_668);
nand U1162 (N_1162,In_167,N_906);
or U1163 (N_1163,N_875,In_2124);
nor U1164 (N_1164,In_1654,N_263);
and U1165 (N_1165,N_731,N_167);
nand U1166 (N_1166,In_571,N_835);
xor U1167 (N_1167,N_360,In_27);
nor U1168 (N_1168,In_2494,N_756);
nand U1169 (N_1169,In_684,In_1728);
or U1170 (N_1170,In_1155,In_1089);
and U1171 (N_1171,In_25,In_910);
and U1172 (N_1172,In_737,N_152);
nor U1173 (N_1173,In_1963,In_2393);
nand U1174 (N_1174,In_226,N_843);
and U1175 (N_1175,In_1105,N_832);
and U1176 (N_1176,In_2250,In_686);
nand U1177 (N_1177,N_891,In_2308);
nor U1178 (N_1178,In_1648,In_1416);
and U1179 (N_1179,N_988,In_1199);
xor U1180 (N_1180,N_948,In_2336);
and U1181 (N_1181,N_528,In_1633);
xor U1182 (N_1182,N_453,In_830);
xor U1183 (N_1183,N_481,In_1635);
xor U1184 (N_1184,N_860,In_15);
and U1185 (N_1185,In_2241,N_349);
nand U1186 (N_1186,In_2389,N_149);
nor U1187 (N_1187,In_1110,N_572);
xnor U1188 (N_1188,In_204,In_1655);
xor U1189 (N_1189,In_1070,In_1826);
and U1190 (N_1190,N_188,In_906);
and U1191 (N_1191,N_965,In_1100);
and U1192 (N_1192,In_290,In_155);
nand U1193 (N_1193,N_786,N_928);
xor U1194 (N_1194,In_1695,N_872);
or U1195 (N_1195,N_394,N_858);
nand U1196 (N_1196,In_1729,N_433);
and U1197 (N_1197,In_527,N_329);
or U1198 (N_1198,N_239,N_958);
and U1199 (N_1199,N_354,In_2304);
nand U1200 (N_1200,In_1411,In_1279);
xnor U1201 (N_1201,N_352,N_1033);
nor U1202 (N_1202,In_104,In_1093);
nand U1203 (N_1203,In_704,N_833);
nor U1204 (N_1204,N_1056,In_1417);
nand U1205 (N_1205,In_1699,In_1726);
and U1206 (N_1206,In_2196,N_1079);
xnor U1207 (N_1207,N_1115,In_1238);
nor U1208 (N_1208,In_21,N_432);
nand U1209 (N_1209,N_400,N_1074);
or U1210 (N_1210,N_451,N_92);
or U1211 (N_1211,In_278,N_599);
nor U1212 (N_1212,N_862,N_537);
and U1213 (N_1213,N_1113,N_74);
nand U1214 (N_1214,In_2180,In_964);
and U1215 (N_1215,In_1310,N_959);
xor U1216 (N_1216,N_1091,N_1145);
or U1217 (N_1217,N_1142,N_890);
nor U1218 (N_1218,In_190,N_659);
and U1219 (N_1219,In_2370,N_667);
nand U1220 (N_1220,In_1079,In_1606);
and U1221 (N_1221,In_2462,N_17);
xor U1222 (N_1222,In_1474,N_330);
xnor U1223 (N_1223,N_1040,In_759);
or U1224 (N_1224,N_887,N_871);
or U1225 (N_1225,N_1029,In_1160);
and U1226 (N_1226,In_1440,N_175);
nor U1227 (N_1227,N_980,In_1116);
nor U1228 (N_1228,In_1288,N_1084);
xor U1229 (N_1229,N_443,N_245);
nor U1230 (N_1230,In_1803,In_587);
or U1231 (N_1231,In_1760,N_683);
or U1232 (N_1232,N_129,N_206);
nand U1233 (N_1233,N_1086,N_1167);
nor U1234 (N_1234,N_1193,N_805);
and U1235 (N_1235,In_2329,In_802);
xnor U1236 (N_1236,N_927,N_723);
nor U1237 (N_1237,N_153,In_909);
or U1238 (N_1238,N_16,N_894);
and U1239 (N_1239,N_602,N_611);
xnor U1240 (N_1240,In_1087,N_933);
xnor U1241 (N_1241,In_1294,In_1143);
and U1242 (N_1242,In_2057,In_1722);
and U1243 (N_1243,N_680,In_2034);
or U1244 (N_1244,N_1041,N_1116);
and U1245 (N_1245,N_1057,N_1011);
and U1246 (N_1246,In_2358,In_1313);
nor U1247 (N_1247,N_259,In_2084);
nand U1248 (N_1248,N_1112,N_252);
or U1249 (N_1249,N_266,In_205);
nand U1250 (N_1250,In_1850,In_2229);
nand U1251 (N_1251,N_134,In_556);
or U1252 (N_1252,N_1004,In_1458);
or U1253 (N_1253,N_1022,In_2067);
or U1254 (N_1254,N_808,N_1003);
xor U1255 (N_1255,N_40,N_1026);
nand U1256 (N_1256,In_1460,N_361);
nand U1257 (N_1257,N_35,N_643);
nor U1258 (N_1258,N_430,In_799);
nand U1259 (N_1259,N_457,In_1887);
or U1260 (N_1260,In_985,N_690);
nand U1261 (N_1261,N_59,In_2429);
nand U1262 (N_1262,In_1599,In_195);
nor U1263 (N_1263,N_800,In_2106);
xor U1264 (N_1264,N_578,N_437);
nor U1265 (N_1265,N_499,N_497);
xor U1266 (N_1266,In_1493,In_1059);
nor U1267 (N_1267,N_714,In_2169);
and U1268 (N_1268,In_1784,In_1549);
and U1269 (N_1269,N_637,N_418);
nor U1270 (N_1270,In_2199,In_1456);
xor U1271 (N_1271,In_2111,N_1085);
xnor U1272 (N_1272,In_67,N_1058);
and U1273 (N_1273,In_1171,N_710);
xor U1274 (N_1274,N_411,N_1078);
xor U1275 (N_1275,In_1837,In_1227);
or U1276 (N_1276,In_1254,N_1059);
nor U1277 (N_1277,N_342,In_43);
or U1278 (N_1278,N_1163,N_1017);
nor U1279 (N_1279,N_986,N_764);
nand U1280 (N_1280,N_592,N_45);
nand U1281 (N_1281,In_1531,In_2050);
xnor U1282 (N_1282,N_979,In_2227);
nor U1283 (N_1283,In_1502,N_628);
xnor U1284 (N_1284,N_345,In_1077);
nand U1285 (N_1285,N_962,N_14);
nand U1286 (N_1286,N_1083,N_938);
and U1287 (N_1287,N_1149,N_283);
or U1288 (N_1288,N_39,In_1516);
nand U1289 (N_1289,N_884,N_522);
and U1290 (N_1290,In_2404,In_1986);
nand U1291 (N_1291,In_1830,N_770);
nand U1292 (N_1292,N_1082,N_994);
xnor U1293 (N_1293,N_1190,N_1125);
nand U1294 (N_1294,In_1685,N_765);
or U1295 (N_1295,N_202,N_1188);
or U1296 (N_1296,N_531,In_1415);
nand U1297 (N_1297,In_2422,In_606);
nand U1298 (N_1298,N_1015,In_1561);
xor U1299 (N_1299,In_680,In_1511);
nor U1300 (N_1300,In_933,N_1053);
nand U1301 (N_1301,In_1807,In_788);
nor U1302 (N_1302,N_1198,In_219);
nor U1303 (N_1303,N_552,N_873);
xnor U1304 (N_1304,N_1080,N_1044);
or U1305 (N_1305,In_580,In_1008);
nand U1306 (N_1306,In_152,In_255);
and U1307 (N_1307,In_2431,In_1323);
nor U1308 (N_1308,In_823,N_431);
nor U1309 (N_1309,In_2112,N_841);
and U1310 (N_1310,N_520,N_692);
xnor U1311 (N_1311,In_555,N_304);
or U1312 (N_1312,N_877,In_230);
or U1313 (N_1313,In_708,In_1533);
or U1314 (N_1314,In_2414,N_880);
nor U1315 (N_1315,N_695,N_929);
nor U1316 (N_1316,N_1036,In_1888);
xnor U1317 (N_1317,In_1033,In_1624);
xor U1318 (N_1318,N_735,In_1137);
nor U1319 (N_1319,In_1282,In_135);
or U1320 (N_1320,In_553,N_274);
nor U1321 (N_1321,N_641,N_234);
or U1322 (N_1322,N_1055,N_27);
nor U1323 (N_1323,In_244,N_26);
nor U1324 (N_1324,In_1675,In_826);
and U1325 (N_1325,In_600,In_793);
or U1326 (N_1326,N_600,N_802);
xor U1327 (N_1327,In_1242,In_2107);
nand U1328 (N_1328,In_1651,N_335);
nor U1329 (N_1329,N_1093,N_893);
or U1330 (N_1330,N_517,In_273);
nand U1331 (N_1331,In_443,N_237);
nand U1332 (N_1332,N_166,N_1136);
nor U1333 (N_1333,In_1970,In_1154);
or U1334 (N_1334,In_877,N_1031);
xor U1335 (N_1335,In_806,In_1472);
nand U1336 (N_1336,N_439,In_1322);
nand U1337 (N_1337,N_332,N_359);
and U1338 (N_1338,N_661,N_993);
nor U1339 (N_1339,N_489,N_1143);
or U1340 (N_1340,N_1178,In_2312);
nor U1341 (N_1341,In_982,N_645);
nor U1342 (N_1342,In_1252,N_1048);
nand U1343 (N_1343,N_1060,In_1500);
nor U1344 (N_1344,In_2238,N_64);
nor U1345 (N_1345,In_120,N_1195);
xnor U1346 (N_1346,In_1424,In_2035);
xor U1347 (N_1347,N_763,In_1512);
nor U1348 (N_1348,N_488,In_938);
or U1349 (N_1349,N_724,In_1625);
and U1350 (N_1350,In_1982,N_784);
nand U1351 (N_1351,N_755,N_720);
and U1352 (N_1352,N_1135,In_643);
and U1353 (N_1353,In_1403,In_512);
or U1354 (N_1354,N_1076,In_248);
xnor U1355 (N_1355,In_1207,In_156);
nor U1356 (N_1356,In_2428,In_2215);
and U1357 (N_1357,In_110,In_2410);
or U1358 (N_1358,N_681,N_1108);
xor U1359 (N_1359,In_1255,In_1369);
xnor U1360 (N_1360,N_684,In_875);
nor U1361 (N_1361,In_1852,N_1121);
nand U1362 (N_1362,In_280,N_144);
or U1363 (N_1363,In_1816,N_1028);
nor U1364 (N_1364,N_544,In_989);
and U1365 (N_1365,N_1182,N_1162);
and U1366 (N_1366,N_66,N_709);
and U1367 (N_1367,In_260,N_865);
nand U1368 (N_1368,In_2262,In_922);
nor U1369 (N_1369,In_1419,N_1009);
xor U1370 (N_1370,N_895,N_1002);
nand U1371 (N_1371,In_1066,In_207);
and U1372 (N_1372,In_927,In_2042);
and U1373 (N_1373,In_550,N_465);
or U1374 (N_1374,N_1124,In_2439);
and U1375 (N_1375,N_982,In_140);
and U1376 (N_1376,In_1078,N_823);
nor U1377 (N_1377,N_194,N_634);
xor U1378 (N_1378,In_2284,N_876);
and U1379 (N_1379,N_1151,In_1035);
nor U1380 (N_1380,N_777,N_1069);
xnor U1381 (N_1381,N_626,N_326);
nor U1382 (N_1382,In_2488,In_1775);
and U1383 (N_1383,N_817,N_631);
and U1384 (N_1384,In_38,In_411);
nor U1385 (N_1385,N_1133,N_353);
and U1386 (N_1386,N_767,N_869);
nand U1387 (N_1387,In_918,In_2256);
or U1388 (N_1388,N_1046,N_700);
nand U1389 (N_1389,N_1132,N_1126);
and U1390 (N_1390,In_1562,In_1190);
nor U1391 (N_1391,N_672,In_459);
nand U1392 (N_1392,N_1019,In_1286);
nor U1393 (N_1393,N_665,N_840);
nand U1394 (N_1394,In_0,N_1166);
or U1395 (N_1395,In_1217,N_417);
and U1396 (N_1396,N_422,In_12);
or U1397 (N_1397,In_1751,N_668);
or U1398 (N_1398,N_744,N_204);
or U1399 (N_1399,N_947,In_391);
nor U1400 (N_1400,In_2390,N_796);
nor U1401 (N_1401,In_454,N_519);
nand U1402 (N_1402,N_847,N_470);
xnor U1403 (N_1403,In_373,In_1938);
nor U1404 (N_1404,N_1240,In_1346);
nand U1405 (N_1405,N_638,N_900);
nand U1406 (N_1406,N_1398,N_1262);
and U1407 (N_1407,N_1281,In_1556);
xor U1408 (N_1408,N_1183,In_1683);
nand U1409 (N_1409,N_693,N_195);
and U1410 (N_1410,N_1154,N_372);
nand U1411 (N_1411,In_233,In_51);
and U1412 (N_1412,N_1228,N_198);
nor U1413 (N_1413,N_381,N_804);
nand U1414 (N_1414,In_1918,N_1327);
and U1415 (N_1415,N_607,In_1570);
nor U1416 (N_1416,N_970,N_581);
xor U1417 (N_1417,N_1035,N_365);
or U1418 (N_1418,In_1890,N_446);
and U1419 (N_1419,N_1043,In_724);
and U1420 (N_1420,In_1216,N_1077);
xor U1421 (N_1421,N_1237,N_1263);
nor U1422 (N_1422,N_621,In_1094);
nor U1423 (N_1423,N_406,N_77);
xor U1424 (N_1424,N_1000,N_1353);
and U1425 (N_1425,N_820,In_320);
xnor U1426 (N_1426,N_945,N_294);
nand U1427 (N_1427,In_1244,In_2222);
and U1428 (N_1428,N_1358,In_1650);
and U1429 (N_1429,In_2175,In_1466);
or U1430 (N_1430,N_1045,N_983);
xor U1431 (N_1431,In_2492,In_2089);
nor U1432 (N_1432,N_1222,N_306);
nand U1433 (N_1433,In_738,In_1914);
or U1434 (N_1434,In_218,In_2476);
or U1435 (N_1435,N_1114,N_826);
or U1436 (N_1436,N_1303,N_1170);
xor U1437 (N_1437,In_1573,In_1659);
or U1438 (N_1438,In_1737,N_1378);
and U1439 (N_1439,In_1798,N_1369);
and U1440 (N_1440,In_577,N_613);
or U1441 (N_1441,In_1124,In_66);
and U1442 (N_1442,N_257,N_317);
or U1443 (N_1443,In_69,In_1902);
xnor U1444 (N_1444,In_317,N_460);
or U1445 (N_1445,In_843,In_2114);
nand U1446 (N_1446,N_1047,N_1309);
or U1447 (N_1447,N_1391,N_728);
and U1448 (N_1448,N_364,In_363);
xnor U1449 (N_1449,N_1130,In_1640);
nor U1450 (N_1450,In_37,In_726);
nor U1451 (N_1451,N_1273,N_705);
nor U1452 (N_1452,N_874,N_1377);
or U1453 (N_1453,N_762,N_727);
nand U1454 (N_1454,N_1230,N_1367);
and U1455 (N_1455,N_1308,N_757);
or U1456 (N_1456,In_2305,N_946);
or U1457 (N_1457,N_1250,N_960);
and U1458 (N_1458,In_627,N_974);
or U1459 (N_1459,N_1209,In_364);
and U1460 (N_1460,N_912,N_790);
nor U1461 (N_1461,N_226,N_1150);
nor U1462 (N_1462,N_913,In_327);
nand U1463 (N_1463,N_1247,N_1204);
or U1464 (N_1464,N_888,In_332);
xnor U1465 (N_1465,N_964,N_656);
and U1466 (N_1466,N_813,In_296);
nor U1467 (N_1467,N_1242,In_2005);
nor U1468 (N_1468,In_1909,N_1334);
and U1469 (N_1469,N_814,In_2296);
or U1470 (N_1470,In_1711,N_1164);
and U1471 (N_1471,N_810,In_2210);
xnor U1472 (N_1472,N_655,N_1386);
nand U1473 (N_1473,In_1036,N_525);
nand U1474 (N_1474,N_1147,N_1236);
nand U1475 (N_1475,N_1052,N_1312);
xnor U1476 (N_1476,N_923,N_1224);
or U1477 (N_1477,In_1999,In_487);
xor U1478 (N_1478,In_834,In_2408);
and U1479 (N_1479,In_581,In_711);
nand U1480 (N_1480,In_456,In_1452);
or U1481 (N_1481,N_1025,In_2348);
xor U1482 (N_1482,N_1089,In_2292);
xor U1483 (N_1483,N_748,In_1652);
nand U1484 (N_1484,In_2211,N_1356);
or U1485 (N_1485,N_1393,N_1300);
nand U1486 (N_1486,N_1324,In_165);
xnor U1487 (N_1487,N_1021,N_1208);
nor U1488 (N_1488,In_1152,N_1368);
or U1489 (N_1489,N_1344,N_1090);
nor U1490 (N_1490,N_1157,N_901);
nand U1491 (N_1491,N_1348,In_2184);
xnor U1492 (N_1492,N_1234,In_1882);
nand U1493 (N_1493,N_1323,In_1583);
nand U1494 (N_1494,N_181,In_2141);
nor U1495 (N_1495,N_1289,In_1463);
nand U1496 (N_1496,N_636,N_33);
and U1497 (N_1497,In_1740,N_1317);
nand U1498 (N_1498,N_972,In_2464);
or U1499 (N_1499,N_1068,N_1279);
or U1500 (N_1500,N_1357,In_714);
xnor U1501 (N_1501,N_1220,In_132);
xor U1502 (N_1502,In_943,N_775);
or U1503 (N_1503,N_1023,N_867);
xnor U1504 (N_1504,N_41,N_1111);
nor U1505 (N_1505,N_557,N_1227);
or U1506 (N_1506,N_1274,N_1128);
nand U1507 (N_1507,N_1148,N_949);
or U1508 (N_1508,N_920,N_269);
xor U1509 (N_1509,N_1229,In_2498);
nor U1510 (N_1510,In_1380,N_1255);
nor U1511 (N_1511,N_65,N_1318);
and U1512 (N_1512,N_1226,N_1319);
nor U1513 (N_1513,N_57,N_1097);
nand U1514 (N_1514,N_936,N_698);
xnor U1515 (N_1515,N_104,In_465);
nand U1516 (N_1516,In_848,In_1339);
nor U1517 (N_1517,N_997,N_1277);
and U1518 (N_1518,N_603,N_58);
nand U1519 (N_1519,In_1704,N_535);
xor U1520 (N_1520,N_47,N_1257);
nand U1521 (N_1521,N_1373,N_1205);
nand U1522 (N_1522,N_857,N_1330);
and U1523 (N_1523,N_586,N_540);
nor U1524 (N_1524,N_1305,N_555);
nor U1525 (N_1525,N_677,In_1284);
and U1526 (N_1526,N_919,In_347);
nor U1527 (N_1527,N_898,N_419);
and U1528 (N_1528,In_1790,N_1248);
xor U1529 (N_1529,In_1109,In_315);
nor U1530 (N_1530,In_1494,N_513);
xor U1531 (N_1531,N_1387,N_1329);
xor U1532 (N_1532,In_1334,In_2450);
or U1533 (N_1533,N_955,N_1217);
or U1534 (N_1534,In_2455,N_1054);
xor U1535 (N_1535,N_951,In_960);
nor U1536 (N_1536,N_109,In_1228);
nand U1537 (N_1537,In_681,N_909);
nor U1538 (N_1538,In_1630,N_1333);
and U1539 (N_1539,N_787,In_232);
and U1540 (N_1540,N_931,N_211);
and U1541 (N_1541,In_498,N_1276);
or U1542 (N_1542,N_984,N_116);
nand U1543 (N_1543,N_454,N_1272);
xnor U1544 (N_1544,N_1337,N_10);
xnor U1545 (N_1545,N_380,In_150);
and U1546 (N_1546,N_1212,In_2466);
xor U1547 (N_1547,In_1506,N_902);
nor U1548 (N_1548,N_1332,N_1020);
and U1549 (N_1549,N_1346,N_323);
or U1550 (N_1550,In_2376,N_1379);
xnor U1551 (N_1551,N_1361,In_2301);
and U1552 (N_1552,N_718,In_2039);
xor U1553 (N_1553,N_1380,N_737);
nand U1554 (N_1554,N_1175,N_1034);
and U1555 (N_1555,In_1637,In_1976);
or U1556 (N_1556,In_2307,In_838);
xor U1557 (N_1557,N_614,In_2367);
and U1558 (N_1558,N_1176,In_1878);
nand U1559 (N_1559,N_1253,N_486);
nor U1560 (N_1560,In_2352,N_620);
nand U1561 (N_1561,In_378,N_989);
or U1562 (N_1562,N_905,In_484);
nor U1563 (N_1563,In_937,N_899);
and U1564 (N_1564,In_773,In_1738);
xor U1565 (N_1565,In_2069,N_1360);
and U1566 (N_1566,N_701,N_89);
or U1567 (N_1567,In_1947,N_246);
nor U1568 (N_1568,In_2061,N_1146);
and U1569 (N_1569,In_125,In_472);
or U1570 (N_1570,In_925,In_886);
nor U1571 (N_1571,N_171,N_1302);
or U1572 (N_1572,N_753,In_551);
nor U1573 (N_1573,N_1328,N_678);
and U1574 (N_1574,In_326,N_1350);
or U1575 (N_1575,In_815,N_1372);
nand U1576 (N_1576,N_1315,In_1062);
or U1577 (N_1577,N_1213,N_1032);
xnor U1578 (N_1578,In_1949,N_1362);
and U1579 (N_1579,In_1927,N_553);
nand U1580 (N_1580,N_184,N_1382);
nor U1581 (N_1581,N_201,N_615);
and U1582 (N_1582,In_1821,N_397);
xnor U1583 (N_1583,N_1061,In_1846);
or U1584 (N_1584,N_1216,In_139);
xor U1585 (N_1585,N_870,N_1005);
and U1586 (N_1586,N_1284,In_1239);
xnor U1587 (N_1587,N_1042,In_2235);
and U1588 (N_1588,N_629,N_815);
or U1589 (N_1589,N_71,N_220);
nand U1590 (N_1590,In_1309,N_1008);
nor U1591 (N_1591,N_940,N_135);
nor U1592 (N_1592,N_1290,In_1131);
nand U1593 (N_1593,N_207,N_62);
nand U1594 (N_1594,N_831,N_382);
xor U1595 (N_1595,N_1160,N_1340);
nand U1596 (N_1596,N_1189,N_1181);
nand U1597 (N_1597,N_533,N_1101);
nand U1598 (N_1598,In_613,N_427);
and U1599 (N_1599,In_501,N_594);
xnor U1600 (N_1600,N_595,N_1286);
nand U1601 (N_1601,N_1428,N_1556);
or U1602 (N_1602,In_1102,N_1285);
and U1603 (N_1603,N_1463,In_1101);
or U1604 (N_1604,N_1480,N_280);
or U1605 (N_1605,N_1409,In_2449);
xnor U1606 (N_1606,In_1672,N_1511);
nand U1607 (N_1607,N_1064,In_2345);
nor U1608 (N_1608,In_735,N_1037);
nand U1609 (N_1609,N_1457,In_595);
nand U1610 (N_1610,N_1464,In_576);
xor U1611 (N_1611,In_2381,N_81);
nor U1612 (N_1612,In_1797,In_2411);
or U1613 (N_1613,N_824,N_1535);
xnor U1614 (N_1614,N_1343,N_1338);
nand U1615 (N_1615,N_1423,N_1313);
or U1616 (N_1616,N_1474,In_780);
or U1617 (N_1617,N_1252,In_1874);
nor U1618 (N_1618,In_1559,In_2425);
xor U1619 (N_1619,N_386,N_1451);
nand U1620 (N_1620,N_1591,N_1172);
and U1621 (N_1621,N_589,N_609);
xnor U1622 (N_1622,N_331,N_1461);
nor U1623 (N_1623,N_1296,N_630);
or U1624 (N_1624,N_1336,In_114);
and U1625 (N_1625,N_1567,N_878);
nand U1626 (N_1626,N_1321,N_1066);
xnor U1627 (N_1627,N_1500,N_1570);
nand U1628 (N_1628,N_1419,In_698);
nand U1629 (N_1629,N_1088,In_525);
xnor U1630 (N_1630,N_1565,In_752);
nand U1631 (N_1631,N_937,In_2373);
and U1632 (N_1632,In_258,N_456);
nand U1633 (N_1633,In_865,N_1030);
or U1634 (N_1634,In_2277,In_879);
nand U1635 (N_1635,N_1203,N_1443);
nor U1636 (N_1636,N_1298,In_56);
xnor U1637 (N_1637,In_124,In_1189);
nor U1638 (N_1638,N_532,In_890);
xnor U1639 (N_1639,In_2136,In_61);
and U1640 (N_1640,In_1266,N_1518);
and U1641 (N_1641,In_1966,N_758);
nor U1642 (N_1642,N_886,N_803);
nor U1643 (N_1643,N_1499,In_70);
nor U1644 (N_1644,N_827,N_1297);
and U1645 (N_1645,N_1425,N_1184);
xnor U1646 (N_1646,N_1445,In_1991);
nor U1647 (N_1647,N_1494,In_439);
nand U1648 (N_1648,N_138,N_1577);
nor U1649 (N_1649,In_22,N_828);
xor U1650 (N_1650,In_50,N_1541);
xnor U1651 (N_1651,N_298,N_567);
and U1652 (N_1652,N_1165,In_1018);
and U1653 (N_1653,N_1013,N_889);
or U1654 (N_1654,In_2090,N_1129);
nand U1655 (N_1655,N_1339,In_2420);
nor U1656 (N_1656,N_1447,N_649);
or U1657 (N_1657,N_1381,N_1524);
or U1658 (N_1658,N_1471,In_1862);
and U1659 (N_1659,In_740,N_1187);
or U1660 (N_1660,N_819,In_142);
xor U1661 (N_1661,N_1588,N_241);
and U1662 (N_1662,N_799,In_176);
and U1663 (N_1663,N_1456,In_287);
nor U1664 (N_1664,N_1374,N_1583);
nor U1665 (N_1665,N_1095,N_284);
or U1666 (N_1666,In_666,In_394);
and U1667 (N_1667,N_1118,N_1210);
nor U1668 (N_1668,In_966,N_740);
xnor U1669 (N_1669,N_1395,In_993);
or U1670 (N_1670,N_530,In_1832);
nor U1671 (N_1671,In_504,N_1192);
nand U1672 (N_1672,N_1572,In_1969);
nor U1673 (N_1673,N_1370,N_1231);
xnor U1674 (N_1674,N_1385,N_1507);
xnor U1675 (N_1675,N_1206,N_648);
nand U1676 (N_1676,N_1530,In_57);
nand U1677 (N_1677,N_738,N_1141);
or U1678 (N_1678,N_772,N_1418);
xnor U1679 (N_1679,N_1410,In_337);
nand U1680 (N_1680,In_76,N_1351);
nand U1681 (N_1681,In_461,N_1554);
xnor U1682 (N_1682,N_1593,N_966);
xor U1683 (N_1683,N_1155,N_117);
xnor U1684 (N_1684,N_812,N_742);
nand U1685 (N_1685,In_2478,In_945);
and U1686 (N_1686,N_848,N_1072);
or U1687 (N_1687,N_518,N_1173);
or U1688 (N_1688,N_1221,N_1412);
or U1689 (N_1689,N_750,N_1075);
and U1690 (N_1690,N_1420,N_1487);
nand U1691 (N_1691,N_1010,N_1437);
nor U1692 (N_1692,N_1516,N_1469);
xnor U1693 (N_1693,N_1441,In_1095);
nor U1694 (N_1694,In_1121,N_1404);
or U1695 (N_1695,N_1589,N_1123);
nor U1696 (N_1696,In_1667,In_371);
nor U1697 (N_1697,In_2243,In_2442);
nand U1698 (N_1698,In_481,N_1103);
nand U1699 (N_1699,N_1552,N_838);
nor U1700 (N_1700,N_1238,N_1014);
nor U1701 (N_1701,In_1283,N_1528);
nand U1702 (N_1702,N_1452,N_1544);
and U1703 (N_1703,N_1269,N_1468);
nor U1704 (N_1704,N_82,N_1239);
and U1705 (N_1705,In_1972,N_1065);
and U1706 (N_1706,In_524,N_1100);
nand U1707 (N_1707,In_601,N_1291);
xnor U1708 (N_1708,N_1522,N_1293);
xor U1709 (N_1709,N_1376,N_538);
and U1710 (N_1710,In_1320,N_1131);
nand U1711 (N_1711,In_950,N_1446);
or U1712 (N_1712,N_1389,In_2299);
xnor U1713 (N_1713,N_1104,N_1051);
or U1714 (N_1714,In_1721,N_1102);
nor U1715 (N_1715,In_2187,N_1062);
nor U1716 (N_1716,N_1159,N_1137);
nor U1717 (N_1717,In_1833,In_2382);
xor U1718 (N_1718,N_569,N_779);
and U1719 (N_1719,N_1388,N_119);
or U1720 (N_1720,N_1557,N_1551);
nor U1721 (N_1721,In_310,In_509);
or U1722 (N_1722,N_968,N_1563);
and U1723 (N_1723,N_1158,In_635);
and U1724 (N_1724,N_1275,In_307);
xor U1725 (N_1725,N_788,N_186);
nor U1726 (N_1726,In_1435,N_549);
nand U1727 (N_1727,In_316,In_1955);
nor U1728 (N_1728,In_2465,N_1363);
nand U1729 (N_1729,In_2132,N_1413);
nor U1730 (N_1730,N_1270,In_35);
or U1731 (N_1731,In_1756,In_1553);
or U1732 (N_1732,N_146,N_1584);
nor U1733 (N_1733,N_293,N_943);
nand U1734 (N_1734,N_1506,In_646);
nor U1735 (N_1735,N_1120,In_904);
or U1736 (N_1736,N_1218,N_903);
and U1737 (N_1737,In_340,N_1523);
nand U1738 (N_1738,N_1287,In_1478);
xor U1739 (N_1739,N_1543,In_97);
nor U1740 (N_1740,N_794,N_1526);
or U1741 (N_1741,N_1199,N_1105);
and U1742 (N_1742,In_1653,N_1405);
or U1743 (N_1743,In_2115,In_891);
or U1744 (N_1744,N_653,In_350);
nor U1745 (N_1745,In_2164,N_987);
or U1746 (N_1746,N_883,In_250);
or U1747 (N_1747,N_1384,In_516);
nand U1748 (N_1748,N_1180,In_1647);
nand U1749 (N_1749,N_1442,N_297);
xnor U1750 (N_1750,N_1512,N_1092);
nand U1751 (N_1751,N_1191,In_2279);
nand U1752 (N_1752,In_2434,N_1449);
xnor U1753 (N_1753,N_1560,N_224);
and U1754 (N_1754,In_1297,N_622);
nor U1755 (N_1755,N_950,N_482);
and U1756 (N_1756,In_2186,N_1169);
or U1757 (N_1757,In_1605,N_1470);
nand U1758 (N_1758,N_1322,N_746);
nor U1759 (N_1759,In_388,In_2354);
nand U1760 (N_1760,N_1585,N_1533);
and U1761 (N_1761,N_825,N_1434);
xor U1762 (N_1762,N_1261,N_911);
or U1763 (N_1763,N_1472,N_892);
and U1764 (N_1764,In_1230,N_669);
or U1765 (N_1765,In_499,N_1549);
and U1766 (N_1766,N_954,N_1219);
or U1767 (N_1767,N_1568,N_1493);
nand U1768 (N_1768,N_1207,N_1415);
xnor U1769 (N_1769,N_1024,In_1619);
and U1770 (N_1770,N_783,In_144);
nand U1771 (N_1771,N_1063,N_442);
or U1772 (N_1772,In_1940,In_240);
nand U1773 (N_1773,N_484,N_1081);
nor U1774 (N_1774,N_1307,N_1525);
and U1775 (N_1775,N_1498,N_1371);
and U1776 (N_1776,N_1027,N_1258);
nor U1777 (N_1777,N_1596,N_921);
or U1778 (N_1778,N_1416,In_1303);
nand U1779 (N_1779,N_1438,N_1260);
nand U1780 (N_1780,In_1631,N_1504);
and U1781 (N_1781,In_1179,N_1430);
or U1782 (N_1782,In_569,N_383);
and U1783 (N_1783,N_1347,In_723);
nand U1784 (N_1784,N_885,N_1495);
nor U1785 (N_1785,N_1482,N_1214);
nor U1786 (N_1786,N_1483,N_1215);
and U1787 (N_1787,N_1590,N_1491);
or U1788 (N_1788,N_1246,In_301);
nand U1789 (N_1789,N_1179,N_1161);
or U1790 (N_1790,In_902,N_1508);
nor U1791 (N_1791,N_1018,In_393);
and U1792 (N_1792,In_2386,In_1773);
or U1793 (N_1793,N_121,In_1185);
xor U1794 (N_1794,N_1454,N_1288);
or U1795 (N_1795,N_1502,N_260);
nand U1796 (N_1796,N_1174,In_1867);
nor U1797 (N_1797,In_2452,N_1197);
xnor U1798 (N_1798,N_1520,N_554);
xor U1799 (N_1799,N_1364,N_852);
and U1800 (N_1800,N_1612,N_161);
nor U1801 (N_1801,In_2168,N_1223);
nand U1802 (N_1802,N_1667,N_1643);
or U1803 (N_1803,In_1396,In_1206);
and U1804 (N_1804,N_1725,N_1467);
nor U1805 (N_1805,N_1266,N_212);
nand U1806 (N_1806,In_2182,N_1631);
xor U1807 (N_1807,N_1440,N_1555);
and U1808 (N_1808,N_156,N_1764);
nand U1809 (N_1809,N_1396,In_46);
xnor U1810 (N_1810,N_324,N_1301);
or U1811 (N_1811,N_1575,N_1649);
xnor U1812 (N_1812,In_1046,In_1815);
nand U1813 (N_1813,In_181,N_1249);
nand U1814 (N_1814,N_1453,N_1012);
nor U1815 (N_1815,In_1483,N_1460);
or U1816 (N_1816,N_1278,In_2176);
nor U1817 (N_1817,N_1657,N_1624);
or U1818 (N_1818,N_1781,N_990);
nand U1819 (N_1819,N_1515,N_1711);
nor U1820 (N_1820,In_2311,N_1784);
nor U1821 (N_1821,N_1519,N_1768);
xnor U1822 (N_1822,N_1618,N_1292);
and U1823 (N_1823,N_1497,In_1831);
nand U1824 (N_1824,N_346,N_1478);
nor U1825 (N_1825,In_1958,N_1345);
and U1826 (N_1826,N_1611,N_1602);
xor U1827 (N_1827,N_633,In_55);
xnor U1828 (N_1828,N_1576,In_2103);
or U1829 (N_1829,N_1196,N_466);
xor U1830 (N_1830,N_1264,N_1320);
nor U1831 (N_1831,N_1772,N_311);
xor U1832 (N_1832,N_1107,N_1539);
xor U1833 (N_1833,N_1673,In_1296);
or U1834 (N_1834,N_1713,N_1786);
and U1835 (N_1835,In_932,In_1895);
and U1836 (N_1836,In_2353,N_1280);
and U1837 (N_1837,N_560,N_561);
and U1838 (N_1838,N_1766,N_1701);
or U1839 (N_1839,In_74,N_1476);
nor U1840 (N_1840,N_1728,N_1626);
nor U1841 (N_1841,In_1327,N_1668);
and U1842 (N_1842,In_2018,N_1406);
or U1843 (N_1843,N_1450,N_1684);
or U1844 (N_1844,N_1734,N_1094);
nand U1845 (N_1845,N_1282,In_419);
nand U1846 (N_1846,N_1407,N_1294);
xor U1847 (N_1847,N_1399,In_644);
or U1848 (N_1848,N_1553,N_1736);
or U1849 (N_1849,N_1299,N_588);
nor U1850 (N_1850,N_1295,N_434);
or U1851 (N_1851,In_1731,In_2402);
or U1852 (N_1852,N_1662,N_1600);
or U1853 (N_1853,In_2493,In_1004);
and U1854 (N_1854,In_2316,N_264);
or U1855 (N_1855,In_2315,N_1746);
or U1856 (N_1856,N_925,N_1201);
nand U1857 (N_1857,N_1194,N_1623);
nor U1858 (N_1858,N_866,N_1375);
xor U1859 (N_1859,N_1202,N_1790);
or U1860 (N_1860,N_1400,N_1411);
and U1861 (N_1861,N_1177,N_1639);
xor U1862 (N_1862,N_1615,In_2);
or U1863 (N_1863,In_276,N_1774);
and U1864 (N_1864,N_1691,N_1743);
or U1865 (N_1865,N_1740,N_1710);
nand U1866 (N_1866,N_1608,N_1752);
nand U1867 (N_1867,In_1697,N_1573);
nand U1868 (N_1868,In_1388,N_1186);
xnor U1869 (N_1869,N_619,In_1978);
xnor U1870 (N_1870,N_1750,N_1007);
or U1871 (N_1871,In_777,N_842);
nand U1872 (N_1872,In_2234,N_1756);
nand U1873 (N_1873,N_1592,N_1049);
or U1874 (N_1874,In_706,N_924);
and U1875 (N_1875,N_1629,N_1598);
and U1876 (N_1876,N_1579,N_1744);
nand U1877 (N_1877,In_599,N_1016);
nand U1878 (N_1878,N_1408,N_1134);
and U1879 (N_1879,N_512,In_1032);
xnor U1880 (N_1880,In_665,N_387);
or U1881 (N_1881,N_1686,N_233);
or U1882 (N_1882,In_1577,N_1473);
nor U1883 (N_1883,N_1696,In_2375);
nor U1884 (N_1884,In_45,N_1661);
xnor U1885 (N_1885,N_1745,N_410);
nor U1886 (N_1886,N_1390,N_1698);
and U1887 (N_1887,N_1316,N_778);
nand U1888 (N_1888,N_1616,N_741);
and U1889 (N_1889,N_1619,In_1973);
nand U1890 (N_1890,In_1361,In_564);
nand U1891 (N_1891,N_1666,N_816);
xnor U1892 (N_1892,N_1505,N_1613);
xor U1893 (N_1893,N_688,N_793);
or U1894 (N_1894,In_325,N_1401);
xor U1895 (N_1895,N_1642,N_416);
and U1896 (N_1896,In_541,N_1271);
or U1897 (N_1897,N_231,In_1793);
nor U1898 (N_1898,N_1098,N_1106);
or U1899 (N_1899,N_642,In_158);
nand U1900 (N_1900,In_2205,N_1352);
and U1901 (N_1901,N_1682,In_172);
nand U1902 (N_1902,N_821,In_178);
and U1903 (N_1903,In_1788,N_1640);
xnor U1904 (N_1904,N_1383,N_1254);
and U1905 (N_1905,N_1233,N_1);
xnor U1906 (N_1906,N_625,N_881);
xor U1907 (N_1907,N_853,N_336);
or U1908 (N_1908,N_491,N_1654);
and U1909 (N_1909,N_1683,In_77);
or U1910 (N_1910,In_1270,N_1751);
and U1911 (N_1911,N_1718,N_1798);
or U1912 (N_1912,N_1672,N_1788);
nand U1913 (N_1913,N_939,N_1564);
nand U1914 (N_1914,In_2457,N_1119);
and U1915 (N_1915,N_216,In_570);
and U1916 (N_1916,N_882,In_1176);
and U1917 (N_1917,N_1704,N_1152);
xor U1918 (N_1918,N_1537,N_1477);
xor U1919 (N_1919,N_1306,In_2062);
nor U1920 (N_1920,In_71,N_1690);
nand U1921 (N_1921,N_1597,N_1601);
or U1922 (N_1922,N_1605,N_1634);
nor U1923 (N_1923,In_842,N_1651);
or U1924 (N_1924,N_1109,N_1444);
or U1925 (N_1925,N_1606,N_1349);
or U1926 (N_1926,N_766,N_1331);
or U1927 (N_1927,In_2298,N_697);
nor U1928 (N_1928,In_206,N_8);
nand U1929 (N_1929,N_563,N_1235);
or U1930 (N_1930,N_1245,N_1426);
nand U1931 (N_1931,In_832,N_1127);
or U1932 (N_1932,N_1628,In_1054);
nand U1933 (N_1933,N_1070,N_1547);
nor U1934 (N_1934,N_1211,N_1436);
nand U1935 (N_1935,In_1710,N_1724);
xor U1936 (N_1936,N_1636,N_1304);
and U1937 (N_1937,N_1765,In_41);
xor U1938 (N_1938,N_405,N_1569);
or U1939 (N_1939,N_1614,N_1748);
or U1940 (N_1940,N_1534,N_1117);
xor U1941 (N_1941,N_1314,N_1087);
or U1942 (N_1942,N_1775,N_1737);
or U1943 (N_1943,N_1785,N_1595);
or U1944 (N_1944,N_1225,N_1168);
and U1945 (N_1945,In_2122,N_205);
nand U1946 (N_1946,N_1342,N_287);
and U1947 (N_1947,In_88,N_1144);
xnor U1948 (N_1948,N_1648,N_420);
and U1949 (N_1949,N_1501,N_296);
xor U1950 (N_1950,In_1893,In_2145);
xnor U1951 (N_1951,In_614,N_854);
nand U1952 (N_1952,N_916,In_1945);
nand U1953 (N_1953,N_953,N_1759);
nor U1954 (N_1954,N_1796,N_1685);
nand U1955 (N_1955,In_1300,N_1599);
or U1956 (N_1956,N_1580,N_1617);
xnor U1957 (N_1957,In_32,N_716);
and U1958 (N_1958,N_829,N_995);
and U1959 (N_1959,In_1813,N_1675);
nor U1960 (N_1960,In_820,N_472);
xnor U1961 (N_1961,In_1034,In_1083);
nor U1962 (N_1962,N_1723,In_1132);
nor U1963 (N_1963,N_1604,N_1659);
nand U1964 (N_1964,N_1753,N_1633);
or U1965 (N_1965,N_1492,N_1514);
nor U1966 (N_1966,N_435,N_1536);
xnor U1967 (N_1967,N_1484,In_1329);
xor U1968 (N_1968,N_1365,N_1665);
nand U1969 (N_1969,N_1663,In_134);
or U1970 (N_1970,N_811,In_1897);
and U1971 (N_1971,N_1767,N_1762);
or U1972 (N_1972,N_1067,N_1758);
xnor U1973 (N_1973,In_1260,In_709);
nor U1974 (N_1974,N_1496,N_373);
nand U1975 (N_1975,N_844,In_813);
and U1976 (N_1976,In_1810,N_1780);
or U1977 (N_1977,In_593,N_1403);
nand U1978 (N_1978,N_1707,In_538);
xor U1979 (N_1979,N_1647,N_412);
xnor U1980 (N_1980,N_1251,N_1283);
or U1981 (N_1981,N_1658,In_931);
and U1982 (N_1982,N_1366,N_932);
xnor U1983 (N_1983,N_1486,N_1587);
xnor U1984 (N_1984,N_1621,N_1709);
xnor U1985 (N_1985,N_255,In_236);
xnor U1986 (N_1986,N_1232,N_806);
nand U1987 (N_1987,N_1326,In_1730);
nand U1988 (N_1988,N_1795,N_1185);
and U1989 (N_1989,N_1637,N_1689);
xnor U1990 (N_1990,N_1038,N_1479);
nor U1991 (N_1991,In_1013,In_1584);
xnor U1992 (N_1992,N_9,In_887);
and U1993 (N_1993,N_1726,In_357);
nand U1994 (N_1994,N_441,N_377);
or U1995 (N_1995,N_1763,N_934);
xnor U1996 (N_1996,In_475,N_897);
or U1997 (N_1997,N_1791,N_685);
nor U1998 (N_1998,N_1669,N_952);
or U1999 (N_1999,N_1676,N_1171);
nor U2000 (N_2000,N_1693,N_1797);
nand U2001 (N_2001,N_1153,N_1848);
xnor U2002 (N_2002,N_1039,N_1895);
nand U2003 (N_2003,N_1439,N_1920);
xor U2004 (N_2004,N_1923,N_1341);
nand U2005 (N_2005,N_1937,In_1898);
nand U2006 (N_2006,N_1993,N_1705);
nand U2007 (N_2007,N_229,N_1972);
nor U2008 (N_2008,In_1824,N_1695);
nor U2009 (N_2009,N_1703,N_1854);
xnor U2010 (N_2010,N_1392,N_1915);
nand U2011 (N_2011,N_1581,N_222);
nand U2012 (N_2012,N_1646,N_1880);
and U2013 (N_2013,N_1858,N_1459);
and U2014 (N_2014,N_1200,N_1842);
or U2015 (N_2015,N_1868,N_1828);
and U2016 (N_2016,In_946,N_1967);
and U2017 (N_2017,N_1894,N_1956);
nor U2018 (N_2018,N_1979,N_1716);
nand U2019 (N_2019,N_845,N_1997);
xor U2020 (N_2020,N_1670,N_1429);
nand U2021 (N_2021,N_1638,N_137);
or U2022 (N_2022,N_1073,N_1903);
xor U2023 (N_2023,N_1870,N_1917);
and U2024 (N_2024,N_1813,N_580);
or U2025 (N_2025,N_624,N_1001);
or U2026 (N_2026,N_1156,In_381);
nand U2027 (N_2027,In_1663,N_1988);
nand U2028 (N_2028,N_1545,N_1964);
or U2029 (N_2029,N_996,N_1462);
or U2030 (N_2030,N_1829,N_1607);
or U2031 (N_2031,N_1538,N_1465);
or U2032 (N_2032,N_1122,N_1980);
xor U2033 (N_2033,N_1966,N_1660);
xor U2034 (N_2034,N_1949,N_523);
nand U2035 (N_2035,N_1991,N_94);
or U2036 (N_2036,N_1945,N_985);
and U2037 (N_2037,N_1717,N_1700);
nor U2038 (N_2038,In_845,In_770);
xor U2039 (N_2039,N_1692,N_1749);
or U2040 (N_2040,N_1632,N_1578);
or U2041 (N_2041,N_1986,In_72);
nand U2042 (N_2042,In_92,N_1906);
nand U2043 (N_2043,N_1973,N_1912);
or U2044 (N_2044,N_1897,N_691);
or U2045 (N_2045,In_1162,N_689);
nor U2046 (N_2046,N_1517,N_1485);
xnor U2047 (N_2047,N_1719,N_1951);
and U2048 (N_2048,N_1708,N_1414);
and U2049 (N_2049,N_1851,In_1395);
xor U2050 (N_2050,N_1856,N_1714);
nand U2051 (N_2051,N_1867,N_1933);
and U2052 (N_2052,N_1812,N_1839);
or U2053 (N_2053,N_1096,N_1489);
nand U2054 (N_2054,N_1747,In_2065);
and U2055 (N_2055,N_1776,N_1397);
nand U2056 (N_2056,N_1926,N_1924);
nand U2057 (N_2057,N_1559,N_1885);
xnor U2058 (N_2058,N_1802,N_1855);
nand U2059 (N_2059,N_978,N_1977);
nor U2060 (N_2060,In_808,N_1849);
xnor U2061 (N_2061,N_1876,In_2409);
and U2062 (N_2062,N_1582,N_1963);
nor U2063 (N_2063,In_1262,N_1907);
and U2064 (N_2064,N_1861,N_1527);
or U2065 (N_2065,N_1981,N_1510);
xnor U2066 (N_2066,N_545,N_1050);
and U2067 (N_2067,N_1422,N_1948);
nand U2068 (N_2068,N_1799,N_309);
and U2069 (N_2069,N_1892,N_1427);
nor U2070 (N_2070,N_1841,N_1878);
xor U2071 (N_2071,N_1845,N_1875);
nand U2072 (N_2072,In_2278,N_1938);
nand U2073 (N_2073,N_1805,N_1139);
nor U2074 (N_2074,N_1941,N_37);
xor U2075 (N_2075,N_1609,N_1687);
nand U2076 (N_2076,N_487,N_1896);
nor U2077 (N_2077,N_1884,N_1729);
or U2078 (N_2078,N_1853,N_1739);
nor U2079 (N_2079,N_769,N_1889);
and U2080 (N_2080,N_1792,N_1819);
xnor U2081 (N_2081,In_1439,N_1241);
or U2082 (N_2082,In_713,N_1838);
nor U2083 (N_2083,N_1417,N_1732);
or U2084 (N_2084,N_1874,N_1866);
or U2085 (N_2085,In_2265,N_1857);
and U2086 (N_2086,N_1432,N_1825);
and U2087 (N_2087,In_2252,N_1140);
xnor U2088 (N_2088,N_1850,N_1099);
xor U2089 (N_2089,In_2319,N_1760);
or U2090 (N_2090,N_103,N_1904);
xor U2091 (N_2091,N_1984,N_1699);
xnor U2092 (N_2092,N_1770,N_1793);
and U2093 (N_2093,N_1550,N_1821);
nor U2094 (N_2094,N_1566,N_1911);
nand U2095 (N_2095,N_1773,In_2337);
xor U2096 (N_2096,N_1914,N_1466);
nor U2097 (N_2097,N_1542,N_1733);
nor U2098 (N_2098,N_1971,N_1778);
and U2099 (N_2099,N_1859,N_1931);
nand U2100 (N_2100,N_1830,N_1843);
nand U2101 (N_2101,N_1893,N_1881);
and U2102 (N_2102,N_1910,N_1735);
xor U2103 (N_2103,N_1138,N_1810);
or U2104 (N_2104,N_1864,N_942);
nor U2105 (N_2105,N_1916,N_1644);
xnor U2106 (N_2106,N_1268,N_1706);
xnor U2107 (N_2107,N_1742,N_1952);
nand U2108 (N_2108,N_1782,N_1877);
and U2109 (N_2109,N_1627,N_837);
xor U2110 (N_2110,N_99,N_1809);
and U2111 (N_2111,In_383,N_1243);
nor U2112 (N_2112,N_1902,N_682);
nand U2113 (N_2113,In_779,N_975);
nand U2114 (N_2114,In_2056,N_1814);
nand U2115 (N_2115,N_68,N_1727);
nand U2116 (N_2116,N_1721,N_1832);
nand U2117 (N_2117,N_863,N_1455);
and U2118 (N_2118,N_1824,N_1521);
or U2119 (N_2119,N_1800,N_1899);
and U2120 (N_2120,N_1831,N_1970);
or U2121 (N_2121,N_1359,N_1652);
nand U2122 (N_2122,N_1987,N_1448);
and U2123 (N_2123,N_1656,In_1844);
or U2124 (N_2124,N_1741,In_2017);
and U2125 (N_2125,N_1930,N_1720);
and U2126 (N_2126,N_1905,N_1887);
nand U2127 (N_2127,N_1594,N_1990);
nand U2128 (N_2128,N_1958,N_1816);
nor U2129 (N_2129,N_1574,N_1653);
or U2130 (N_2130,N_424,N_1908);
xor U2131 (N_2131,In_1782,N_1561);
xnor U2132 (N_2132,N_1837,N_1900);
nand U2133 (N_2133,N_1840,N_1818);
xnor U2134 (N_2134,N_1962,N_1531);
nand U2135 (N_2135,N_1994,N_1421);
nor U2136 (N_2136,In_585,N_1942);
or U2137 (N_2137,N_1974,N_1940);
xor U2138 (N_2138,In_285,In_1674);
and U2139 (N_2139,N_671,In_1537);
nor U2140 (N_2140,In_2060,N_1808);
and U2141 (N_2141,In_2055,N_1833);
nor U2142 (N_2142,In_1060,N_1622);
nand U2143 (N_2143,N_1803,N_1674);
and U2144 (N_2144,N_1562,N_1655);
xnor U2145 (N_2145,N_1688,N_1757);
xnor U2146 (N_2146,N_1955,N_1935);
nor U2147 (N_2147,N_1925,N_1969);
or U2148 (N_2148,N_1540,N_1960);
nand U2149 (N_2149,N_248,In_133);
nand U2150 (N_2150,N_1730,N_1789);
and U2151 (N_2151,N_1806,N_1978);
or U2152 (N_2152,N_1548,In_1754);
xnor U2153 (N_2153,N_1815,N_1603);
and U2154 (N_2154,N_855,N_1256);
xor U2155 (N_2155,N_1625,N_1712);
or U2156 (N_2156,N_1481,In_1962);
xnor U2157 (N_2157,N_1879,N_1823);
nor U2158 (N_2158,N_1424,N_1834);
nand U2159 (N_2159,In_2351,N_1883);
xnor U2160 (N_2160,N_1355,N_1431);
nand U2161 (N_2161,N_1976,N_1811);
and U2162 (N_2162,N_1650,N_1836);
or U2163 (N_2163,N_1865,N_839);
and U2164 (N_2164,N_1999,N_1961);
nor U2165 (N_2165,N_1909,N_1996);
and U2166 (N_2166,N_617,N_1433);
or U2167 (N_2167,N_1928,N_1671);
xor U2168 (N_2168,N_918,N_1913);
nand U2169 (N_2169,N_1265,N_1532);
or U2170 (N_2170,N_830,N_1947);
nor U2171 (N_2171,N_1769,N_1738);
and U2172 (N_2172,N_1939,N_1968);
nand U2173 (N_2173,N_1965,N_768);
xnor U2174 (N_2174,N_1959,N_496);
nor U2175 (N_2175,N_1620,N_1694);
nor U2176 (N_2176,N_1847,In_1540);
and U2177 (N_2177,N_1863,N_1677);
nand U2178 (N_2178,N_1954,N_1957);
and U2179 (N_2179,N_1641,N_1860);
and U2180 (N_2180,N_1558,N_961);
xor U2181 (N_2181,In_109,N_1804);
or U2182 (N_2182,In_1716,N_1898);
and U2183 (N_2183,N_1513,N_1890);
nand U2184 (N_2184,N_60,N_1529);
xor U2185 (N_2185,In_962,N_1681);
xnor U2186 (N_2186,In_2049,In_2228);
xnor U2187 (N_2187,N_1310,N_1771);
nand U2188 (N_2188,In_765,N_1715);
xor U2189 (N_2189,N_1503,N_1754);
nor U2190 (N_2190,In_407,N_1918);
xnor U2191 (N_2191,N_449,N_1995);
or U2192 (N_2192,N_1794,N_1458);
or U2193 (N_2193,N_1932,N_1801);
nor U2194 (N_2194,N_1755,N_448);
xor U2195 (N_2195,N_1946,N_1852);
nor U2196 (N_2196,N_1927,In_2063);
nand U2197 (N_2197,In_1662,N_1846);
or U2198 (N_2198,N_1871,N_461);
and U2199 (N_2199,N_967,N_850);
nand U2200 (N_2200,N_2039,N_2084);
nor U2201 (N_2201,N_2165,N_2027);
nor U2202 (N_2202,N_1998,N_2146);
or U2203 (N_2203,N_2154,N_1787);
nor U2204 (N_2204,N_2003,N_2071);
or U2205 (N_2205,N_2096,N_2133);
nor U2206 (N_2206,N_2193,N_2016);
or U2207 (N_2207,N_2194,N_2181);
nand U2208 (N_2208,N_2189,N_2175);
xnor U2209 (N_2209,N_1817,N_2184);
or U2210 (N_2210,N_2017,N_2088);
nand U2211 (N_2211,N_2187,N_356);
nand U2212 (N_2212,N_2191,N_2123);
and U2213 (N_2213,N_2002,In_814);
or U2214 (N_2214,N_1402,N_2135);
or U2215 (N_2215,N_2035,N_2190);
nand U2216 (N_2216,N_56,In_312);
xnor U2217 (N_2217,N_2049,N_861);
nor U2218 (N_2218,N_849,N_2130);
xnor U2219 (N_2219,N_2060,N_1807);
nand U2220 (N_2220,N_956,N_2119);
or U2221 (N_2221,N_2058,N_2050);
nor U2222 (N_2222,N_2083,N_1731);
nor U2223 (N_2223,In_2320,N_1872);
xnor U2224 (N_2224,N_2104,N_2177);
nand U2225 (N_2225,N_2073,In_1360);
and U2226 (N_2226,N_2033,N_2167);
xor U2227 (N_2227,N_2069,N_2090);
xor U2228 (N_2228,N_2009,N_2155);
xor U2229 (N_2229,N_2005,N_2097);
nor U2230 (N_2230,N_2185,N_2140);
or U2231 (N_2231,N_1509,N_2172);
nor U2232 (N_2232,N_2196,N_2080);
nand U2233 (N_2233,N_2137,N_2077);
or U2234 (N_2234,N_2007,N_2173);
or U2235 (N_2235,N_2015,N_1950);
or U2236 (N_2236,N_1680,N_2106);
or U2237 (N_2237,N_1325,N_2041);
or U2238 (N_2238,N_2149,N_2051);
xor U2239 (N_2239,N_2108,N_2101);
or U2240 (N_2240,N_1610,N_2112);
and U2241 (N_2241,N_2004,N_2166);
and U2242 (N_2242,N_2110,N_907);
or U2243 (N_2243,N_2078,N_2021);
xnor U2244 (N_2244,N_2195,N_1944);
or U2245 (N_2245,N_1697,N_1983);
or U2246 (N_2246,N_2019,N_1886);
or U2247 (N_2247,N_2114,N_1953);
or U2248 (N_2248,N_2075,N_2192);
or U2249 (N_2249,N_797,N_2043);
nand U2250 (N_2250,N_2199,N_1311);
nor U2251 (N_2251,N_2001,N_2044);
or U2252 (N_2252,N_2063,N_1936);
or U2253 (N_2253,N_2030,N_2098);
nor U2254 (N_2254,N_501,N_2126);
xnor U2255 (N_2255,N_2198,N_2006);
nor U2256 (N_2256,In_1222,N_2168);
xor U2257 (N_2257,N_2047,N_2131);
and U2258 (N_2258,N_1888,N_2176);
xnor U2259 (N_2259,N_1982,N_2120);
and U2260 (N_2260,N_1354,N_1635);
nor U2261 (N_2261,N_2170,N_1862);
xor U2262 (N_2262,N_2145,N_1586);
nand U2263 (N_2263,N_1761,N_2152);
and U2264 (N_2264,N_2142,N_2139);
and U2265 (N_2265,N_1820,N_2150);
nor U2266 (N_2266,N_1490,N_2138);
or U2267 (N_2267,N_1678,N_2086);
nor U2268 (N_2268,N_590,N_2032);
nand U2269 (N_2269,N_2031,N_706);
or U2270 (N_2270,N_1435,N_2188);
and U2271 (N_2271,N_2113,N_1488);
and U2272 (N_2272,N_2111,N_1071);
and U2273 (N_2273,In_745,N_2008);
and U2274 (N_2274,N_2029,N_1989);
and U2275 (N_2275,N_1645,N_725);
or U2276 (N_2276,N_2055,N_2020);
nand U2277 (N_2277,N_1630,N_2100);
nor U2278 (N_2278,N_2057,N_2143);
nor U2279 (N_2279,N_2064,N_1919);
nor U2280 (N_2280,N_2085,N_2115);
nand U2281 (N_2281,N_1922,N_2136);
and U2282 (N_2282,N_2014,N_1869);
or U2283 (N_2283,N_1571,N_2182);
and U2284 (N_2284,N_1259,N_2065);
nand U2285 (N_2285,N_1244,N_2067);
and U2286 (N_2286,N_2128,N_904);
or U2287 (N_2287,N_675,N_2162);
xnor U2288 (N_2288,N_2107,N_2070);
nor U2289 (N_2289,N_1702,N_2116);
and U2290 (N_2290,N_2074,N_2072);
nand U2291 (N_2291,N_2186,N_2062);
xor U2292 (N_2292,In_1291,N_2164);
nor U2293 (N_2293,N_2151,N_2028);
nor U2294 (N_2294,N_2183,N_2056);
nand U2295 (N_2295,N_1929,N_2091);
and U2296 (N_2296,N_2180,N_1394);
nor U2297 (N_2297,N_1835,N_2082);
or U2298 (N_2298,N_2054,N_1934);
xor U2299 (N_2299,N_2109,N_1975);
xnor U2300 (N_2300,N_2025,N_2171);
or U2301 (N_2301,N_2079,N_1779);
nand U2302 (N_2302,N_2037,N_2105);
xor U2303 (N_2303,N_2157,N_2087);
xor U2304 (N_2304,In_451,N_1992);
nor U2305 (N_2305,N_1985,N_2178);
and U2306 (N_2306,N_2034,N_2144);
nor U2307 (N_2307,N_2132,N_1844);
and U2308 (N_2308,N_2048,N_2129);
xnor U2309 (N_2309,N_2024,N_1679);
xnor U2310 (N_2310,N_1827,N_2068);
or U2311 (N_2311,N_2169,In_558);
nor U2312 (N_2312,N_1826,N_495);
and U2313 (N_2313,N_1475,N_2125);
nand U2314 (N_2314,N_1722,N_2158);
xnor U2315 (N_2315,N_2042,N_2038);
nand U2316 (N_2316,N_2018,In_786);
nor U2317 (N_2317,N_1783,N_2121);
xnor U2318 (N_2318,N_2197,N_2141);
nand U2319 (N_2319,N_2023,N_2012);
nor U2320 (N_2320,N_2163,In_2028);
nand U2321 (N_2321,N_2093,N_2174);
and U2322 (N_2322,N_1006,N_2026);
and U2323 (N_2323,In_284,N_1882);
xnor U2324 (N_2324,N_2103,N_1822);
or U2325 (N_2325,N_2000,N_2127);
or U2326 (N_2326,N_2095,N_2122);
nor U2327 (N_2327,N_2053,N_2179);
nor U2328 (N_2328,N_2153,N_1901);
and U2329 (N_2329,N_2052,N_2092);
nand U2330 (N_2330,N_2094,N_2118);
or U2331 (N_2331,N_2059,N_1921);
or U2332 (N_2332,N_1943,N_2066);
and U2333 (N_2333,N_2081,In_2128);
and U2334 (N_2334,N_1546,N_2160);
or U2335 (N_2335,N_2013,N_2156);
nand U2336 (N_2336,N_2046,N_991);
xor U2337 (N_2337,N_1777,N_2159);
or U2338 (N_2338,N_2117,N_2036);
or U2339 (N_2339,N_1873,N_2134);
nand U2340 (N_2340,N_1891,N_2124);
and U2341 (N_2341,N_2148,N_2040);
nand U2342 (N_2342,N_2011,N_2045);
nor U2343 (N_2343,N_593,N_1335);
xor U2344 (N_2344,N_2102,N_2161);
nor U2345 (N_2345,N_1664,N_2061);
and U2346 (N_2346,N_2099,N_2147);
or U2347 (N_2347,N_1110,N_2022);
nand U2348 (N_2348,N_2076,N_1267);
nand U2349 (N_2349,N_2010,N_2089);
xnor U2350 (N_2350,In_2320,N_1919);
xor U2351 (N_2351,N_904,N_2190);
nand U2352 (N_2352,N_2003,N_2093);
nand U2353 (N_2353,N_2088,N_1325);
and U2354 (N_2354,N_1664,N_1586);
and U2355 (N_2355,N_2194,N_1950);
nand U2356 (N_2356,N_2049,N_2168);
nand U2357 (N_2357,N_1982,N_2038);
and U2358 (N_2358,N_2067,N_2056);
or U2359 (N_2359,N_2089,N_2087);
xnor U2360 (N_2360,N_2142,N_2199);
nor U2361 (N_2361,N_2043,N_2038);
xnor U2362 (N_2362,N_2158,N_2068);
xnor U2363 (N_2363,N_2084,N_2126);
xnor U2364 (N_2364,N_2008,N_2093);
and U2365 (N_2365,N_501,N_2072);
and U2366 (N_2366,N_2199,N_2184);
and U2367 (N_2367,N_1919,N_2179);
or U2368 (N_2368,N_2140,N_1944);
nand U2369 (N_2369,N_2176,N_2113);
and U2370 (N_2370,N_2176,N_2064);
and U2371 (N_2371,N_904,N_1998);
and U2372 (N_2372,N_2165,N_1862);
nor U2373 (N_2373,N_1901,N_2024);
nand U2374 (N_2374,N_2044,N_861);
and U2375 (N_2375,N_2060,N_1929);
nand U2376 (N_2376,N_1822,N_2097);
nor U2377 (N_2377,N_2084,N_2041);
nand U2378 (N_2378,N_2197,N_1820);
and U2379 (N_2379,N_2096,N_2094);
nor U2380 (N_2380,N_2116,N_2158);
and U2381 (N_2381,N_2015,N_2095);
or U2382 (N_2382,N_1998,N_2165);
nand U2383 (N_2383,N_2159,N_2103);
nand U2384 (N_2384,N_2132,N_1731);
nand U2385 (N_2385,N_1869,N_1827);
nand U2386 (N_2386,N_2147,N_2092);
xnor U2387 (N_2387,In_284,N_2126);
nand U2388 (N_2388,N_2072,N_2037);
and U2389 (N_2389,N_1335,N_2191);
nand U2390 (N_2390,N_1936,N_1680);
or U2391 (N_2391,N_1827,N_501);
xnor U2392 (N_2392,N_1645,N_2154);
or U2393 (N_2393,N_2039,N_1901);
or U2394 (N_2394,In_1222,N_1777);
or U2395 (N_2395,N_1488,N_2001);
nand U2396 (N_2396,N_2168,N_2036);
xor U2397 (N_2397,N_2011,N_2091);
or U2398 (N_2398,N_2085,In_2320);
xnor U2399 (N_2399,N_2033,N_1944);
or U2400 (N_2400,N_2283,N_2366);
and U2401 (N_2401,N_2386,N_2271);
or U2402 (N_2402,N_2258,N_2262);
nand U2403 (N_2403,N_2268,N_2310);
and U2404 (N_2404,N_2218,N_2249);
nor U2405 (N_2405,N_2321,N_2213);
nor U2406 (N_2406,N_2395,N_2375);
nor U2407 (N_2407,N_2287,N_2254);
nor U2408 (N_2408,N_2306,N_2270);
nor U2409 (N_2409,N_2320,N_2274);
or U2410 (N_2410,N_2316,N_2233);
and U2411 (N_2411,N_2279,N_2288);
nor U2412 (N_2412,N_2391,N_2383);
nand U2413 (N_2413,N_2337,N_2392);
and U2414 (N_2414,N_2236,N_2245);
xor U2415 (N_2415,N_2368,N_2294);
xnor U2416 (N_2416,N_2393,N_2250);
xor U2417 (N_2417,N_2353,N_2315);
nand U2418 (N_2418,N_2220,N_2342);
nor U2419 (N_2419,N_2360,N_2277);
nor U2420 (N_2420,N_2215,N_2361);
and U2421 (N_2421,N_2272,N_2334);
nor U2422 (N_2422,N_2354,N_2370);
and U2423 (N_2423,N_2265,N_2255);
and U2424 (N_2424,N_2308,N_2327);
and U2425 (N_2425,N_2344,N_2292);
nor U2426 (N_2426,N_2303,N_2323);
nand U2427 (N_2427,N_2256,N_2318);
nand U2428 (N_2428,N_2253,N_2299);
xnor U2429 (N_2429,N_2244,N_2397);
or U2430 (N_2430,N_2248,N_2351);
xor U2431 (N_2431,N_2398,N_2309);
nand U2432 (N_2432,N_2227,N_2399);
or U2433 (N_2433,N_2359,N_2263);
or U2434 (N_2434,N_2210,N_2295);
or U2435 (N_2435,N_2385,N_2281);
nand U2436 (N_2436,N_2242,N_2211);
nand U2437 (N_2437,N_2269,N_2201);
or U2438 (N_2438,N_2203,N_2297);
and U2439 (N_2439,N_2300,N_2214);
xor U2440 (N_2440,N_2241,N_2280);
or U2441 (N_2441,N_2205,N_2243);
and U2442 (N_2442,N_2212,N_2276);
or U2443 (N_2443,N_2379,N_2330);
and U2444 (N_2444,N_2314,N_2208);
and U2445 (N_2445,N_2313,N_2225);
nor U2446 (N_2446,N_2356,N_2217);
or U2447 (N_2447,N_2260,N_2329);
or U2448 (N_2448,N_2322,N_2289);
and U2449 (N_2449,N_2264,N_2317);
nor U2450 (N_2450,N_2387,N_2349);
nor U2451 (N_2451,N_2219,N_2372);
or U2452 (N_2452,N_2257,N_2298);
nor U2453 (N_2453,N_2363,N_2305);
and U2454 (N_2454,N_2286,N_2296);
nand U2455 (N_2455,N_2350,N_2396);
nor U2456 (N_2456,N_2346,N_2369);
and U2457 (N_2457,N_2378,N_2340);
or U2458 (N_2458,N_2324,N_2348);
or U2459 (N_2459,N_2278,N_2240);
nor U2460 (N_2460,N_2332,N_2234);
xor U2461 (N_2461,N_2216,N_2358);
nand U2462 (N_2462,N_2222,N_2290);
xnor U2463 (N_2463,N_2252,N_2377);
and U2464 (N_2464,N_2311,N_2284);
nor U2465 (N_2465,N_2221,N_2293);
xnor U2466 (N_2466,N_2231,N_2237);
nand U2467 (N_2467,N_2376,N_2247);
nor U2468 (N_2468,N_2335,N_2206);
nand U2469 (N_2469,N_2246,N_2302);
or U2470 (N_2470,N_2235,N_2259);
or U2471 (N_2471,N_2204,N_2390);
nand U2472 (N_2472,N_2261,N_2336);
xor U2473 (N_2473,N_2338,N_2365);
or U2474 (N_2474,N_2364,N_2223);
xor U2475 (N_2475,N_2226,N_2239);
nand U2476 (N_2476,N_2251,N_2357);
and U2477 (N_2477,N_2267,N_2367);
nand U2478 (N_2478,N_2200,N_2238);
and U2479 (N_2479,N_2373,N_2394);
and U2480 (N_2480,N_2347,N_2333);
or U2481 (N_2481,N_2339,N_2266);
nor U2482 (N_2482,N_2312,N_2328);
nand U2483 (N_2483,N_2389,N_2343);
xnor U2484 (N_2484,N_2229,N_2362);
nand U2485 (N_2485,N_2352,N_2380);
or U2486 (N_2486,N_2374,N_2273);
and U2487 (N_2487,N_2291,N_2228);
or U2488 (N_2488,N_2388,N_2371);
or U2489 (N_2489,N_2355,N_2326);
or U2490 (N_2490,N_2209,N_2232);
nor U2491 (N_2491,N_2224,N_2382);
nor U2492 (N_2492,N_2304,N_2341);
nand U2493 (N_2493,N_2202,N_2230);
and U2494 (N_2494,N_2275,N_2345);
nand U2495 (N_2495,N_2384,N_2381);
xor U2496 (N_2496,N_2307,N_2331);
and U2497 (N_2497,N_2319,N_2282);
nand U2498 (N_2498,N_2285,N_2301);
nor U2499 (N_2499,N_2325,N_2207);
nand U2500 (N_2500,N_2376,N_2339);
nand U2501 (N_2501,N_2326,N_2324);
or U2502 (N_2502,N_2327,N_2250);
nand U2503 (N_2503,N_2253,N_2215);
nand U2504 (N_2504,N_2357,N_2303);
and U2505 (N_2505,N_2379,N_2345);
nor U2506 (N_2506,N_2216,N_2378);
nand U2507 (N_2507,N_2227,N_2395);
and U2508 (N_2508,N_2231,N_2352);
nand U2509 (N_2509,N_2324,N_2277);
nor U2510 (N_2510,N_2268,N_2291);
nor U2511 (N_2511,N_2223,N_2387);
or U2512 (N_2512,N_2376,N_2336);
and U2513 (N_2513,N_2226,N_2295);
nand U2514 (N_2514,N_2209,N_2301);
or U2515 (N_2515,N_2238,N_2346);
and U2516 (N_2516,N_2364,N_2235);
nor U2517 (N_2517,N_2298,N_2394);
xnor U2518 (N_2518,N_2272,N_2318);
and U2519 (N_2519,N_2266,N_2210);
nor U2520 (N_2520,N_2327,N_2388);
nand U2521 (N_2521,N_2260,N_2310);
and U2522 (N_2522,N_2359,N_2393);
and U2523 (N_2523,N_2257,N_2314);
xnor U2524 (N_2524,N_2323,N_2216);
nor U2525 (N_2525,N_2274,N_2397);
and U2526 (N_2526,N_2374,N_2202);
nor U2527 (N_2527,N_2263,N_2266);
xor U2528 (N_2528,N_2334,N_2309);
xnor U2529 (N_2529,N_2311,N_2382);
nand U2530 (N_2530,N_2281,N_2374);
and U2531 (N_2531,N_2297,N_2204);
nor U2532 (N_2532,N_2226,N_2257);
or U2533 (N_2533,N_2280,N_2335);
and U2534 (N_2534,N_2366,N_2398);
nand U2535 (N_2535,N_2214,N_2301);
nor U2536 (N_2536,N_2344,N_2367);
nand U2537 (N_2537,N_2256,N_2227);
nand U2538 (N_2538,N_2370,N_2387);
xnor U2539 (N_2539,N_2336,N_2241);
or U2540 (N_2540,N_2230,N_2290);
nor U2541 (N_2541,N_2327,N_2284);
xnor U2542 (N_2542,N_2261,N_2308);
or U2543 (N_2543,N_2247,N_2241);
xnor U2544 (N_2544,N_2364,N_2241);
and U2545 (N_2545,N_2247,N_2222);
xnor U2546 (N_2546,N_2276,N_2273);
and U2547 (N_2547,N_2289,N_2245);
xor U2548 (N_2548,N_2213,N_2364);
nor U2549 (N_2549,N_2382,N_2278);
xor U2550 (N_2550,N_2341,N_2324);
nor U2551 (N_2551,N_2320,N_2235);
xnor U2552 (N_2552,N_2294,N_2315);
nor U2553 (N_2553,N_2202,N_2385);
and U2554 (N_2554,N_2347,N_2204);
or U2555 (N_2555,N_2272,N_2325);
xor U2556 (N_2556,N_2213,N_2204);
and U2557 (N_2557,N_2292,N_2317);
nor U2558 (N_2558,N_2215,N_2228);
xor U2559 (N_2559,N_2381,N_2399);
and U2560 (N_2560,N_2341,N_2274);
nand U2561 (N_2561,N_2210,N_2373);
nor U2562 (N_2562,N_2386,N_2286);
nor U2563 (N_2563,N_2321,N_2334);
nor U2564 (N_2564,N_2217,N_2366);
xor U2565 (N_2565,N_2296,N_2270);
nand U2566 (N_2566,N_2259,N_2324);
and U2567 (N_2567,N_2214,N_2314);
or U2568 (N_2568,N_2353,N_2330);
xnor U2569 (N_2569,N_2303,N_2343);
and U2570 (N_2570,N_2259,N_2243);
nor U2571 (N_2571,N_2294,N_2299);
and U2572 (N_2572,N_2215,N_2218);
nor U2573 (N_2573,N_2351,N_2315);
xor U2574 (N_2574,N_2398,N_2323);
nand U2575 (N_2575,N_2245,N_2323);
nand U2576 (N_2576,N_2346,N_2215);
nor U2577 (N_2577,N_2269,N_2299);
nand U2578 (N_2578,N_2226,N_2212);
nand U2579 (N_2579,N_2210,N_2255);
or U2580 (N_2580,N_2273,N_2294);
or U2581 (N_2581,N_2356,N_2292);
nor U2582 (N_2582,N_2274,N_2254);
nand U2583 (N_2583,N_2267,N_2381);
nor U2584 (N_2584,N_2274,N_2217);
xnor U2585 (N_2585,N_2294,N_2364);
nor U2586 (N_2586,N_2221,N_2339);
nor U2587 (N_2587,N_2307,N_2209);
and U2588 (N_2588,N_2275,N_2386);
xor U2589 (N_2589,N_2212,N_2269);
nand U2590 (N_2590,N_2207,N_2200);
and U2591 (N_2591,N_2249,N_2352);
nor U2592 (N_2592,N_2315,N_2318);
xor U2593 (N_2593,N_2248,N_2266);
or U2594 (N_2594,N_2239,N_2235);
and U2595 (N_2595,N_2232,N_2267);
nand U2596 (N_2596,N_2360,N_2212);
nor U2597 (N_2597,N_2300,N_2362);
nand U2598 (N_2598,N_2389,N_2303);
nor U2599 (N_2599,N_2229,N_2347);
and U2600 (N_2600,N_2436,N_2523);
or U2601 (N_2601,N_2484,N_2576);
xor U2602 (N_2602,N_2459,N_2432);
xor U2603 (N_2603,N_2567,N_2411);
nor U2604 (N_2604,N_2513,N_2535);
nand U2605 (N_2605,N_2511,N_2497);
or U2606 (N_2606,N_2556,N_2549);
xor U2607 (N_2607,N_2444,N_2597);
nand U2608 (N_2608,N_2595,N_2572);
and U2609 (N_2609,N_2467,N_2435);
nor U2610 (N_2610,N_2558,N_2583);
xor U2611 (N_2611,N_2538,N_2580);
or U2612 (N_2612,N_2550,N_2562);
and U2613 (N_2613,N_2448,N_2500);
or U2614 (N_2614,N_2574,N_2417);
and U2615 (N_2615,N_2437,N_2494);
nand U2616 (N_2616,N_2464,N_2402);
and U2617 (N_2617,N_2489,N_2461);
nand U2618 (N_2618,N_2483,N_2468);
and U2619 (N_2619,N_2530,N_2531);
nor U2620 (N_2620,N_2554,N_2537);
nor U2621 (N_2621,N_2557,N_2462);
and U2622 (N_2622,N_2482,N_2487);
and U2623 (N_2623,N_2569,N_2443);
or U2624 (N_2624,N_2427,N_2424);
and U2625 (N_2625,N_2493,N_2454);
or U2626 (N_2626,N_2564,N_2519);
nand U2627 (N_2627,N_2582,N_2544);
xnor U2628 (N_2628,N_2496,N_2401);
nand U2629 (N_2629,N_2520,N_2423);
and U2630 (N_2630,N_2472,N_2490);
nand U2631 (N_2631,N_2488,N_2566);
nor U2632 (N_2632,N_2473,N_2452);
nand U2633 (N_2633,N_2475,N_2471);
nand U2634 (N_2634,N_2598,N_2503);
nand U2635 (N_2635,N_2455,N_2505);
nand U2636 (N_2636,N_2545,N_2457);
or U2637 (N_2637,N_2438,N_2413);
nor U2638 (N_2638,N_2477,N_2546);
nand U2639 (N_2639,N_2409,N_2529);
and U2640 (N_2640,N_2516,N_2465);
nand U2641 (N_2641,N_2495,N_2573);
or U2642 (N_2642,N_2585,N_2589);
nand U2643 (N_2643,N_2508,N_2577);
nor U2644 (N_2644,N_2446,N_2591);
nand U2645 (N_2645,N_2506,N_2414);
and U2646 (N_2646,N_2474,N_2415);
nand U2647 (N_2647,N_2479,N_2555);
and U2648 (N_2648,N_2400,N_2469);
xor U2649 (N_2649,N_2407,N_2594);
and U2650 (N_2650,N_2571,N_2560);
and U2651 (N_2651,N_2426,N_2451);
nor U2652 (N_2652,N_2463,N_2596);
nor U2653 (N_2653,N_2449,N_2552);
xor U2654 (N_2654,N_2532,N_2551);
nand U2655 (N_2655,N_2416,N_2460);
and U2656 (N_2656,N_2439,N_2581);
nand U2657 (N_2657,N_2445,N_2470);
or U2658 (N_2658,N_2434,N_2450);
nand U2659 (N_2659,N_2502,N_2534);
or U2660 (N_2660,N_2579,N_2515);
xnor U2661 (N_2661,N_2441,N_2425);
xor U2662 (N_2662,N_2447,N_2418);
nor U2663 (N_2663,N_2561,N_2584);
xor U2664 (N_2664,N_2476,N_2403);
xnor U2665 (N_2665,N_2547,N_2570);
nand U2666 (N_2666,N_2412,N_2420);
xnor U2667 (N_2667,N_2518,N_2599);
nor U2668 (N_2668,N_2406,N_2575);
nand U2669 (N_2669,N_2528,N_2428);
xnor U2670 (N_2670,N_2410,N_2499);
nor U2671 (N_2671,N_2404,N_2536);
or U2672 (N_2672,N_2512,N_2429);
xor U2673 (N_2673,N_2517,N_2480);
nand U2674 (N_2674,N_2501,N_2542);
and U2675 (N_2675,N_2478,N_2588);
nand U2676 (N_2676,N_2559,N_2543);
and U2677 (N_2677,N_2408,N_2548);
nand U2678 (N_2678,N_2458,N_2421);
nand U2679 (N_2679,N_2540,N_2533);
or U2680 (N_2680,N_2592,N_2525);
xnor U2681 (N_2681,N_2527,N_2422);
nand U2682 (N_2682,N_2586,N_2453);
or U2683 (N_2683,N_2553,N_2509);
nand U2684 (N_2684,N_2433,N_2442);
or U2685 (N_2685,N_2524,N_2431);
nand U2686 (N_2686,N_2440,N_2522);
and U2687 (N_2687,N_2578,N_2539);
nand U2688 (N_2688,N_2521,N_2430);
and U2689 (N_2689,N_2568,N_2466);
or U2690 (N_2690,N_2507,N_2514);
nand U2691 (N_2691,N_2481,N_2485);
xor U2692 (N_2692,N_2419,N_2565);
or U2693 (N_2693,N_2593,N_2405);
nand U2694 (N_2694,N_2541,N_2504);
nor U2695 (N_2695,N_2456,N_2510);
or U2696 (N_2696,N_2491,N_2498);
or U2697 (N_2697,N_2486,N_2526);
and U2698 (N_2698,N_2492,N_2590);
nand U2699 (N_2699,N_2563,N_2587);
nor U2700 (N_2700,N_2455,N_2521);
and U2701 (N_2701,N_2565,N_2599);
and U2702 (N_2702,N_2467,N_2492);
xor U2703 (N_2703,N_2577,N_2569);
nand U2704 (N_2704,N_2409,N_2540);
nand U2705 (N_2705,N_2436,N_2482);
xnor U2706 (N_2706,N_2441,N_2440);
and U2707 (N_2707,N_2593,N_2542);
nand U2708 (N_2708,N_2458,N_2467);
nor U2709 (N_2709,N_2568,N_2553);
xnor U2710 (N_2710,N_2504,N_2555);
and U2711 (N_2711,N_2568,N_2413);
xor U2712 (N_2712,N_2531,N_2566);
nor U2713 (N_2713,N_2473,N_2482);
xnor U2714 (N_2714,N_2401,N_2430);
nor U2715 (N_2715,N_2482,N_2508);
xnor U2716 (N_2716,N_2480,N_2587);
or U2717 (N_2717,N_2592,N_2585);
xor U2718 (N_2718,N_2570,N_2543);
nor U2719 (N_2719,N_2450,N_2590);
xnor U2720 (N_2720,N_2557,N_2592);
or U2721 (N_2721,N_2540,N_2588);
nand U2722 (N_2722,N_2596,N_2470);
xor U2723 (N_2723,N_2414,N_2478);
nand U2724 (N_2724,N_2540,N_2593);
nand U2725 (N_2725,N_2487,N_2410);
nor U2726 (N_2726,N_2440,N_2500);
and U2727 (N_2727,N_2477,N_2560);
xnor U2728 (N_2728,N_2458,N_2580);
and U2729 (N_2729,N_2432,N_2560);
xor U2730 (N_2730,N_2407,N_2512);
and U2731 (N_2731,N_2434,N_2533);
xnor U2732 (N_2732,N_2441,N_2487);
xnor U2733 (N_2733,N_2494,N_2452);
nor U2734 (N_2734,N_2402,N_2401);
nand U2735 (N_2735,N_2593,N_2407);
xor U2736 (N_2736,N_2477,N_2552);
xor U2737 (N_2737,N_2447,N_2445);
or U2738 (N_2738,N_2538,N_2577);
and U2739 (N_2739,N_2408,N_2509);
and U2740 (N_2740,N_2467,N_2597);
nor U2741 (N_2741,N_2490,N_2486);
or U2742 (N_2742,N_2480,N_2427);
and U2743 (N_2743,N_2555,N_2548);
xnor U2744 (N_2744,N_2533,N_2415);
nand U2745 (N_2745,N_2562,N_2450);
nand U2746 (N_2746,N_2465,N_2417);
nand U2747 (N_2747,N_2463,N_2503);
nand U2748 (N_2748,N_2441,N_2520);
xor U2749 (N_2749,N_2496,N_2423);
and U2750 (N_2750,N_2412,N_2465);
nand U2751 (N_2751,N_2433,N_2405);
or U2752 (N_2752,N_2536,N_2598);
and U2753 (N_2753,N_2493,N_2535);
nor U2754 (N_2754,N_2500,N_2446);
xor U2755 (N_2755,N_2500,N_2544);
nor U2756 (N_2756,N_2466,N_2440);
or U2757 (N_2757,N_2419,N_2545);
nand U2758 (N_2758,N_2421,N_2496);
or U2759 (N_2759,N_2411,N_2456);
or U2760 (N_2760,N_2537,N_2449);
or U2761 (N_2761,N_2409,N_2473);
or U2762 (N_2762,N_2585,N_2479);
nand U2763 (N_2763,N_2516,N_2571);
nor U2764 (N_2764,N_2497,N_2471);
xnor U2765 (N_2765,N_2459,N_2473);
or U2766 (N_2766,N_2462,N_2543);
and U2767 (N_2767,N_2424,N_2488);
or U2768 (N_2768,N_2592,N_2437);
and U2769 (N_2769,N_2449,N_2491);
and U2770 (N_2770,N_2535,N_2599);
nand U2771 (N_2771,N_2455,N_2553);
xnor U2772 (N_2772,N_2532,N_2580);
xor U2773 (N_2773,N_2473,N_2595);
nor U2774 (N_2774,N_2483,N_2459);
xnor U2775 (N_2775,N_2566,N_2471);
nor U2776 (N_2776,N_2509,N_2574);
and U2777 (N_2777,N_2571,N_2460);
nand U2778 (N_2778,N_2520,N_2471);
nor U2779 (N_2779,N_2443,N_2582);
nand U2780 (N_2780,N_2502,N_2437);
and U2781 (N_2781,N_2432,N_2566);
nand U2782 (N_2782,N_2414,N_2442);
or U2783 (N_2783,N_2417,N_2436);
xnor U2784 (N_2784,N_2455,N_2478);
nor U2785 (N_2785,N_2553,N_2567);
nand U2786 (N_2786,N_2520,N_2466);
or U2787 (N_2787,N_2563,N_2470);
nand U2788 (N_2788,N_2573,N_2568);
and U2789 (N_2789,N_2599,N_2428);
nand U2790 (N_2790,N_2482,N_2452);
nand U2791 (N_2791,N_2417,N_2443);
nand U2792 (N_2792,N_2496,N_2435);
xnor U2793 (N_2793,N_2496,N_2475);
nand U2794 (N_2794,N_2456,N_2579);
and U2795 (N_2795,N_2467,N_2502);
or U2796 (N_2796,N_2421,N_2485);
nand U2797 (N_2797,N_2436,N_2598);
nand U2798 (N_2798,N_2576,N_2489);
nand U2799 (N_2799,N_2474,N_2477);
nand U2800 (N_2800,N_2635,N_2662);
nor U2801 (N_2801,N_2748,N_2674);
xor U2802 (N_2802,N_2756,N_2622);
or U2803 (N_2803,N_2728,N_2755);
xnor U2804 (N_2804,N_2694,N_2619);
nor U2805 (N_2805,N_2772,N_2659);
xor U2806 (N_2806,N_2722,N_2610);
and U2807 (N_2807,N_2676,N_2734);
and U2808 (N_2808,N_2654,N_2727);
or U2809 (N_2809,N_2784,N_2679);
xor U2810 (N_2810,N_2758,N_2737);
and U2811 (N_2811,N_2718,N_2702);
nor U2812 (N_2812,N_2708,N_2765);
and U2813 (N_2813,N_2785,N_2740);
nand U2814 (N_2814,N_2751,N_2775);
or U2815 (N_2815,N_2717,N_2613);
xnor U2816 (N_2816,N_2744,N_2675);
xnor U2817 (N_2817,N_2642,N_2766);
nand U2818 (N_2818,N_2787,N_2617);
nor U2819 (N_2819,N_2652,N_2670);
xnor U2820 (N_2820,N_2738,N_2600);
nor U2821 (N_2821,N_2671,N_2754);
and U2822 (N_2822,N_2774,N_2649);
nand U2823 (N_2823,N_2624,N_2742);
nor U2824 (N_2824,N_2614,N_2672);
nor U2825 (N_2825,N_2690,N_2605);
and U2826 (N_2826,N_2630,N_2776);
and U2827 (N_2827,N_2777,N_2746);
xor U2828 (N_2828,N_2680,N_2745);
xor U2829 (N_2829,N_2608,N_2711);
nor U2830 (N_2830,N_2601,N_2645);
xnor U2831 (N_2831,N_2759,N_2706);
nand U2832 (N_2832,N_2730,N_2664);
and U2833 (N_2833,N_2701,N_2604);
nor U2834 (N_2834,N_2636,N_2696);
nand U2835 (N_2835,N_2697,N_2749);
nand U2836 (N_2836,N_2723,N_2692);
or U2837 (N_2837,N_2797,N_2793);
or U2838 (N_2838,N_2716,N_2733);
nor U2839 (N_2839,N_2673,N_2799);
nand U2840 (N_2840,N_2623,N_2705);
nand U2841 (N_2841,N_2731,N_2781);
nand U2842 (N_2842,N_2620,N_2648);
and U2843 (N_2843,N_2631,N_2661);
and U2844 (N_2844,N_2660,N_2655);
or U2845 (N_2845,N_2780,N_2720);
nor U2846 (N_2846,N_2750,N_2669);
nor U2847 (N_2847,N_2668,N_2699);
or U2848 (N_2848,N_2704,N_2741);
xnor U2849 (N_2849,N_2689,N_2687);
xor U2850 (N_2850,N_2770,N_2753);
and U2851 (N_2851,N_2710,N_2633);
or U2852 (N_2852,N_2663,N_2693);
nand U2853 (N_2853,N_2651,N_2795);
nand U2854 (N_2854,N_2621,N_2713);
and U2855 (N_2855,N_2752,N_2681);
or U2856 (N_2856,N_2653,N_2739);
xor U2857 (N_2857,N_2762,N_2606);
nor U2858 (N_2858,N_2644,N_2714);
and U2859 (N_2859,N_2779,N_2732);
xnor U2860 (N_2860,N_2771,N_2626);
and U2861 (N_2861,N_2667,N_2647);
nand U2862 (N_2862,N_2629,N_2643);
nor U2863 (N_2863,N_2627,N_2700);
nor U2864 (N_2864,N_2725,N_2682);
or U2865 (N_2865,N_2794,N_2639);
and U2866 (N_2866,N_2736,N_2703);
nand U2867 (N_2867,N_2789,N_2640);
nand U2868 (N_2868,N_2603,N_2609);
nand U2869 (N_2869,N_2625,N_2783);
nor U2870 (N_2870,N_2729,N_2641);
or U2871 (N_2871,N_2657,N_2735);
and U2872 (N_2872,N_2616,N_2684);
xnor U2873 (N_2873,N_2782,N_2637);
and U2874 (N_2874,N_2658,N_2666);
or U2875 (N_2875,N_2677,N_2778);
or U2876 (N_2876,N_2724,N_2747);
and U2877 (N_2877,N_2791,N_2761);
nor U2878 (N_2878,N_2615,N_2683);
xor U2879 (N_2879,N_2796,N_2691);
and U2880 (N_2880,N_2618,N_2790);
or U2881 (N_2881,N_2611,N_2678);
or U2882 (N_2882,N_2686,N_2665);
and U2883 (N_2883,N_2612,N_2602);
and U2884 (N_2884,N_2688,N_2646);
or U2885 (N_2885,N_2788,N_2638);
xor U2886 (N_2886,N_2760,N_2656);
nor U2887 (N_2887,N_2768,N_2786);
or U2888 (N_2888,N_2764,N_2773);
and U2889 (N_2889,N_2767,N_2634);
nand U2890 (N_2890,N_2607,N_2769);
and U2891 (N_2891,N_2726,N_2743);
nor U2892 (N_2892,N_2707,N_2798);
xor U2893 (N_2893,N_2650,N_2763);
nor U2894 (N_2894,N_2719,N_2685);
and U2895 (N_2895,N_2695,N_2757);
nor U2896 (N_2896,N_2721,N_2712);
or U2897 (N_2897,N_2709,N_2698);
xnor U2898 (N_2898,N_2632,N_2792);
or U2899 (N_2899,N_2628,N_2715);
nand U2900 (N_2900,N_2655,N_2630);
or U2901 (N_2901,N_2646,N_2719);
nand U2902 (N_2902,N_2784,N_2730);
nand U2903 (N_2903,N_2701,N_2693);
xor U2904 (N_2904,N_2663,N_2787);
and U2905 (N_2905,N_2751,N_2757);
nor U2906 (N_2906,N_2670,N_2790);
nand U2907 (N_2907,N_2769,N_2612);
nand U2908 (N_2908,N_2669,N_2651);
xor U2909 (N_2909,N_2782,N_2736);
xnor U2910 (N_2910,N_2714,N_2705);
nor U2911 (N_2911,N_2685,N_2632);
and U2912 (N_2912,N_2759,N_2608);
nor U2913 (N_2913,N_2765,N_2659);
nand U2914 (N_2914,N_2625,N_2672);
or U2915 (N_2915,N_2780,N_2679);
nand U2916 (N_2916,N_2688,N_2677);
or U2917 (N_2917,N_2600,N_2612);
and U2918 (N_2918,N_2755,N_2679);
and U2919 (N_2919,N_2648,N_2691);
or U2920 (N_2920,N_2605,N_2736);
nor U2921 (N_2921,N_2610,N_2697);
nor U2922 (N_2922,N_2640,N_2645);
and U2923 (N_2923,N_2670,N_2798);
nor U2924 (N_2924,N_2753,N_2613);
and U2925 (N_2925,N_2636,N_2760);
or U2926 (N_2926,N_2770,N_2670);
or U2927 (N_2927,N_2631,N_2690);
nor U2928 (N_2928,N_2642,N_2693);
xnor U2929 (N_2929,N_2600,N_2602);
or U2930 (N_2930,N_2779,N_2745);
and U2931 (N_2931,N_2622,N_2780);
or U2932 (N_2932,N_2719,N_2622);
nor U2933 (N_2933,N_2747,N_2648);
nor U2934 (N_2934,N_2748,N_2630);
nand U2935 (N_2935,N_2691,N_2749);
or U2936 (N_2936,N_2717,N_2618);
nand U2937 (N_2937,N_2626,N_2777);
xnor U2938 (N_2938,N_2707,N_2749);
nand U2939 (N_2939,N_2671,N_2791);
or U2940 (N_2940,N_2665,N_2606);
nand U2941 (N_2941,N_2732,N_2614);
xor U2942 (N_2942,N_2637,N_2722);
nand U2943 (N_2943,N_2764,N_2790);
xnor U2944 (N_2944,N_2738,N_2779);
and U2945 (N_2945,N_2784,N_2777);
xor U2946 (N_2946,N_2756,N_2772);
xor U2947 (N_2947,N_2602,N_2725);
or U2948 (N_2948,N_2765,N_2616);
or U2949 (N_2949,N_2785,N_2670);
nor U2950 (N_2950,N_2704,N_2723);
and U2951 (N_2951,N_2653,N_2616);
nor U2952 (N_2952,N_2679,N_2685);
nand U2953 (N_2953,N_2657,N_2645);
nor U2954 (N_2954,N_2688,N_2609);
and U2955 (N_2955,N_2657,N_2630);
or U2956 (N_2956,N_2760,N_2702);
xnor U2957 (N_2957,N_2793,N_2680);
or U2958 (N_2958,N_2790,N_2619);
and U2959 (N_2959,N_2752,N_2618);
nand U2960 (N_2960,N_2799,N_2658);
nand U2961 (N_2961,N_2778,N_2796);
nand U2962 (N_2962,N_2685,N_2714);
and U2963 (N_2963,N_2694,N_2737);
xor U2964 (N_2964,N_2677,N_2655);
nor U2965 (N_2965,N_2754,N_2644);
and U2966 (N_2966,N_2635,N_2717);
or U2967 (N_2967,N_2695,N_2686);
or U2968 (N_2968,N_2725,N_2723);
nand U2969 (N_2969,N_2628,N_2773);
nand U2970 (N_2970,N_2646,N_2701);
nand U2971 (N_2971,N_2771,N_2753);
nand U2972 (N_2972,N_2632,N_2743);
and U2973 (N_2973,N_2669,N_2749);
or U2974 (N_2974,N_2780,N_2778);
and U2975 (N_2975,N_2728,N_2652);
or U2976 (N_2976,N_2751,N_2768);
and U2977 (N_2977,N_2799,N_2748);
xnor U2978 (N_2978,N_2750,N_2749);
xnor U2979 (N_2979,N_2707,N_2688);
nand U2980 (N_2980,N_2717,N_2641);
nor U2981 (N_2981,N_2698,N_2694);
nor U2982 (N_2982,N_2682,N_2705);
or U2983 (N_2983,N_2793,N_2759);
nor U2984 (N_2984,N_2794,N_2630);
or U2985 (N_2985,N_2764,N_2794);
xor U2986 (N_2986,N_2673,N_2715);
xnor U2987 (N_2987,N_2624,N_2728);
or U2988 (N_2988,N_2664,N_2776);
and U2989 (N_2989,N_2651,N_2741);
xnor U2990 (N_2990,N_2774,N_2671);
xnor U2991 (N_2991,N_2614,N_2725);
and U2992 (N_2992,N_2640,N_2750);
nor U2993 (N_2993,N_2733,N_2652);
or U2994 (N_2994,N_2721,N_2791);
xnor U2995 (N_2995,N_2773,N_2703);
or U2996 (N_2996,N_2761,N_2756);
xnor U2997 (N_2997,N_2780,N_2662);
and U2998 (N_2998,N_2784,N_2749);
xor U2999 (N_2999,N_2780,N_2716);
nor U3000 (N_3000,N_2875,N_2862);
and U3001 (N_3001,N_2884,N_2878);
and U3002 (N_3002,N_2869,N_2906);
xor U3003 (N_3003,N_2907,N_2966);
and U3004 (N_3004,N_2913,N_2924);
xor U3005 (N_3005,N_2822,N_2929);
nor U3006 (N_3006,N_2898,N_2986);
nand U3007 (N_3007,N_2838,N_2904);
nand U3008 (N_3008,N_2815,N_2810);
and U3009 (N_3009,N_2902,N_2811);
xor U3010 (N_3010,N_2874,N_2819);
and U3011 (N_3011,N_2813,N_2958);
and U3012 (N_3012,N_2814,N_2826);
and U3013 (N_3013,N_2859,N_2877);
nor U3014 (N_3014,N_2899,N_2962);
nor U3015 (N_3015,N_2833,N_2892);
or U3016 (N_3016,N_2837,N_2854);
nand U3017 (N_3017,N_2809,N_2827);
nor U3018 (N_3018,N_2805,N_2903);
and U3019 (N_3019,N_2823,N_2952);
or U3020 (N_3020,N_2830,N_2896);
nor U3021 (N_3021,N_2840,N_2905);
nor U3022 (N_3022,N_2974,N_2982);
nand U3023 (N_3023,N_2939,N_2856);
nand U3024 (N_3024,N_2825,N_2973);
nand U3025 (N_3025,N_2941,N_2940);
xnor U3026 (N_3026,N_2953,N_2914);
xnor U3027 (N_3027,N_2866,N_2992);
xor U3028 (N_3028,N_2891,N_2926);
and U3029 (N_3029,N_2967,N_2820);
xnor U3030 (N_3030,N_2969,N_2872);
and U3031 (N_3031,N_2976,N_2829);
nor U3032 (N_3032,N_2945,N_2812);
nor U3033 (N_3033,N_2930,N_2909);
or U3034 (N_3034,N_2870,N_2994);
or U3035 (N_3035,N_2828,N_2844);
and U3036 (N_3036,N_2916,N_2954);
nand U3037 (N_3037,N_2951,N_2804);
or U3038 (N_3038,N_2818,N_2927);
and U3039 (N_3039,N_2993,N_2988);
and U3040 (N_3040,N_2831,N_2853);
xor U3041 (N_3041,N_2880,N_2843);
xor U3042 (N_3042,N_2855,N_2981);
and U3043 (N_3043,N_2824,N_2996);
and U3044 (N_3044,N_2802,N_2922);
and U3045 (N_3045,N_2890,N_2889);
and U3046 (N_3046,N_2895,N_2979);
and U3047 (N_3047,N_2997,N_2999);
xor U3048 (N_3048,N_2871,N_2832);
nand U3049 (N_3049,N_2955,N_2977);
xnor U3050 (N_3050,N_2876,N_2942);
nand U3051 (N_3051,N_2918,N_2821);
or U3052 (N_3052,N_2842,N_2881);
nand U3053 (N_3053,N_2946,N_2852);
or U3054 (N_3054,N_2816,N_2975);
xnor U3055 (N_3055,N_2925,N_2964);
nor U3056 (N_3056,N_2801,N_2841);
and U3057 (N_3057,N_2860,N_2873);
nand U3058 (N_3058,N_2806,N_2868);
or U3059 (N_3059,N_2901,N_2935);
xnor U3060 (N_3060,N_2919,N_2894);
nor U3061 (N_3061,N_2836,N_2947);
xor U3062 (N_3062,N_2960,N_2938);
and U3063 (N_3063,N_2845,N_2949);
xor U3064 (N_3064,N_2835,N_2972);
and U3065 (N_3065,N_2934,N_2839);
and U3066 (N_3066,N_2879,N_2915);
nand U3067 (N_3067,N_2849,N_2937);
or U3068 (N_3068,N_2932,N_2931);
nor U3069 (N_3069,N_2920,N_2912);
nand U3070 (N_3070,N_2923,N_2908);
xnor U3071 (N_3071,N_2957,N_2987);
nor U3072 (N_3072,N_2961,N_2959);
nand U3073 (N_3073,N_2995,N_2897);
nand U3074 (N_3074,N_2864,N_2850);
nand U3075 (N_3075,N_2956,N_2867);
nand U3076 (N_3076,N_2863,N_2989);
xor U3077 (N_3077,N_2968,N_2834);
and U3078 (N_3078,N_2803,N_2808);
xor U3079 (N_3079,N_2985,N_2800);
or U3080 (N_3080,N_2893,N_2921);
xor U3081 (N_3081,N_2851,N_2865);
and U3082 (N_3082,N_2983,N_2943);
and U3083 (N_3083,N_2886,N_2963);
and U3084 (N_3084,N_2882,N_2984);
or U3085 (N_3085,N_2933,N_2928);
nand U3086 (N_3086,N_2980,N_2888);
or U3087 (N_3087,N_2965,N_2971);
xnor U3088 (N_3088,N_2911,N_2936);
xor U3089 (N_3089,N_2846,N_2991);
and U3090 (N_3090,N_2950,N_2944);
nand U3091 (N_3091,N_2887,N_2978);
nor U3092 (N_3092,N_2998,N_2917);
nand U3093 (N_3093,N_2885,N_2948);
xor U3094 (N_3094,N_2858,N_2990);
nor U3095 (N_3095,N_2848,N_2900);
nor U3096 (N_3096,N_2861,N_2883);
or U3097 (N_3097,N_2807,N_2970);
nand U3098 (N_3098,N_2857,N_2847);
nor U3099 (N_3099,N_2910,N_2817);
or U3100 (N_3100,N_2934,N_2941);
nand U3101 (N_3101,N_2970,N_2948);
xnor U3102 (N_3102,N_2960,N_2991);
nor U3103 (N_3103,N_2875,N_2801);
nand U3104 (N_3104,N_2986,N_2846);
and U3105 (N_3105,N_2833,N_2926);
nor U3106 (N_3106,N_2985,N_2993);
and U3107 (N_3107,N_2806,N_2814);
xnor U3108 (N_3108,N_2955,N_2897);
nor U3109 (N_3109,N_2827,N_2916);
nor U3110 (N_3110,N_2824,N_2937);
or U3111 (N_3111,N_2982,N_2856);
and U3112 (N_3112,N_2942,N_2862);
nand U3113 (N_3113,N_2868,N_2949);
nor U3114 (N_3114,N_2979,N_2961);
or U3115 (N_3115,N_2879,N_2894);
xnor U3116 (N_3116,N_2910,N_2997);
and U3117 (N_3117,N_2991,N_2840);
xor U3118 (N_3118,N_2830,N_2839);
or U3119 (N_3119,N_2911,N_2934);
nor U3120 (N_3120,N_2881,N_2871);
or U3121 (N_3121,N_2867,N_2984);
or U3122 (N_3122,N_2960,N_2802);
or U3123 (N_3123,N_2978,N_2800);
and U3124 (N_3124,N_2849,N_2855);
and U3125 (N_3125,N_2845,N_2873);
nor U3126 (N_3126,N_2917,N_2849);
xnor U3127 (N_3127,N_2874,N_2890);
and U3128 (N_3128,N_2841,N_2976);
and U3129 (N_3129,N_2955,N_2823);
nor U3130 (N_3130,N_2954,N_2908);
nand U3131 (N_3131,N_2824,N_2883);
nand U3132 (N_3132,N_2850,N_2870);
and U3133 (N_3133,N_2987,N_2896);
nand U3134 (N_3134,N_2959,N_2868);
and U3135 (N_3135,N_2833,N_2855);
or U3136 (N_3136,N_2886,N_2935);
xor U3137 (N_3137,N_2976,N_2804);
nor U3138 (N_3138,N_2854,N_2870);
xnor U3139 (N_3139,N_2890,N_2911);
or U3140 (N_3140,N_2861,N_2863);
and U3141 (N_3141,N_2909,N_2869);
xor U3142 (N_3142,N_2830,N_2924);
or U3143 (N_3143,N_2957,N_2811);
and U3144 (N_3144,N_2947,N_2936);
and U3145 (N_3145,N_2895,N_2905);
nor U3146 (N_3146,N_2961,N_2945);
or U3147 (N_3147,N_2960,N_2865);
xor U3148 (N_3148,N_2801,N_2944);
or U3149 (N_3149,N_2954,N_2992);
xnor U3150 (N_3150,N_2930,N_2826);
or U3151 (N_3151,N_2986,N_2992);
nand U3152 (N_3152,N_2835,N_2994);
and U3153 (N_3153,N_2801,N_2971);
or U3154 (N_3154,N_2859,N_2856);
or U3155 (N_3155,N_2869,N_2849);
xor U3156 (N_3156,N_2865,N_2919);
and U3157 (N_3157,N_2874,N_2981);
and U3158 (N_3158,N_2867,N_2949);
or U3159 (N_3159,N_2977,N_2938);
nor U3160 (N_3160,N_2986,N_2825);
or U3161 (N_3161,N_2865,N_2843);
nor U3162 (N_3162,N_2860,N_2994);
xnor U3163 (N_3163,N_2801,N_2910);
nand U3164 (N_3164,N_2846,N_2964);
nor U3165 (N_3165,N_2909,N_2908);
xor U3166 (N_3166,N_2980,N_2854);
or U3167 (N_3167,N_2931,N_2848);
or U3168 (N_3168,N_2868,N_2881);
xnor U3169 (N_3169,N_2814,N_2991);
nor U3170 (N_3170,N_2983,N_2992);
and U3171 (N_3171,N_2872,N_2828);
xnor U3172 (N_3172,N_2985,N_2988);
and U3173 (N_3173,N_2924,N_2951);
and U3174 (N_3174,N_2842,N_2896);
xnor U3175 (N_3175,N_2902,N_2804);
nand U3176 (N_3176,N_2808,N_2846);
or U3177 (N_3177,N_2808,N_2996);
nand U3178 (N_3178,N_2859,N_2825);
nand U3179 (N_3179,N_2945,N_2920);
nor U3180 (N_3180,N_2854,N_2888);
xor U3181 (N_3181,N_2854,N_2920);
and U3182 (N_3182,N_2922,N_2907);
or U3183 (N_3183,N_2924,N_2997);
nand U3184 (N_3184,N_2906,N_2989);
or U3185 (N_3185,N_2985,N_2959);
nand U3186 (N_3186,N_2836,N_2843);
nand U3187 (N_3187,N_2816,N_2934);
xor U3188 (N_3188,N_2815,N_2987);
nor U3189 (N_3189,N_2809,N_2966);
and U3190 (N_3190,N_2990,N_2971);
xnor U3191 (N_3191,N_2959,N_2963);
nor U3192 (N_3192,N_2958,N_2959);
xnor U3193 (N_3193,N_2963,N_2866);
xor U3194 (N_3194,N_2980,N_2878);
or U3195 (N_3195,N_2902,N_2968);
nor U3196 (N_3196,N_2929,N_2842);
nand U3197 (N_3197,N_2848,N_2857);
xnor U3198 (N_3198,N_2859,N_2981);
nand U3199 (N_3199,N_2911,N_2854);
nand U3200 (N_3200,N_3030,N_3144);
and U3201 (N_3201,N_3015,N_3155);
and U3202 (N_3202,N_3073,N_3056);
nor U3203 (N_3203,N_3069,N_3041);
or U3204 (N_3204,N_3016,N_3079);
or U3205 (N_3205,N_3173,N_3191);
and U3206 (N_3206,N_3168,N_3060);
nand U3207 (N_3207,N_3190,N_3031);
nor U3208 (N_3208,N_3006,N_3127);
and U3209 (N_3209,N_3166,N_3120);
xnor U3210 (N_3210,N_3178,N_3121);
and U3211 (N_3211,N_3078,N_3038);
nor U3212 (N_3212,N_3167,N_3068);
nand U3213 (N_3213,N_3087,N_3081);
xor U3214 (N_3214,N_3109,N_3074);
nor U3215 (N_3215,N_3021,N_3125);
and U3216 (N_3216,N_3008,N_3054);
nor U3217 (N_3217,N_3010,N_3142);
xor U3218 (N_3218,N_3149,N_3072);
or U3219 (N_3219,N_3018,N_3089);
nor U3220 (N_3220,N_3161,N_3138);
nand U3221 (N_3221,N_3132,N_3196);
xor U3222 (N_3222,N_3172,N_3082);
nand U3223 (N_3223,N_3098,N_3176);
nor U3224 (N_3224,N_3184,N_3195);
and U3225 (N_3225,N_3177,N_3123);
nor U3226 (N_3226,N_3198,N_3034);
nand U3227 (N_3227,N_3174,N_3063);
nand U3228 (N_3228,N_3017,N_3092);
xnor U3229 (N_3229,N_3066,N_3111);
nor U3230 (N_3230,N_3024,N_3146);
and U3231 (N_3231,N_3171,N_3106);
nor U3232 (N_3232,N_3045,N_3085);
nor U3233 (N_3233,N_3137,N_3160);
or U3234 (N_3234,N_3004,N_3185);
xor U3235 (N_3235,N_3107,N_3152);
xnor U3236 (N_3236,N_3105,N_3165);
or U3237 (N_3237,N_3032,N_3150);
nand U3238 (N_3238,N_3128,N_3169);
nand U3239 (N_3239,N_3058,N_3181);
nand U3240 (N_3240,N_3187,N_3023);
nor U3241 (N_3241,N_3156,N_3000);
xor U3242 (N_3242,N_3026,N_3100);
nand U3243 (N_3243,N_3099,N_3055);
and U3244 (N_3244,N_3094,N_3005);
and U3245 (N_3245,N_3151,N_3158);
nand U3246 (N_3246,N_3014,N_3022);
nor U3247 (N_3247,N_3076,N_3130);
xor U3248 (N_3248,N_3065,N_3129);
or U3249 (N_3249,N_3180,N_3194);
nand U3250 (N_3250,N_3095,N_3011);
or U3251 (N_3251,N_3117,N_3003);
nand U3252 (N_3252,N_3153,N_3088);
nor U3253 (N_3253,N_3103,N_3020);
nand U3254 (N_3254,N_3157,N_3053);
xor U3255 (N_3255,N_3007,N_3080);
nand U3256 (N_3256,N_3002,N_3119);
nand U3257 (N_3257,N_3019,N_3083);
xnor U3258 (N_3258,N_3159,N_3182);
nor U3259 (N_3259,N_3048,N_3001);
nand U3260 (N_3260,N_3049,N_3009);
and U3261 (N_3261,N_3090,N_3122);
nor U3262 (N_3262,N_3039,N_3114);
or U3263 (N_3263,N_3064,N_3179);
nor U3264 (N_3264,N_3037,N_3136);
and U3265 (N_3265,N_3025,N_3046);
or U3266 (N_3266,N_3110,N_3145);
or U3267 (N_3267,N_3044,N_3051);
or U3268 (N_3268,N_3047,N_3108);
nand U3269 (N_3269,N_3084,N_3050);
xor U3270 (N_3270,N_3141,N_3036);
nand U3271 (N_3271,N_3101,N_3183);
xor U3272 (N_3272,N_3131,N_3189);
nor U3273 (N_3273,N_3188,N_3112);
nand U3274 (N_3274,N_3086,N_3013);
nand U3275 (N_3275,N_3134,N_3097);
nand U3276 (N_3276,N_3040,N_3075);
and U3277 (N_3277,N_3139,N_3140);
nor U3278 (N_3278,N_3096,N_3012);
and U3279 (N_3279,N_3028,N_3148);
or U3280 (N_3280,N_3033,N_3070);
or U3281 (N_3281,N_3052,N_3133);
nand U3282 (N_3282,N_3035,N_3126);
nand U3283 (N_3283,N_3091,N_3118);
nand U3284 (N_3284,N_3062,N_3059);
nand U3285 (N_3285,N_3170,N_3186);
nor U3286 (N_3286,N_3192,N_3147);
nor U3287 (N_3287,N_3113,N_3027);
and U3288 (N_3288,N_3042,N_3143);
nand U3289 (N_3289,N_3067,N_3124);
or U3290 (N_3290,N_3164,N_3193);
or U3291 (N_3291,N_3102,N_3197);
nand U3292 (N_3292,N_3057,N_3043);
nor U3293 (N_3293,N_3163,N_3154);
xnor U3294 (N_3294,N_3162,N_3077);
and U3295 (N_3295,N_3199,N_3029);
nor U3296 (N_3296,N_3093,N_3104);
and U3297 (N_3297,N_3071,N_3175);
or U3298 (N_3298,N_3116,N_3115);
nand U3299 (N_3299,N_3061,N_3135);
and U3300 (N_3300,N_3098,N_3083);
nand U3301 (N_3301,N_3132,N_3141);
nand U3302 (N_3302,N_3009,N_3128);
or U3303 (N_3303,N_3163,N_3188);
nand U3304 (N_3304,N_3166,N_3113);
nor U3305 (N_3305,N_3117,N_3104);
xor U3306 (N_3306,N_3184,N_3062);
nor U3307 (N_3307,N_3068,N_3045);
xnor U3308 (N_3308,N_3075,N_3173);
nor U3309 (N_3309,N_3143,N_3121);
and U3310 (N_3310,N_3073,N_3179);
and U3311 (N_3311,N_3107,N_3007);
nand U3312 (N_3312,N_3039,N_3008);
or U3313 (N_3313,N_3162,N_3161);
nor U3314 (N_3314,N_3114,N_3115);
or U3315 (N_3315,N_3086,N_3111);
or U3316 (N_3316,N_3075,N_3030);
nand U3317 (N_3317,N_3164,N_3194);
or U3318 (N_3318,N_3047,N_3096);
and U3319 (N_3319,N_3157,N_3049);
or U3320 (N_3320,N_3048,N_3119);
nand U3321 (N_3321,N_3114,N_3197);
xnor U3322 (N_3322,N_3029,N_3059);
or U3323 (N_3323,N_3137,N_3184);
xnor U3324 (N_3324,N_3000,N_3097);
nand U3325 (N_3325,N_3123,N_3150);
nor U3326 (N_3326,N_3030,N_3014);
nand U3327 (N_3327,N_3168,N_3038);
nor U3328 (N_3328,N_3189,N_3101);
and U3329 (N_3329,N_3151,N_3165);
xnor U3330 (N_3330,N_3158,N_3065);
and U3331 (N_3331,N_3130,N_3077);
nor U3332 (N_3332,N_3123,N_3015);
nor U3333 (N_3333,N_3025,N_3065);
xor U3334 (N_3334,N_3098,N_3034);
xnor U3335 (N_3335,N_3046,N_3177);
or U3336 (N_3336,N_3166,N_3107);
xnor U3337 (N_3337,N_3127,N_3087);
nor U3338 (N_3338,N_3181,N_3180);
nor U3339 (N_3339,N_3090,N_3129);
nand U3340 (N_3340,N_3123,N_3143);
xor U3341 (N_3341,N_3000,N_3063);
or U3342 (N_3342,N_3182,N_3061);
nand U3343 (N_3343,N_3052,N_3073);
nand U3344 (N_3344,N_3131,N_3052);
xnor U3345 (N_3345,N_3084,N_3137);
nor U3346 (N_3346,N_3047,N_3168);
or U3347 (N_3347,N_3175,N_3166);
and U3348 (N_3348,N_3119,N_3055);
nor U3349 (N_3349,N_3125,N_3072);
or U3350 (N_3350,N_3036,N_3153);
nand U3351 (N_3351,N_3048,N_3128);
xnor U3352 (N_3352,N_3028,N_3123);
or U3353 (N_3353,N_3130,N_3120);
nand U3354 (N_3354,N_3052,N_3031);
or U3355 (N_3355,N_3033,N_3099);
or U3356 (N_3356,N_3120,N_3058);
nand U3357 (N_3357,N_3039,N_3145);
xor U3358 (N_3358,N_3075,N_3099);
or U3359 (N_3359,N_3061,N_3086);
nor U3360 (N_3360,N_3067,N_3033);
nand U3361 (N_3361,N_3020,N_3030);
and U3362 (N_3362,N_3095,N_3105);
nand U3363 (N_3363,N_3059,N_3078);
or U3364 (N_3364,N_3104,N_3034);
nand U3365 (N_3365,N_3044,N_3182);
or U3366 (N_3366,N_3190,N_3180);
nand U3367 (N_3367,N_3055,N_3180);
or U3368 (N_3368,N_3123,N_3011);
and U3369 (N_3369,N_3115,N_3096);
or U3370 (N_3370,N_3075,N_3048);
nor U3371 (N_3371,N_3074,N_3165);
and U3372 (N_3372,N_3081,N_3040);
and U3373 (N_3373,N_3048,N_3087);
nand U3374 (N_3374,N_3085,N_3027);
nand U3375 (N_3375,N_3028,N_3031);
nor U3376 (N_3376,N_3112,N_3132);
nand U3377 (N_3377,N_3143,N_3061);
nor U3378 (N_3378,N_3095,N_3142);
nand U3379 (N_3379,N_3148,N_3195);
or U3380 (N_3380,N_3115,N_3180);
nand U3381 (N_3381,N_3172,N_3062);
nand U3382 (N_3382,N_3007,N_3047);
or U3383 (N_3383,N_3163,N_3127);
or U3384 (N_3384,N_3118,N_3187);
or U3385 (N_3385,N_3193,N_3082);
and U3386 (N_3386,N_3180,N_3006);
xnor U3387 (N_3387,N_3000,N_3172);
nand U3388 (N_3388,N_3143,N_3063);
nor U3389 (N_3389,N_3004,N_3027);
xor U3390 (N_3390,N_3038,N_3099);
nand U3391 (N_3391,N_3004,N_3020);
and U3392 (N_3392,N_3014,N_3150);
xor U3393 (N_3393,N_3019,N_3165);
xnor U3394 (N_3394,N_3134,N_3152);
and U3395 (N_3395,N_3024,N_3137);
or U3396 (N_3396,N_3191,N_3009);
and U3397 (N_3397,N_3113,N_3155);
nand U3398 (N_3398,N_3128,N_3096);
and U3399 (N_3399,N_3136,N_3107);
nand U3400 (N_3400,N_3378,N_3216);
and U3401 (N_3401,N_3208,N_3236);
or U3402 (N_3402,N_3224,N_3337);
nand U3403 (N_3403,N_3373,N_3345);
xnor U3404 (N_3404,N_3235,N_3308);
nand U3405 (N_3405,N_3259,N_3312);
and U3406 (N_3406,N_3269,N_3324);
nor U3407 (N_3407,N_3205,N_3281);
nand U3408 (N_3408,N_3255,N_3207);
nor U3409 (N_3409,N_3364,N_3361);
nor U3410 (N_3410,N_3356,N_3202);
nor U3411 (N_3411,N_3241,N_3365);
xnor U3412 (N_3412,N_3382,N_3334);
nor U3413 (N_3413,N_3239,N_3222);
or U3414 (N_3414,N_3232,N_3354);
xnor U3415 (N_3415,N_3260,N_3328);
nor U3416 (N_3416,N_3227,N_3340);
or U3417 (N_3417,N_3242,N_3321);
xnor U3418 (N_3418,N_3371,N_3355);
or U3419 (N_3419,N_3266,N_3213);
and U3420 (N_3420,N_3295,N_3217);
and U3421 (N_3421,N_3284,N_3200);
nand U3422 (N_3422,N_3368,N_3268);
nand U3423 (N_3423,N_3301,N_3313);
nand U3424 (N_3424,N_3351,N_3293);
or U3425 (N_3425,N_3325,N_3370);
xor U3426 (N_3426,N_3289,N_3349);
or U3427 (N_3427,N_3316,N_3342);
nor U3428 (N_3428,N_3362,N_3240);
nand U3429 (N_3429,N_3258,N_3294);
xor U3430 (N_3430,N_3393,N_3226);
nor U3431 (N_3431,N_3347,N_3306);
or U3432 (N_3432,N_3244,N_3253);
xor U3433 (N_3433,N_3265,N_3336);
or U3434 (N_3434,N_3237,N_3302);
nand U3435 (N_3435,N_3287,N_3267);
and U3436 (N_3436,N_3288,N_3383);
or U3437 (N_3437,N_3204,N_3249);
nand U3438 (N_3438,N_3214,N_3327);
nand U3439 (N_3439,N_3344,N_3298);
and U3440 (N_3440,N_3212,N_3329);
xnor U3441 (N_3441,N_3272,N_3391);
xnor U3442 (N_3442,N_3320,N_3206);
xnor U3443 (N_3443,N_3300,N_3231);
nor U3444 (N_3444,N_3264,N_3238);
or U3445 (N_3445,N_3395,N_3397);
and U3446 (N_3446,N_3396,N_3201);
xnor U3447 (N_3447,N_3379,N_3219);
nand U3448 (N_3448,N_3210,N_3292);
nand U3449 (N_3449,N_3353,N_3317);
nor U3450 (N_3450,N_3277,N_3352);
nand U3451 (N_3451,N_3311,N_3233);
xnor U3452 (N_3452,N_3279,N_3338);
xnor U3453 (N_3453,N_3282,N_3384);
nor U3454 (N_3454,N_3263,N_3322);
xnor U3455 (N_3455,N_3331,N_3399);
nor U3456 (N_3456,N_3385,N_3250);
nand U3457 (N_3457,N_3394,N_3375);
nand U3458 (N_3458,N_3341,N_3376);
or U3459 (N_3459,N_3230,N_3234);
nand U3460 (N_3460,N_3304,N_3330);
nor U3461 (N_3461,N_3366,N_3203);
nor U3462 (N_3462,N_3286,N_3318);
or U3463 (N_3463,N_3276,N_3339);
nor U3464 (N_3464,N_3346,N_3254);
nor U3465 (N_3465,N_3248,N_3392);
nand U3466 (N_3466,N_3319,N_3297);
and U3467 (N_3467,N_3220,N_3315);
or U3468 (N_3468,N_3299,N_3332);
xor U3469 (N_3469,N_3246,N_3314);
or U3470 (N_3470,N_3273,N_3228);
xnor U3471 (N_3471,N_3271,N_3398);
or U3472 (N_3472,N_3360,N_3247);
or U3473 (N_3473,N_3305,N_3257);
xnor U3474 (N_3474,N_3215,N_3218);
or U3475 (N_3475,N_3358,N_3291);
and U3476 (N_3476,N_3221,N_3296);
nand U3477 (N_3477,N_3283,N_3323);
nand U3478 (N_3478,N_3388,N_3251);
nor U3479 (N_3479,N_3369,N_3389);
or U3480 (N_3480,N_3367,N_3387);
or U3481 (N_3481,N_3278,N_3380);
nor U3482 (N_3482,N_3343,N_3211);
xnor U3483 (N_3483,N_3270,N_3348);
or U3484 (N_3484,N_3209,N_3274);
nor U3485 (N_3485,N_3229,N_3290);
nor U3486 (N_3486,N_3310,N_3377);
or U3487 (N_3487,N_3333,N_3252);
nor U3488 (N_3488,N_3381,N_3223);
nand U3489 (N_3489,N_3256,N_3280);
nor U3490 (N_3490,N_3261,N_3307);
xor U3491 (N_3491,N_3363,N_3285);
and U3492 (N_3492,N_3245,N_3326);
and U3493 (N_3493,N_3374,N_3262);
xor U3494 (N_3494,N_3309,N_3243);
xor U3495 (N_3495,N_3350,N_3335);
or U3496 (N_3496,N_3225,N_3386);
nor U3497 (N_3497,N_3372,N_3359);
nor U3498 (N_3498,N_3275,N_3357);
xor U3499 (N_3499,N_3390,N_3303);
xnor U3500 (N_3500,N_3340,N_3394);
xnor U3501 (N_3501,N_3364,N_3365);
nand U3502 (N_3502,N_3284,N_3348);
and U3503 (N_3503,N_3345,N_3299);
and U3504 (N_3504,N_3340,N_3330);
xor U3505 (N_3505,N_3394,N_3216);
xnor U3506 (N_3506,N_3306,N_3370);
nand U3507 (N_3507,N_3308,N_3288);
nand U3508 (N_3508,N_3298,N_3354);
nor U3509 (N_3509,N_3253,N_3393);
or U3510 (N_3510,N_3345,N_3262);
or U3511 (N_3511,N_3294,N_3226);
nor U3512 (N_3512,N_3268,N_3309);
nor U3513 (N_3513,N_3250,N_3238);
and U3514 (N_3514,N_3202,N_3204);
and U3515 (N_3515,N_3272,N_3373);
nand U3516 (N_3516,N_3345,N_3342);
nor U3517 (N_3517,N_3229,N_3227);
or U3518 (N_3518,N_3265,N_3255);
nor U3519 (N_3519,N_3348,N_3299);
nand U3520 (N_3520,N_3280,N_3334);
or U3521 (N_3521,N_3253,N_3254);
and U3522 (N_3522,N_3299,N_3352);
nor U3523 (N_3523,N_3231,N_3333);
nand U3524 (N_3524,N_3224,N_3340);
nor U3525 (N_3525,N_3344,N_3369);
xnor U3526 (N_3526,N_3396,N_3388);
or U3527 (N_3527,N_3220,N_3394);
or U3528 (N_3528,N_3253,N_3350);
and U3529 (N_3529,N_3301,N_3232);
nand U3530 (N_3530,N_3386,N_3312);
nor U3531 (N_3531,N_3364,N_3316);
nand U3532 (N_3532,N_3244,N_3258);
nand U3533 (N_3533,N_3379,N_3306);
or U3534 (N_3534,N_3302,N_3259);
xor U3535 (N_3535,N_3311,N_3313);
nor U3536 (N_3536,N_3270,N_3327);
xnor U3537 (N_3537,N_3338,N_3202);
and U3538 (N_3538,N_3308,N_3368);
and U3539 (N_3539,N_3204,N_3326);
or U3540 (N_3540,N_3264,N_3236);
nor U3541 (N_3541,N_3366,N_3251);
nor U3542 (N_3542,N_3240,N_3365);
nand U3543 (N_3543,N_3326,N_3220);
nand U3544 (N_3544,N_3267,N_3356);
nand U3545 (N_3545,N_3213,N_3247);
xor U3546 (N_3546,N_3297,N_3391);
xnor U3547 (N_3547,N_3332,N_3251);
xnor U3548 (N_3548,N_3234,N_3367);
xnor U3549 (N_3549,N_3358,N_3377);
and U3550 (N_3550,N_3235,N_3267);
and U3551 (N_3551,N_3319,N_3314);
and U3552 (N_3552,N_3214,N_3227);
nor U3553 (N_3553,N_3276,N_3344);
nor U3554 (N_3554,N_3233,N_3388);
xnor U3555 (N_3555,N_3386,N_3251);
nand U3556 (N_3556,N_3342,N_3376);
nand U3557 (N_3557,N_3306,N_3212);
and U3558 (N_3558,N_3325,N_3230);
nand U3559 (N_3559,N_3353,N_3212);
xnor U3560 (N_3560,N_3388,N_3294);
and U3561 (N_3561,N_3238,N_3391);
and U3562 (N_3562,N_3397,N_3278);
or U3563 (N_3563,N_3351,N_3342);
and U3564 (N_3564,N_3239,N_3211);
or U3565 (N_3565,N_3209,N_3359);
nor U3566 (N_3566,N_3221,N_3213);
and U3567 (N_3567,N_3234,N_3220);
or U3568 (N_3568,N_3269,N_3206);
and U3569 (N_3569,N_3349,N_3254);
xor U3570 (N_3570,N_3212,N_3352);
xor U3571 (N_3571,N_3380,N_3291);
xor U3572 (N_3572,N_3301,N_3346);
or U3573 (N_3573,N_3320,N_3221);
nor U3574 (N_3574,N_3268,N_3336);
xor U3575 (N_3575,N_3243,N_3375);
and U3576 (N_3576,N_3337,N_3259);
nand U3577 (N_3577,N_3273,N_3333);
or U3578 (N_3578,N_3238,N_3281);
nand U3579 (N_3579,N_3378,N_3322);
and U3580 (N_3580,N_3291,N_3334);
and U3581 (N_3581,N_3203,N_3387);
nor U3582 (N_3582,N_3301,N_3350);
xor U3583 (N_3583,N_3319,N_3347);
or U3584 (N_3584,N_3276,N_3329);
or U3585 (N_3585,N_3383,N_3313);
and U3586 (N_3586,N_3261,N_3242);
and U3587 (N_3587,N_3313,N_3241);
nor U3588 (N_3588,N_3351,N_3200);
nand U3589 (N_3589,N_3203,N_3398);
xor U3590 (N_3590,N_3277,N_3381);
nor U3591 (N_3591,N_3223,N_3360);
and U3592 (N_3592,N_3311,N_3396);
nand U3593 (N_3593,N_3211,N_3272);
and U3594 (N_3594,N_3207,N_3339);
or U3595 (N_3595,N_3298,N_3367);
and U3596 (N_3596,N_3231,N_3270);
and U3597 (N_3597,N_3334,N_3287);
xor U3598 (N_3598,N_3271,N_3323);
xor U3599 (N_3599,N_3392,N_3310);
and U3600 (N_3600,N_3532,N_3449);
nor U3601 (N_3601,N_3442,N_3470);
or U3602 (N_3602,N_3543,N_3491);
nand U3603 (N_3603,N_3411,N_3569);
nand U3604 (N_3604,N_3483,N_3472);
xor U3605 (N_3605,N_3594,N_3534);
nor U3606 (N_3606,N_3447,N_3456);
or U3607 (N_3607,N_3413,N_3476);
xor U3608 (N_3608,N_3509,N_3469);
and U3609 (N_3609,N_3558,N_3530);
or U3610 (N_3610,N_3497,N_3460);
nand U3611 (N_3611,N_3599,N_3478);
nor U3612 (N_3612,N_3550,N_3523);
xor U3613 (N_3613,N_3482,N_3495);
and U3614 (N_3614,N_3420,N_3492);
nor U3615 (N_3615,N_3416,N_3572);
xnor U3616 (N_3616,N_3508,N_3443);
nor U3617 (N_3617,N_3562,N_3405);
or U3618 (N_3618,N_3598,N_3500);
nand U3619 (N_3619,N_3518,N_3587);
xnor U3620 (N_3620,N_3404,N_3526);
and U3621 (N_3621,N_3506,N_3560);
or U3622 (N_3622,N_3589,N_3593);
or U3623 (N_3623,N_3512,N_3474);
or U3624 (N_3624,N_3540,N_3503);
nand U3625 (N_3625,N_3584,N_3490);
nand U3626 (N_3626,N_3477,N_3453);
xnor U3627 (N_3627,N_3513,N_3432);
nand U3628 (N_3628,N_3410,N_3402);
xnor U3629 (N_3629,N_3465,N_3583);
nor U3630 (N_3630,N_3457,N_3585);
nand U3631 (N_3631,N_3450,N_3564);
and U3632 (N_3632,N_3507,N_3535);
or U3633 (N_3633,N_3570,N_3521);
and U3634 (N_3634,N_3438,N_3592);
nor U3635 (N_3635,N_3496,N_3554);
nor U3636 (N_3636,N_3529,N_3525);
and U3637 (N_3637,N_3423,N_3544);
nand U3638 (N_3638,N_3458,N_3439);
nor U3639 (N_3639,N_3557,N_3537);
nor U3640 (N_3640,N_3577,N_3546);
nor U3641 (N_3641,N_3571,N_3579);
nand U3642 (N_3642,N_3552,N_3510);
or U3643 (N_3643,N_3556,N_3433);
nand U3644 (N_3644,N_3517,N_3549);
and U3645 (N_3645,N_3454,N_3436);
or U3646 (N_3646,N_3418,N_3417);
nand U3647 (N_3647,N_3565,N_3446);
and U3648 (N_3648,N_3504,N_3515);
or U3649 (N_3649,N_3441,N_3553);
nand U3650 (N_3650,N_3555,N_3547);
and U3651 (N_3651,N_3488,N_3591);
nor U3652 (N_3652,N_3498,N_3561);
xor U3653 (N_3653,N_3581,N_3461);
or U3654 (N_3654,N_3573,N_3580);
nor U3655 (N_3655,N_3464,N_3401);
nand U3656 (N_3656,N_3480,N_3596);
and U3657 (N_3657,N_3516,N_3493);
or U3658 (N_3658,N_3531,N_3429);
and U3659 (N_3659,N_3473,N_3533);
or U3660 (N_3660,N_3536,N_3566);
nand U3661 (N_3661,N_3479,N_3403);
nand U3662 (N_3662,N_3568,N_3582);
or U3663 (N_3663,N_3485,N_3514);
nand U3664 (N_3664,N_3430,N_3407);
xnor U3665 (N_3665,N_3501,N_3511);
nor U3666 (N_3666,N_3467,N_3426);
and U3667 (N_3667,N_3445,N_3588);
xor U3668 (N_3668,N_3428,N_3538);
nand U3669 (N_3669,N_3412,N_3595);
nand U3670 (N_3670,N_3471,N_3578);
xor U3671 (N_3671,N_3466,N_3419);
nor U3672 (N_3672,N_3425,N_3431);
or U3673 (N_3673,N_3437,N_3539);
nand U3674 (N_3674,N_3400,N_3590);
nor U3675 (N_3675,N_3559,N_3484);
nor U3676 (N_3676,N_3487,N_3434);
or U3677 (N_3677,N_3597,N_3586);
xnor U3678 (N_3678,N_3415,N_3422);
and U3679 (N_3679,N_3494,N_3452);
and U3680 (N_3680,N_3421,N_3448);
and U3681 (N_3681,N_3455,N_3567);
xnor U3682 (N_3682,N_3489,N_3427);
xor U3683 (N_3683,N_3406,N_3459);
or U3684 (N_3684,N_3575,N_3424);
or U3685 (N_3685,N_3520,N_3527);
or U3686 (N_3686,N_3409,N_3542);
and U3687 (N_3687,N_3475,N_3541);
and U3688 (N_3688,N_3444,N_3414);
xnor U3689 (N_3689,N_3528,N_3548);
xnor U3690 (N_3690,N_3502,N_3524);
or U3691 (N_3691,N_3451,N_3499);
nor U3692 (N_3692,N_3563,N_3522);
nand U3693 (N_3693,N_3462,N_3505);
or U3694 (N_3694,N_3576,N_3486);
xnor U3695 (N_3695,N_3463,N_3468);
nor U3696 (N_3696,N_3574,N_3440);
nand U3697 (N_3697,N_3435,N_3551);
xor U3698 (N_3698,N_3408,N_3545);
xnor U3699 (N_3699,N_3519,N_3481);
nand U3700 (N_3700,N_3416,N_3534);
and U3701 (N_3701,N_3472,N_3440);
xnor U3702 (N_3702,N_3450,N_3536);
nand U3703 (N_3703,N_3595,N_3445);
nand U3704 (N_3704,N_3521,N_3481);
xor U3705 (N_3705,N_3511,N_3463);
xnor U3706 (N_3706,N_3449,N_3484);
nand U3707 (N_3707,N_3509,N_3529);
xor U3708 (N_3708,N_3569,N_3446);
nor U3709 (N_3709,N_3525,N_3460);
nand U3710 (N_3710,N_3589,N_3505);
or U3711 (N_3711,N_3466,N_3447);
nand U3712 (N_3712,N_3433,N_3555);
xnor U3713 (N_3713,N_3577,N_3475);
and U3714 (N_3714,N_3569,N_3421);
and U3715 (N_3715,N_3487,N_3514);
or U3716 (N_3716,N_3473,N_3434);
and U3717 (N_3717,N_3595,N_3442);
and U3718 (N_3718,N_3404,N_3462);
and U3719 (N_3719,N_3529,N_3514);
nand U3720 (N_3720,N_3549,N_3485);
xor U3721 (N_3721,N_3511,N_3428);
and U3722 (N_3722,N_3414,N_3564);
xor U3723 (N_3723,N_3444,N_3437);
nand U3724 (N_3724,N_3444,N_3463);
or U3725 (N_3725,N_3429,N_3514);
nor U3726 (N_3726,N_3425,N_3406);
xor U3727 (N_3727,N_3463,N_3493);
or U3728 (N_3728,N_3494,N_3582);
nand U3729 (N_3729,N_3471,N_3430);
nor U3730 (N_3730,N_3585,N_3405);
nand U3731 (N_3731,N_3436,N_3555);
and U3732 (N_3732,N_3491,N_3582);
nand U3733 (N_3733,N_3587,N_3467);
nand U3734 (N_3734,N_3462,N_3439);
nand U3735 (N_3735,N_3591,N_3549);
nand U3736 (N_3736,N_3567,N_3542);
and U3737 (N_3737,N_3425,N_3554);
or U3738 (N_3738,N_3589,N_3420);
or U3739 (N_3739,N_3414,N_3529);
xor U3740 (N_3740,N_3475,N_3486);
nand U3741 (N_3741,N_3488,N_3564);
nor U3742 (N_3742,N_3400,N_3493);
nand U3743 (N_3743,N_3486,N_3562);
xor U3744 (N_3744,N_3481,N_3518);
nor U3745 (N_3745,N_3403,N_3532);
and U3746 (N_3746,N_3592,N_3425);
nor U3747 (N_3747,N_3510,N_3501);
or U3748 (N_3748,N_3475,N_3436);
xnor U3749 (N_3749,N_3435,N_3511);
nor U3750 (N_3750,N_3423,N_3453);
or U3751 (N_3751,N_3587,N_3479);
nor U3752 (N_3752,N_3415,N_3588);
or U3753 (N_3753,N_3546,N_3519);
nor U3754 (N_3754,N_3411,N_3429);
nand U3755 (N_3755,N_3489,N_3440);
xnor U3756 (N_3756,N_3574,N_3527);
nor U3757 (N_3757,N_3405,N_3448);
and U3758 (N_3758,N_3406,N_3469);
xnor U3759 (N_3759,N_3538,N_3560);
and U3760 (N_3760,N_3585,N_3598);
nor U3761 (N_3761,N_3536,N_3571);
nor U3762 (N_3762,N_3453,N_3435);
and U3763 (N_3763,N_3547,N_3595);
or U3764 (N_3764,N_3518,N_3580);
xor U3765 (N_3765,N_3439,N_3486);
xor U3766 (N_3766,N_3585,N_3590);
nor U3767 (N_3767,N_3462,N_3598);
and U3768 (N_3768,N_3426,N_3436);
xnor U3769 (N_3769,N_3536,N_3487);
nand U3770 (N_3770,N_3551,N_3505);
and U3771 (N_3771,N_3553,N_3538);
nor U3772 (N_3772,N_3506,N_3500);
and U3773 (N_3773,N_3419,N_3562);
and U3774 (N_3774,N_3568,N_3559);
or U3775 (N_3775,N_3416,N_3503);
nand U3776 (N_3776,N_3494,N_3414);
nand U3777 (N_3777,N_3586,N_3463);
nand U3778 (N_3778,N_3590,N_3408);
nor U3779 (N_3779,N_3445,N_3479);
xor U3780 (N_3780,N_3424,N_3585);
and U3781 (N_3781,N_3582,N_3570);
nor U3782 (N_3782,N_3557,N_3490);
xor U3783 (N_3783,N_3526,N_3486);
xnor U3784 (N_3784,N_3547,N_3590);
nand U3785 (N_3785,N_3433,N_3483);
nand U3786 (N_3786,N_3557,N_3416);
xnor U3787 (N_3787,N_3557,N_3508);
and U3788 (N_3788,N_3458,N_3533);
nor U3789 (N_3789,N_3488,N_3461);
and U3790 (N_3790,N_3518,N_3529);
nand U3791 (N_3791,N_3562,N_3533);
nor U3792 (N_3792,N_3456,N_3409);
nor U3793 (N_3793,N_3475,N_3449);
xnor U3794 (N_3794,N_3425,N_3545);
xor U3795 (N_3795,N_3564,N_3535);
xor U3796 (N_3796,N_3438,N_3455);
xor U3797 (N_3797,N_3555,N_3503);
or U3798 (N_3798,N_3461,N_3414);
nand U3799 (N_3799,N_3419,N_3539);
nor U3800 (N_3800,N_3683,N_3756);
nor U3801 (N_3801,N_3650,N_3717);
xnor U3802 (N_3802,N_3671,N_3730);
xnor U3803 (N_3803,N_3727,N_3762);
and U3804 (N_3804,N_3697,N_3720);
and U3805 (N_3805,N_3644,N_3773);
xnor U3806 (N_3806,N_3696,N_3793);
and U3807 (N_3807,N_3783,N_3654);
nor U3808 (N_3808,N_3629,N_3739);
and U3809 (N_3809,N_3675,N_3797);
nand U3810 (N_3810,N_3642,N_3602);
nor U3811 (N_3811,N_3663,N_3632);
or U3812 (N_3812,N_3687,N_3798);
nand U3813 (N_3813,N_3634,N_3627);
nor U3814 (N_3814,N_3630,N_3778);
xor U3815 (N_3815,N_3626,N_3685);
nand U3816 (N_3816,N_3728,N_3677);
or U3817 (N_3817,N_3693,N_3624);
xnor U3818 (N_3818,N_3600,N_3708);
nand U3819 (N_3819,N_3705,N_3787);
nor U3820 (N_3820,N_3726,N_3615);
nor U3821 (N_3821,N_3784,N_3755);
and U3822 (N_3822,N_3741,N_3712);
nor U3823 (N_3823,N_3698,N_3651);
nor U3824 (N_3824,N_3733,N_3790);
nand U3825 (N_3825,N_3657,N_3635);
xor U3826 (N_3826,N_3640,N_3611);
and U3827 (N_3827,N_3767,N_3723);
or U3828 (N_3828,N_3788,N_3659);
nand U3829 (N_3829,N_3606,N_3758);
nand U3830 (N_3830,N_3732,N_3740);
or U3831 (N_3831,N_3751,N_3777);
or U3832 (N_3832,N_3770,N_3753);
xnor U3833 (N_3833,N_3669,N_3704);
nor U3834 (N_3834,N_3625,N_3795);
nor U3835 (N_3835,N_3769,N_3631);
nor U3836 (N_3836,N_3721,N_3713);
xnor U3837 (N_3837,N_3614,N_3724);
nor U3838 (N_3838,N_3765,N_3668);
or U3839 (N_3839,N_3662,N_3621);
nand U3840 (N_3840,N_3707,N_3716);
and U3841 (N_3841,N_3672,N_3792);
xnor U3842 (N_3842,N_3609,N_3676);
nor U3843 (N_3843,N_3618,N_3749);
xor U3844 (N_3844,N_3619,N_3620);
or U3845 (N_3845,N_3617,N_3735);
xor U3846 (N_3846,N_3737,N_3639);
xnor U3847 (N_3847,N_3745,N_3791);
and U3848 (N_3848,N_3776,N_3694);
and U3849 (N_3849,N_3743,N_3691);
and U3850 (N_3850,N_3695,N_3628);
nor U3851 (N_3851,N_3763,N_3656);
nor U3852 (N_3852,N_3768,N_3718);
or U3853 (N_3853,N_3796,N_3710);
or U3854 (N_3854,N_3754,N_3670);
xnor U3855 (N_3855,N_3766,N_3667);
nand U3856 (N_3856,N_3701,N_3623);
nand U3857 (N_3857,N_3722,N_3771);
nand U3858 (N_3858,N_3608,N_3750);
nor U3859 (N_3859,N_3633,N_3719);
xor U3860 (N_3860,N_3780,N_3748);
nor U3861 (N_3861,N_3782,N_3605);
nand U3862 (N_3862,N_3799,N_3781);
and U3863 (N_3863,N_3764,N_3616);
xnor U3864 (N_3864,N_3678,N_3655);
xnor U3865 (N_3865,N_3729,N_3636);
nor U3866 (N_3866,N_3752,N_3702);
nor U3867 (N_3867,N_3774,N_3607);
or U3868 (N_3868,N_3610,N_3658);
and U3869 (N_3869,N_3601,N_3686);
nor U3870 (N_3870,N_3637,N_3690);
and U3871 (N_3871,N_3736,N_3674);
nand U3872 (N_3872,N_3692,N_3638);
xor U3873 (N_3873,N_3664,N_3682);
and U3874 (N_3874,N_3738,N_3785);
or U3875 (N_3875,N_3725,N_3703);
nand U3876 (N_3876,N_3714,N_3789);
nand U3877 (N_3877,N_3652,N_3679);
and U3878 (N_3878,N_3731,N_3734);
and U3879 (N_3879,N_3760,N_3715);
nor U3880 (N_3880,N_3794,N_3747);
nand U3881 (N_3881,N_3680,N_3706);
and U3882 (N_3882,N_3757,N_3648);
nand U3883 (N_3883,N_3761,N_3673);
nor U3884 (N_3884,N_3688,N_3689);
and U3885 (N_3885,N_3645,N_3775);
xor U3886 (N_3886,N_3699,N_3613);
or U3887 (N_3887,N_3684,N_3661);
and U3888 (N_3888,N_3603,N_3660);
nand U3889 (N_3889,N_3746,N_3759);
xor U3890 (N_3890,N_3709,N_3786);
nor U3891 (N_3891,N_3711,N_3612);
nor U3892 (N_3892,N_3653,N_3649);
nor U3893 (N_3893,N_3779,N_3641);
or U3894 (N_3894,N_3647,N_3744);
or U3895 (N_3895,N_3666,N_3604);
nor U3896 (N_3896,N_3665,N_3772);
or U3897 (N_3897,N_3646,N_3622);
xnor U3898 (N_3898,N_3681,N_3643);
xnor U3899 (N_3899,N_3700,N_3742);
or U3900 (N_3900,N_3613,N_3671);
xnor U3901 (N_3901,N_3622,N_3674);
and U3902 (N_3902,N_3734,N_3697);
xnor U3903 (N_3903,N_3601,N_3637);
nor U3904 (N_3904,N_3684,N_3721);
or U3905 (N_3905,N_3787,N_3724);
or U3906 (N_3906,N_3788,N_3744);
and U3907 (N_3907,N_3728,N_3710);
nor U3908 (N_3908,N_3736,N_3763);
and U3909 (N_3909,N_3641,N_3759);
xnor U3910 (N_3910,N_3773,N_3616);
or U3911 (N_3911,N_3662,N_3632);
or U3912 (N_3912,N_3698,N_3799);
nand U3913 (N_3913,N_3647,N_3621);
or U3914 (N_3914,N_3752,N_3739);
nor U3915 (N_3915,N_3713,N_3707);
or U3916 (N_3916,N_3787,N_3659);
nor U3917 (N_3917,N_3790,N_3723);
and U3918 (N_3918,N_3652,N_3630);
nand U3919 (N_3919,N_3669,N_3637);
and U3920 (N_3920,N_3671,N_3708);
and U3921 (N_3921,N_3737,N_3759);
xnor U3922 (N_3922,N_3680,N_3641);
xnor U3923 (N_3923,N_3782,N_3637);
nand U3924 (N_3924,N_3781,N_3674);
and U3925 (N_3925,N_3602,N_3638);
or U3926 (N_3926,N_3627,N_3715);
xor U3927 (N_3927,N_3770,N_3701);
or U3928 (N_3928,N_3776,N_3714);
xnor U3929 (N_3929,N_3600,N_3710);
nor U3930 (N_3930,N_3711,N_3607);
xnor U3931 (N_3931,N_3669,N_3732);
nor U3932 (N_3932,N_3779,N_3685);
or U3933 (N_3933,N_3726,N_3646);
xnor U3934 (N_3934,N_3696,N_3678);
or U3935 (N_3935,N_3761,N_3611);
nor U3936 (N_3936,N_3678,N_3756);
or U3937 (N_3937,N_3724,N_3768);
and U3938 (N_3938,N_3798,N_3651);
xnor U3939 (N_3939,N_3665,N_3674);
and U3940 (N_3940,N_3710,N_3726);
or U3941 (N_3941,N_3785,N_3755);
xnor U3942 (N_3942,N_3709,N_3633);
nand U3943 (N_3943,N_3729,N_3671);
xnor U3944 (N_3944,N_3623,N_3799);
nand U3945 (N_3945,N_3745,N_3603);
nor U3946 (N_3946,N_3674,N_3663);
nand U3947 (N_3947,N_3636,N_3717);
nand U3948 (N_3948,N_3725,N_3710);
nand U3949 (N_3949,N_3653,N_3705);
nand U3950 (N_3950,N_3747,N_3705);
nand U3951 (N_3951,N_3603,N_3627);
or U3952 (N_3952,N_3718,N_3726);
and U3953 (N_3953,N_3664,N_3636);
or U3954 (N_3954,N_3730,N_3694);
and U3955 (N_3955,N_3785,N_3631);
nand U3956 (N_3956,N_3656,N_3698);
or U3957 (N_3957,N_3676,N_3770);
nor U3958 (N_3958,N_3732,N_3624);
and U3959 (N_3959,N_3774,N_3716);
and U3960 (N_3960,N_3630,N_3690);
nand U3961 (N_3961,N_3709,N_3624);
or U3962 (N_3962,N_3606,N_3627);
xor U3963 (N_3963,N_3796,N_3714);
xnor U3964 (N_3964,N_3613,N_3774);
and U3965 (N_3965,N_3655,N_3646);
and U3966 (N_3966,N_3666,N_3791);
and U3967 (N_3967,N_3759,N_3610);
nor U3968 (N_3968,N_3693,N_3742);
or U3969 (N_3969,N_3695,N_3618);
nor U3970 (N_3970,N_3784,N_3604);
or U3971 (N_3971,N_3733,N_3747);
nor U3972 (N_3972,N_3751,N_3768);
nor U3973 (N_3973,N_3743,N_3625);
nand U3974 (N_3974,N_3712,N_3748);
xor U3975 (N_3975,N_3674,N_3779);
nor U3976 (N_3976,N_3720,N_3610);
and U3977 (N_3977,N_3739,N_3691);
xnor U3978 (N_3978,N_3603,N_3615);
and U3979 (N_3979,N_3628,N_3663);
or U3980 (N_3980,N_3736,N_3774);
or U3981 (N_3981,N_3648,N_3713);
nand U3982 (N_3982,N_3733,N_3766);
and U3983 (N_3983,N_3770,N_3602);
and U3984 (N_3984,N_3624,N_3741);
or U3985 (N_3985,N_3786,N_3604);
xor U3986 (N_3986,N_3720,N_3712);
xor U3987 (N_3987,N_3738,N_3643);
xor U3988 (N_3988,N_3755,N_3667);
nand U3989 (N_3989,N_3758,N_3728);
nor U3990 (N_3990,N_3715,N_3757);
nor U3991 (N_3991,N_3783,N_3630);
or U3992 (N_3992,N_3783,N_3784);
nand U3993 (N_3993,N_3614,N_3633);
nand U3994 (N_3994,N_3739,N_3725);
or U3995 (N_3995,N_3728,N_3683);
or U3996 (N_3996,N_3650,N_3655);
or U3997 (N_3997,N_3674,N_3724);
xnor U3998 (N_3998,N_3643,N_3665);
and U3999 (N_3999,N_3684,N_3743);
or U4000 (N_4000,N_3877,N_3976);
nor U4001 (N_4001,N_3853,N_3991);
nand U4002 (N_4002,N_3829,N_3827);
nor U4003 (N_4003,N_3905,N_3859);
nor U4004 (N_4004,N_3898,N_3843);
nor U4005 (N_4005,N_3884,N_3803);
xnor U4006 (N_4006,N_3917,N_3994);
and U4007 (N_4007,N_3927,N_3995);
nand U4008 (N_4008,N_3990,N_3825);
nor U4009 (N_4009,N_3801,N_3894);
nand U4010 (N_4010,N_3868,N_3960);
nor U4011 (N_4011,N_3914,N_3890);
or U4012 (N_4012,N_3984,N_3831);
and U4013 (N_4013,N_3924,N_3883);
and U4014 (N_4014,N_3922,N_3981);
nor U4015 (N_4015,N_3849,N_3959);
or U4016 (N_4016,N_3904,N_3919);
or U4017 (N_4017,N_3972,N_3806);
nor U4018 (N_4018,N_3968,N_3974);
xnor U4019 (N_4019,N_3839,N_3891);
xnor U4020 (N_4020,N_3973,N_3941);
and U4021 (N_4021,N_3886,N_3881);
and U4022 (N_4022,N_3808,N_3841);
nand U4023 (N_4023,N_3949,N_3889);
and U4024 (N_4024,N_3809,N_3888);
nor U4025 (N_4025,N_3899,N_3921);
or U4026 (N_4026,N_3817,N_3937);
or U4027 (N_4027,N_3842,N_3856);
nand U4028 (N_4028,N_3908,N_3854);
xnor U4029 (N_4029,N_3861,N_3875);
nor U4030 (N_4030,N_3804,N_3978);
nand U4031 (N_4031,N_3931,N_3869);
xnor U4032 (N_4032,N_3837,N_3951);
nand U4033 (N_4033,N_3851,N_3993);
or U4034 (N_4034,N_3961,N_3985);
nand U4035 (N_4035,N_3900,N_3971);
nor U4036 (N_4036,N_3925,N_3999);
xnor U4037 (N_4037,N_3812,N_3935);
and U4038 (N_4038,N_3864,N_3838);
or U4039 (N_4039,N_3977,N_3901);
nor U4040 (N_4040,N_3873,N_3880);
or U4041 (N_4041,N_3997,N_3926);
and U4042 (N_4042,N_3895,N_3975);
nand U4043 (N_4043,N_3858,N_3867);
nand U4044 (N_4044,N_3987,N_3848);
or U4045 (N_4045,N_3818,N_3969);
and U4046 (N_4046,N_3957,N_3950);
nor U4047 (N_4047,N_3844,N_3902);
nor U4048 (N_4048,N_3930,N_3852);
or U4049 (N_4049,N_3915,N_3826);
nand U4050 (N_4050,N_3910,N_3810);
nand U4051 (N_4051,N_3966,N_3821);
nor U4052 (N_4052,N_3982,N_3897);
nand U4053 (N_4053,N_3929,N_3815);
nor U4054 (N_4054,N_3836,N_3862);
xor U4055 (N_4055,N_3923,N_3807);
xnor U4056 (N_4056,N_3948,N_3980);
xnor U4057 (N_4057,N_3952,N_3866);
xnor U4058 (N_4058,N_3823,N_3945);
and U4059 (N_4059,N_3805,N_3892);
and U4060 (N_4060,N_3824,N_3903);
and U4061 (N_4061,N_3955,N_3863);
nor U4062 (N_4062,N_3833,N_3847);
nand U4063 (N_4063,N_3846,N_3964);
xnor U4064 (N_4064,N_3814,N_3947);
xor U4065 (N_4065,N_3800,N_3822);
nor U4066 (N_4066,N_3944,N_3860);
or U4067 (N_4067,N_3954,N_3970);
xor U4068 (N_4068,N_3936,N_3958);
or U4069 (N_4069,N_3934,N_3878);
nor U4070 (N_4070,N_3988,N_3992);
or U4071 (N_4071,N_3946,N_3874);
and U4072 (N_4072,N_3855,N_3893);
nor U4073 (N_4073,N_3835,N_3906);
or U4074 (N_4074,N_3940,N_3870);
nand U4075 (N_4075,N_3820,N_3998);
or U4076 (N_4076,N_3965,N_3887);
and U4077 (N_4077,N_3996,N_3879);
xor U4078 (N_4078,N_3967,N_3933);
and U4079 (N_4079,N_3909,N_3896);
nand U4080 (N_4080,N_3850,N_3939);
nand U4081 (N_4081,N_3865,N_3832);
and U4082 (N_4082,N_3962,N_3907);
or U4083 (N_4083,N_3834,N_3885);
or U4084 (N_4084,N_3912,N_3871);
xor U4085 (N_4085,N_3811,N_3918);
nor U4086 (N_4086,N_3857,N_3956);
nand U4087 (N_4087,N_3989,N_3943);
nor U4088 (N_4088,N_3942,N_3845);
or U4089 (N_4089,N_3979,N_3816);
or U4090 (N_4090,N_3876,N_3840);
nor U4091 (N_4091,N_3963,N_3938);
or U4092 (N_4092,N_3986,N_3911);
and U4093 (N_4093,N_3819,N_3882);
and U4094 (N_4094,N_3916,N_3813);
or U4095 (N_4095,N_3828,N_3932);
or U4096 (N_4096,N_3928,N_3913);
and U4097 (N_4097,N_3920,N_3872);
xnor U4098 (N_4098,N_3802,N_3830);
nand U4099 (N_4099,N_3953,N_3983);
nand U4100 (N_4100,N_3933,N_3982);
nand U4101 (N_4101,N_3988,N_3872);
nor U4102 (N_4102,N_3906,N_3905);
and U4103 (N_4103,N_3922,N_3990);
nor U4104 (N_4104,N_3997,N_3915);
or U4105 (N_4105,N_3803,N_3950);
nand U4106 (N_4106,N_3905,N_3860);
and U4107 (N_4107,N_3891,N_3985);
and U4108 (N_4108,N_3948,N_3999);
nor U4109 (N_4109,N_3962,N_3958);
nor U4110 (N_4110,N_3825,N_3979);
and U4111 (N_4111,N_3929,N_3908);
and U4112 (N_4112,N_3957,N_3922);
and U4113 (N_4113,N_3948,N_3818);
xor U4114 (N_4114,N_3956,N_3901);
nor U4115 (N_4115,N_3884,N_3975);
xnor U4116 (N_4116,N_3827,N_3944);
and U4117 (N_4117,N_3801,N_3980);
nor U4118 (N_4118,N_3960,N_3917);
xnor U4119 (N_4119,N_3994,N_3901);
and U4120 (N_4120,N_3931,N_3811);
or U4121 (N_4121,N_3816,N_3872);
nand U4122 (N_4122,N_3950,N_3921);
and U4123 (N_4123,N_3881,N_3893);
nor U4124 (N_4124,N_3904,N_3906);
xnor U4125 (N_4125,N_3813,N_3957);
or U4126 (N_4126,N_3805,N_3821);
xor U4127 (N_4127,N_3982,N_3996);
nor U4128 (N_4128,N_3992,N_3828);
or U4129 (N_4129,N_3923,N_3904);
nand U4130 (N_4130,N_3961,N_3998);
or U4131 (N_4131,N_3925,N_3857);
nand U4132 (N_4132,N_3950,N_3859);
and U4133 (N_4133,N_3958,N_3881);
nand U4134 (N_4134,N_3976,N_3806);
and U4135 (N_4135,N_3911,N_3865);
and U4136 (N_4136,N_3936,N_3978);
nor U4137 (N_4137,N_3995,N_3875);
xor U4138 (N_4138,N_3994,N_3836);
and U4139 (N_4139,N_3853,N_3940);
nand U4140 (N_4140,N_3803,N_3998);
and U4141 (N_4141,N_3904,N_3841);
and U4142 (N_4142,N_3909,N_3820);
or U4143 (N_4143,N_3961,N_3831);
nand U4144 (N_4144,N_3934,N_3914);
xor U4145 (N_4145,N_3909,N_3836);
and U4146 (N_4146,N_3858,N_3893);
and U4147 (N_4147,N_3990,N_3811);
xor U4148 (N_4148,N_3977,N_3984);
and U4149 (N_4149,N_3960,N_3944);
nor U4150 (N_4150,N_3917,N_3885);
nor U4151 (N_4151,N_3927,N_3810);
and U4152 (N_4152,N_3961,N_3860);
or U4153 (N_4153,N_3891,N_3972);
xor U4154 (N_4154,N_3928,N_3979);
nand U4155 (N_4155,N_3928,N_3898);
or U4156 (N_4156,N_3843,N_3890);
nor U4157 (N_4157,N_3929,N_3894);
xor U4158 (N_4158,N_3827,N_3973);
nand U4159 (N_4159,N_3822,N_3977);
and U4160 (N_4160,N_3980,N_3878);
and U4161 (N_4161,N_3912,N_3973);
and U4162 (N_4162,N_3867,N_3971);
or U4163 (N_4163,N_3994,N_3835);
and U4164 (N_4164,N_3903,N_3835);
nand U4165 (N_4165,N_3837,N_3807);
and U4166 (N_4166,N_3850,N_3847);
and U4167 (N_4167,N_3991,N_3983);
xor U4168 (N_4168,N_3809,N_3814);
and U4169 (N_4169,N_3883,N_3984);
xnor U4170 (N_4170,N_3889,N_3930);
or U4171 (N_4171,N_3883,N_3843);
or U4172 (N_4172,N_3849,N_3917);
xnor U4173 (N_4173,N_3800,N_3959);
nor U4174 (N_4174,N_3909,N_3920);
nor U4175 (N_4175,N_3954,N_3887);
xnor U4176 (N_4176,N_3849,N_3998);
nand U4177 (N_4177,N_3953,N_3851);
nor U4178 (N_4178,N_3879,N_3881);
xor U4179 (N_4179,N_3914,N_3989);
and U4180 (N_4180,N_3883,N_3818);
or U4181 (N_4181,N_3846,N_3851);
or U4182 (N_4182,N_3829,N_3812);
nor U4183 (N_4183,N_3877,N_3871);
and U4184 (N_4184,N_3994,N_3980);
or U4185 (N_4185,N_3953,N_3934);
nor U4186 (N_4186,N_3911,N_3993);
nand U4187 (N_4187,N_3876,N_3915);
nor U4188 (N_4188,N_3957,N_3823);
nor U4189 (N_4189,N_3873,N_3980);
and U4190 (N_4190,N_3905,N_3977);
nor U4191 (N_4191,N_3837,N_3966);
nor U4192 (N_4192,N_3820,N_3852);
nand U4193 (N_4193,N_3813,N_3935);
xnor U4194 (N_4194,N_3983,N_3920);
xnor U4195 (N_4195,N_3988,N_3931);
nand U4196 (N_4196,N_3996,N_3914);
xor U4197 (N_4197,N_3808,N_3899);
nor U4198 (N_4198,N_3828,N_3841);
or U4199 (N_4199,N_3809,N_3874);
nand U4200 (N_4200,N_4019,N_4029);
nor U4201 (N_4201,N_4174,N_4152);
nor U4202 (N_4202,N_4132,N_4162);
nand U4203 (N_4203,N_4054,N_4065);
nand U4204 (N_4204,N_4072,N_4192);
nor U4205 (N_4205,N_4038,N_4058);
nand U4206 (N_4206,N_4000,N_4002);
nor U4207 (N_4207,N_4024,N_4083);
nor U4208 (N_4208,N_4167,N_4067);
nor U4209 (N_4209,N_4124,N_4149);
and U4210 (N_4210,N_4120,N_4033);
nand U4211 (N_4211,N_4096,N_4143);
xnor U4212 (N_4212,N_4118,N_4094);
nor U4213 (N_4213,N_4056,N_4111);
or U4214 (N_4214,N_4112,N_4098);
and U4215 (N_4215,N_4077,N_4177);
nand U4216 (N_4216,N_4106,N_4166);
or U4217 (N_4217,N_4133,N_4171);
or U4218 (N_4218,N_4046,N_4031);
xnor U4219 (N_4219,N_4105,N_4178);
or U4220 (N_4220,N_4059,N_4087);
and U4221 (N_4221,N_4146,N_4119);
xnor U4222 (N_4222,N_4104,N_4006);
nand U4223 (N_4223,N_4023,N_4176);
and U4224 (N_4224,N_4041,N_4088);
xor U4225 (N_4225,N_4109,N_4130);
or U4226 (N_4226,N_4020,N_4183);
nor U4227 (N_4227,N_4026,N_4122);
xor U4228 (N_4228,N_4001,N_4062);
and U4229 (N_4229,N_4158,N_4060);
and U4230 (N_4230,N_4103,N_4173);
nand U4231 (N_4231,N_4199,N_4147);
nand U4232 (N_4232,N_4014,N_4057);
nor U4233 (N_4233,N_4049,N_4193);
nor U4234 (N_4234,N_4125,N_4044);
or U4235 (N_4235,N_4194,N_4078);
nor U4236 (N_4236,N_4101,N_4117);
nor U4237 (N_4237,N_4074,N_4114);
nor U4238 (N_4238,N_4028,N_4022);
and U4239 (N_4239,N_4195,N_4172);
nand U4240 (N_4240,N_4186,N_4136);
nand U4241 (N_4241,N_4076,N_4090);
nor U4242 (N_4242,N_4055,N_4005);
nor U4243 (N_4243,N_4003,N_4021);
and U4244 (N_4244,N_4126,N_4017);
or U4245 (N_4245,N_4196,N_4155);
nand U4246 (N_4246,N_4025,N_4018);
or U4247 (N_4247,N_4154,N_4053);
nor U4248 (N_4248,N_4165,N_4036);
nand U4249 (N_4249,N_4063,N_4181);
and U4250 (N_4250,N_4160,N_4068);
nand U4251 (N_4251,N_4004,N_4008);
or U4252 (N_4252,N_4045,N_4188);
nor U4253 (N_4253,N_4108,N_4048);
nand U4254 (N_4254,N_4051,N_4140);
and U4255 (N_4255,N_4086,N_4010);
nor U4256 (N_4256,N_4157,N_4121);
xor U4257 (N_4257,N_4137,N_4161);
xnor U4258 (N_4258,N_4159,N_4082);
nand U4259 (N_4259,N_4070,N_4073);
or U4260 (N_4260,N_4071,N_4189);
or U4261 (N_4261,N_4131,N_4197);
nand U4262 (N_4262,N_4135,N_4097);
or U4263 (N_4263,N_4035,N_4179);
xnor U4264 (N_4264,N_4175,N_4061);
nand U4265 (N_4265,N_4148,N_4011);
xnor U4266 (N_4266,N_4156,N_4037);
and U4267 (N_4267,N_4184,N_4187);
nand U4268 (N_4268,N_4050,N_4134);
nand U4269 (N_4269,N_4182,N_4151);
and U4270 (N_4270,N_4030,N_4039);
nor U4271 (N_4271,N_4169,N_4064);
and U4272 (N_4272,N_4084,N_4142);
or U4273 (N_4273,N_4127,N_4081);
nand U4274 (N_4274,N_4040,N_4164);
or U4275 (N_4275,N_4091,N_4047);
and U4276 (N_4276,N_4027,N_4052);
nand U4277 (N_4277,N_4123,N_4128);
nand U4278 (N_4278,N_4163,N_4190);
nor U4279 (N_4279,N_4080,N_4107);
nand U4280 (N_4280,N_4069,N_4079);
or U4281 (N_4281,N_4042,N_4099);
xor U4282 (N_4282,N_4145,N_4129);
nor U4283 (N_4283,N_4113,N_4141);
and U4284 (N_4284,N_4102,N_4150);
or U4285 (N_4285,N_4092,N_4180);
and U4286 (N_4286,N_4144,N_4115);
xor U4287 (N_4287,N_4153,N_4093);
nand U4288 (N_4288,N_4013,N_4009);
nor U4289 (N_4289,N_4116,N_4085);
nor U4290 (N_4290,N_4032,N_4015);
or U4291 (N_4291,N_4138,N_4016);
or U4292 (N_4292,N_4100,N_4191);
nor U4293 (N_4293,N_4198,N_4095);
nand U4294 (N_4294,N_4007,N_4110);
and U4295 (N_4295,N_4139,N_4066);
or U4296 (N_4296,N_4089,N_4034);
or U4297 (N_4297,N_4043,N_4185);
or U4298 (N_4298,N_4170,N_4168);
nor U4299 (N_4299,N_4012,N_4075);
and U4300 (N_4300,N_4180,N_4046);
xnor U4301 (N_4301,N_4180,N_4045);
nand U4302 (N_4302,N_4031,N_4028);
nor U4303 (N_4303,N_4145,N_4070);
xnor U4304 (N_4304,N_4115,N_4197);
nor U4305 (N_4305,N_4124,N_4074);
or U4306 (N_4306,N_4056,N_4093);
nor U4307 (N_4307,N_4129,N_4038);
nor U4308 (N_4308,N_4188,N_4110);
and U4309 (N_4309,N_4028,N_4122);
nand U4310 (N_4310,N_4083,N_4053);
or U4311 (N_4311,N_4139,N_4163);
and U4312 (N_4312,N_4029,N_4063);
and U4313 (N_4313,N_4101,N_4150);
xor U4314 (N_4314,N_4179,N_4119);
and U4315 (N_4315,N_4131,N_4186);
xnor U4316 (N_4316,N_4062,N_4104);
xnor U4317 (N_4317,N_4034,N_4039);
and U4318 (N_4318,N_4132,N_4024);
nor U4319 (N_4319,N_4047,N_4176);
nor U4320 (N_4320,N_4186,N_4110);
or U4321 (N_4321,N_4191,N_4085);
xnor U4322 (N_4322,N_4011,N_4049);
nand U4323 (N_4323,N_4141,N_4190);
and U4324 (N_4324,N_4016,N_4090);
nor U4325 (N_4325,N_4029,N_4163);
nor U4326 (N_4326,N_4078,N_4099);
nor U4327 (N_4327,N_4165,N_4091);
and U4328 (N_4328,N_4041,N_4195);
nor U4329 (N_4329,N_4197,N_4129);
nor U4330 (N_4330,N_4179,N_4070);
or U4331 (N_4331,N_4175,N_4142);
and U4332 (N_4332,N_4156,N_4086);
or U4333 (N_4333,N_4000,N_4117);
xnor U4334 (N_4334,N_4061,N_4051);
or U4335 (N_4335,N_4049,N_4051);
nor U4336 (N_4336,N_4160,N_4138);
and U4337 (N_4337,N_4126,N_4016);
or U4338 (N_4338,N_4160,N_4019);
nor U4339 (N_4339,N_4016,N_4150);
xnor U4340 (N_4340,N_4085,N_4163);
nand U4341 (N_4341,N_4027,N_4000);
or U4342 (N_4342,N_4109,N_4145);
and U4343 (N_4343,N_4057,N_4146);
xnor U4344 (N_4344,N_4151,N_4064);
and U4345 (N_4345,N_4130,N_4125);
or U4346 (N_4346,N_4030,N_4014);
and U4347 (N_4347,N_4024,N_4115);
and U4348 (N_4348,N_4156,N_4059);
and U4349 (N_4349,N_4152,N_4117);
xor U4350 (N_4350,N_4015,N_4133);
nor U4351 (N_4351,N_4016,N_4160);
nor U4352 (N_4352,N_4161,N_4006);
or U4353 (N_4353,N_4178,N_4180);
xor U4354 (N_4354,N_4066,N_4046);
and U4355 (N_4355,N_4075,N_4010);
nor U4356 (N_4356,N_4075,N_4143);
and U4357 (N_4357,N_4018,N_4031);
xnor U4358 (N_4358,N_4038,N_4116);
nor U4359 (N_4359,N_4168,N_4119);
or U4360 (N_4360,N_4013,N_4143);
nand U4361 (N_4361,N_4058,N_4096);
and U4362 (N_4362,N_4062,N_4170);
or U4363 (N_4363,N_4152,N_4123);
nor U4364 (N_4364,N_4156,N_4094);
and U4365 (N_4365,N_4072,N_4146);
or U4366 (N_4366,N_4089,N_4168);
and U4367 (N_4367,N_4139,N_4116);
xnor U4368 (N_4368,N_4080,N_4015);
or U4369 (N_4369,N_4132,N_4198);
nor U4370 (N_4370,N_4165,N_4093);
nor U4371 (N_4371,N_4063,N_4159);
xor U4372 (N_4372,N_4084,N_4196);
nor U4373 (N_4373,N_4102,N_4125);
or U4374 (N_4374,N_4171,N_4100);
nor U4375 (N_4375,N_4018,N_4070);
or U4376 (N_4376,N_4123,N_4074);
nor U4377 (N_4377,N_4104,N_4093);
nor U4378 (N_4378,N_4175,N_4171);
xnor U4379 (N_4379,N_4002,N_4182);
and U4380 (N_4380,N_4151,N_4032);
and U4381 (N_4381,N_4017,N_4187);
and U4382 (N_4382,N_4154,N_4036);
and U4383 (N_4383,N_4099,N_4197);
xor U4384 (N_4384,N_4073,N_4055);
and U4385 (N_4385,N_4090,N_4195);
nor U4386 (N_4386,N_4137,N_4086);
nor U4387 (N_4387,N_4160,N_4141);
xnor U4388 (N_4388,N_4094,N_4022);
xor U4389 (N_4389,N_4090,N_4132);
and U4390 (N_4390,N_4187,N_4118);
and U4391 (N_4391,N_4151,N_4149);
nor U4392 (N_4392,N_4019,N_4012);
or U4393 (N_4393,N_4031,N_4016);
and U4394 (N_4394,N_4132,N_4026);
or U4395 (N_4395,N_4030,N_4150);
or U4396 (N_4396,N_4053,N_4162);
or U4397 (N_4397,N_4166,N_4062);
nand U4398 (N_4398,N_4006,N_4119);
nand U4399 (N_4399,N_4120,N_4129);
or U4400 (N_4400,N_4372,N_4221);
xor U4401 (N_4401,N_4252,N_4293);
xnor U4402 (N_4402,N_4310,N_4202);
and U4403 (N_4403,N_4235,N_4318);
xnor U4404 (N_4404,N_4374,N_4237);
and U4405 (N_4405,N_4383,N_4268);
nor U4406 (N_4406,N_4258,N_4327);
or U4407 (N_4407,N_4342,N_4377);
xor U4408 (N_4408,N_4204,N_4364);
and U4409 (N_4409,N_4236,N_4322);
nor U4410 (N_4410,N_4270,N_4307);
xor U4411 (N_4411,N_4203,N_4287);
nand U4412 (N_4412,N_4304,N_4217);
xor U4413 (N_4413,N_4321,N_4314);
or U4414 (N_4414,N_4373,N_4345);
nor U4415 (N_4415,N_4295,N_4357);
and U4416 (N_4416,N_4256,N_4257);
nand U4417 (N_4417,N_4246,N_4389);
nor U4418 (N_4418,N_4245,N_4278);
and U4419 (N_4419,N_4382,N_4206);
and U4420 (N_4420,N_4209,N_4396);
and U4421 (N_4421,N_4264,N_4296);
nand U4422 (N_4422,N_4274,N_4326);
nor U4423 (N_4423,N_4343,N_4335);
nand U4424 (N_4424,N_4338,N_4341);
nor U4425 (N_4425,N_4375,N_4255);
nor U4426 (N_4426,N_4360,N_4240);
or U4427 (N_4427,N_4228,N_4350);
xor U4428 (N_4428,N_4398,N_4379);
and U4429 (N_4429,N_4297,N_4356);
nand U4430 (N_4430,N_4311,N_4312);
xor U4431 (N_4431,N_4349,N_4271);
or U4432 (N_4432,N_4239,N_4336);
xor U4433 (N_4433,N_4220,N_4390);
nor U4434 (N_4434,N_4251,N_4242);
nor U4435 (N_4435,N_4368,N_4201);
xor U4436 (N_4436,N_4225,N_4316);
nor U4437 (N_4437,N_4254,N_4320);
and U4438 (N_4438,N_4393,N_4354);
and U4439 (N_4439,N_4391,N_4294);
nor U4440 (N_4440,N_4285,N_4283);
or U4441 (N_4441,N_4248,N_4230);
xor U4442 (N_4442,N_4244,N_4232);
nor U4443 (N_4443,N_4308,N_4234);
nor U4444 (N_4444,N_4212,N_4381);
nor U4445 (N_4445,N_4331,N_4333);
nor U4446 (N_4446,N_4284,N_4323);
and U4447 (N_4447,N_4369,N_4250);
nor U4448 (N_4448,N_4395,N_4227);
nor U4449 (N_4449,N_4328,N_4309);
or U4450 (N_4450,N_4371,N_4388);
xnor U4451 (N_4451,N_4306,N_4397);
and U4452 (N_4452,N_4200,N_4215);
or U4453 (N_4453,N_4226,N_4213);
and U4454 (N_4454,N_4365,N_4280);
xnor U4455 (N_4455,N_4399,N_4261);
and U4456 (N_4456,N_4359,N_4394);
xor U4457 (N_4457,N_4259,N_4224);
xnor U4458 (N_4458,N_4355,N_4288);
nor U4459 (N_4459,N_4281,N_4231);
or U4460 (N_4460,N_4247,N_4214);
nor U4461 (N_4461,N_4313,N_4299);
or U4462 (N_4462,N_4292,N_4253);
nor U4463 (N_4463,N_4301,N_4273);
xnor U4464 (N_4464,N_4269,N_4208);
nand U4465 (N_4465,N_4210,N_4303);
nand U4466 (N_4466,N_4305,N_4367);
nand U4467 (N_4467,N_4218,N_4380);
xor U4468 (N_4468,N_4386,N_4263);
and U4469 (N_4469,N_4222,N_4219);
nand U4470 (N_4470,N_4233,N_4286);
and U4471 (N_4471,N_4358,N_4211);
xor U4472 (N_4472,N_4347,N_4229);
and U4473 (N_4473,N_4366,N_4339);
xnor U4474 (N_4474,N_4262,N_4282);
nor U4475 (N_4475,N_4291,N_4329);
xnor U4476 (N_4476,N_4376,N_4205);
xor U4477 (N_4477,N_4385,N_4249);
nand U4478 (N_4478,N_4279,N_4351);
xor U4479 (N_4479,N_4216,N_4241);
nand U4480 (N_4480,N_4207,N_4378);
nand U4481 (N_4481,N_4277,N_4346);
nor U4482 (N_4482,N_4289,N_4265);
and U4483 (N_4483,N_4272,N_4266);
nor U4484 (N_4484,N_4317,N_4392);
and U4485 (N_4485,N_4330,N_4223);
and U4486 (N_4486,N_4324,N_4325);
nand U4487 (N_4487,N_4275,N_4298);
and U4488 (N_4488,N_4363,N_4353);
or U4489 (N_4489,N_4238,N_4260);
nand U4490 (N_4490,N_4319,N_4348);
or U4491 (N_4491,N_4387,N_4315);
and U4492 (N_4492,N_4300,N_4340);
xnor U4493 (N_4493,N_4243,N_4362);
nor U4494 (N_4494,N_4352,N_4276);
nor U4495 (N_4495,N_4361,N_4332);
and U4496 (N_4496,N_4370,N_4334);
nor U4497 (N_4497,N_4267,N_4290);
nand U4498 (N_4498,N_4302,N_4337);
xnor U4499 (N_4499,N_4344,N_4384);
and U4500 (N_4500,N_4240,N_4290);
nand U4501 (N_4501,N_4331,N_4261);
or U4502 (N_4502,N_4265,N_4201);
xor U4503 (N_4503,N_4395,N_4397);
and U4504 (N_4504,N_4330,N_4356);
xor U4505 (N_4505,N_4337,N_4324);
or U4506 (N_4506,N_4348,N_4261);
and U4507 (N_4507,N_4289,N_4331);
or U4508 (N_4508,N_4294,N_4375);
nand U4509 (N_4509,N_4234,N_4261);
nor U4510 (N_4510,N_4360,N_4378);
nand U4511 (N_4511,N_4269,N_4363);
or U4512 (N_4512,N_4330,N_4335);
and U4513 (N_4513,N_4255,N_4309);
nor U4514 (N_4514,N_4343,N_4257);
xor U4515 (N_4515,N_4267,N_4291);
nor U4516 (N_4516,N_4225,N_4228);
nor U4517 (N_4517,N_4314,N_4223);
and U4518 (N_4518,N_4273,N_4337);
nand U4519 (N_4519,N_4229,N_4352);
nor U4520 (N_4520,N_4365,N_4287);
nand U4521 (N_4521,N_4297,N_4204);
xor U4522 (N_4522,N_4375,N_4336);
and U4523 (N_4523,N_4228,N_4229);
nand U4524 (N_4524,N_4245,N_4281);
and U4525 (N_4525,N_4233,N_4216);
nor U4526 (N_4526,N_4380,N_4347);
xnor U4527 (N_4527,N_4354,N_4283);
xor U4528 (N_4528,N_4309,N_4241);
nor U4529 (N_4529,N_4284,N_4254);
nand U4530 (N_4530,N_4318,N_4250);
and U4531 (N_4531,N_4254,N_4396);
xnor U4532 (N_4532,N_4273,N_4278);
nand U4533 (N_4533,N_4217,N_4338);
xor U4534 (N_4534,N_4208,N_4329);
xnor U4535 (N_4535,N_4207,N_4375);
nand U4536 (N_4536,N_4231,N_4334);
nor U4537 (N_4537,N_4336,N_4380);
xnor U4538 (N_4538,N_4218,N_4328);
nor U4539 (N_4539,N_4273,N_4256);
and U4540 (N_4540,N_4318,N_4305);
or U4541 (N_4541,N_4316,N_4219);
and U4542 (N_4542,N_4364,N_4253);
nand U4543 (N_4543,N_4340,N_4236);
or U4544 (N_4544,N_4398,N_4233);
and U4545 (N_4545,N_4240,N_4308);
and U4546 (N_4546,N_4310,N_4331);
xnor U4547 (N_4547,N_4251,N_4360);
or U4548 (N_4548,N_4331,N_4270);
xnor U4549 (N_4549,N_4241,N_4277);
nand U4550 (N_4550,N_4270,N_4382);
xor U4551 (N_4551,N_4381,N_4392);
nand U4552 (N_4552,N_4231,N_4261);
and U4553 (N_4553,N_4282,N_4277);
nor U4554 (N_4554,N_4378,N_4290);
nor U4555 (N_4555,N_4245,N_4316);
and U4556 (N_4556,N_4373,N_4355);
nor U4557 (N_4557,N_4340,N_4215);
or U4558 (N_4558,N_4333,N_4365);
and U4559 (N_4559,N_4365,N_4236);
xnor U4560 (N_4560,N_4208,N_4299);
nor U4561 (N_4561,N_4365,N_4242);
and U4562 (N_4562,N_4372,N_4362);
and U4563 (N_4563,N_4355,N_4222);
xnor U4564 (N_4564,N_4257,N_4236);
and U4565 (N_4565,N_4254,N_4228);
and U4566 (N_4566,N_4298,N_4389);
xnor U4567 (N_4567,N_4262,N_4224);
nand U4568 (N_4568,N_4319,N_4399);
and U4569 (N_4569,N_4362,N_4341);
nor U4570 (N_4570,N_4329,N_4287);
and U4571 (N_4571,N_4310,N_4391);
or U4572 (N_4572,N_4271,N_4306);
nand U4573 (N_4573,N_4356,N_4325);
xnor U4574 (N_4574,N_4231,N_4206);
nor U4575 (N_4575,N_4312,N_4318);
nand U4576 (N_4576,N_4311,N_4264);
nor U4577 (N_4577,N_4207,N_4315);
nor U4578 (N_4578,N_4252,N_4257);
or U4579 (N_4579,N_4368,N_4355);
or U4580 (N_4580,N_4278,N_4264);
xor U4581 (N_4581,N_4367,N_4206);
xor U4582 (N_4582,N_4355,N_4369);
or U4583 (N_4583,N_4211,N_4250);
or U4584 (N_4584,N_4269,N_4392);
nand U4585 (N_4585,N_4397,N_4283);
nand U4586 (N_4586,N_4348,N_4239);
xnor U4587 (N_4587,N_4282,N_4244);
nor U4588 (N_4588,N_4273,N_4288);
xor U4589 (N_4589,N_4390,N_4213);
xnor U4590 (N_4590,N_4337,N_4331);
nor U4591 (N_4591,N_4223,N_4382);
nand U4592 (N_4592,N_4213,N_4229);
and U4593 (N_4593,N_4379,N_4282);
and U4594 (N_4594,N_4327,N_4232);
nand U4595 (N_4595,N_4379,N_4318);
xnor U4596 (N_4596,N_4379,N_4244);
and U4597 (N_4597,N_4360,N_4242);
or U4598 (N_4598,N_4238,N_4285);
or U4599 (N_4599,N_4303,N_4397);
xnor U4600 (N_4600,N_4522,N_4523);
xnor U4601 (N_4601,N_4549,N_4457);
or U4602 (N_4602,N_4443,N_4459);
or U4603 (N_4603,N_4560,N_4486);
nand U4604 (N_4604,N_4594,N_4592);
and U4605 (N_4605,N_4510,N_4422);
nor U4606 (N_4606,N_4526,N_4585);
or U4607 (N_4607,N_4410,N_4438);
nand U4608 (N_4608,N_4559,N_4403);
nand U4609 (N_4609,N_4516,N_4412);
and U4610 (N_4610,N_4495,N_4404);
and U4611 (N_4611,N_4481,N_4458);
or U4612 (N_4612,N_4416,N_4465);
xor U4613 (N_4613,N_4553,N_4448);
xnor U4614 (N_4614,N_4445,N_4565);
xor U4615 (N_4615,N_4597,N_4451);
nand U4616 (N_4616,N_4596,N_4591);
nand U4617 (N_4617,N_4444,N_4562);
nand U4618 (N_4618,N_4479,N_4543);
nand U4619 (N_4619,N_4478,N_4452);
or U4620 (N_4620,N_4497,N_4508);
and U4621 (N_4621,N_4558,N_4456);
or U4622 (N_4622,N_4521,N_4493);
and U4623 (N_4623,N_4477,N_4476);
nand U4624 (N_4624,N_4460,N_4566);
and U4625 (N_4625,N_4402,N_4574);
xor U4626 (N_4626,N_4466,N_4506);
nor U4627 (N_4627,N_4524,N_4432);
nand U4628 (N_4628,N_4496,N_4442);
xor U4629 (N_4629,N_4586,N_4408);
or U4630 (N_4630,N_4469,N_4428);
nor U4631 (N_4631,N_4419,N_4576);
xor U4632 (N_4632,N_4482,N_4461);
xor U4633 (N_4633,N_4545,N_4421);
nor U4634 (N_4634,N_4575,N_4552);
xor U4635 (N_4635,N_4449,N_4595);
xor U4636 (N_4636,N_4563,N_4587);
and U4637 (N_4637,N_4401,N_4531);
and U4638 (N_4638,N_4498,N_4567);
or U4639 (N_4639,N_4472,N_4453);
xor U4640 (N_4640,N_4436,N_4546);
xor U4641 (N_4641,N_4499,N_4420);
nand U4642 (N_4642,N_4467,N_4534);
and U4643 (N_4643,N_4581,N_4547);
xnor U4644 (N_4644,N_4409,N_4470);
nand U4645 (N_4645,N_4474,N_4503);
and U4646 (N_4646,N_4429,N_4414);
or U4647 (N_4647,N_4505,N_4431);
and U4648 (N_4648,N_4583,N_4555);
nor U4649 (N_4649,N_4532,N_4441);
nand U4650 (N_4650,N_4550,N_4568);
or U4651 (N_4651,N_4439,N_4484);
xnor U4652 (N_4652,N_4489,N_4570);
and U4653 (N_4653,N_4572,N_4535);
xnor U4654 (N_4654,N_4485,N_4454);
or U4655 (N_4655,N_4541,N_4538);
and U4656 (N_4656,N_4582,N_4415);
nand U4657 (N_4657,N_4598,N_4475);
xnor U4658 (N_4658,N_4539,N_4517);
nand U4659 (N_4659,N_4500,N_4492);
xnor U4660 (N_4660,N_4557,N_4400);
and U4661 (N_4661,N_4571,N_4514);
nand U4662 (N_4662,N_4446,N_4490);
xor U4663 (N_4663,N_4556,N_4440);
xor U4664 (N_4664,N_4544,N_4520);
xnor U4665 (N_4665,N_4483,N_4424);
and U4666 (N_4666,N_4464,N_4513);
xnor U4667 (N_4667,N_4588,N_4488);
nor U4668 (N_4668,N_4406,N_4507);
nand U4669 (N_4669,N_4504,N_4512);
and U4670 (N_4670,N_4437,N_4423);
nor U4671 (N_4671,N_4533,N_4589);
xor U4672 (N_4672,N_4599,N_4471);
nand U4673 (N_4673,N_4468,N_4536);
nor U4674 (N_4674,N_4417,N_4593);
or U4675 (N_4675,N_4501,N_4430);
xnor U4676 (N_4676,N_4425,N_4426);
nor U4677 (N_4677,N_4542,N_4502);
nor U4678 (N_4678,N_4434,N_4515);
or U4679 (N_4679,N_4418,N_4411);
nand U4680 (N_4680,N_4554,N_4527);
xnor U4681 (N_4681,N_4511,N_4573);
or U4682 (N_4682,N_4525,N_4528);
nand U4683 (N_4683,N_4580,N_4433);
xnor U4684 (N_4684,N_4450,N_4530);
or U4685 (N_4685,N_4435,N_4564);
nor U4686 (N_4686,N_4463,N_4462);
xor U4687 (N_4687,N_4561,N_4491);
xor U4688 (N_4688,N_4413,N_4509);
or U4689 (N_4689,N_4579,N_4487);
or U4690 (N_4690,N_4494,N_4405);
or U4691 (N_4691,N_4569,N_4427);
and U4692 (N_4692,N_4529,N_4578);
xor U4693 (N_4693,N_4519,N_4447);
and U4694 (N_4694,N_4584,N_4540);
xor U4695 (N_4695,N_4473,N_4518);
nand U4696 (N_4696,N_4407,N_4551);
and U4697 (N_4697,N_4455,N_4480);
xor U4698 (N_4698,N_4577,N_4537);
and U4699 (N_4699,N_4590,N_4548);
nand U4700 (N_4700,N_4419,N_4400);
and U4701 (N_4701,N_4585,N_4560);
nand U4702 (N_4702,N_4487,N_4495);
xnor U4703 (N_4703,N_4552,N_4464);
or U4704 (N_4704,N_4519,N_4444);
xnor U4705 (N_4705,N_4560,N_4404);
or U4706 (N_4706,N_4481,N_4425);
and U4707 (N_4707,N_4481,N_4436);
nand U4708 (N_4708,N_4433,N_4574);
or U4709 (N_4709,N_4537,N_4488);
nand U4710 (N_4710,N_4583,N_4433);
xnor U4711 (N_4711,N_4469,N_4403);
or U4712 (N_4712,N_4479,N_4574);
or U4713 (N_4713,N_4588,N_4524);
xor U4714 (N_4714,N_4570,N_4482);
xnor U4715 (N_4715,N_4430,N_4482);
and U4716 (N_4716,N_4535,N_4520);
or U4717 (N_4717,N_4521,N_4465);
nor U4718 (N_4718,N_4590,N_4489);
or U4719 (N_4719,N_4475,N_4495);
xnor U4720 (N_4720,N_4454,N_4506);
xnor U4721 (N_4721,N_4564,N_4551);
xor U4722 (N_4722,N_4559,N_4521);
and U4723 (N_4723,N_4592,N_4597);
nor U4724 (N_4724,N_4597,N_4511);
nor U4725 (N_4725,N_4465,N_4404);
xor U4726 (N_4726,N_4474,N_4414);
and U4727 (N_4727,N_4515,N_4415);
xnor U4728 (N_4728,N_4478,N_4457);
nand U4729 (N_4729,N_4561,N_4595);
nand U4730 (N_4730,N_4422,N_4400);
and U4731 (N_4731,N_4544,N_4527);
or U4732 (N_4732,N_4471,N_4511);
xnor U4733 (N_4733,N_4555,N_4546);
nand U4734 (N_4734,N_4571,N_4547);
and U4735 (N_4735,N_4483,N_4506);
or U4736 (N_4736,N_4569,N_4542);
xnor U4737 (N_4737,N_4504,N_4479);
nand U4738 (N_4738,N_4486,N_4445);
nand U4739 (N_4739,N_4525,N_4447);
and U4740 (N_4740,N_4464,N_4403);
and U4741 (N_4741,N_4482,N_4489);
and U4742 (N_4742,N_4568,N_4599);
nand U4743 (N_4743,N_4523,N_4599);
or U4744 (N_4744,N_4471,N_4477);
or U4745 (N_4745,N_4591,N_4451);
xnor U4746 (N_4746,N_4566,N_4569);
and U4747 (N_4747,N_4555,N_4440);
and U4748 (N_4748,N_4596,N_4527);
or U4749 (N_4749,N_4584,N_4509);
xor U4750 (N_4750,N_4558,N_4423);
and U4751 (N_4751,N_4571,N_4502);
xnor U4752 (N_4752,N_4522,N_4546);
and U4753 (N_4753,N_4438,N_4539);
nand U4754 (N_4754,N_4481,N_4525);
and U4755 (N_4755,N_4485,N_4547);
nand U4756 (N_4756,N_4446,N_4591);
nand U4757 (N_4757,N_4456,N_4465);
xnor U4758 (N_4758,N_4426,N_4491);
or U4759 (N_4759,N_4480,N_4404);
nor U4760 (N_4760,N_4592,N_4588);
and U4761 (N_4761,N_4540,N_4468);
xnor U4762 (N_4762,N_4476,N_4492);
nor U4763 (N_4763,N_4534,N_4517);
nor U4764 (N_4764,N_4574,N_4491);
and U4765 (N_4765,N_4531,N_4430);
nor U4766 (N_4766,N_4488,N_4420);
nand U4767 (N_4767,N_4423,N_4537);
xnor U4768 (N_4768,N_4544,N_4543);
xor U4769 (N_4769,N_4468,N_4544);
and U4770 (N_4770,N_4554,N_4411);
or U4771 (N_4771,N_4504,N_4559);
nand U4772 (N_4772,N_4536,N_4484);
xnor U4773 (N_4773,N_4558,N_4458);
nand U4774 (N_4774,N_4487,N_4553);
xor U4775 (N_4775,N_4461,N_4567);
or U4776 (N_4776,N_4572,N_4447);
nand U4777 (N_4777,N_4408,N_4432);
xnor U4778 (N_4778,N_4409,N_4596);
xor U4779 (N_4779,N_4402,N_4555);
nand U4780 (N_4780,N_4544,N_4450);
nor U4781 (N_4781,N_4405,N_4465);
xor U4782 (N_4782,N_4540,N_4479);
nand U4783 (N_4783,N_4451,N_4458);
xor U4784 (N_4784,N_4558,N_4518);
xnor U4785 (N_4785,N_4425,N_4496);
xnor U4786 (N_4786,N_4529,N_4548);
nor U4787 (N_4787,N_4442,N_4492);
or U4788 (N_4788,N_4454,N_4492);
nand U4789 (N_4789,N_4558,N_4533);
and U4790 (N_4790,N_4480,N_4517);
xor U4791 (N_4791,N_4423,N_4424);
xor U4792 (N_4792,N_4445,N_4444);
nor U4793 (N_4793,N_4562,N_4580);
nand U4794 (N_4794,N_4408,N_4587);
nand U4795 (N_4795,N_4518,N_4427);
xnor U4796 (N_4796,N_4512,N_4558);
or U4797 (N_4797,N_4573,N_4496);
xor U4798 (N_4798,N_4521,N_4458);
nor U4799 (N_4799,N_4587,N_4480);
xnor U4800 (N_4800,N_4705,N_4631);
and U4801 (N_4801,N_4713,N_4608);
nand U4802 (N_4802,N_4621,N_4738);
and U4803 (N_4803,N_4798,N_4796);
nand U4804 (N_4804,N_4782,N_4750);
or U4805 (N_4805,N_4716,N_4693);
and U4806 (N_4806,N_4775,N_4799);
nor U4807 (N_4807,N_4648,N_4629);
nor U4808 (N_4808,N_4725,N_4615);
xnor U4809 (N_4809,N_4737,N_4707);
xor U4810 (N_4810,N_4771,N_4718);
nand U4811 (N_4811,N_4640,N_4745);
nand U4812 (N_4812,N_4724,N_4690);
and U4813 (N_4813,N_4671,N_4754);
xor U4814 (N_4814,N_4676,N_4632);
and U4815 (N_4815,N_4670,N_4624);
or U4816 (N_4816,N_4768,N_4647);
and U4817 (N_4817,N_4669,N_4781);
xnor U4818 (N_4818,N_4739,N_4733);
nor U4819 (N_4819,N_4712,N_4762);
and U4820 (N_4820,N_4607,N_4744);
nand U4821 (N_4821,N_4665,N_4740);
xnor U4822 (N_4822,N_4625,N_4653);
and U4823 (N_4823,N_4643,N_4779);
nor U4824 (N_4824,N_4635,N_4763);
and U4825 (N_4825,N_4777,N_4756);
xor U4826 (N_4826,N_4715,N_4675);
xor U4827 (N_4827,N_4746,N_4674);
or U4828 (N_4828,N_4680,N_4612);
or U4829 (N_4829,N_4797,N_4658);
nor U4830 (N_4830,N_4641,N_4776);
nor U4831 (N_4831,N_4691,N_4664);
and U4832 (N_4832,N_4759,N_4787);
xnor U4833 (N_4833,N_4668,N_4736);
xnor U4834 (N_4834,N_4619,N_4684);
nand U4835 (N_4835,N_4679,N_4678);
and U4836 (N_4836,N_4644,N_4639);
or U4837 (N_4837,N_4789,N_4741);
xnor U4838 (N_4838,N_4758,N_4623);
nor U4839 (N_4839,N_4645,N_4720);
and U4840 (N_4840,N_4732,N_4666);
nand U4841 (N_4841,N_4618,N_4651);
nand U4842 (N_4842,N_4654,N_4634);
nor U4843 (N_4843,N_4793,N_4726);
xnor U4844 (N_4844,N_4774,N_4614);
nand U4845 (N_4845,N_4613,N_4620);
nand U4846 (N_4846,N_4687,N_4714);
xnor U4847 (N_4847,N_4711,N_4660);
xor U4848 (N_4848,N_4742,N_4765);
nor U4849 (N_4849,N_4766,N_4761);
nand U4850 (N_4850,N_4609,N_4760);
xor U4851 (N_4851,N_4785,N_4702);
and U4852 (N_4852,N_4650,N_4734);
xnor U4853 (N_4853,N_4611,N_4661);
xor U4854 (N_4854,N_4637,N_4704);
and U4855 (N_4855,N_4795,N_4681);
xor U4856 (N_4856,N_4723,N_4752);
nor U4857 (N_4857,N_4659,N_4706);
xor U4858 (N_4858,N_4603,N_4667);
xor U4859 (N_4859,N_4694,N_4672);
nor U4860 (N_4860,N_4717,N_4788);
nor U4861 (N_4861,N_4606,N_4682);
nor U4862 (N_4862,N_4626,N_4686);
nor U4863 (N_4863,N_4722,N_4767);
or U4864 (N_4864,N_4772,N_4698);
or U4865 (N_4865,N_4770,N_4710);
nand U4866 (N_4866,N_4656,N_4757);
nor U4867 (N_4867,N_4735,N_4688);
or U4868 (N_4868,N_4792,N_4700);
or U4869 (N_4869,N_4683,N_4778);
and U4870 (N_4870,N_4692,N_4604);
nand U4871 (N_4871,N_4689,N_4638);
nand U4872 (N_4872,N_4673,N_4655);
nand U4873 (N_4873,N_4780,N_4794);
xor U4874 (N_4874,N_4791,N_4703);
or U4875 (N_4875,N_4605,N_4790);
xor U4876 (N_4876,N_4753,N_4748);
and U4877 (N_4877,N_4657,N_4749);
nor U4878 (N_4878,N_4628,N_4642);
or U4879 (N_4879,N_4731,N_4636);
nor U4880 (N_4880,N_4677,N_4747);
nand U4881 (N_4881,N_4743,N_4646);
nor U4882 (N_4882,N_4783,N_4764);
or U4883 (N_4883,N_4719,N_4695);
or U4884 (N_4884,N_4685,N_4610);
or U4885 (N_4885,N_4730,N_4630);
and U4886 (N_4886,N_4727,N_4649);
nand U4887 (N_4887,N_4617,N_4699);
nor U4888 (N_4888,N_4709,N_4697);
nand U4889 (N_4889,N_4786,N_4729);
and U4890 (N_4890,N_4616,N_4663);
nor U4891 (N_4891,N_4600,N_4601);
or U4892 (N_4892,N_4622,N_4696);
nor U4893 (N_4893,N_4708,N_4784);
nor U4894 (N_4894,N_4701,N_4633);
or U4895 (N_4895,N_4627,N_4652);
and U4896 (N_4896,N_4773,N_4728);
or U4897 (N_4897,N_4751,N_4602);
and U4898 (N_4898,N_4755,N_4769);
and U4899 (N_4899,N_4662,N_4721);
and U4900 (N_4900,N_4764,N_4706);
nand U4901 (N_4901,N_4783,N_4653);
or U4902 (N_4902,N_4773,N_4772);
nor U4903 (N_4903,N_4655,N_4738);
nand U4904 (N_4904,N_4656,N_4630);
xnor U4905 (N_4905,N_4716,N_4772);
nand U4906 (N_4906,N_4763,N_4634);
or U4907 (N_4907,N_4618,N_4661);
nand U4908 (N_4908,N_4615,N_4774);
or U4909 (N_4909,N_4653,N_4674);
xnor U4910 (N_4910,N_4795,N_4788);
xnor U4911 (N_4911,N_4641,N_4730);
nand U4912 (N_4912,N_4777,N_4699);
or U4913 (N_4913,N_4621,N_4601);
nand U4914 (N_4914,N_4772,N_4780);
nand U4915 (N_4915,N_4773,N_4693);
xnor U4916 (N_4916,N_4640,N_4695);
nand U4917 (N_4917,N_4715,N_4756);
nor U4918 (N_4918,N_4707,N_4628);
and U4919 (N_4919,N_4669,N_4607);
or U4920 (N_4920,N_4778,N_4641);
xnor U4921 (N_4921,N_4753,N_4687);
nand U4922 (N_4922,N_4739,N_4635);
nand U4923 (N_4923,N_4688,N_4663);
and U4924 (N_4924,N_4736,N_4682);
nand U4925 (N_4925,N_4601,N_4797);
nand U4926 (N_4926,N_4759,N_4792);
xnor U4927 (N_4927,N_4604,N_4744);
nor U4928 (N_4928,N_4647,N_4740);
or U4929 (N_4929,N_4684,N_4717);
nor U4930 (N_4930,N_4762,N_4765);
xor U4931 (N_4931,N_4609,N_4754);
and U4932 (N_4932,N_4612,N_4675);
nand U4933 (N_4933,N_4665,N_4791);
xor U4934 (N_4934,N_4686,N_4780);
xnor U4935 (N_4935,N_4758,N_4709);
and U4936 (N_4936,N_4788,N_4608);
or U4937 (N_4937,N_4784,N_4753);
and U4938 (N_4938,N_4748,N_4789);
or U4939 (N_4939,N_4725,N_4691);
xnor U4940 (N_4940,N_4691,N_4659);
nand U4941 (N_4941,N_4622,N_4667);
xnor U4942 (N_4942,N_4609,N_4696);
xor U4943 (N_4943,N_4651,N_4658);
or U4944 (N_4944,N_4749,N_4694);
xnor U4945 (N_4945,N_4755,N_4739);
nor U4946 (N_4946,N_4763,N_4756);
xor U4947 (N_4947,N_4666,N_4707);
nor U4948 (N_4948,N_4616,N_4736);
and U4949 (N_4949,N_4690,N_4765);
nand U4950 (N_4950,N_4694,N_4636);
nor U4951 (N_4951,N_4652,N_4692);
xor U4952 (N_4952,N_4637,N_4730);
xor U4953 (N_4953,N_4699,N_4723);
nor U4954 (N_4954,N_4743,N_4645);
nor U4955 (N_4955,N_4633,N_4671);
or U4956 (N_4956,N_4660,N_4763);
nand U4957 (N_4957,N_4730,N_4626);
nand U4958 (N_4958,N_4744,N_4749);
nor U4959 (N_4959,N_4715,N_4749);
or U4960 (N_4960,N_4774,N_4673);
and U4961 (N_4961,N_4752,N_4725);
or U4962 (N_4962,N_4780,N_4656);
xor U4963 (N_4963,N_4784,N_4788);
xor U4964 (N_4964,N_4629,N_4742);
xnor U4965 (N_4965,N_4745,N_4795);
or U4966 (N_4966,N_4704,N_4705);
nor U4967 (N_4967,N_4615,N_4699);
or U4968 (N_4968,N_4733,N_4639);
and U4969 (N_4969,N_4711,N_4682);
xnor U4970 (N_4970,N_4691,N_4721);
or U4971 (N_4971,N_4767,N_4675);
or U4972 (N_4972,N_4666,N_4636);
nand U4973 (N_4973,N_4663,N_4635);
and U4974 (N_4974,N_4720,N_4787);
nor U4975 (N_4975,N_4623,N_4796);
xnor U4976 (N_4976,N_4713,N_4605);
nand U4977 (N_4977,N_4799,N_4603);
or U4978 (N_4978,N_4717,N_4626);
and U4979 (N_4979,N_4760,N_4671);
nand U4980 (N_4980,N_4627,N_4721);
and U4981 (N_4981,N_4791,N_4788);
or U4982 (N_4982,N_4621,N_4619);
or U4983 (N_4983,N_4644,N_4617);
xnor U4984 (N_4984,N_4739,N_4724);
nor U4985 (N_4985,N_4656,N_4746);
nand U4986 (N_4986,N_4787,N_4629);
nor U4987 (N_4987,N_4734,N_4753);
nor U4988 (N_4988,N_4740,N_4624);
or U4989 (N_4989,N_4609,N_4777);
or U4990 (N_4990,N_4736,N_4634);
nor U4991 (N_4991,N_4786,N_4760);
or U4992 (N_4992,N_4615,N_4771);
and U4993 (N_4993,N_4796,N_4777);
or U4994 (N_4994,N_4600,N_4689);
xor U4995 (N_4995,N_4602,N_4791);
nand U4996 (N_4996,N_4764,N_4784);
nand U4997 (N_4997,N_4729,N_4681);
and U4998 (N_4998,N_4751,N_4631);
or U4999 (N_4999,N_4691,N_4662);
xor U5000 (N_5000,N_4873,N_4827);
nand U5001 (N_5001,N_4911,N_4884);
xor U5002 (N_5002,N_4852,N_4988);
xnor U5003 (N_5003,N_4981,N_4935);
or U5004 (N_5004,N_4917,N_4947);
xnor U5005 (N_5005,N_4913,N_4956);
xnor U5006 (N_5006,N_4848,N_4963);
xnor U5007 (N_5007,N_4928,N_4991);
nor U5008 (N_5008,N_4909,N_4934);
xnor U5009 (N_5009,N_4892,N_4970);
xnor U5010 (N_5010,N_4898,N_4978);
and U5011 (N_5011,N_4811,N_4916);
nand U5012 (N_5012,N_4835,N_4983);
nor U5013 (N_5013,N_4859,N_4942);
nor U5014 (N_5014,N_4986,N_4843);
nand U5015 (N_5015,N_4851,N_4918);
xor U5016 (N_5016,N_4854,N_4940);
or U5017 (N_5017,N_4887,N_4922);
and U5018 (N_5018,N_4954,N_4992);
and U5019 (N_5019,N_4905,N_4869);
nor U5020 (N_5020,N_4958,N_4828);
xor U5021 (N_5021,N_4872,N_4876);
xnor U5022 (N_5022,N_4894,N_4987);
and U5023 (N_5023,N_4858,N_4800);
nor U5024 (N_5024,N_4865,N_4816);
nor U5025 (N_5025,N_4930,N_4932);
nor U5026 (N_5026,N_4857,N_4860);
nor U5027 (N_5027,N_4994,N_4867);
xor U5028 (N_5028,N_4814,N_4920);
xor U5029 (N_5029,N_4946,N_4919);
and U5030 (N_5030,N_4964,N_4822);
nand U5031 (N_5031,N_4912,N_4999);
and U5032 (N_5032,N_4863,N_4808);
xor U5033 (N_5033,N_4925,N_4823);
nand U5034 (N_5034,N_4955,N_4997);
xnor U5035 (N_5035,N_4837,N_4907);
and U5036 (N_5036,N_4924,N_4976);
xnor U5037 (N_5037,N_4874,N_4980);
nand U5038 (N_5038,N_4906,N_4806);
xor U5039 (N_5039,N_4923,N_4952);
or U5040 (N_5040,N_4805,N_4965);
nor U5041 (N_5041,N_4998,N_4902);
nor U5042 (N_5042,N_4943,N_4996);
xnor U5043 (N_5043,N_4836,N_4972);
and U5044 (N_5044,N_4871,N_4853);
or U5045 (N_5045,N_4929,N_4937);
nand U5046 (N_5046,N_4830,N_4927);
nand U5047 (N_5047,N_4888,N_4815);
nand U5048 (N_5048,N_4977,N_4961);
or U5049 (N_5049,N_4801,N_4804);
and U5050 (N_5050,N_4939,N_4969);
xnor U5051 (N_5051,N_4862,N_4866);
nor U5052 (N_5052,N_4834,N_4844);
or U5053 (N_5053,N_4826,N_4810);
xnor U5054 (N_5054,N_4879,N_4832);
nand U5055 (N_5055,N_4861,N_4901);
xor U5056 (N_5056,N_4985,N_4819);
and U5057 (N_5057,N_4921,N_4842);
and U5058 (N_5058,N_4829,N_4979);
and U5059 (N_5059,N_4938,N_4973);
and U5060 (N_5060,N_4893,N_4974);
and U5061 (N_5061,N_4885,N_4936);
or U5062 (N_5062,N_4941,N_4850);
nand U5063 (N_5063,N_4926,N_4877);
and U5064 (N_5064,N_4904,N_4864);
or U5065 (N_5065,N_4899,N_4812);
nand U5066 (N_5066,N_4802,N_4957);
nor U5067 (N_5067,N_4838,N_4914);
or U5068 (N_5068,N_4856,N_4881);
nand U5069 (N_5069,N_4984,N_4945);
or U5070 (N_5070,N_4831,N_4990);
nor U5071 (N_5071,N_4908,N_4896);
xor U5072 (N_5072,N_4966,N_4845);
and U5073 (N_5073,N_4949,N_4891);
or U5074 (N_5074,N_4933,N_4890);
xnor U5075 (N_5075,N_4989,N_4951);
nor U5076 (N_5076,N_4818,N_4882);
xor U5077 (N_5077,N_4821,N_4968);
and U5078 (N_5078,N_4875,N_4982);
nor U5079 (N_5079,N_4971,N_4960);
and U5080 (N_5080,N_4833,N_4895);
nand U5081 (N_5081,N_4903,N_4878);
nand U5082 (N_5082,N_4993,N_4975);
nand U5083 (N_5083,N_4995,N_4855);
and U5084 (N_5084,N_4870,N_4944);
xnor U5085 (N_5085,N_4948,N_4915);
nor U5086 (N_5086,N_4967,N_4897);
nand U5087 (N_5087,N_4813,N_4886);
and U5088 (N_5088,N_4847,N_4910);
and U5089 (N_5089,N_4880,N_4868);
nor U5090 (N_5090,N_4824,N_4809);
and U5091 (N_5091,N_4817,N_4803);
nor U5092 (N_5092,N_4950,N_4839);
nor U5093 (N_5093,N_4841,N_4883);
nand U5094 (N_5094,N_4900,N_4931);
xor U5095 (N_5095,N_4889,N_4962);
nand U5096 (N_5096,N_4849,N_4953);
and U5097 (N_5097,N_4846,N_4840);
or U5098 (N_5098,N_4820,N_4825);
xor U5099 (N_5099,N_4959,N_4807);
nand U5100 (N_5100,N_4818,N_4814);
or U5101 (N_5101,N_4904,N_4839);
nand U5102 (N_5102,N_4949,N_4870);
and U5103 (N_5103,N_4882,N_4961);
xor U5104 (N_5104,N_4939,N_4841);
nand U5105 (N_5105,N_4826,N_4951);
xor U5106 (N_5106,N_4830,N_4925);
nor U5107 (N_5107,N_4897,N_4802);
or U5108 (N_5108,N_4902,N_4939);
nor U5109 (N_5109,N_4985,N_4967);
or U5110 (N_5110,N_4945,N_4879);
and U5111 (N_5111,N_4800,N_4832);
nand U5112 (N_5112,N_4854,N_4989);
xnor U5113 (N_5113,N_4897,N_4926);
or U5114 (N_5114,N_4999,N_4937);
or U5115 (N_5115,N_4839,N_4971);
nor U5116 (N_5116,N_4899,N_4924);
and U5117 (N_5117,N_4979,N_4981);
and U5118 (N_5118,N_4908,N_4910);
and U5119 (N_5119,N_4849,N_4934);
xor U5120 (N_5120,N_4904,N_4983);
nor U5121 (N_5121,N_4942,N_4965);
and U5122 (N_5122,N_4915,N_4933);
nor U5123 (N_5123,N_4916,N_4893);
or U5124 (N_5124,N_4856,N_4911);
xnor U5125 (N_5125,N_4968,N_4949);
xnor U5126 (N_5126,N_4993,N_4932);
xor U5127 (N_5127,N_4858,N_4840);
or U5128 (N_5128,N_4987,N_4864);
and U5129 (N_5129,N_4837,N_4875);
and U5130 (N_5130,N_4834,N_4928);
xor U5131 (N_5131,N_4989,N_4844);
xor U5132 (N_5132,N_4808,N_4947);
nor U5133 (N_5133,N_4959,N_4869);
nand U5134 (N_5134,N_4832,N_4899);
and U5135 (N_5135,N_4816,N_4822);
and U5136 (N_5136,N_4888,N_4988);
and U5137 (N_5137,N_4980,N_4903);
and U5138 (N_5138,N_4800,N_4895);
nand U5139 (N_5139,N_4997,N_4832);
and U5140 (N_5140,N_4978,N_4847);
xor U5141 (N_5141,N_4810,N_4827);
xnor U5142 (N_5142,N_4897,N_4893);
nor U5143 (N_5143,N_4876,N_4931);
nand U5144 (N_5144,N_4924,N_4839);
and U5145 (N_5145,N_4854,N_4897);
xor U5146 (N_5146,N_4939,N_4844);
nand U5147 (N_5147,N_4935,N_4802);
and U5148 (N_5148,N_4819,N_4855);
or U5149 (N_5149,N_4831,N_4884);
xnor U5150 (N_5150,N_4836,N_4898);
and U5151 (N_5151,N_4840,N_4893);
and U5152 (N_5152,N_4931,N_4875);
and U5153 (N_5153,N_4870,N_4912);
nor U5154 (N_5154,N_4996,N_4935);
nand U5155 (N_5155,N_4896,N_4903);
and U5156 (N_5156,N_4867,N_4841);
xor U5157 (N_5157,N_4848,N_4921);
xnor U5158 (N_5158,N_4814,N_4915);
or U5159 (N_5159,N_4977,N_4866);
or U5160 (N_5160,N_4916,N_4868);
xnor U5161 (N_5161,N_4859,N_4939);
and U5162 (N_5162,N_4846,N_4854);
and U5163 (N_5163,N_4935,N_4805);
and U5164 (N_5164,N_4810,N_4956);
and U5165 (N_5165,N_4990,N_4877);
nor U5166 (N_5166,N_4863,N_4864);
xor U5167 (N_5167,N_4817,N_4836);
and U5168 (N_5168,N_4806,N_4896);
xnor U5169 (N_5169,N_4873,N_4973);
xor U5170 (N_5170,N_4824,N_4901);
xor U5171 (N_5171,N_4837,N_4995);
nor U5172 (N_5172,N_4961,N_4831);
and U5173 (N_5173,N_4828,N_4868);
xor U5174 (N_5174,N_4995,N_4984);
and U5175 (N_5175,N_4854,N_4876);
nor U5176 (N_5176,N_4946,N_4956);
or U5177 (N_5177,N_4811,N_4945);
or U5178 (N_5178,N_4886,N_4939);
or U5179 (N_5179,N_4956,N_4986);
xor U5180 (N_5180,N_4904,N_4857);
or U5181 (N_5181,N_4821,N_4933);
or U5182 (N_5182,N_4940,N_4868);
and U5183 (N_5183,N_4920,N_4941);
nand U5184 (N_5184,N_4816,N_4844);
nor U5185 (N_5185,N_4880,N_4833);
nor U5186 (N_5186,N_4984,N_4871);
and U5187 (N_5187,N_4820,N_4887);
or U5188 (N_5188,N_4970,N_4998);
nand U5189 (N_5189,N_4957,N_4961);
nand U5190 (N_5190,N_4841,N_4854);
and U5191 (N_5191,N_4867,N_4959);
nor U5192 (N_5192,N_4890,N_4978);
nor U5193 (N_5193,N_4847,N_4900);
or U5194 (N_5194,N_4881,N_4925);
nand U5195 (N_5195,N_4831,N_4912);
nand U5196 (N_5196,N_4880,N_4983);
and U5197 (N_5197,N_4921,N_4873);
xnor U5198 (N_5198,N_4826,N_4975);
nor U5199 (N_5199,N_4854,N_4947);
or U5200 (N_5200,N_5070,N_5166);
and U5201 (N_5201,N_5179,N_5152);
nand U5202 (N_5202,N_5130,N_5011);
nor U5203 (N_5203,N_5085,N_5171);
or U5204 (N_5204,N_5073,N_5198);
and U5205 (N_5205,N_5149,N_5056);
nand U5206 (N_5206,N_5163,N_5119);
or U5207 (N_5207,N_5050,N_5048);
nor U5208 (N_5208,N_5147,N_5187);
xnor U5209 (N_5209,N_5021,N_5041);
xnor U5210 (N_5210,N_5156,N_5093);
and U5211 (N_5211,N_5110,N_5026);
nand U5212 (N_5212,N_5078,N_5057);
nor U5213 (N_5213,N_5135,N_5023);
xnor U5214 (N_5214,N_5067,N_5003);
xor U5215 (N_5215,N_5175,N_5060);
and U5216 (N_5216,N_5063,N_5064);
or U5217 (N_5217,N_5183,N_5189);
nand U5218 (N_5218,N_5049,N_5127);
or U5219 (N_5219,N_5062,N_5009);
or U5220 (N_5220,N_5168,N_5154);
nor U5221 (N_5221,N_5027,N_5020);
nor U5222 (N_5222,N_5172,N_5106);
xnor U5223 (N_5223,N_5108,N_5001);
and U5224 (N_5224,N_5145,N_5014);
or U5225 (N_5225,N_5055,N_5019);
and U5226 (N_5226,N_5118,N_5116);
and U5227 (N_5227,N_5104,N_5142);
nand U5228 (N_5228,N_5046,N_5131);
or U5229 (N_5229,N_5177,N_5159);
xnor U5230 (N_5230,N_5109,N_5160);
nand U5231 (N_5231,N_5071,N_5059);
and U5232 (N_5232,N_5080,N_5047);
nor U5233 (N_5233,N_5005,N_5045);
nand U5234 (N_5234,N_5065,N_5165);
or U5235 (N_5235,N_5138,N_5068);
and U5236 (N_5236,N_5195,N_5044);
nor U5237 (N_5237,N_5174,N_5030);
xnor U5238 (N_5238,N_5040,N_5033);
xor U5239 (N_5239,N_5101,N_5006);
and U5240 (N_5240,N_5117,N_5148);
nand U5241 (N_5241,N_5182,N_5096);
nand U5242 (N_5242,N_5042,N_5105);
nor U5243 (N_5243,N_5146,N_5089);
xnor U5244 (N_5244,N_5140,N_5025);
nand U5245 (N_5245,N_5024,N_5144);
or U5246 (N_5246,N_5029,N_5169);
xnor U5247 (N_5247,N_5010,N_5188);
xnor U5248 (N_5248,N_5120,N_5113);
nor U5249 (N_5249,N_5186,N_5121);
nand U5250 (N_5250,N_5132,N_5091);
or U5251 (N_5251,N_5061,N_5137);
xnor U5252 (N_5252,N_5155,N_5015);
nand U5253 (N_5253,N_5087,N_5141);
nand U5254 (N_5254,N_5150,N_5007);
xor U5255 (N_5255,N_5051,N_5128);
or U5256 (N_5256,N_5129,N_5158);
nand U5257 (N_5257,N_5196,N_5094);
and U5258 (N_5258,N_5016,N_5054);
and U5259 (N_5259,N_5170,N_5000);
nor U5260 (N_5260,N_5157,N_5036);
xor U5261 (N_5261,N_5122,N_5066);
and U5262 (N_5262,N_5034,N_5018);
nor U5263 (N_5263,N_5004,N_5114);
nor U5264 (N_5264,N_5176,N_5095);
xor U5265 (N_5265,N_5008,N_5125);
nand U5266 (N_5266,N_5102,N_5037);
nor U5267 (N_5267,N_5035,N_5192);
and U5268 (N_5268,N_5185,N_5022);
and U5269 (N_5269,N_5123,N_5002);
nand U5270 (N_5270,N_5112,N_5076);
nand U5271 (N_5271,N_5190,N_5180);
and U5272 (N_5272,N_5058,N_5098);
nor U5273 (N_5273,N_5031,N_5139);
nor U5274 (N_5274,N_5100,N_5017);
xor U5275 (N_5275,N_5092,N_5153);
and U5276 (N_5276,N_5084,N_5097);
nor U5277 (N_5277,N_5115,N_5083);
xor U5278 (N_5278,N_5103,N_5124);
or U5279 (N_5279,N_5082,N_5181);
and U5280 (N_5280,N_5013,N_5074);
nand U5281 (N_5281,N_5032,N_5081);
nand U5282 (N_5282,N_5167,N_5143);
nand U5283 (N_5283,N_5012,N_5126);
and U5284 (N_5284,N_5086,N_5039);
and U5285 (N_5285,N_5194,N_5053);
and U5286 (N_5286,N_5164,N_5072);
nor U5287 (N_5287,N_5043,N_5038);
and U5288 (N_5288,N_5184,N_5151);
nand U5289 (N_5289,N_5199,N_5079);
nor U5290 (N_5290,N_5090,N_5133);
nand U5291 (N_5291,N_5077,N_5111);
xor U5292 (N_5292,N_5069,N_5173);
nand U5293 (N_5293,N_5193,N_5099);
nand U5294 (N_5294,N_5088,N_5107);
xor U5295 (N_5295,N_5178,N_5161);
and U5296 (N_5296,N_5197,N_5191);
nand U5297 (N_5297,N_5075,N_5162);
nor U5298 (N_5298,N_5052,N_5134);
or U5299 (N_5299,N_5136,N_5028);
or U5300 (N_5300,N_5072,N_5173);
nor U5301 (N_5301,N_5099,N_5181);
nor U5302 (N_5302,N_5078,N_5070);
or U5303 (N_5303,N_5154,N_5121);
xor U5304 (N_5304,N_5119,N_5083);
nand U5305 (N_5305,N_5095,N_5186);
nor U5306 (N_5306,N_5140,N_5048);
xor U5307 (N_5307,N_5184,N_5034);
and U5308 (N_5308,N_5075,N_5065);
and U5309 (N_5309,N_5128,N_5076);
nor U5310 (N_5310,N_5114,N_5031);
and U5311 (N_5311,N_5003,N_5013);
or U5312 (N_5312,N_5149,N_5140);
and U5313 (N_5313,N_5069,N_5116);
xor U5314 (N_5314,N_5156,N_5077);
xor U5315 (N_5315,N_5138,N_5110);
nand U5316 (N_5316,N_5101,N_5062);
nand U5317 (N_5317,N_5015,N_5039);
and U5318 (N_5318,N_5044,N_5024);
xnor U5319 (N_5319,N_5026,N_5076);
or U5320 (N_5320,N_5128,N_5152);
or U5321 (N_5321,N_5077,N_5193);
xnor U5322 (N_5322,N_5019,N_5063);
nor U5323 (N_5323,N_5165,N_5043);
xor U5324 (N_5324,N_5024,N_5157);
and U5325 (N_5325,N_5186,N_5066);
or U5326 (N_5326,N_5107,N_5121);
nand U5327 (N_5327,N_5147,N_5003);
or U5328 (N_5328,N_5099,N_5147);
xor U5329 (N_5329,N_5150,N_5085);
or U5330 (N_5330,N_5138,N_5043);
and U5331 (N_5331,N_5113,N_5188);
nand U5332 (N_5332,N_5168,N_5063);
nand U5333 (N_5333,N_5190,N_5020);
or U5334 (N_5334,N_5089,N_5165);
nand U5335 (N_5335,N_5130,N_5003);
xor U5336 (N_5336,N_5038,N_5003);
xor U5337 (N_5337,N_5088,N_5008);
or U5338 (N_5338,N_5099,N_5013);
nor U5339 (N_5339,N_5077,N_5135);
and U5340 (N_5340,N_5195,N_5037);
or U5341 (N_5341,N_5109,N_5042);
xnor U5342 (N_5342,N_5002,N_5075);
nor U5343 (N_5343,N_5068,N_5170);
nor U5344 (N_5344,N_5033,N_5097);
nor U5345 (N_5345,N_5117,N_5040);
and U5346 (N_5346,N_5036,N_5167);
xnor U5347 (N_5347,N_5045,N_5033);
xnor U5348 (N_5348,N_5116,N_5109);
nor U5349 (N_5349,N_5196,N_5144);
nand U5350 (N_5350,N_5166,N_5127);
nor U5351 (N_5351,N_5141,N_5126);
or U5352 (N_5352,N_5075,N_5177);
xnor U5353 (N_5353,N_5156,N_5121);
and U5354 (N_5354,N_5108,N_5178);
xnor U5355 (N_5355,N_5112,N_5035);
xor U5356 (N_5356,N_5006,N_5171);
or U5357 (N_5357,N_5117,N_5180);
and U5358 (N_5358,N_5135,N_5095);
nand U5359 (N_5359,N_5086,N_5145);
or U5360 (N_5360,N_5092,N_5171);
xnor U5361 (N_5361,N_5103,N_5170);
nor U5362 (N_5362,N_5098,N_5121);
or U5363 (N_5363,N_5002,N_5157);
and U5364 (N_5364,N_5060,N_5063);
nand U5365 (N_5365,N_5199,N_5024);
and U5366 (N_5366,N_5087,N_5104);
nand U5367 (N_5367,N_5057,N_5129);
nand U5368 (N_5368,N_5102,N_5018);
nor U5369 (N_5369,N_5046,N_5154);
or U5370 (N_5370,N_5024,N_5185);
or U5371 (N_5371,N_5142,N_5080);
xnor U5372 (N_5372,N_5039,N_5005);
xor U5373 (N_5373,N_5033,N_5147);
xnor U5374 (N_5374,N_5087,N_5161);
or U5375 (N_5375,N_5173,N_5075);
and U5376 (N_5376,N_5093,N_5133);
nand U5377 (N_5377,N_5051,N_5082);
nand U5378 (N_5378,N_5040,N_5047);
nand U5379 (N_5379,N_5039,N_5167);
or U5380 (N_5380,N_5097,N_5186);
xnor U5381 (N_5381,N_5103,N_5117);
nand U5382 (N_5382,N_5153,N_5028);
xnor U5383 (N_5383,N_5191,N_5054);
xnor U5384 (N_5384,N_5051,N_5009);
xnor U5385 (N_5385,N_5177,N_5076);
xnor U5386 (N_5386,N_5192,N_5174);
nor U5387 (N_5387,N_5068,N_5093);
and U5388 (N_5388,N_5092,N_5023);
or U5389 (N_5389,N_5113,N_5114);
xnor U5390 (N_5390,N_5179,N_5116);
nor U5391 (N_5391,N_5190,N_5058);
nand U5392 (N_5392,N_5031,N_5044);
nand U5393 (N_5393,N_5023,N_5139);
nand U5394 (N_5394,N_5073,N_5054);
and U5395 (N_5395,N_5189,N_5007);
nor U5396 (N_5396,N_5099,N_5121);
xnor U5397 (N_5397,N_5017,N_5087);
and U5398 (N_5398,N_5078,N_5092);
nor U5399 (N_5399,N_5143,N_5010);
nor U5400 (N_5400,N_5298,N_5240);
and U5401 (N_5401,N_5201,N_5225);
nor U5402 (N_5402,N_5301,N_5333);
and U5403 (N_5403,N_5370,N_5250);
nand U5404 (N_5404,N_5362,N_5203);
nor U5405 (N_5405,N_5294,N_5359);
xor U5406 (N_5406,N_5227,N_5205);
and U5407 (N_5407,N_5356,N_5316);
or U5408 (N_5408,N_5334,N_5255);
nand U5409 (N_5409,N_5273,N_5383);
xor U5410 (N_5410,N_5235,N_5239);
and U5411 (N_5411,N_5322,N_5393);
nand U5412 (N_5412,N_5207,N_5284);
nor U5413 (N_5413,N_5305,N_5204);
and U5414 (N_5414,N_5303,N_5267);
xnor U5415 (N_5415,N_5283,N_5200);
or U5416 (N_5416,N_5378,N_5296);
xor U5417 (N_5417,N_5248,N_5319);
xor U5418 (N_5418,N_5350,N_5249);
nand U5419 (N_5419,N_5368,N_5245);
nor U5420 (N_5420,N_5339,N_5399);
and U5421 (N_5421,N_5282,N_5244);
and U5422 (N_5422,N_5338,N_5254);
and U5423 (N_5423,N_5261,N_5398);
nand U5424 (N_5424,N_5340,N_5327);
and U5425 (N_5425,N_5358,N_5387);
nand U5426 (N_5426,N_5324,N_5347);
nor U5427 (N_5427,N_5236,N_5367);
nor U5428 (N_5428,N_5260,N_5252);
nor U5429 (N_5429,N_5384,N_5394);
or U5430 (N_5430,N_5262,N_5277);
xor U5431 (N_5431,N_5314,N_5330);
nor U5432 (N_5432,N_5247,N_5288);
and U5433 (N_5433,N_5234,N_5208);
and U5434 (N_5434,N_5269,N_5263);
and U5435 (N_5435,N_5373,N_5286);
nor U5436 (N_5436,N_5326,N_5361);
nor U5437 (N_5437,N_5376,N_5329);
and U5438 (N_5438,N_5352,N_5279);
xor U5439 (N_5439,N_5274,N_5251);
and U5440 (N_5440,N_5278,N_5275);
xnor U5441 (N_5441,N_5217,N_5337);
xor U5442 (N_5442,N_5232,N_5320);
nand U5443 (N_5443,N_5349,N_5342);
xor U5444 (N_5444,N_5310,N_5391);
nor U5445 (N_5445,N_5224,N_5295);
nand U5446 (N_5446,N_5315,N_5307);
and U5447 (N_5447,N_5229,N_5377);
and U5448 (N_5448,N_5243,N_5335);
nand U5449 (N_5449,N_5202,N_5292);
xnor U5450 (N_5450,N_5276,N_5233);
nor U5451 (N_5451,N_5346,N_5385);
xnor U5452 (N_5452,N_5375,N_5213);
and U5453 (N_5453,N_5231,N_5280);
and U5454 (N_5454,N_5364,N_5325);
nand U5455 (N_5455,N_5369,N_5285);
nor U5456 (N_5456,N_5268,N_5311);
xnor U5457 (N_5457,N_5223,N_5281);
and U5458 (N_5458,N_5230,N_5341);
nand U5459 (N_5459,N_5271,N_5293);
nand U5460 (N_5460,N_5287,N_5308);
and U5461 (N_5461,N_5366,N_5216);
nand U5462 (N_5462,N_5343,N_5211);
or U5463 (N_5463,N_5246,N_5379);
nand U5464 (N_5464,N_5300,N_5360);
and U5465 (N_5465,N_5210,N_5270);
or U5466 (N_5466,N_5218,N_5266);
or U5467 (N_5467,N_5272,N_5212);
and U5468 (N_5468,N_5354,N_5392);
and U5469 (N_5469,N_5220,N_5332);
xnor U5470 (N_5470,N_5257,N_5289);
xnor U5471 (N_5471,N_5253,N_5265);
and U5472 (N_5472,N_5323,N_5336);
nand U5473 (N_5473,N_5299,N_5363);
nor U5474 (N_5474,N_5264,N_5388);
or U5475 (N_5475,N_5317,N_5222);
xnor U5476 (N_5476,N_5389,N_5221);
xnor U5477 (N_5477,N_5215,N_5302);
or U5478 (N_5478,N_5258,N_5290);
nor U5479 (N_5479,N_5331,N_5355);
xor U5480 (N_5480,N_5371,N_5238);
or U5481 (N_5481,N_5242,N_5321);
xnor U5482 (N_5482,N_5386,N_5226);
and U5483 (N_5483,N_5365,N_5328);
xnor U5484 (N_5484,N_5374,N_5382);
xnor U5485 (N_5485,N_5318,N_5256);
or U5486 (N_5486,N_5297,N_5380);
nor U5487 (N_5487,N_5344,N_5237);
xor U5488 (N_5488,N_5241,N_5312);
xor U5489 (N_5489,N_5397,N_5351);
nand U5490 (N_5490,N_5306,N_5206);
xnor U5491 (N_5491,N_5381,N_5395);
and U5492 (N_5492,N_5396,N_5214);
xnor U5493 (N_5493,N_5219,N_5304);
nor U5494 (N_5494,N_5390,N_5309);
nor U5495 (N_5495,N_5313,N_5209);
or U5496 (N_5496,N_5345,N_5291);
or U5497 (N_5497,N_5259,N_5348);
and U5498 (N_5498,N_5357,N_5228);
or U5499 (N_5499,N_5372,N_5353);
nand U5500 (N_5500,N_5357,N_5382);
and U5501 (N_5501,N_5372,N_5338);
nor U5502 (N_5502,N_5204,N_5335);
nor U5503 (N_5503,N_5305,N_5340);
nor U5504 (N_5504,N_5265,N_5372);
nor U5505 (N_5505,N_5381,N_5294);
nor U5506 (N_5506,N_5345,N_5249);
and U5507 (N_5507,N_5386,N_5325);
or U5508 (N_5508,N_5389,N_5304);
nand U5509 (N_5509,N_5218,N_5353);
or U5510 (N_5510,N_5280,N_5347);
or U5511 (N_5511,N_5286,N_5251);
or U5512 (N_5512,N_5283,N_5275);
xor U5513 (N_5513,N_5385,N_5366);
or U5514 (N_5514,N_5363,N_5284);
and U5515 (N_5515,N_5318,N_5244);
or U5516 (N_5516,N_5218,N_5327);
or U5517 (N_5517,N_5312,N_5348);
xnor U5518 (N_5518,N_5328,N_5336);
and U5519 (N_5519,N_5286,N_5337);
and U5520 (N_5520,N_5396,N_5389);
or U5521 (N_5521,N_5234,N_5328);
and U5522 (N_5522,N_5374,N_5245);
xnor U5523 (N_5523,N_5287,N_5283);
xnor U5524 (N_5524,N_5281,N_5399);
xor U5525 (N_5525,N_5222,N_5261);
and U5526 (N_5526,N_5340,N_5364);
nand U5527 (N_5527,N_5281,N_5236);
nand U5528 (N_5528,N_5241,N_5209);
and U5529 (N_5529,N_5364,N_5388);
nor U5530 (N_5530,N_5322,N_5299);
nor U5531 (N_5531,N_5355,N_5378);
nor U5532 (N_5532,N_5275,N_5217);
or U5533 (N_5533,N_5256,N_5268);
or U5534 (N_5534,N_5308,N_5265);
nand U5535 (N_5535,N_5326,N_5362);
nor U5536 (N_5536,N_5323,N_5303);
nor U5537 (N_5537,N_5320,N_5288);
nand U5538 (N_5538,N_5313,N_5361);
xor U5539 (N_5539,N_5353,N_5399);
or U5540 (N_5540,N_5357,N_5270);
xnor U5541 (N_5541,N_5233,N_5318);
nand U5542 (N_5542,N_5276,N_5328);
and U5543 (N_5543,N_5217,N_5347);
or U5544 (N_5544,N_5350,N_5231);
nor U5545 (N_5545,N_5242,N_5387);
and U5546 (N_5546,N_5325,N_5388);
and U5547 (N_5547,N_5237,N_5347);
nand U5548 (N_5548,N_5279,N_5210);
nand U5549 (N_5549,N_5208,N_5207);
xnor U5550 (N_5550,N_5303,N_5217);
nand U5551 (N_5551,N_5268,N_5372);
and U5552 (N_5552,N_5220,N_5372);
nor U5553 (N_5553,N_5367,N_5359);
xor U5554 (N_5554,N_5215,N_5348);
nand U5555 (N_5555,N_5266,N_5312);
nand U5556 (N_5556,N_5208,N_5209);
or U5557 (N_5557,N_5399,N_5318);
xnor U5558 (N_5558,N_5275,N_5206);
and U5559 (N_5559,N_5215,N_5225);
or U5560 (N_5560,N_5279,N_5286);
or U5561 (N_5561,N_5314,N_5307);
nand U5562 (N_5562,N_5209,N_5262);
xor U5563 (N_5563,N_5204,N_5356);
nor U5564 (N_5564,N_5385,N_5237);
xnor U5565 (N_5565,N_5222,N_5239);
or U5566 (N_5566,N_5306,N_5355);
xnor U5567 (N_5567,N_5399,N_5251);
xnor U5568 (N_5568,N_5266,N_5399);
or U5569 (N_5569,N_5323,N_5223);
xor U5570 (N_5570,N_5276,N_5266);
or U5571 (N_5571,N_5390,N_5305);
nor U5572 (N_5572,N_5279,N_5313);
nor U5573 (N_5573,N_5308,N_5330);
or U5574 (N_5574,N_5334,N_5230);
nor U5575 (N_5575,N_5337,N_5383);
xor U5576 (N_5576,N_5200,N_5211);
nand U5577 (N_5577,N_5336,N_5324);
xnor U5578 (N_5578,N_5360,N_5201);
nand U5579 (N_5579,N_5254,N_5303);
nand U5580 (N_5580,N_5313,N_5386);
nand U5581 (N_5581,N_5273,N_5225);
nor U5582 (N_5582,N_5213,N_5206);
nor U5583 (N_5583,N_5325,N_5297);
nor U5584 (N_5584,N_5220,N_5294);
or U5585 (N_5585,N_5252,N_5331);
nand U5586 (N_5586,N_5247,N_5282);
nor U5587 (N_5587,N_5308,N_5348);
nand U5588 (N_5588,N_5282,N_5377);
or U5589 (N_5589,N_5362,N_5338);
xnor U5590 (N_5590,N_5344,N_5332);
and U5591 (N_5591,N_5336,N_5270);
nor U5592 (N_5592,N_5305,N_5213);
xor U5593 (N_5593,N_5363,N_5208);
or U5594 (N_5594,N_5313,N_5302);
xor U5595 (N_5595,N_5308,N_5342);
xnor U5596 (N_5596,N_5277,N_5230);
or U5597 (N_5597,N_5377,N_5345);
nand U5598 (N_5598,N_5274,N_5372);
or U5599 (N_5599,N_5211,N_5354);
and U5600 (N_5600,N_5567,N_5440);
or U5601 (N_5601,N_5474,N_5593);
or U5602 (N_5602,N_5491,N_5461);
and U5603 (N_5603,N_5577,N_5548);
nor U5604 (N_5604,N_5546,N_5404);
and U5605 (N_5605,N_5464,N_5459);
or U5606 (N_5606,N_5592,N_5597);
and U5607 (N_5607,N_5498,N_5494);
nor U5608 (N_5608,N_5415,N_5478);
nor U5609 (N_5609,N_5535,N_5420);
or U5610 (N_5610,N_5559,N_5504);
xor U5611 (N_5611,N_5574,N_5564);
and U5612 (N_5612,N_5471,N_5545);
and U5613 (N_5613,N_5455,N_5492);
xnor U5614 (N_5614,N_5448,N_5534);
nand U5615 (N_5615,N_5562,N_5523);
xnor U5616 (N_5616,N_5553,N_5516);
nor U5617 (N_5617,N_5473,N_5527);
or U5618 (N_5618,N_5457,N_5525);
nand U5619 (N_5619,N_5490,N_5583);
and U5620 (N_5620,N_5401,N_5449);
nand U5621 (N_5621,N_5513,N_5596);
and U5622 (N_5622,N_5419,N_5454);
or U5623 (N_5623,N_5453,N_5495);
xnor U5624 (N_5624,N_5555,N_5486);
xnor U5625 (N_5625,N_5496,N_5536);
nand U5626 (N_5626,N_5407,N_5552);
nand U5627 (N_5627,N_5432,N_5443);
and U5628 (N_5628,N_5417,N_5410);
and U5629 (N_5629,N_5437,N_5469);
nand U5630 (N_5630,N_5507,N_5537);
or U5631 (N_5631,N_5585,N_5547);
and U5632 (N_5632,N_5423,N_5533);
nor U5633 (N_5633,N_5581,N_5460);
nand U5634 (N_5634,N_5430,N_5402);
xnor U5635 (N_5635,N_5502,N_5493);
nand U5636 (N_5636,N_5556,N_5403);
nand U5637 (N_5637,N_5406,N_5515);
nor U5638 (N_5638,N_5595,N_5436);
and U5639 (N_5639,N_5450,N_5598);
xnor U5640 (N_5640,N_5451,N_5447);
nand U5641 (N_5641,N_5517,N_5586);
nor U5642 (N_5642,N_5499,N_5569);
or U5643 (N_5643,N_5488,N_5505);
and U5644 (N_5644,N_5442,N_5560);
nor U5645 (N_5645,N_5429,N_5518);
or U5646 (N_5646,N_5412,N_5572);
nand U5647 (N_5647,N_5416,N_5508);
and U5648 (N_5648,N_5409,N_5418);
or U5649 (N_5649,N_5514,N_5489);
xor U5650 (N_5650,N_5421,N_5479);
and U5651 (N_5651,N_5456,N_5541);
nor U5652 (N_5652,N_5438,N_5511);
nor U5653 (N_5653,N_5590,N_5468);
or U5654 (N_5654,N_5475,N_5529);
or U5655 (N_5655,N_5582,N_5462);
xor U5656 (N_5656,N_5483,N_5446);
and U5657 (N_5657,N_5414,N_5543);
and U5658 (N_5658,N_5441,N_5571);
nand U5659 (N_5659,N_5465,N_5522);
nand U5660 (N_5660,N_5424,N_5466);
xor U5661 (N_5661,N_5472,N_5463);
and U5662 (N_5662,N_5530,N_5487);
nand U5663 (N_5663,N_5578,N_5554);
or U5664 (N_5664,N_5444,N_5563);
and U5665 (N_5665,N_5550,N_5549);
nand U5666 (N_5666,N_5579,N_5539);
or U5667 (N_5667,N_5480,N_5566);
or U5668 (N_5668,N_5427,N_5576);
nand U5669 (N_5669,N_5557,N_5520);
and U5670 (N_5670,N_5551,N_5526);
nor U5671 (N_5671,N_5580,N_5408);
nand U5672 (N_5672,N_5599,N_5524);
or U5673 (N_5673,N_5411,N_5484);
nand U5674 (N_5674,N_5570,N_5594);
or U5675 (N_5675,N_5568,N_5400);
nand U5676 (N_5676,N_5542,N_5512);
nand U5677 (N_5677,N_5509,N_5428);
nand U5678 (N_5678,N_5497,N_5470);
and U5679 (N_5679,N_5573,N_5503);
and U5680 (N_5680,N_5422,N_5538);
or U5681 (N_5681,N_5561,N_5519);
and U5682 (N_5682,N_5477,N_5435);
or U5683 (N_5683,N_5467,N_5425);
nand U5684 (N_5684,N_5485,N_5500);
nor U5685 (N_5685,N_5584,N_5458);
nand U5686 (N_5686,N_5506,N_5540);
xor U5687 (N_5687,N_5413,N_5591);
or U5688 (N_5688,N_5544,N_5532);
nand U5689 (N_5689,N_5589,N_5433);
and U5690 (N_5690,N_5531,N_5439);
nor U5691 (N_5691,N_5431,N_5510);
xor U5692 (N_5692,N_5405,N_5575);
nand U5693 (N_5693,N_5426,N_5528);
nand U5694 (N_5694,N_5565,N_5445);
nand U5695 (N_5695,N_5482,N_5452);
nor U5696 (N_5696,N_5481,N_5587);
or U5697 (N_5697,N_5521,N_5558);
or U5698 (N_5698,N_5476,N_5588);
nand U5699 (N_5699,N_5434,N_5501);
and U5700 (N_5700,N_5427,N_5459);
nand U5701 (N_5701,N_5433,N_5458);
xor U5702 (N_5702,N_5586,N_5590);
and U5703 (N_5703,N_5429,N_5519);
xor U5704 (N_5704,N_5415,N_5580);
nand U5705 (N_5705,N_5542,N_5487);
xor U5706 (N_5706,N_5516,N_5559);
nand U5707 (N_5707,N_5543,N_5555);
and U5708 (N_5708,N_5573,N_5438);
and U5709 (N_5709,N_5433,N_5464);
nor U5710 (N_5710,N_5580,N_5593);
or U5711 (N_5711,N_5508,N_5521);
nor U5712 (N_5712,N_5483,N_5525);
xor U5713 (N_5713,N_5596,N_5583);
nand U5714 (N_5714,N_5527,N_5493);
and U5715 (N_5715,N_5501,N_5458);
and U5716 (N_5716,N_5410,N_5543);
and U5717 (N_5717,N_5512,N_5436);
or U5718 (N_5718,N_5415,N_5542);
or U5719 (N_5719,N_5508,N_5589);
or U5720 (N_5720,N_5525,N_5441);
nand U5721 (N_5721,N_5550,N_5448);
xnor U5722 (N_5722,N_5412,N_5454);
nor U5723 (N_5723,N_5425,N_5498);
xnor U5724 (N_5724,N_5479,N_5505);
nor U5725 (N_5725,N_5497,N_5407);
nand U5726 (N_5726,N_5403,N_5589);
xnor U5727 (N_5727,N_5524,N_5490);
nor U5728 (N_5728,N_5416,N_5592);
or U5729 (N_5729,N_5466,N_5471);
xnor U5730 (N_5730,N_5483,N_5449);
nor U5731 (N_5731,N_5563,N_5489);
xnor U5732 (N_5732,N_5495,N_5598);
xor U5733 (N_5733,N_5539,N_5529);
and U5734 (N_5734,N_5567,N_5502);
and U5735 (N_5735,N_5412,N_5410);
xor U5736 (N_5736,N_5563,N_5570);
nand U5737 (N_5737,N_5538,N_5529);
or U5738 (N_5738,N_5596,N_5421);
nand U5739 (N_5739,N_5475,N_5464);
nor U5740 (N_5740,N_5549,N_5412);
xnor U5741 (N_5741,N_5468,N_5565);
nand U5742 (N_5742,N_5407,N_5501);
or U5743 (N_5743,N_5468,N_5494);
nor U5744 (N_5744,N_5466,N_5421);
nand U5745 (N_5745,N_5480,N_5419);
xor U5746 (N_5746,N_5565,N_5498);
nand U5747 (N_5747,N_5572,N_5465);
and U5748 (N_5748,N_5405,N_5417);
nand U5749 (N_5749,N_5489,N_5502);
nand U5750 (N_5750,N_5594,N_5578);
xor U5751 (N_5751,N_5589,N_5425);
nor U5752 (N_5752,N_5505,N_5515);
nor U5753 (N_5753,N_5481,N_5478);
and U5754 (N_5754,N_5418,N_5510);
xnor U5755 (N_5755,N_5454,N_5555);
xor U5756 (N_5756,N_5533,N_5406);
or U5757 (N_5757,N_5428,N_5568);
and U5758 (N_5758,N_5418,N_5544);
nor U5759 (N_5759,N_5584,N_5538);
nor U5760 (N_5760,N_5466,N_5478);
and U5761 (N_5761,N_5466,N_5411);
nand U5762 (N_5762,N_5456,N_5591);
xnor U5763 (N_5763,N_5583,N_5422);
and U5764 (N_5764,N_5493,N_5536);
or U5765 (N_5765,N_5410,N_5562);
or U5766 (N_5766,N_5415,N_5416);
xnor U5767 (N_5767,N_5483,N_5464);
xnor U5768 (N_5768,N_5486,N_5569);
nand U5769 (N_5769,N_5423,N_5450);
nor U5770 (N_5770,N_5485,N_5522);
nand U5771 (N_5771,N_5578,N_5512);
and U5772 (N_5772,N_5451,N_5535);
xor U5773 (N_5773,N_5556,N_5489);
and U5774 (N_5774,N_5402,N_5525);
nor U5775 (N_5775,N_5502,N_5475);
and U5776 (N_5776,N_5599,N_5525);
nand U5777 (N_5777,N_5527,N_5410);
or U5778 (N_5778,N_5515,N_5513);
and U5779 (N_5779,N_5532,N_5481);
nand U5780 (N_5780,N_5542,N_5413);
xnor U5781 (N_5781,N_5492,N_5457);
nand U5782 (N_5782,N_5470,N_5504);
and U5783 (N_5783,N_5502,N_5588);
and U5784 (N_5784,N_5566,N_5547);
and U5785 (N_5785,N_5518,N_5584);
xnor U5786 (N_5786,N_5569,N_5507);
nor U5787 (N_5787,N_5468,N_5589);
xnor U5788 (N_5788,N_5557,N_5554);
xnor U5789 (N_5789,N_5589,N_5551);
nand U5790 (N_5790,N_5415,N_5401);
nand U5791 (N_5791,N_5522,N_5479);
and U5792 (N_5792,N_5508,N_5450);
xnor U5793 (N_5793,N_5593,N_5482);
nor U5794 (N_5794,N_5569,N_5594);
xor U5795 (N_5795,N_5447,N_5438);
nor U5796 (N_5796,N_5533,N_5547);
or U5797 (N_5797,N_5562,N_5457);
nor U5798 (N_5798,N_5592,N_5485);
xor U5799 (N_5799,N_5507,N_5535);
xnor U5800 (N_5800,N_5682,N_5778);
nor U5801 (N_5801,N_5662,N_5741);
and U5802 (N_5802,N_5645,N_5796);
and U5803 (N_5803,N_5616,N_5607);
xor U5804 (N_5804,N_5679,N_5769);
nor U5805 (N_5805,N_5759,N_5749);
nor U5806 (N_5806,N_5795,N_5736);
nor U5807 (N_5807,N_5617,N_5794);
nor U5808 (N_5808,N_5764,N_5687);
or U5809 (N_5809,N_5601,N_5709);
and U5810 (N_5810,N_5746,N_5660);
nand U5811 (N_5811,N_5638,N_5781);
nor U5812 (N_5812,N_5658,N_5694);
xnor U5813 (N_5813,N_5791,N_5716);
xnor U5814 (N_5814,N_5634,N_5783);
xnor U5815 (N_5815,N_5792,N_5632);
or U5816 (N_5816,N_5624,N_5717);
nor U5817 (N_5817,N_5665,N_5603);
xnor U5818 (N_5818,N_5748,N_5643);
nor U5819 (N_5819,N_5644,N_5674);
nand U5820 (N_5820,N_5788,N_5630);
nor U5821 (N_5821,N_5712,N_5670);
xnor U5822 (N_5822,N_5691,N_5787);
nand U5823 (N_5823,N_5742,N_5752);
xor U5824 (N_5824,N_5680,N_5790);
xor U5825 (N_5825,N_5744,N_5641);
or U5826 (N_5826,N_5618,N_5668);
and U5827 (N_5827,N_5753,N_5614);
or U5828 (N_5828,N_5775,N_5779);
xor U5829 (N_5829,N_5755,N_5737);
and U5830 (N_5830,N_5667,N_5719);
xnor U5831 (N_5831,N_5689,N_5756);
nand U5832 (N_5832,N_5653,N_5705);
nand U5833 (N_5833,N_5762,N_5777);
and U5834 (N_5834,N_5728,N_5707);
and U5835 (N_5835,N_5743,N_5760);
or U5836 (N_5836,N_5609,N_5798);
or U5837 (N_5837,N_5782,N_5715);
xnor U5838 (N_5838,N_5718,N_5704);
nor U5839 (N_5839,N_5612,N_5771);
and U5840 (N_5840,N_5686,N_5611);
or U5841 (N_5841,N_5730,N_5710);
nand U5842 (N_5842,N_5797,N_5733);
nand U5843 (N_5843,N_5692,N_5640);
nor U5844 (N_5844,N_5786,N_5672);
nand U5845 (N_5845,N_5620,N_5697);
xor U5846 (N_5846,N_5745,N_5631);
or U5847 (N_5847,N_5673,N_5659);
nor U5848 (N_5848,N_5669,N_5766);
or U5849 (N_5849,N_5608,N_5765);
and U5850 (N_5850,N_5642,N_5625);
nor U5851 (N_5851,N_5636,N_5706);
and U5852 (N_5852,N_5734,N_5610);
nand U5853 (N_5853,N_5619,N_5780);
xor U5854 (N_5854,N_5681,N_5621);
nand U5855 (N_5855,N_5700,N_5626);
nor U5856 (N_5856,N_5684,N_5725);
or U5857 (N_5857,N_5649,N_5683);
nor U5858 (N_5858,N_5648,N_5677);
or U5859 (N_5859,N_5713,N_5761);
and U5860 (N_5860,N_5767,N_5637);
nand U5861 (N_5861,N_5664,N_5652);
xnor U5862 (N_5862,N_5678,N_5747);
xor U5863 (N_5863,N_5639,N_5606);
nor U5864 (N_5864,N_5785,N_5698);
or U5865 (N_5865,N_5774,N_5615);
nand U5866 (N_5866,N_5789,N_5655);
nor U5867 (N_5867,N_5758,N_5699);
nand U5868 (N_5868,N_5726,N_5627);
or U5869 (N_5869,N_5666,N_5635);
nand U5870 (N_5870,N_5754,N_5696);
and U5871 (N_5871,N_5708,N_5629);
nand U5872 (N_5872,N_5602,N_5732);
nand U5873 (N_5873,N_5628,N_5757);
nand U5874 (N_5874,N_5650,N_5651);
xor U5875 (N_5875,N_5770,N_5695);
and U5876 (N_5876,N_5722,N_5661);
or U5877 (N_5877,N_5702,N_5711);
nand U5878 (N_5878,N_5654,N_5772);
nor U5879 (N_5879,N_5776,N_5633);
xnor U5880 (N_5880,N_5671,N_5693);
nand U5881 (N_5881,N_5723,N_5721);
nand U5882 (N_5882,N_5604,N_5729);
nor U5883 (N_5883,N_5793,N_5646);
or U5884 (N_5884,N_5663,N_5688);
nor U5885 (N_5885,N_5763,N_5685);
nand U5886 (N_5886,N_5720,N_5600);
and U5887 (N_5887,N_5724,N_5703);
nor U5888 (N_5888,N_5799,N_5605);
and U5889 (N_5889,N_5751,N_5701);
nor U5890 (N_5890,N_5613,N_5676);
nand U5891 (N_5891,N_5675,N_5623);
nand U5892 (N_5892,N_5740,N_5690);
nand U5893 (N_5893,N_5750,N_5714);
or U5894 (N_5894,N_5739,N_5768);
nor U5895 (N_5895,N_5773,N_5622);
or U5896 (N_5896,N_5784,N_5731);
nor U5897 (N_5897,N_5735,N_5647);
nor U5898 (N_5898,N_5738,N_5656);
nor U5899 (N_5899,N_5657,N_5727);
nand U5900 (N_5900,N_5630,N_5697);
xnor U5901 (N_5901,N_5661,N_5670);
or U5902 (N_5902,N_5788,N_5741);
nand U5903 (N_5903,N_5798,N_5702);
and U5904 (N_5904,N_5742,N_5725);
nand U5905 (N_5905,N_5742,N_5627);
and U5906 (N_5906,N_5603,N_5790);
nand U5907 (N_5907,N_5734,N_5716);
nor U5908 (N_5908,N_5693,N_5660);
and U5909 (N_5909,N_5760,N_5642);
nand U5910 (N_5910,N_5652,N_5704);
and U5911 (N_5911,N_5644,N_5684);
nor U5912 (N_5912,N_5607,N_5680);
nor U5913 (N_5913,N_5760,N_5679);
nand U5914 (N_5914,N_5761,N_5736);
or U5915 (N_5915,N_5654,N_5684);
xnor U5916 (N_5916,N_5643,N_5731);
or U5917 (N_5917,N_5781,N_5615);
nor U5918 (N_5918,N_5667,N_5712);
or U5919 (N_5919,N_5664,N_5714);
or U5920 (N_5920,N_5798,N_5727);
and U5921 (N_5921,N_5766,N_5790);
nand U5922 (N_5922,N_5646,N_5764);
xnor U5923 (N_5923,N_5677,N_5664);
or U5924 (N_5924,N_5784,N_5725);
nor U5925 (N_5925,N_5669,N_5653);
nand U5926 (N_5926,N_5649,N_5715);
nor U5927 (N_5927,N_5756,N_5688);
xor U5928 (N_5928,N_5739,N_5659);
xnor U5929 (N_5929,N_5772,N_5609);
and U5930 (N_5930,N_5662,N_5695);
and U5931 (N_5931,N_5698,N_5741);
nor U5932 (N_5932,N_5723,N_5630);
xnor U5933 (N_5933,N_5659,N_5705);
or U5934 (N_5934,N_5626,N_5748);
or U5935 (N_5935,N_5770,N_5727);
xnor U5936 (N_5936,N_5794,N_5696);
or U5937 (N_5937,N_5667,N_5650);
and U5938 (N_5938,N_5798,N_5790);
xor U5939 (N_5939,N_5632,N_5645);
xnor U5940 (N_5940,N_5694,N_5634);
and U5941 (N_5941,N_5739,N_5762);
nand U5942 (N_5942,N_5686,N_5630);
xnor U5943 (N_5943,N_5648,N_5688);
xnor U5944 (N_5944,N_5704,N_5716);
nor U5945 (N_5945,N_5786,N_5766);
nand U5946 (N_5946,N_5616,N_5767);
xnor U5947 (N_5947,N_5775,N_5703);
and U5948 (N_5948,N_5610,N_5611);
xnor U5949 (N_5949,N_5701,N_5672);
nand U5950 (N_5950,N_5664,N_5706);
and U5951 (N_5951,N_5683,N_5666);
nor U5952 (N_5952,N_5645,N_5649);
or U5953 (N_5953,N_5766,N_5796);
nor U5954 (N_5954,N_5690,N_5758);
xnor U5955 (N_5955,N_5789,N_5762);
and U5956 (N_5956,N_5626,N_5661);
xor U5957 (N_5957,N_5624,N_5766);
and U5958 (N_5958,N_5672,N_5663);
nor U5959 (N_5959,N_5702,N_5743);
and U5960 (N_5960,N_5676,N_5733);
and U5961 (N_5961,N_5698,N_5772);
nor U5962 (N_5962,N_5701,N_5788);
and U5963 (N_5963,N_5671,N_5707);
or U5964 (N_5964,N_5745,N_5711);
or U5965 (N_5965,N_5792,N_5674);
xor U5966 (N_5966,N_5726,N_5777);
xnor U5967 (N_5967,N_5669,N_5697);
and U5968 (N_5968,N_5768,N_5726);
xor U5969 (N_5969,N_5798,N_5688);
and U5970 (N_5970,N_5695,N_5683);
and U5971 (N_5971,N_5628,N_5703);
nand U5972 (N_5972,N_5789,N_5792);
nor U5973 (N_5973,N_5624,N_5633);
xor U5974 (N_5974,N_5743,N_5765);
nor U5975 (N_5975,N_5659,N_5754);
or U5976 (N_5976,N_5787,N_5758);
nor U5977 (N_5977,N_5712,N_5761);
or U5978 (N_5978,N_5681,N_5646);
and U5979 (N_5979,N_5739,N_5774);
nand U5980 (N_5980,N_5769,N_5685);
nand U5981 (N_5981,N_5795,N_5739);
nand U5982 (N_5982,N_5792,N_5658);
nor U5983 (N_5983,N_5624,N_5736);
nand U5984 (N_5984,N_5775,N_5630);
nor U5985 (N_5985,N_5675,N_5619);
or U5986 (N_5986,N_5607,N_5760);
nor U5987 (N_5987,N_5611,N_5626);
nor U5988 (N_5988,N_5736,N_5645);
nand U5989 (N_5989,N_5769,N_5745);
nor U5990 (N_5990,N_5782,N_5794);
nor U5991 (N_5991,N_5766,N_5602);
or U5992 (N_5992,N_5772,N_5758);
and U5993 (N_5993,N_5761,N_5730);
nand U5994 (N_5994,N_5732,N_5775);
nor U5995 (N_5995,N_5787,N_5745);
xnor U5996 (N_5996,N_5725,N_5606);
nor U5997 (N_5997,N_5613,N_5687);
xnor U5998 (N_5998,N_5728,N_5731);
nor U5999 (N_5999,N_5705,N_5707);
nand U6000 (N_6000,N_5929,N_5856);
and U6001 (N_6001,N_5881,N_5967);
or U6002 (N_6002,N_5859,N_5830);
or U6003 (N_6003,N_5957,N_5923);
nor U6004 (N_6004,N_5840,N_5991);
and U6005 (N_6005,N_5926,N_5836);
nand U6006 (N_6006,N_5997,N_5839);
nor U6007 (N_6007,N_5925,N_5921);
and U6008 (N_6008,N_5936,N_5828);
nand U6009 (N_6009,N_5905,N_5998);
nand U6010 (N_6010,N_5949,N_5866);
or U6011 (N_6011,N_5910,N_5976);
and U6012 (N_6012,N_5847,N_5915);
and U6013 (N_6013,N_5906,N_5927);
and U6014 (N_6014,N_5803,N_5988);
xnor U6015 (N_6015,N_5911,N_5950);
or U6016 (N_6016,N_5855,N_5874);
and U6017 (N_6017,N_5885,N_5817);
xor U6018 (N_6018,N_5992,N_5939);
nor U6019 (N_6019,N_5888,N_5959);
or U6020 (N_6020,N_5878,N_5909);
or U6021 (N_6021,N_5889,N_5837);
xor U6022 (N_6022,N_5989,N_5864);
and U6023 (N_6023,N_5970,N_5971);
xor U6024 (N_6024,N_5984,N_5813);
or U6025 (N_6025,N_5882,N_5816);
and U6026 (N_6026,N_5850,N_5987);
and U6027 (N_6027,N_5823,N_5873);
and U6028 (N_6028,N_5933,N_5819);
and U6029 (N_6029,N_5846,N_5952);
nor U6030 (N_6030,N_5996,N_5809);
and U6031 (N_6031,N_5938,N_5831);
xor U6032 (N_6032,N_5886,N_5972);
xnor U6033 (N_6033,N_5969,N_5851);
or U6034 (N_6034,N_5835,N_5807);
and U6035 (N_6035,N_5993,N_5907);
and U6036 (N_6036,N_5951,N_5860);
xor U6037 (N_6037,N_5867,N_5812);
nand U6038 (N_6038,N_5872,N_5948);
nand U6039 (N_6039,N_5945,N_5980);
and U6040 (N_6040,N_5820,N_5887);
nor U6041 (N_6041,N_5919,N_5917);
or U6042 (N_6042,N_5838,N_5894);
xnor U6043 (N_6043,N_5897,N_5883);
and U6044 (N_6044,N_5893,N_5900);
nor U6045 (N_6045,N_5833,N_5901);
nor U6046 (N_6046,N_5953,N_5822);
xnor U6047 (N_6047,N_5814,N_5958);
nand U6048 (N_6048,N_5890,N_5986);
nand U6049 (N_6049,N_5841,N_5918);
or U6050 (N_6050,N_5931,N_5818);
xor U6051 (N_6051,N_5962,N_5990);
nand U6052 (N_6052,N_5854,N_5960);
nor U6053 (N_6053,N_5937,N_5827);
nor U6054 (N_6054,N_5832,N_5963);
or U6055 (N_6055,N_5943,N_5928);
nor U6056 (N_6056,N_5935,N_5940);
xnor U6057 (N_6057,N_5876,N_5930);
or U6058 (N_6058,N_5995,N_5942);
nor U6059 (N_6059,N_5973,N_5974);
and U6060 (N_6060,N_5824,N_5884);
nor U6061 (N_6061,N_5826,N_5898);
or U6062 (N_6062,N_5869,N_5810);
xor U6063 (N_6063,N_5868,N_5982);
xor U6064 (N_6064,N_5983,N_5999);
or U6065 (N_6065,N_5896,N_5870);
and U6066 (N_6066,N_5922,N_5968);
nor U6067 (N_6067,N_5857,N_5956);
or U6068 (N_6068,N_5975,N_5863);
and U6069 (N_6069,N_5802,N_5892);
or U6070 (N_6070,N_5912,N_5964);
nand U6071 (N_6071,N_5934,N_5804);
and U6072 (N_6072,N_5916,N_5902);
xor U6073 (N_6073,N_5941,N_5944);
xor U6074 (N_6074,N_5852,N_5899);
xnor U6075 (N_6075,N_5806,N_5924);
or U6076 (N_6076,N_5853,N_5801);
and U6077 (N_6077,N_5811,N_5877);
or U6078 (N_6078,N_5842,N_5932);
nor U6079 (N_6079,N_5848,N_5844);
or U6080 (N_6080,N_5977,N_5808);
xnor U6081 (N_6081,N_5834,N_5845);
nor U6082 (N_6082,N_5805,N_5843);
nor U6083 (N_6083,N_5829,N_5880);
nor U6084 (N_6084,N_5815,N_5965);
xnor U6085 (N_6085,N_5849,N_5947);
or U6086 (N_6086,N_5979,N_5861);
and U6087 (N_6087,N_5800,N_5821);
xnor U6088 (N_6088,N_5920,N_5862);
nand U6089 (N_6089,N_5994,N_5946);
and U6090 (N_6090,N_5891,N_5985);
or U6091 (N_6091,N_5978,N_5966);
and U6092 (N_6092,N_5913,N_5908);
xnor U6093 (N_6093,N_5895,N_5981);
nand U6094 (N_6094,N_5865,N_5903);
or U6095 (N_6095,N_5954,N_5825);
or U6096 (N_6096,N_5914,N_5904);
xnor U6097 (N_6097,N_5961,N_5955);
nor U6098 (N_6098,N_5858,N_5879);
and U6099 (N_6099,N_5875,N_5871);
nand U6100 (N_6100,N_5824,N_5948);
or U6101 (N_6101,N_5904,N_5819);
nor U6102 (N_6102,N_5840,N_5819);
xnor U6103 (N_6103,N_5894,N_5947);
nand U6104 (N_6104,N_5963,N_5931);
nor U6105 (N_6105,N_5811,N_5839);
or U6106 (N_6106,N_5811,N_5821);
and U6107 (N_6107,N_5809,N_5992);
or U6108 (N_6108,N_5874,N_5959);
or U6109 (N_6109,N_5827,N_5907);
and U6110 (N_6110,N_5961,N_5883);
nand U6111 (N_6111,N_5835,N_5883);
or U6112 (N_6112,N_5976,N_5926);
and U6113 (N_6113,N_5959,N_5923);
xnor U6114 (N_6114,N_5803,N_5835);
xor U6115 (N_6115,N_5830,N_5856);
nor U6116 (N_6116,N_5943,N_5947);
and U6117 (N_6117,N_5987,N_5965);
nand U6118 (N_6118,N_5878,N_5854);
xnor U6119 (N_6119,N_5995,N_5973);
nor U6120 (N_6120,N_5810,N_5948);
xor U6121 (N_6121,N_5906,N_5950);
nor U6122 (N_6122,N_5949,N_5946);
nand U6123 (N_6123,N_5892,N_5848);
or U6124 (N_6124,N_5927,N_5973);
nand U6125 (N_6125,N_5943,N_5944);
and U6126 (N_6126,N_5919,N_5861);
or U6127 (N_6127,N_5974,N_5975);
nor U6128 (N_6128,N_5859,N_5815);
nor U6129 (N_6129,N_5931,N_5895);
or U6130 (N_6130,N_5959,N_5977);
and U6131 (N_6131,N_5978,N_5841);
and U6132 (N_6132,N_5837,N_5810);
xor U6133 (N_6133,N_5869,N_5881);
and U6134 (N_6134,N_5875,N_5967);
nor U6135 (N_6135,N_5983,N_5980);
and U6136 (N_6136,N_5840,N_5877);
xor U6137 (N_6137,N_5803,N_5987);
nand U6138 (N_6138,N_5938,N_5954);
and U6139 (N_6139,N_5983,N_5824);
nor U6140 (N_6140,N_5932,N_5943);
or U6141 (N_6141,N_5829,N_5918);
nand U6142 (N_6142,N_5990,N_5953);
nor U6143 (N_6143,N_5832,N_5885);
xor U6144 (N_6144,N_5993,N_5875);
nor U6145 (N_6145,N_5938,N_5902);
nand U6146 (N_6146,N_5927,N_5805);
nor U6147 (N_6147,N_5991,N_5974);
xnor U6148 (N_6148,N_5943,N_5861);
xor U6149 (N_6149,N_5939,N_5894);
nor U6150 (N_6150,N_5858,N_5856);
nand U6151 (N_6151,N_5808,N_5811);
or U6152 (N_6152,N_5885,N_5853);
and U6153 (N_6153,N_5833,N_5967);
xnor U6154 (N_6154,N_5829,N_5953);
nand U6155 (N_6155,N_5962,N_5860);
nor U6156 (N_6156,N_5875,N_5807);
or U6157 (N_6157,N_5840,N_5805);
or U6158 (N_6158,N_5814,N_5874);
or U6159 (N_6159,N_5971,N_5812);
xnor U6160 (N_6160,N_5919,N_5853);
nand U6161 (N_6161,N_5943,N_5904);
and U6162 (N_6162,N_5827,N_5995);
nand U6163 (N_6163,N_5889,N_5806);
and U6164 (N_6164,N_5858,N_5863);
nor U6165 (N_6165,N_5934,N_5970);
or U6166 (N_6166,N_5873,N_5929);
and U6167 (N_6167,N_5854,N_5813);
and U6168 (N_6168,N_5993,N_5944);
and U6169 (N_6169,N_5801,N_5877);
and U6170 (N_6170,N_5997,N_5841);
or U6171 (N_6171,N_5914,N_5890);
xor U6172 (N_6172,N_5913,N_5988);
xor U6173 (N_6173,N_5814,N_5824);
and U6174 (N_6174,N_5984,N_5936);
xnor U6175 (N_6175,N_5816,N_5958);
nand U6176 (N_6176,N_5913,N_5876);
xor U6177 (N_6177,N_5945,N_5850);
nor U6178 (N_6178,N_5856,N_5885);
xor U6179 (N_6179,N_5960,N_5972);
and U6180 (N_6180,N_5966,N_5980);
nand U6181 (N_6181,N_5975,N_5930);
and U6182 (N_6182,N_5800,N_5890);
nand U6183 (N_6183,N_5983,N_5876);
and U6184 (N_6184,N_5835,N_5831);
nor U6185 (N_6185,N_5808,N_5917);
nor U6186 (N_6186,N_5815,N_5881);
or U6187 (N_6187,N_5878,N_5960);
nor U6188 (N_6188,N_5803,N_5888);
nor U6189 (N_6189,N_5896,N_5846);
nor U6190 (N_6190,N_5926,N_5848);
nor U6191 (N_6191,N_5962,N_5811);
or U6192 (N_6192,N_5933,N_5944);
nand U6193 (N_6193,N_5918,N_5866);
nor U6194 (N_6194,N_5803,N_5869);
and U6195 (N_6195,N_5911,N_5997);
nor U6196 (N_6196,N_5824,N_5892);
xor U6197 (N_6197,N_5973,N_5904);
and U6198 (N_6198,N_5846,N_5863);
and U6199 (N_6199,N_5810,N_5842);
xor U6200 (N_6200,N_6028,N_6034);
nor U6201 (N_6201,N_6086,N_6142);
xor U6202 (N_6202,N_6174,N_6193);
nand U6203 (N_6203,N_6137,N_6003);
or U6204 (N_6204,N_6143,N_6195);
nand U6205 (N_6205,N_6103,N_6129);
nor U6206 (N_6206,N_6116,N_6110);
or U6207 (N_6207,N_6097,N_6173);
nor U6208 (N_6208,N_6198,N_6049);
xor U6209 (N_6209,N_6043,N_6088);
xor U6210 (N_6210,N_6172,N_6082);
nor U6211 (N_6211,N_6163,N_6153);
xor U6212 (N_6212,N_6108,N_6022);
xor U6213 (N_6213,N_6181,N_6117);
nand U6214 (N_6214,N_6111,N_6178);
nor U6215 (N_6215,N_6096,N_6112);
or U6216 (N_6216,N_6199,N_6044);
and U6217 (N_6217,N_6139,N_6134);
and U6218 (N_6218,N_6125,N_6026);
xnor U6219 (N_6219,N_6128,N_6188);
xnor U6220 (N_6220,N_6085,N_6042);
or U6221 (N_6221,N_6063,N_6057);
nand U6222 (N_6222,N_6030,N_6098);
nor U6223 (N_6223,N_6033,N_6020);
nor U6224 (N_6224,N_6152,N_6005);
and U6225 (N_6225,N_6048,N_6131);
nor U6226 (N_6226,N_6038,N_6056);
nand U6227 (N_6227,N_6079,N_6169);
and U6228 (N_6228,N_6059,N_6055);
and U6229 (N_6229,N_6120,N_6018);
nand U6230 (N_6230,N_6100,N_6076);
xor U6231 (N_6231,N_6113,N_6000);
nand U6232 (N_6232,N_6095,N_6107);
or U6233 (N_6233,N_6104,N_6035);
or U6234 (N_6234,N_6058,N_6187);
and U6235 (N_6235,N_6092,N_6122);
xnor U6236 (N_6236,N_6151,N_6023);
or U6237 (N_6237,N_6166,N_6191);
nor U6238 (N_6238,N_6062,N_6013);
or U6239 (N_6239,N_6135,N_6007);
nand U6240 (N_6240,N_6154,N_6075);
and U6241 (N_6241,N_6155,N_6146);
and U6242 (N_6242,N_6010,N_6041);
and U6243 (N_6243,N_6133,N_6051);
or U6244 (N_6244,N_6066,N_6077);
and U6245 (N_6245,N_6127,N_6150);
nor U6246 (N_6246,N_6024,N_6118);
or U6247 (N_6247,N_6130,N_6064);
nor U6248 (N_6248,N_6138,N_6185);
or U6249 (N_6249,N_6012,N_6084);
xnor U6250 (N_6250,N_6186,N_6016);
nand U6251 (N_6251,N_6065,N_6194);
or U6252 (N_6252,N_6109,N_6009);
xor U6253 (N_6253,N_6053,N_6080);
and U6254 (N_6254,N_6196,N_6072);
and U6255 (N_6255,N_6180,N_6037);
xnor U6256 (N_6256,N_6182,N_6011);
and U6257 (N_6257,N_6078,N_6147);
nand U6258 (N_6258,N_6145,N_6074);
nand U6259 (N_6259,N_6031,N_6073);
nand U6260 (N_6260,N_6175,N_6019);
nor U6261 (N_6261,N_6148,N_6170);
or U6262 (N_6262,N_6017,N_6032);
nand U6263 (N_6263,N_6156,N_6021);
nor U6264 (N_6264,N_6114,N_6036);
xnor U6265 (N_6265,N_6029,N_6069);
or U6266 (N_6266,N_6183,N_6008);
and U6267 (N_6267,N_6162,N_6083);
or U6268 (N_6268,N_6046,N_6165);
xnor U6269 (N_6269,N_6071,N_6039);
nand U6270 (N_6270,N_6176,N_6171);
or U6271 (N_6271,N_6192,N_6106);
nor U6272 (N_6272,N_6091,N_6050);
nand U6273 (N_6273,N_6157,N_6115);
or U6274 (N_6274,N_6102,N_6070);
xor U6275 (N_6275,N_6159,N_6184);
xor U6276 (N_6276,N_6126,N_6067);
and U6277 (N_6277,N_6167,N_6094);
and U6278 (N_6278,N_6087,N_6006);
xnor U6279 (N_6279,N_6132,N_6015);
nor U6280 (N_6280,N_6144,N_6001);
or U6281 (N_6281,N_6052,N_6141);
xor U6282 (N_6282,N_6179,N_6124);
xor U6283 (N_6283,N_6197,N_6123);
nand U6284 (N_6284,N_6045,N_6158);
or U6285 (N_6285,N_6160,N_6025);
nand U6286 (N_6286,N_6149,N_6168);
nand U6287 (N_6287,N_6054,N_6121);
nor U6288 (N_6288,N_6089,N_6004);
nand U6289 (N_6289,N_6136,N_6090);
nor U6290 (N_6290,N_6164,N_6119);
or U6291 (N_6291,N_6081,N_6047);
and U6292 (N_6292,N_6027,N_6061);
nor U6293 (N_6293,N_6105,N_6099);
nor U6294 (N_6294,N_6093,N_6189);
nand U6295 (N_6295,N_6002,N_6177);
or U6296 (N_6296,N_6068,N_6014);
and U6297 (N_6297,N_6060,N_6161);
and U6298 (N_6298,N_6040,N_6190);
or U6299 (N_6299,N_6140,N_6101);
nor U6300 (N_6300,N_6135,N_6177);
or U6301 (N_6301,N_6166,N_6110);
xnor U6302 (N_6302,N_6177,N_6150);
nor U6303 (N_6303,N_6054,N_6050);
nand U6304 (N_6304,N_6087,N_6163);
nor U6305 (N_6305,N_6179,N_6027);
nor U6306 (N_6306,N_6028,N_6136);
or U6307 (N_6307,N_6031,N_6128);
nand U6308 (N_6308,N_6062,N_6042);
xor U6309 (N_6309,N_6109,N_6105);
nand U6310 (N_6310,N_6127,N_6176);
nand U6311 (N_6311,N_6177,N_6075);
or U6312 (N_6312,N_6181,N_6054);
nor U6313 (N_6313,N_6168,N_6017);
xnor U6314 (N_6314,N_6112,N_6013);
nand U6315 (N_6315,N_6122,N_6159);
or U6316 (N_6316,N_6000,N_6055);
nor U6317 (N_6317,N_6132,N_6060);
or U6318 (N_6318,N_6123,N_6162);
nor U6319 (N_6319,N_6140,N_6019);
xor U6320 (N_6320,N_6123,N_6071);
or U6321 (N_6321,N_6167,N_6189);
nand U6322 (N_6322,N_6042,N_6097);
or U6323 (N_6323,N_6028,N_6129);
nand U6324 (N_6324,N_6173,N_6153);
and U6325 (N_6325,N_6107,N_6166);
nand U6326 (N_6326,N_6056,N_6009);
or U6327 (N_6327,N_6003,N_6193);
xor U6328 (N_6328,N_6047,N_6065);
nor U6329 (N_6329,N_6162,N_6011);
or U6330 (N_6330,N_6097,N_6091);
nand U6331 (N_6331,N_6107,N_6021);
nor U6332 (N_6332,N_6164,N_6141);
xor U6333 (N_6333,N_6007,N_6027);
or U6334 (N_6334,N_6106,N_6172);
or U6335 (N_6335,N_6192,N_6102);
or U6336 (N_6336,N_6043,N_6038);
and U6337 (N_6337,N_6146,N_6101);
or U6338 (N_6338,N_6003,N_6141);
or U6339 (N_6339,N_6194,N_6051);
nor U6340 (N_6340,N_6060,N_6089);
nor U6341 (N_6341,N_6127,N_6080);
nand U6342 (N_6342,N_6008,N_6140);
or U6343 (N_6343,N_6034,N_6062);
nand U6344 (N_6344,N_6178,N_6146);
nand U6345 (N_6345,N_6060,N_6155);
and U6346 (N_6346,N_6111,N_6017);
and U6347 (N_6347,N_6172,N_6080);
nand U6348 (N_6348,N_6068,N_6049);
and U6349 (N_6349,N_6063,N_6008);
nand U6350 (N_6350,N_6145,N_6118);
nand U6351 (N_6351,N_6023,N_6061);
nand U6352 (N_6352,N_6101,N_6061);
nand U6353 (N_6353,N_6168,N_6101);
nor U6354 (N_6354,N_6076,N_6043);
or U6355 (N_6355,N_6115,N_6165);
and U6356 (N_6356,N_6109,N_6036);
xor U6357 (N_6357,N_6170,N_6166);
and U6358 (N_6358,N_6176,N_6032);
or U6359 (N_6359,N_6038,N_6103);
xor U6360 (N_6360,N_6134,N_6197);
or U6361 (N_6361,N_6043,N_6065);
nor U6362 (N_6362,N_6055,N_6198);
or U6363 (N_6363,N_6094,N_6190);
and U6364 (N_6364,N_6067,N_6071);
nand U6365 (N_6365,N_6040,N_6004);
nor U6366 (N_6366,N_6143,N_6132);
xor U6367 (N_6367,N_6167,N_6149);
or U6368 (N_6368,N_6157,N_6173);
nand U6369 (N_6369,N_6125,N_6035);
nor U6370 (N_6370,N_6185,N_6036);
nand U6371 (N_6371,N_6117,N_6046);
nor U6372 (N_6372,N_6121,N_6197);
and U6373 (N_6373,N_6098,N_6125);
xor U6374 (N_6374,N_6050,N_6133);
nand U6375 (N_6375,N_6143,N_6007);
xnor U6376 (N_6376,N_6033,N_6162);
nand U6377 (N_6377,N_6051,N_6108);
and U6378 (N_6378,N_6003,N_6185);
nor U6379 (N_6379,N_6008,N_6079);
nand U6380 (N_6380,N_6100,N_6159);
or U6381 (N_6381,N_6007,N_6127);
or U6382 (N_6382,N_6004,N_6172);
and U6383 (N_6383,N_6176,N_6116);
xor U6384 (N_6384,N_6113,N_6046);
nor U6385 (N_6385,N_6056,N_6030);
nand U6386 (N_6386,N_6143,N_6070);
xnor U6387 (N_6387,N_6166,N_6009);
or U6388 (N_6388,N_6154,N_6014);
and U6389 (N_6389,N_6055,N_6083);
nor U6390 (N_6390,N_6045,N_6165);
nand U6391 (N_6391,N_6068,N_6156);
nand U6392 (N_6392,N_6089,N_6061);
nor U6393 (N_6393,N_6045,N_6055);
xnor U6394 (N_6394,N_6037,N_6072);
and U6395 (N_6395,N_6172,N_6126);
and U6396 (N_6396,N_6189,N_6133);
nor U6397 (N_6397,N_6010,N_6178);
or U6398 (N_6398,N_6071,N_6183);
xor U6399 (N_6399,N_6057,N_6027);
or U6400 (N_6400,N_6323,N_6303);
nor U6401 (N_6401,N_6343,N_6265);
nand U6402 (N_6402,N_6273,N_6249);
and U6403 (N_6403,N_6298,N_6350);
nor U6404 (N_6404,N_6378,N_6375);
nor U6405 (N_6405,N_6299,N_6367);
nand U6406 (N_6406,N_6397,N_6208);
or U6407 (N_6407,N_6221,N_6382);
nor U6408 (N_6408,N_6234,N_6289);
xnor U6409 (N_6409,N_6260,N_6347);
nor U6410 (N_6410,N_6241,N_6227);
xnor U6411 (N_6411,N_6387,N_6339);
nand U6412 (N_6412,N_6261,N_6225);
nor U6413 (N_6413,N_6229,N_6310);
nand U6414 (N_6414,N_6304,N_6292);
nor U6415 (N_6415,N_6243,N_6256);
xor U6416 (N_6416,N_6263,N_6270);
nand U6417 (N_6417,N_6223,N_6251);
or U6418 (N_6418,N_6207,N_6321);
nand U6419 (N_6419,N_6317,N_6385);
xnor U6420 (N_6420,N_6202,N_6365);
and U6421 (N_6421,N_6334,N_6286);
xnor U6422 (N_6422,N_6236,N_6340);
nor U6423 (N_6423,N_6253,N_6337);
and U6424 (N_6424,N_6277,N_6248);
nor U6425 (N_6425,N_6206,N_6250);
and U6426 (N_6426,N_6259,N_6362);
nand U6427 (N_6427,N_6266,N_6305);
and U6428 (N_6428,N_6246,N_6281);
and U6429 (N_6429,N_6214,N_6373);
and U6430 (N_6430,N_6218,N_6237);
xnor U6431 (N_6431,N_6257,N_6293);
nor U6432 (N_6432,N_6247,N_6344);
or U6433 (N_6433,N_6242,N_6336);
xor U6434 (N_6434,N_6228,N_6363);
xor U6435 (N_6435,N_6395,N_6268);
or U6436 (N_6436,N_6216,N_6325);
nand U6437 (N_6437,N_6296,N_6307);
xnor U6438 (N_6438,N_6329,N_6211);
or U6439 (N_6439,N_6383,N_6276);
xnor U6440 (N_6440,N_6391,N_6215);
and U6441 (N_6441,N_6244,N_6379);
and U6442 (N_6442,N_6287,N_6278);
and U6443 (N_6443,N_6330,N_6342);
or U6444 (N_6444,N_6275,N_6272);
nor U6445 (N_6445,N_6357,N_6369);
xor U6446 (N_6446,N_6280,N_6359);
or U6447 (N_6447,N_6230,N_6254);
nand U6448 (N_6448,N_6346,N_6291);
nor U6449 (N_6449,N_6302,N_6209);
or U6450 (N_6450,N_6290,N_6399);
nor U6451 (N_6451,N_6376,N_6239);
or U6452 (N_6452,N_6312,N_6372);
nand U6453 (N_6453,N_6220,N_6213);
xnor U6454 (N_6454,N_6233,N_6394);
and U6455 (N_6455,N_6271,N_6327);
xor U6456 (N_6456,N_6390,N_6356);
nand U6457 (N_6457,N_6301,N_6267);
xnor U6458 (N_6458,N_6258,N_6348);
and U6459 (N_6459,N_6354,N_6279);
and U6460 (N_6460,N_6335,N_6297);
or U6461 (N_6461,N_6324,N_6316);
xor U6462 (N_6462,N_6349,N_6288);
nor U6463 (N_6463,N_6381,N_6224);
or U6464 (N_6464,N_6205,N_6384);
and U6465 (N_6465,N_6300,N_6235);
xor U6466 (N_6466,N_6204,N_6283);
nor U6467 (N_6467,N_6309,N_6201);
xnor U6468 (N_6468,N_6351,N_6358);
and U6469 (N_6469,N_6315,N_6360);
or U6470 (N_6470,N_6217,N_6274);
xnor U6471 (N_6471,N_6322,N_6386);
nor U6472 (N_6472,N_6308,N_6314);
nor U6473 (N_6473,N_6313,N_6231);
xnor U6474 (N_6474,N_6238,N_6341);
nand U6475 (N_6475,N_6252,N_6264);
xor U6476 (N_6476,N_6338,N_6388);
xnor U6477 (N_6477,N_6262,N_6232);
nor U6478 (N_6478,N_6226,N_6219);
xor U6479 (N_6479,N_6355,N_6200);
nand U6480 (N_6480,N_6240,N_6212);
nor U6481 (N_6481,N_6245,N_6295);
or U6482 (N_6482,N_6282,N_6396);
nand U6483 (N_6483,N_6326,N_6345);
xor U6484 (N_6484,N_6371,N_6377);
xnor U6485 (N_6485,N_6392,N_6210);
xnor U6486 (N_6486,N_6333,N_6222);
and U6487 (N_6487,N_6368,N_6389);
nand U6488 (N_6488,N_6255,N_6320);
and U6489 (N_6489,N_6328,N_6364);
or U6490 (N_6490,N_6318,N_6374);
nor U6491 (N_6491,N_6366,N_6311);
xnor U6492 (N_6492,N_6361,N_6294);
or U6493 (N_6493,N_6284,N_6352);
or U6494 (N_6494,N_6353,N_6370);
and U6495 (N_6495,N_6331,N_6285);
nor U6496 (N_6496,N_6203,N_6380);
and U6497 (N_6497,N_6269,N_6393);
xnor U6498 (N_6498,N_6398,N_6306);
nand U6499 (N_6499,N_6319,N_6332);
nor U6500 (N_6500,N_6241,N_6263);
or U6501 (N_6501,N_6323,N_6210);
or U6502 (N_6502,N_6374,N_6373);
and U6503 (N_6503,N_6354,N_6272);
and U6504 (N_6504,N_6343,N_6246);
xnor U6505 (N_6505,N_6341,N_6388);
or U6506 (N_6506,N_6230,N_6343);
or U6507 (N_6507,N_6378,N_6350);
nor U6508 (N_6508,N_6255,N_6253);
or U6509 (N_6509,N_6251,N_6397);
and U6510 (N_6510,N_6241,N_6239);
nand U6511 (N_6511,N_6311,N_6261);
xor U6512 (N_6512,N_6232,N_6367);
or U6513 (N_6513,N_6349,N_6386);
and U6514 (N_6514,N_6248,N_6206);
or U6515 (N_6515,N_6204,N_6235);
or U6516 (N_6516,N_6322,N_6397);
xnor U6517 (N_6517,N_6254,N_6375);
or U6518 (N_6518,N_6316,N_6230);
and U6519 (N_6519,N_6317,N_6344);
nand U6520 (N_6520,N_6243,N_6388);
nand U6521 (N_6521,N_6330,N_6344);
xor U6522 (N_6522,N_6242,N_6312);
nand U6523 (N_6523,N_6209,N_6326);
xnor U6524 (N_6524,N_6359,N_6395);
and U6525 (N_6525,N_6300,N_6203);
xnor U6526 (N_6526,N_6203,N_6218);
nand U6527 (N_6527,N_6203,N_6204);
xor U6528 (N_6528,N_6258,N_6256);
xnor U6529 (N_6529,N_6228,N_6350);
or U6530 (N_6530,N_6272,N_6319);
nand U6531 (N_6531,N_6334,N_6339);
or U6532 (N_6532,N_6326,N_6253);
nor U6533 (N_6533,N_6256,N_6222);
and U6534 (N_6534,N_6218,N_6236);
and U6535 (N_6535,N_6395,N_6255);
xor U6536 (N_6536,N_6307,N_6289);
nand U6537 (N_6537,N_6267,N_6379);
nor U6538 (N_6538,N_6319,N_6230);
or U6539 (N_6539,N_6286,N_6230);
nor U6540 (N_6540,N_6263,N_6249);
nand U6541 (N_6541,N_6314,N_6239);
and U6542 (N_6542,N_6300,N_6222);
or U6543 (N_6543,N_6355,N_6243);
nand U6544 (N_6544,N_6337,N_6345);
and U6545 (N_6545,N_6390,N_6344);
and U6546 (N_6546,N_6209,N_6394);
nand U6547 (N_6547,N_6205,N_6329);
or U6548 (N_6548,N_6382,N_6236);
xnor U6549 (N_6549,N_6390,N_6352);
nor U6550 (N_6550,N_6205,N_6382);
nand U6551 (N_6551,N_6203,N_6282);
and U6552 (N_6552,N_6328,N_6359);
or U6553 (N_6553,N_6364,N_6319);
nor U6554 (N_6554,N_6303,N_6206);
and U6555 (N_6555,N_6219,N_6217);
nor U6556 (N_6556,N_6268,N_6238);
nor U6557 (N_6557,N_6348,N_6242);
and U6558 (N_6558,N_6311,N_6309);
nand U6559 (N_6559,N_6270,N_6311);
nor U6560 (N_6560,N_6369,N_6249);
xnor U6561 (N_6561,N_6239,N_6328);
and U6562 (N_6562,N_6324,N_6332);
nand U6563 (N_6563,N_6280,N_6346);
xor U6564 (N_6564,N_6380,N_6233);
xor U6565 (N_6565,N_6274,N_6367);
nand U6566 (N_6566,N_6243,N_6284);
xor U6567 (N_6567,N_6281,N_6308);
and U6568 (N_6568,N_6291,N_6361);
or U6569 (N_6569,N_6269,N_6257);
nand U6570 (N_6570,N_6291,N_6311);
nor U6571 (N_6571,N_6310,N_6372);
nand U6572 (N_6572,N_6214,N_6255);
xor U6573 (N_6573,N_6352,N_6321);
or U6574 (N_6574,N_6324,N_6395);
nor U6575 (N_6575,N_6276,N_6290);
nor U6576 (N_6576,N_6241,N_6382);
and U6577 (N_6577,N_6270,N_6386);
nand U6578 (N_6578,N_6305,N_6272);
xnor U6579 (N_6579,N_6241,N_6262);
nand U6580 (N_6580,N_6283,N_6398);
nor U6581 (N_6581,N_6277,N_6235);
and U6582 (N_6582,N_6266,N_6220);
nand U6583 (N_6583,N_6343,N_6284);
xor U6584 (N_6584,N_6236,N_6310);
nand U6585 (N_6585,N_6277,N_6372);
xnor U6586 (N_6586,N_6385,N_6395);
nor U6587 (N_6587,N_6285,N_6293);
xnor U6588 (N_6588,N_6293,N_6366);
or U6589 (N_6589,N_6384,N_6392);
or U6590 (N_6590,N_6200,N_6239);
nand U6591 (N_6591,N_6309,N_6230);
xnor U6592 (N_6592,N_6284,N_6224);
xnor U6593 (N_6593,N_6216,N_6296);
nand U6594 (N_6594,N_6330,N_6206);
or U6595 (N_6595,N_6382,N_6230);
xor U6596 (N_6596,N_6217,N_6364);
nor U6597 (N_6597,N_6200,N_6284);
nor U6598 (N_6598,N_6200,N_6300);
xnor U6599 (N_6599,N_6375,N_6251);
nand U6600 (N_6600,N_6421,N_6411);
and U6601 (N_6601,N_6414,N_6463);
or U6602 (N_6602,N_6523,N_6549);
and U6603 (N_6603,N_6489,N_6532);
nand U6604 (N_6604,N_6587,N_6468);
and U6605 (N_6605,N_6426,N_6545);
xor U6606 (N_6606,N_6454,N_6563);
or U6607 (N_6607,N_6579,N_6483);
nor U6608 (N_6608,N_6445,N_6435);
and U6609 (N_6609,N_6437,N_6491);
nor U6610 (N_6610,N_6560,N_6590);
or U6611 (N_6611,N_6462,N_6588);
nor U6612 (N_6612,N_6420,N_6510);
xnor U6613 (N_6613,N_6527,N_6548);
nor U6614 (N_6614,N_6551,N_6596);
xnor U6615 (N_6615,N_6506,N_6458);
and U6616 (N_6616,N_6429,N_6584);
nand U6617 (N_6617,N_6474,N_6475);
xor U6618 (N_6618,N_6511,N_6504);
nand U6619 (N_6619,N_6413,N_6455);
or U6620 (N_6620,N_6485,N_6519);
nor U6621 (N_6621,N_6405,N_6492);
or U6622 (N_6622,N_6419,N_6573);
xnor U6623 (N_6623,N_6409,N_6477);
nand U6624 (N_6624,N_6521,N_6503);
xnor U6625 (N_6625,N_6571,N_6402);
nor U6626 (N_6626,N_6577,N_6481);
and U6627 (N_6627,N_6518,N_6436);
and U6628 (N_6628,N_6514,N_6517);
xor U6629 (N_6629,N_6494,N_6479);
xor U6630 (N_6630,N_6448,N_6499);
or U6631 (N_6631,N_6407,N_6487);
xnor U6632 (N_6632,N_6582,N_6403);
nand U6633 (N_6633,N_6442,N_6476);
nand U6634 (N_6634,N_6439,N_6469);
nor U6635 (N_6635,N_6418,N_6456);
and U6636 (N_6636,N_6593,N_6546);
and U6637 (N_6637,N_6417,N_6501);
xnor U6638 (N_6638,N_6452,N_6460);
nor U6639 (N_6639,N_6516,N_6533);
nand U6640 (N_6640,N_6561,N_6470);
nor U6641 (N_6641,N_6430,N_6453);
xnor U6642 (N_6642,N_6434,N_6500);
nand U6643 (N_6643,N_6482,N_6581);
nor U6644 (N_6644,N_6594,N_6423);
or U6645 (N_6645,N_6424,N_6558);
or U6646 (N_6646,N_6450,N_6406);
nor U6647 (N_6647,N_6446,N_6520);
xnor U6648 (N_6648,N_6565,N_6473);
xnor U6649 (N_6649,N_6449,N_6562);
and U6650 (N_6650,N_6459,N_6515);
or U6651 (N_6651,N_6490,N_6444);
xnor U6652 (N_6652,N_6525,N_6522);
nor U6653 (N_6653,N_6583,N_6538);
nand U6654 (N_6654,N_6537,N_6451);
nor U6655 (N_6655,N_6478,N_6528);
and U6656 (N_6656,N_6567,N_6544);
or U6657 (N_6657,N_6438,N_6597);
or U6658 (N_6658,N_6591,N_6440);
and U6659 (N_6659,N_6566,N_6578);
nor U6660 (N_6660,N_6529,N_6472);
nand U6661 (N_6661,N_6592,N_6447);
or U6662 (N_6662,N_6461,N_6428);
nor U6663 (N_6663,N_6408,N_6598);
xor U6664 (N_6664,N_6498,N_6552);
xor U6665 (N_6665,N_6556,N_6540);
nand U6666 (N_6666,N_6502,N_6569);
xor U6667 (N_6667,N_6585,N_6547);
nor U6668 (N_6668,N_6484,N_6572);
nand U6669 (N_6669,N_6542,N_6534);
nand U6670 (N_6670,N_6466,N_6404);
nand U6671 (N_6671,N_6480,N_6550);
nand U6672 (N_6672,N_6557,N_6431);
xnor U6673 (N_6673,N_6559,N_6535);
nand U6674 (N_6674,N_6543,N_6570);
or U6675 (N_6675,N_6495,N_6422);
nor U6676 (N_6676,N_6576,N_6496);
nand U6677 (N_6677,N_6513,N_6505);
xor U6678 (N_6678,N_6531,N_6416);
and U6679 (N_6679,N_6589,N_6465);
xnor U6680 (N_6680,N_6553,N_6574);
or U6681 (N_6681,N_6526,N_6595);
nand U6682 (N_6682,N_6493,N_6539);
and U6683 (N_6683,N_6425,N_6443);
and U6684 (N_6684,N_6568,N_6412);
nand U6685 (N_6685,N_6400,N_6564);
and U6686 (N_6686,N_6586,N_6457);
nand U6687 (N_6687,N_6410,N_6554);
xor U6688 (N_6688,N_6524,N_6467);
xor U6689 (N_6689,N_6486,N_6541);
nor U6690 (N_6690,N_6464,N_6415);
nand U6691 (N_6691,N_6575,N_6488);
xor U6692 (N_6692,N_6427,N_6599);
nor U6693 (N_6693,N_6497,N_6509);
xor U6694 (N_6694,N_6433,N_6580);
xnor U6695 (N_6695,N_6530,N_6512);
nand U6696 (N_6696,N_6441,N_6507);
and U6697 (N_6697,N_6432,N_6471);
xnor U6698 (N_6698,N_6536,N_6508);
or U6699 (N_6699,N_6401,N_6555);
xnor U6700 (N_6700,N_6421,N_6466);
nor U6701 (N_6701,N_6472,N_6560);
and U6702 (N_6702,N_6518,N_6543);
xor U6703 (N_6703,N_6442,N_6413);
nor U6704 (N_6704,N_6472,N_6535);
xor U6705 (N_6705,N_6402,N_6575);
nor U6706 (N_6706,N_6437,N_6507);
nor U6707 (N_6707,N_6472,N_6577);
and U6708 (N_6708,N_6562,N_6461);
and U6709 (N_6709,N_6567,N_6517);
and U6710 (N_6710,N_6520,N_6439);
or U6711 (N_6711,N_6533,N_6596);
xor U6712 (N_6712,N_6437,N_6573);
xor U6713 (N_6713,N_6470,N_6474);
nand U6714 (N_6714,N_6533,N_6446);
nand U6715 (N_6715,N_6533,N_6430);
and U6716 (N_6716,N_6452,N_6561);
xor U6717 (N_6717,N_6451,N_6524);
nand U6718 (N_6718,N_6553,N_6529);
and U6719 (N_6719,N_6473,N_6498);
nand U6720 (N_6720,N_6592,N_6502);
or U6721 (N_6721,N_6504,N_6559);
nor U6722 (N_6722,N_6570,N_6485);
nor U6723 (N_6723,N_6455,N_6597);
xor U6724 (N_6724,N_6546,N_6517);
and U6725 (N_6725,N_6461,N_6490);
xor U6726 (N_6726,N_6447,N_6577);
nor U6727 (N_6727,N_6500,N_6498);
xnor U6728 (N_6728,N_6549,N_6419);
nand U6729 (N_6729,N_6459,N_6562);
xor U6730 (N_6730,N_6552,N_6439);
nor U6731 (N_6731,N_6554,N_6535);
nand U6732 (N_6732,N_6506,N_6431);
nor U6733 (N_6733,N_6423,N_6452);
nor U6734 (N_6734,N_6454,N_6470);
nor U6735 (N_6735,N_6583,N_6455);
or U6736 (N_6736,N_6454,N_6556);
xor U6737 (N_6737,N_6402,N_6576);
and U6738 (N_6738,N_6431,N_6555);
nor U6739 (N_6739,N_6497,N_6447);
nand U6740 (N_6740,N_6471,N_6578);
nand U6741 (N_6741,N_6494,N_6428);
xnor U6742 (N_6742,N_6402,N_6462);
xor U6743 (N_6743,N_6527,N_6509);
nand U6744 (N_6744,N_6557,N_6512);
and U6745 (N_6745,N_6597,N_6506);
nor U6746 (N_6746,N_6545,N_6508);
nor U6747 (N_6747,N_6400,N_6437);
nand U6748 (N_6748,N_6595,N_6579);
nor U6749 (N_6749,N_6554,N_6508);
xnor U6750 (N_6750,N_6510,N_6520);
xor U6751 (N_6751,N_6497,N_6466);
nand U6752 (N_6752,N_6572,N_6433);
xor U6753 (N_6753,N_6406,N_6490);
nand U6754 (N_6754,N_6519,N_6570);
or U6755 (N_6755,N_6565,N_6490);
nand U6756 (N_6756,N_6405,N_6475);
nand U6757 (N_6757,N_6593,N_6428);
and U6758 (N_6758,N_6599,N_6426);
nand U6759 (N_6759,N_6578,N_6473);
nor U6760 (N_6760,N_6429,N_6423);
nor U6761 (N_6761,N_6505,N_6587);
xor U6762 (N_6762,N_6428,N_6503);
nor U6763 (N_6763,N_6590,N_6407);
or U6764 (N_6764,N_6492,N_6545);
or U6765 (N_6765,N_6574,N_6534);
xor U6766 (N_6766,N_6595,N_6403);
and U6767 (N_6767,N_6490,N_6429);
and U6768 (N_6768,N_6415,N_6420);
nor U6769 (N_6769,N_6427,N_6445);
nand U6770 (N_6770,N_6504,N_6537);
nor U6771 (N_6771,N_6513,N_6416);
or U6772 (N_6772,N_6568,N_6480);
nor U6773 (N_6773,N_6588,N_6476);
or U6774 (N_6774,N_6519,N_6560);
nor U6775 (N_6775,N_6464,N_6413);
and U6776 (N_6776,N_6518,N_6434);
xor U6777 (N_6777,N_6576,N_6431);
xnor U6778 (N_6778,N_6550,N_6535);
nand U6779 (N_6779,N_6437,N_6482);
nor U6780 (N_6780,N_6469,N_6416);
or U6781 (N_6781,N_6485,N_6446);
and U6782 (N_6782,N_6477,N_6540);
nand U6783 (N_6783,N_6489,N_6555);
nor U6784 (N_6784,N_6424,N_6487);
nand U6785 (N_6785,N_6418,N_6491);
or U6786 (N_6786,N_6526,N_6599);
nor U6787 (N_6787,N_6503,N_6552);
or U6788 (N_6788,N_6422,N_6536);
nand U6789 (N_6789,N_6585,N_6432);
nand U6790 (N_6790,N_6595,N_6443);
or U6791 (N_6791,N_6460,N_6471);
or U6792 (N_6792,N_6413,N_6559);
and U6793 (N_6793,N_6404,N_6570);
nor U6794 (N_6794,N_6421,N_6413);
or U6795 (N_6795,N_6566,N_6589);
or U6796 (N_6796,N_6495,N_6598);
nor U6797 (N_6797,N_6489,N_6420);
nor U6798 (N_6798,N_6576,N_6427);
nor U6799 (N_6799,N_6540,N_6497);
xnor U6800 (N_6800,N_6618,N_6605);
or U6801 (N_6801,N_6634,N_6650);
or U6802 (N_6802,N_6694,N_6771);
nor U6803 (N_6803,N_6705,N_6672);
xor U6804 (N_6804,N_6777,N_6722);
or U6805 (N_6805,N_6749,N_6610);
xor U6806 (N_6806,N_6666,N_6641);
nor U6807 (N_6807,N_6730,N_6715);
xor U6808 (N_6808,N_6619,N_6707);
nand U6809 (N_6809,N_6796,N_6698);
or U6810 (N_6810,N_6688,N_6713);
or U6811 (N_6811,N_6752,N_6778);
nor U6812 (N_6812,N_6792,N_6660);
xnor U6813 (N_6813,N_6620,N_6714);
xnor U6814 (N_6814,N_6682,N_6793);
nor U6815 (N_6815,N_6656,N_6668);
nand U6816 (N_6816,N_6644,N_6766);
or U6817 (N_6817,N_6731,N_6667);
nand U6818 (N_6818,N_6700,N_6652);
or U6819 (N_6819,N_6779,N_6763);
xor U6820 (N_6820,N_6745,N_6612);
xor U6821 (N_6821,N_6699,N_6642);
xnor U6822 (N_6822,N_6638,N_6692);
or U6823 (N_6823,N_6647,N_6753);
nor U6824 (N_6824,N_6783,N_6616);
nand U6825 (N_6825,N_6720,N_6795);
and U6826 (N_6826,N_6636,N_6663);
and U6827 (N_6827,N_6750,N_6633);
nor U6828 (N_6828,N_6628,N_6780);
or U6829 (N_6829,N_6625,N_6611);
or U6830 (N_6830,N_6737,N_6629);
nor U6831 (N_6831,N_6623,N_6600);
or U6832 (N_6832,N_6704,N_6691);
and U6833 (N_6833,N_6748,N_6662);
nor U6834 (N_6834,N_6751,N_6676);
nor U6835 (N_6835,N_6710,N_6759);
or U6836 (N_6836,N_6643,N_6728);
and U6837 (N_6837,N_6739,N_6788);
xor U6838 (N_6838,N_6661,N_6614);
xnor U6839 (N_6839,N_6635,N_6673);
xor U6840 (N_6840,N_6740,N_6613);
or U6841 (N_6841,N_6726,N_6712);
nor U6842 (N_6842,N_6741,N_6653);
or U6843 (N_6843,N_6729,N_6622);
and U6844 (N_6844,N_6743,N_6790);
xnor U6845 (N_6845,N_6708,N_6786);
nor U6846 (N_6846,N_6669,N_6703);
and U6847 (N_6847,N_6646,N_6723);
xnor U6848 (N_6848,N_6655,N_6609);
nand U6849 (N_6849,N_6761,N_6727);
or U6850 (N_6850,N_6735,N_6794);
nand U6851 (N_6851,N_6626,N_6683);
xor U6852 (N_6852,N_6709,N_6665);
xor U6853 (N_6853,N_6657,N_6744);
xor U6854 (N_6854,N_6798,N_6760);
xnor U6855 (N_6855,N_6640,N_6639);
nor U6856 (N_6856,N_6770,N_6670);
or U6857 (N_6857,N_6637,N_6658);
nand U6858 (N_6858,N_6690,N_6606);
and U6859 (N_6859,N_6717,N_6687);
and U6860 (N_6860,N_6725,N_6696);
or U6861 (N_6861,N_6689,N_6651);
xnor U6862 (N_6862,N_6695,N_6756);
nand U6863 (N_6863,N_6732,N_6724);
or U6864 (N_6864,N_6615,N_6706);
xor U6865 (N_6865,N_6604,N_6603);
or U6866 (N_6866,N_6686,N_6654);
or U6867 (N_6867,N_6693,N_6697);
nor U6868 (N_6868,N_6632,N_6675);
or U6869 (N_6869,N_6601,N_6762);
or U6870 (N_6870,N_6674,N_6701);
or U6871 (N_6871,N_6734,N_6621);
nand U6872 (N_6872,N_6624,N_6738);
nor U6873 (N_6873,N_6671,N_6630);
nor U6874 (N_6874,N_6773,N_6681);
nand U6875 (N_6875,N_6719,N_6765);
and U6876 (N_6876,N_6767,N_6789);
nor U6877 (N_6877,N_6677,N_6742);
xnor U6878 (N_6878,N_6631,N_6608);
or U6879 (N_6879,N_6799,N_6797);
and U6880 (N_6880,N_6758,N_6721);
and U6881 (N_6881,N_6664,N_6781);
and U6882 (N_6882,N_6659,N_6775);
xor U6883 (N_6883,N_6774,N_6736);
nor U6884 (N_6884,N_6702,N_6772);
nand U6885 (N_6885,N_6684,N_6768);
nand U6886 (N_6886,N_6787,N_6648);
xnor U6887 (N_6887,N_6678,N_6685);
and U6888 (N_6888,N_6791,N_6680);
or U6889 (N_6889,N_6782,N_6764);
or U6890 (N_6890,N_6776,N_6711);
nand U6891 (N_6891,N_6716,N_6769);
nor U6892 (N_6892,N_6607,N_6649);
nor U6893 (N_6893,N_6617,N_6718);
and U6894 (N_6894,N_6757,N_6733);
nor U6895 (N_6895,N_6785,N_6746);
xor U6896 (N_6896,N_6747,N_6602);
nand U6897 (N_6897,N_6784,N_6679);
nor U6898 (N_6898,N_6627,N_6755);
nor U6899 (N_6899,N_6645,N_6754);
and U6900 (N_6900,N_6668,N_6696);
and U6901 (N_6901,N_6659,N_6607);
nand U6902 (N_6902,N_6713,N_6762);
nand U6903 (N_6903,N_6694,N_6696);
nand U6904 (N_6904,N_6690,N_6701);
nand U6905 (N_6905,N_6636,N_6773);
and U6906 (N_6906,N_6672,N_6786);
xnor U6907 (N_6907,N_6783,N_6744);
or U6908 (N_6908,N_6714,N_6618);
and U6909 (N_6909,N_6741,N_6755);
and U6910 (N_6910,N_6753,N_6645);
xnor U6911 (N_6911,N_6620,N_6633);
xnor U6912 (N_6912,N_6714,N_6685);
xnor U6913 (N_6913,N_6600,N_6787);
xor U6914 (N_6914,N_6655,N_6723);
xnor U6915 (N_6915,N_6779,N_6764);
nor U6916 (N_6916,N_6786,N_6718);
nand U6917 (N_6917,N_6707,N_6663);
nor U6918 (N_6918,N_6608,N_6741);
or U6919 (N_6919,N_6696,N_6655);
nand U6920 (N_6920,N_6608,N_6693);
xor U6921 (N_6921,N_6763,N_6690);
xor U6922 (N_6922,N_6622,N_6666);
nor U6923 (N_6923,N_6730,N_6793);
and U6924 (N_6924,N_6764,N_6742);
xor U6925 (N_6925,N_6718,N_6621);
nand U6926 (N_6926,N_6748,N_6703);
nand U6927 (N_6927,N_6761,N_6728);
and U6928 (N_6928,N_6659,N_6762);
nand U6929 (N_6929,N_6651,N_6664);
and U6930 (N_6930,N_6784,N_6722);
xnor U6931 (N_6931,N_6640,N_6744);
xnor U6932 (N_6932,N_6650,N_6729);
nor U6933 (N_6933,N_6622,N_6751);
nand U6934 (N_6934,N_6693,N_6768);
xnor U6935 (N_6935,N_6798,N_6666);
xor U6936 (N_6936,N_6688,N_6696);
nand U6937 (N_6937,N_6746,N_6799);
and U6938 (N_6938,N_6661,N_6635);
and U6939 (N_6939,N_6682,N_6622);
nand U6940 (N_6940,N_6701,N_6620);
and U6941 (N_6941,N_6795,N_6670);
or U6942 (N_6942,N_6787,N_6757);
nand U6943 (N_6943,N_6737,N_6780);
xnor U6944 (N_6944,N_6709,N_6694);
and U6945 (N_6945,N_6615,N_6658);
nand U6946 (N_6946,N_6782,N_6747);
and U6947 (N_6947,N_6728,N_6776);
nand U6948 (N_6948,N_6651,N_6743);
nor U6949 (N_6949,N_6754,N_6646);
and U6950 (N_6950,N_6728,N_6733);
or U6951 (N_6951,N_6754,N_6618);
nand U6952 (N_6952,N_6692,N_6787);
nand U6953 (N_6953,N_6607,N_6787);
xor U6954 (N_6954,N_6731,N_6668);
or U6955 (N_6955,N_6745,N_6665);
nand U6956 (N_6956,N_6799,N_6675);
nor U6957 (N_6957,N_6714,N_6791);
xor U6958 (N_6958,N_6644,N_6705);
and U6959 (N_6959,N_6679,N_6666);
nor U6960 (N_6960,N_6698,N_6626);
xor U6961 (N_6961,N_6643,N_6678);
nor U6962 (N_6962,N_6795,N_6757);
and U6963 (N_6963,N_6668,N_6699);
xnor U6964 (N_6964,N_6717,N_6726);
or U6965 (N_6965,N_6607,N_6608);
or U6966 (N_6966,N_6798,N_6604);
and U6967 (N_6967,N_6612,N_6643);
and U6968 (N_6968,N_6662,N_6753);
or U6969 (N_6969,N_6761,N_6662);
nand U6970 (N_6970,N_6757,N_6745);
xor U6971 (N_6971,N_6752,N_6610);
xnor U6972 (N_6972,N_6767,N_6658);
nor U6973 (N_6973,N_6667,N_6790);
and U6974 (N_6974,N_6773,N_6745);
or U6975 (N_6975,N_6700,N_6689);
nand U6976 (N_6976,N_6688,N_6706);
and U6977 (N_6977,N_6616,N_6660);
or U6978 (N_6978,N_6649,N_6666);
and U6979 (N_6979,N_6773,N_6797);
nor U6980 (N_6980,N_6706,N_6691);
or U6981 (N_6981,N_6663,N_6625);
xnor U6982 (N_6982,N_6724,N_6699);
and U6983 (N_6983,N_6682,N_6725);
xor U6984 (N_6984,N_6690,N_6653);
nor U6985 (N_6985,N_6703,N_6698);
nand U6986 (N_6986,N_6726,N_6729);
nor U6987 (N_6987,N_6730,N_6659);
xnor U6988 (N_6988,N_6764,N_6658);
nand U6989 (N_6989,N_6749,N_6778);
xnor U6990 (N_6990,N_6702,N_6727);
and U6991 (N_6991,N_6755,N_6667);
nand U6992 (N_6992,N_6687,N_6766);
and U6993 (N_6993,N_6767,N_6703);
xor U6994 (N_6994,N_6710,N_6608);
xor U6995 (N_6995,N_6618,N_6682);
xnor U6996 (N_6996,N_6782,N_6718);
xnor U6997 (N_6997,N_6643,N_6628);
or U6998 (N_6998,N_6713,N_6731);
and U6999 (N_6999,N_6736,N_6745);
or U7000 (N_7000,N_6963,N_6978);
xnor U7001 (N_7001,N_6883,N_6938);
nand U7002 (N_7002,N_6936,N_6828);
nor U7003 (N_7003,N_6994,N_6998);
or U7004 (N_7004,N_6966,N_6809);
nor U7005 (N_7005,N_6988,N_6950);
nand U7006 (N_7006,N_6992,N_6852);
xnor U7007 (N_7007,N_6801,N_6807);
or U7008 (N_7008,N_6908,N_6831);
nor U7009 (N_7009,N_6848,N_6878);
and U7010 (N_7010,N_6941,N_6960);
nor U7011 (N_7011,N_6884,N_6811);
xor U7012 (N_7012,N_6979,N_6923);
or U7013 (N_7013,N_6949,N_6971);
xor U7014 (N_7014,N_6913,N_6866);
or U7015 (N_7015,N_6974,N_6862);
and U7016 (N_7016,N_6850,N_6969);
or U7017 (N_7017,N_6934,N_6871);
nor U7018 (N_7018,N_6898,N_6910);
nor U7019 (N_7019,N_6912,N_6944);
xor U7020 (N_7020,N_6815,N_6926);
nand U7021 (N_7021,N_6854,N_6967);
nor U7022 (N_7022,N_6847,N_6834);
nand U7023 (N_7023,N_6805,N_6835);
or U7024 (N_7024,N_6858,N_6890);
nand U7025 (N_7025,N_6980,N_6970);
and U7026 (N_7026,N_6906,N_6867);
nand U7027 (N_7027,N_6822,N_6911);
and U7028 (N_7028,N_6940,N_6957);
xor U7029 (N_7029,N_6881,N_6958);
nand U7030 (N_7030,N_6841,N_6899);
nor U7031 (N_7031,N_6845,N_6943);
nor U7032 (N_7032,N_6997,N_6996);
nor U7033 (N_7033,N_6985,N_6942);
nand U7034 (N_7034,N_6977,N_6932);
or U7035 (N_7035,N_6951,N_6909);
or U7036 (N_7036,N_6916,N_6843);
xnor U7037 (N_7037,N_6856,N_6863);
xor U7038 (N_7038,N_6816,N_6893);
nand U7039 (N_7039,N_6823,N_6917);
xnor U7040 (N_7040,N_6982,N_6990);
xor U7041 (N_7041,N_6861,N_6902);
or U7042 (N_7042,N_6879,N_6891);
nand U7043 (N_7043,N_6993,N_6933);
or U7044 (N_7044,N_6973,N_6839);
and U7045 (N_7045,N_6922,N_6824);
and U7046 (N_7046,N_6952,N_6872);
or U7047 (N_7047,N_6851,N_6897);
and U7048 (N_7048,N_6842,N_6888);
nor U7049 (N_7049,N_6868,N_6864);
or U7050 (N_7050,N_6929,N_6935);
xnor U7051 (N_7051,N_6976,N_6875);
xor U7052 (N_7052,N_6876,N_6959);
xor U7053 (N_7053,N_6921,N_6900);
nand U7054 (N_7054,N_6968,N_6873);
xnor U7055 (N_7055,N_6999,N_6955);
xnor U7056 (N_7056,N_6972,N_6846);
nor U7057 (N_7057,N_6844,N_6887);
nand U7058 (N_7058,N_6826,N_6810);
and U7059 (N_7059,N_6849,N_6914);
nand U7060 (N_7060,N_6825,N_6987);
nand U7061 (N_7061,N_6857,N_6855);
nor U7062 (N_7062,N_6975,N_6814);
xnor U7063 (N_7063,N_6837,N_6803);
or U7064 (N_7064,N_6925,N_6865);
xnor U7065 (N_7065,N_6838,N_6802);
xor U7066 (N_7066,N_6896,N_6986);
nand U7067 (N_7067,N_6927,N_6808);
and U7068 (N_7068,N_6915,N_6924);
xor U7069 (N_7069,N_6829,N_6953);
nand U7070 (N_7070,N_6836,N_6947);
nor U7071 (N_7071,N_6946,N_6859);
nand U7072 (N_7072,N_6901,N_6882);
nand U7073 (N_7073,N_6903,N_6930);
and U7074 (N_7074,N_6919,N_6833);
or U7075 (N_7075,N_6821,N_6869);
and U7076 (N_7076,N_6870,N_6981);
xor U7077 (N_7077,N_6813,N_6892);
and U7078 (N_7078,N_6956,N_6948);
or U7079 (N_7079,N_6918,N_6937);
xor U7080 (N_7080,N_6830,N_6961);
nor U7081 (N_7081,N_6832,N_6800);
or U7082 (N_7082,N_6954,N_6989);
and U7083 (N_7083,N_6984,N_6818);
and U7084 (N_7084,N_6886,N_6991);
or U7085 (N_7085,N_6804,N_6874);
nand U7086 (N_7086,N_6905,N_6840);
nor U7087 (N_7087,N_6920,N_6820);
nor U7088 (N_7088,N_6928,N_6962);
and U7089 (N_7089,N_6894,N_6827);
nand U7090 (N_7090,N_6895,N_6860);
nand U7091 (N_7091,N_6995,N_6812);
or U7092 (N_7092,N_6939,N_6945);
nand U7093 (N_7093,N_6817,N_6885);
xnor U7094 (N_7094,N_6880,N_6877);
nor U7095 (N_7095,N_6931,N_6819);
nand U7096 (N_7096,N_6964,N_6889);
or U7097 (N_7097,N_6983,N_6965);
xnor U7098 (N_7098,N_6904,N_6853);
and U7099 (N_7099,N_6806,N_6907);
and U7100 (N_7100,N_6840,N_6950);
and U7101 (N_7101,N_6874,N_6986);
or U7102 (N_7102,N_6928,N_6889);
and U7103 (N_7103,N_6927,N_6815);
and U7104 (N_7104,N_6855,N_6868);
or U7105 (N_7105,N_6980,N_6951);
nand U7106 (N_7106,N_6831,N_6987);
xnor U7107 (N_7107,N_6920,N_6823);
nand U7108 (N_7108,N_6816,N_6920);
and U7109 (N_7109,N_6972,N_6808);
or U7110 (N_7110,N_6920,N_6849);
nand U7111 (N_7111,N_6837,N_6809);
or U7112 (N_7112,N_6884,N_6852);
nor U7113 (N_7113,N_6986,N_6869);
and U7114 (N_7114,N_6824,N_6916);
xnor U7115 (N_7115,N_6966,N_6870);
and U7116 (N_7116,N_6812,N_6898);
nand U7117 (N_7117,N_6943,N_6834);
or U7118 (N_7118,N_6806,N_6950);
nand U7119 (N_7119,N_6963,N_6936);
xor U7120 (N_7120,N_6913,N_6821);
nand U7121 (N_7121,N_6949,N_6939);
nand U7122 (N_7122,N_6837,N_6976);
xnor U7123 (N_7123,N_6853,N_6872);
xor U7124 (N_7124,N_6956,N_6813);
nand U7125 (N_7125,N_6934,N_6915);
and U7126 (N_7126,N_6907,N_6811);
nand U7127 (N_7127,N_6853,N_6876);
nand U7128 (N_7128,N_6852,N_6831);
nor U7129 (N_7129,N_6838,N_6836);
xor U7130 (N_7130,N_6904,N_6869);
nor U7131 (N_7131,N_6940,N_6952);
nand U7132 (N_7132,N_6882,N_6801);
and U7133 (N_7133,N_6884,N_6878);
and U7134 (N_7134,N_6996,N_6886);
xnor U7135 (N_7135,N_6807,N_6978);
or U7136 (N_7136,N_6845,N_6985);
or U7137 (N_7137,N_6939,N_6824);
or U7138 (N_7138,N_6871,N_6848);
nor U7139 (N_7139,N_6803,N_6993);
and U7140 (N_7140,N_6849,N_6813);
nand U7141 (N_7141,N_6997,N_6970);
nand U7142 (N_7142,N_6921,N_6836);
or U7143 (N_7143,N_6930,N_6956);
nand U7144 (N_7144,N_6847,N_6931);
or U7145 (N_7145,N_6925,N_6937);
or U7146 (N_7146,N_6819,N_6994);
xnor U7147 (N_7147,N_6859,N_6854);
nor U7148 (N_7148,N_6946,N_6867);
or U7149 (N_7149,N_6995,N_6981);
xnor U7150 (N_7150,N_6968,N_6851);
and U7151 (N_7151,N_6848,N_6846);
nor U7152 (N_7152,N_6801,N_6991);
nand U7153 (N_7153,N_6981,N_6976);
xnor U7154 (N_7154,N_6990,N_6998);
and U7155 (N_7155,N_6955,N_6839);
nand U7156 (N_7156,N_6872,N_6997);
and U7157 (N_7157,N_6851,N_6827);
or U7158 (N_7158,N_6998,N_6809);
xnor U7159 (N_7159,N_6934,N_6869);
nor U7160 (N_7160,N_6817,N_6851);
xnor U7161 (N_7161,N_6868,N_6878);
or U7162 (N_7162,N_6806,N_6998);
and U7163 (N_7163,N_6947,N_6990);
or U7164 (N_7164,N_6897,N_6954);
and U7165 (N_7165,N_6969,N_6933);
or U7166 (N_7166,N_6944,N_6849);
nor U7167 (N_7167,N_6912,N_6803);
nor U7168 (N_7168,N_6863,N_6855);
nand U7169 (N_7169,N_6863,N_6908);
nand U7170 (N_7170,N_6872,N_6915);
or U7171 (N_7171,N_6854,N_6825);
nand U7172 (N_7172,N_6865,N_6864);
and U7173 (N_7173,N_6944,N_6958);
or U7174 (N_7174,N_6852,N_6903);
xnor U7175 (N_7175,N_6995,N_6828);
or U7176 (N_7176,N_6847,N_6855);
and U7177 (N_7177,N_6886,N_6849);
or U7178 (N_7178,N_6811,N_6827);
and U7179 (N_7179,N_6929,N_6808);
nor U7180 (N_7180,N_6961,N_6855);
and U7181 (N_7181,N_6961,N_6818);
and U7182 (N_7182,N_6929,N_6812);
xor U7183 (N_7183,N_6945,N_6993);
nor U7184 (N_7184,N_6972,N_6850);
or U7185 (N_7185,N_6969,N_6908);
xor U7186 (N_7186,N_6873,N_6808);
nand U7187 (N_7187,N_6863,N_6893);
nor U7188 (N_7188,N_6869,N_6876);
xnor U7189 (N_7189,N_6906,N_6915);
and U7190 (N_7190,N_6910,N_6850);
xor U7191 (N_7191,N_6958,N_6820);
xnor U7192 (N_7192,N_6969,N_6938);
nor U7193 (N_7193,N_6987,N_6864);
nand U7194 (N_7194,N_6947,N_6800);
nand U7195 (N_7195,N_6935,N_6914);
nand U7196 (N_7196,N_6802,N_6979);
and U7197 (N_7197,N_6873,N_6908);
nor U7198 (N_7198,N_6940,N_6994);
nor U7199 (N_7199,N_6918,N_6829);
xnor U7200 (N_7200,N_7168,N_7119);
nand U7201 (N_7201,N_7063,N_7005);
nor U7202 (N_7202,N_7157,N_7175);
and U7203 (N_7203,N_7142,N_7122);
nor U7204 (N_7204,N_7037,N_7174);
nand U7205 (N_7205,N_7112,N_7128);
xor U7206 (N_7206,N_7177,N_7064);
nor U7207 (N_7207,N_7066,N_7199);
xor U7208 (N_7208,N_7072,N_7051);
or U7209 (N_7209,N_7137,N_7023);
and U7210 (N_7210,N_7116,N_7166);
nand U7211 (N_7211,N_7082,N_7036);
nor U7212 (N_7212,N_7086,N_7053);
nand U7213 (N_7213,N_7096,N_7004);
nand U7214 (N_7214,N_7045,N_7031);
or U7215 (N_7215,N_7007,N_7078);
nand U7216 (N_7216,N_7021,N_7011);
xnor U7217 (N_7217,N_7077,N_7092);
or U7218 (N_7218,N_7149,N_7041);
and U7219 (N_7219,N_7093,N_7145);
or U7220 (N_7220,N_7020,N_7016);
xnor U7221 (N_7221,N_7181,N_7131);
or U7222 (N_7222,N_7187,N_7067);
or U7223 (N_7223,N_7167,N_7173);
nand U7224 (N_7224,N_7030,N_7069);
or U7225 (N_7225,N_7024,N_7022);
nand U7226 (N_7226,N_7099,N_7121);
nor U7227 (N_7227,N_7110,N_7098);
nand U7228 (N_7228,N_7114,N_7068);
and U7229 (N_7229,N_7097,N_7115);
or U7230 (N_7230,N_7192,N_7136);
or U7231 (N_7231,N_7188,N_7140);
or U7232 (N_7232,N_7026,N_7184);
nor U7233 (N_7233,N_7125,N_7002);
xor U7234 (N_7234,N_7159,N_7001);
xor U7235 (N_7235,N_7034,N_7139);
xnor U7236 (N_7236,N_7176,N_7084);
xor U7237 (N_7237,N_7025,N_7038);
and U7238 (N_7238,N_7183,N_7010);
nor U7239 (N_7239,N_7169,N_7126);
nand U7240 (N_7240,N_7057,N_7150);
xor U7241 (N_7241,N_7155,N_7158);
nor U7242 (N_7242,N_7132,N_7154);
nand U7243 (N_7243,N_7029,N_7056);
nor U7244 (N_7244,N_7135,N_7180);
nand U7245 (N_7245,N_7087,N_7091);
nand U7246 (N_7246,N_7081,N_7039);
or U7247 (N_7247,N_7108,N_7151);
nor U7248 (N_7248,N_7111,N_7117);
nand U7249 (N_7249,N_7042,N_7171);
or U7250 (N_7250,N_7165,N_7172);
nand U7251 (N_7251,N_7133,N_7073);
nand U7252 (N_7252,N_7054,N_7161);
and U7253 (N_7253,N_7058,N_7185);
nor U7254 (N_7254,N_7196,N_7090);
or U7255 (N_7255,N_7198,N_7040);
nor U7256 (N_7256,N_7074,N_7178);
nand U7257 (N_7257,N_7003,N_7044);
or U7258 (N_7258,N_7160,N_7052);
nor U7259 (N_7259,N_7000,N_7018);
or U7260 (N_7260,N_7153,N_7028);
or U7261 (N_7261,N_7075,N_7027);
nor U7262 (N_7262,N_7047,N_7013);
or U7263 (N_7263,N_7144,N_7106);
and U7264 (N_7264,N_7130,N_7162);
and U7265 (N_7265,N_7102,N_7186);
nor U7266 (N_7266,N_7197,N_7035);
or U7267 (N_7267,N_7109,N_7046);
xnor U7268 (N_7268,N_7061,N_7118);
and U7269 (N_7269,N_7089,N_7182);
xor U7270 (N_7270,N_7017,N_7095);
nor U7271 (N_7271,N_7146,N_7138);
xnor U7272 (N_7272,N_7164,N_7148);
nand U7273 (N_7273,N_7195,N_7123);
nor U7274 (N_7274,N_7059,N_7170);
nor U7275 (N_7275,N_7062,N_7085);
or U7276 (N_7276,N_7152,N_7179);
nand U7277 (N_7277,N_7088,N_7033);
xnor U7278 (N_7278,N_7083,N_7079);
nor U7279 (N_7279,N_7107,N_7009);
and U7280 (N_7280,N_7141,N_7124);
or U7281 (N_7281,N_7050,N_7094);
or U7282 (N_7282,N_7076,N_7019);
and U7283 (N_7283,N_7015,N_7101);
nand U7284 (N_7284,N_7127,N_7048);
and U7285 (N_7285,N_7100,N_7194);
nand U7286 (N_7286,N_7113,N_7032);
nand U7287 (N_7287,N_7134,N_7190);
nor U7288 (N_7288,N_7156,N_7012);
nand U7289 (N_7289,N_7070,N_7080);
nor U7290 (N_7290,N_7014,N_7065);
nand U7291 (N_7291,N_7163,N_7071);
or U7292 (N_7292,N_7055,N_7189);
nor U7293 (N_7293,N_7143,N_7103);
or U7294 (N_7294,N_7060,N_7049);
nor U7295 (N_7295,N_7193,N_7129);
nand U7296 (N_7296,N_7043,N_7008);
xnor U7297 (N_7297,N_7006,N_7120);
nand U7298 (N_7298,N_7105,N_7104);
nor U7299 (N_7299,N_7191,N_7147);
and U7300 (N_7300,N_7001,N_7154);
nor U7301 (N_7301,N_7022,N_7000);
and U7302 (N_7302,N_7031,N_7163);
and U7303 (N_7303,N_7049,N_7179);
xor U7304 (N_7304,N_7062,N_7023);
and U7305 (N_7305,N_7032,N_7098);
and U7306 (N_7306,N_7092,N_7142);
and U7307 (N_7307,N_7136,N_7000);
or U7308 (N_7308,N_7131,N_7012);
or U7309 (N_7309,N_7158,N_7092);
or U7310 (N_7310,N_7047,N_7073);
nand U7311 (N_7311,N_7105,N_7121);
and U7312 (N_7312,N_7019,N_7173);
nand U7313 (N_7313,N_7195,N_7104);
xnor U7314 (N_7314,N_7085,N_7001);
xor U7315 (N_7315,N_7110,N_7051);
or U7316 (N_7316,N_7041,N_7133);
nand U7317 (N_7317,N_7043,N_7190);
and U7318 (N_7318,N_7118,N_7077);
xnor U7319 (N_7319,N_7079,N_7142);
nor U7320 (N_7320,N_7197,N_7136);
nand U7321 (N_7321,N_7176,N_7086);
nor U7322 (N_7322,N_7069,N_7147);
nand U7323 (N_7323,N_7144,N_7140);
or U7324 (N_7324,N_7145,N_7166);
nor U7325 (N_7325,N_7088,N_7133);
or U7326 (N_7326,N_7022,N_7088);
xnor U7327 (N_7327,N_7074,N_7106);
nor U7328 (N_7328,N_7074,N_7198);
and U7329 (N_7329,N_7106,N_7035);
or U7330 (N_7330,N_7127,N_7178);
nand U7331 (N_7331,N_7103,N_7028);
xnor U7332 (N_7332,N_7123,N_7117);
nand U7333 (N_7333,N_7121,N_7170);
nand U7334 (N_7334,N_7005,N_7190);
nor U7335 (N_7335,N_7035,N_7145);
and U7336 (N_7336,N_7162,N_7108);
xnor U7337 (N_7337,N_7190,N_7035);
nor U7338 (N_7338,N_7029,N_7182);
nand U7339 (N_7339,N_7194,N_7011);
xor U7340 (N_7340,N_7190,N_7072);
nor U7341 (N_7341,N_7178,N_7175);
nor U7342 (N_7342,N_7013,N_7129);
or U7343 (N_7343,N_7117,N_7023);
nor U7344 (N_7344,N_7025,N_7071);
nand U7345 (N_7345,N_7042,N_7067);
xnor U7346 (N_7346,N_7180,N_7079);
nor U7347 (N_7347,N_7038,N_7032);
or U7348 (N_7348,N_7170,N_7197);
or U7349 (N_7349,N_7067,N_7146);
nand U7350 (N_7350,N_7068,N_7076);
nand U7351 (N_7351,N_7198,N_7137);
and U7352 (N_7352,N_7199,N_7133);
xor U7353 (N_7353,N_7005,N_7060);
xnor U7354 (N_7354,N_7107,N_7001);
xnor U7355 (N_7355,N_7008,N_7007);
nor U7356 (N_7356,N_7030,N_7019);
nor U7357 (N_7357,N_7034,N_7156);
nor U7358 (N_7358,N_7161,N_7078);
nand U7359 (N_7359,N_7171,N_7081);
xnor U7360 (N_7360,N_7170,N_7153);
xor U7361 (N_7361,N_7062,N_7199);
or U7362 (N_7362,N_7188,N_7172);
xnor U7363 (N_7363,N_7094,N_7161);
and U7364 (N_7364,N_7058,N_7189);
or U7365 (N_7365,N_7002,N_7059);
nor U7366 (N_7366,N_7145,N_7045);
or U7367 (N_7367,N_7161,N_7061);
xor U7368 (N_7368,N_7084,N_7098);
and U7369 (N_7369,N_7140,N_7104);
or U7370 (N_7370,N_7014,N_7172);
xnor U7371 (N_7371,N_7166,N_7164);
nand U7372 (N_7372,N_7049,N_7126);
and U7373 (N_7373,N_7171,N_7190);
nor U7374 (N_7374,N_7174,N_7107);
and U7375 (N_7375,N_7141,N_7179);
nand U7376 (N_7376,N_7011,N_7085);
nor U7377 (N_7377,N_7114,N_7121);
nand U7378 (N_7378,N_7159,N_7179);
or U7379 (N_7379,N_7057,N_7198);
xor U7380 (N_7380,N_7187,N_7026);
or U7381 (N_7381,N_7156,N_7084);
nor U7382 (N_7382,N_7062,N_7079);
xor U7383 (N_7383,N_7025,N_7181);
and U7384 (N_7384,N_7143,N_7159);
and U7385 (N_7385,N_7127,N_7037);
xnor U7386 (N_7386,N_7080,N_7035);
xnor U7387 (N_7387,N_7060,N_7051);
nand U7388 (N_7388,N_7171,N_7131);
xor U7389 (N_7389,N_7037,N_7125);
nor U7390 (N_7390,N_7127,N_7049);
nor U7391 (N_7391,N_7184,N_7162);
xnor U7392 (N_7392,N_7024,N_7107);
and U7393 (N_7393,N_7048,N_7045);
xor U7394 (N_7394,N_7169,N_7196);
nor U7395 (N_7395,N_7022,N_7104);
nor U7396 (N_7396,N_7118,N_7124);
or U7397 (N_7397,N_7165,N_7108);
nand U7398 (N_7398,N_7000,N_7042);
or U7399 (N_7399,N_7049,N_7029);
xnor U7400 (N_7400,N_7244,N_7341);
nor U7401 (N_7401,N_7246,N_7370);
nor U7402 (N_7402,N_7282,N_7249);
nand U7403 (N_7403,N_7360,N_7220);
xor U7404 (N_7404,N_7335,N_7237);
xnor U7405 (N_7405,N_7343,N_7269);
or U7406 (N_7406,N_7375,N_7298);
xnor U7407 (N_7407,N_7262,N_7297);
nand U7408 (N_7408,N_7231,N_7272);
or U7409 (N_7409,N_7353,N_7386);
nand U7410 (N_7410,N_7257,N_7385);
nor U7411 (N_7411,N_7234,N_7252);
xnor U7412 (N_7412,N_7296,N_7273);
or U7413 (N_7413,N_7278,N_7317);
nor U7414 (N_7414,N_7392,N_7293);
and U7415 (N_7415,N_7329,N_7376);
and U7416 (N_7416,N_7202,N_7387);
or U7417 (N_7417,N_7280,N_7215);
and U7418 (N_7418,N_7213,N_7345);
nor U7419 (N_7419,N_7359,N_7292);
and U7420 (N_7420,N_7340,N_7286);
and U7421 (N_7421,N_7396,N_7330);
xor U7422 (N_7422,N_7325,N_7238);
nand U7423 (N_7423,N_7263,N_7253);
xnor U7424 (N_7424,N_7354,N_7367);
or U7425 (N_7425,N_7362,N_7261);
nand U7426 (N_7426,N_7274,N_7245);
and U7427 (N_7427,N_7356,N_7208);
xnor U7428 (N_7428,N_7332,N_7346);
and U7429 (N_7429,N_7328,N_7352);
nand U7430 (N_7430,N_7259,N_7247);
nor U7431 (N_7431,N_7344,N_7336);
xor U7432 (N_7432,N_7368,N_7290);
and U7433 (N_7433,N_7326,N_7222);
nand U7434 (N_7434,N_7209,N_7369);
xnor U7435 (N_7435,N_7337,N_7397);
or U7436 (N_7436,N_7279,N_7363);
and U7437 (N_7437,N_7393,N_7289);
nand U7438 (N_7438,N_7384,N_7364);
xnor U7439 (N_7439,N_7226,N_7255);
nor U7440 (N_7440,N_7240,N_7235);
or U7441 (N_7441,N_7260,N_7207);
nor U7442 (N_7442,N_7324,N_7301);
and U7443 (N_7443,N_7258,N_7294);
nand U7444 (N_7444,N_7312,N_7378);
nand U7445 (N_7445,N_7311,N_7270);
nor U7446 (N_7446,N_7204,N_7358);
xor U7447 (N_7447,N_7266,N_7327);
nor U7448 (N_7448,N_7214,N_7374);
or U7449 (N_7449,N_7239,N_7265);
nor U7450 (N_7450,N_7224,N_7276);
and U7451 (N_7451,N_7373,N_7366);
nand U7452 (N_7452,N_7212,N_7306);
or U7453 (N_7453,N_7355,N_7281);
or U7454 (N_7454,N_7395,N_7251);
or U7455 (N_7455,N_7284,N_7242);
xor U7456 (N_7456,N_7236,N_7219);
nor U7457 (N_7457,N_7203,N_7267);
xor U7458 (N_7458,N_7342,N_7241);
nor U7459 (N_7459,N_7377,N_7394);
nor U7460 (N_7460,N_7268,N_7216);
or U7461 (N_7461,N_7264,N_7308);
or U7462 (N_7462,N_7254,N_7210);
xnor U7463 (N_7463,N_7200,N_7232);
xnor U7464 (N_7464,N_7307,N_7229);
xnor U7465 (N_7465,N_7304,N_7217);
xnor U7466 (N_7466,N_7361,N_7365);
nand U7467 (N_7467,N_7382,N_7250);
xor U7468 (N_7468,N_7201,N_7357);
or U7469 (N_7469,N_7338,N_7379);
or U7470 (N_7470,N_7228,N_7218);
xnor U7471 (N_7471,N_7390,N_7313);
and U7472 (N_7472,N_7322,N_7287);
nand U7473 (N_7473,N_7399,N_7320);
and U7474 (N_7474,N_7333,N_7302);
xnor U7475 (N_7475,N_7248,N_7211);
xnor U7476 (N_7476,N_7380,N_7398);
and U7477 (N_7477,N_7275,N_7319);
and U7478 (N_7478,N_7303,N_7314);
nor U7479 (N_7479,N_7389,N_7309);
and U7480 (N_7480,N_7300,N_7388);
nand U7481 (N_7481,N_7233,N_7295);
and U7482 (N_7482,N_7288,N_7323);
nor U7483 (N_7483,N_7383,N_7347);
or U7484 (N_7484,N_7277,N_7283);
or U7485 (N_7485,N_7256,N_7305);
and U7486 (N_7486,N_7243,N_7371);
and U7487 (N_7487,N_7372,N_7227);
xnor U7488 (N_7488,N_7315,N_7316);
nor U7489 (N_7489,N_7221,N_7349);
xor U7490 (N_7490,N_7351,N_7350);
and U7491 (N_7491,N_7205,N_7318);
or U7492 (N_7492,N_7391,N_7321);
or U7493 (N_7493,N_7271,N_7334);
and U7494 (N_7494,N_7223,N_7291);
nand U7495 (N_7495,N_7225,N_7339);
xor U7496 (N_7496,N_7299,N_7310);
nor U7497 (N_7497,N_7331,N_7230);
nor U7498 (N_7498,N_7285,N_7381);
nor U7499 (N_7499,N_7206,N_7348);
nand U7500 (N_7500,N_7232,N_7227);
xnor U7501 (N_7501,N_7323,N_7236);
and U7502 (N_7502,N_7395,N_7261);
nor U7503 (N_7503,N_7209,N_7218);
nand U7504 (N_7504,N_7311,N_7361);
and U7505 (N_7505,N_7369,N_7273);
and U7506 (N_7506,N_7310,N_7354);
nor U7507 (N_7507,N_7387,N_7381);
xor U7508 (N_7508,N_7304,N_7242);
or U7509 (N_7509,N_7311,N_7343);
xnor U7510 (N_7510,N_7308,N_7224);
nor U7511 (N_7511,N_7281,N_7298);
or U7512 (N_7512,N_7391,N_7315);
xor U7513 (N_7513,N_7241,N_7316);
or U7514 (N_7514,N_7207,N_7213);
nor U7515 (N_7515,N_7343,N_7339);
xor U7516 (N_7516,N_7328,N_7216);
nand U7517 (N_7517,N_7341,N_7368);
xnor U7518 (N_7518,N_7366,N_7305);
nand U7519 (N_7519,N_7343,N_7321);
nor U7520 (N_7520,N_7356,N_7322);
and U7521 (N_7521,N_7330,N_7399);
and U7522 (N_7522,N_7354,N_7323);
nor U7523 (N_7523,N_7265,N_7340);
xor U7524 (N_7524,N_7212,N_7201);
nor U7525 (N_7525,N_7393,N_7257);
and U7526 (N_7526,N_7366,N_7206);
and U7527 (N_7527,N_7294,N_7399);
nor U7528 (N_7528,N_7221,N_7388);
or U7529 (N_7529,N_7240,N_7227);
nor U7530 (N_7530,N_7243,N_7211);
xnor U7531 (N_7531,N_7243,N_7389);
or U7532 (N_7532,N_7251,N_7312);
nand U7533 (N_7533,N_7307,N_7396);
nand U7534 (N_7534,N_7202,N_7239);
and U7535 (N_7535,N_7278,N_7202);
or U7536 (N_7536,N_7292,N_7261);
and U7537 (N_7537,N_7353,N_7381);
or U7538 (N_7538,N_7372,N_7255);
and U7539 (N_7539,N_7371,N_7280);
nor U7540 (N_7540,N_7221,N_7322);
xor U7541 (N_7541,N_7399,N_7264);
and U7542 (N_7542,N_7334,N_7353);
nand U7543 (N_7543,N_7265,N_7367);
nor U7544 (N_7544,N_7223,N_7320);
nor U7545 (N_7545,N_7364,N_7378);
nand U7546 (N_7546,N_7307,N_7298);
nand U7547 (N_7547,N_7245,N_7394);
or U7548 (N_7548,N_7342,N_7323);
or U7549 (N_7549,N_7352,N_7309);
xnor U7550 (N_7550,N_7311,N_7367);
nor U7551 (N_7551,N_7342,N_7207);
or U7552 (N_7552,N_7291,N_7230);
nor U7553 (N_7553,N_7227,N_7388);
nand U7554 (N_7554,N_7315,N_7205);
nor U7555 (N_7555,N_7209,N_7339);
nand U7556 (N_7556,N_7374,N_7364);
or U7557 (N_7557,N_7353,N_7233);
nand U7558 (N_7558,N_7207,N_7340);
nor U7559 (N_7559,N_7317,N_7215);
or U7560 (N_7560,N_7314,N_7321);
or U7561 (N_7561,N_7201,N_7276);
or U7562 (N_7562,N_7212,N_7206);
or U7563 (N_7563,N_7365,N_7252);
nand U7564 (N_7564,N_7234,N_7390);
or U7565 (N_7565,N_7361,N_7310);
or U7566 (N_7566,N_7298,N_7268);
and U7567 (N_7567,N_7287,N_7344);
nor U7568 (N_7568,N_7223,N_7290);
and U7569 (N_7569,N_7306,N_7372);
or U7570 (N_7570,N_7352,N_7224);
and U7571 (N_7571,N_7367,N_7270);
and U7572 (N_7572,N_7393,N_7367);
nand U7573 (N_7573,N_7278,N_7214);
or U7574 (N_7574,N_7378,N_7282);
nor U7575 (N_7575,N_7256,N_7226);
or U7576 (N_7576,N_7264,N_7202);
nor U7577 (N_7577,N_7387,N_7362);
and U7578 (N_7578,N_7273,N_7269);
and U7579 (N_7579,N_7323,N_7345);
nor U7580 (N_7580,N_7328,N_7214);
or U7581 (N_7581,N_7365,N_7380);
xnor U7582 (N_7582,N_7355,N_7325);
xnor U7583 (N_7583,N_7354,N_7307);
nand U7584 (N_7584,N_7244,N_7268);
nand U7585 (N_7585,N_7306,N_7282);
nand U7586 (N_7586,N_7380,N_7314);
xor U7587 (N_7587,N_7372,N_7245);
and U7588 (N_7588,N_7274,N_7344);
and U7589 (N_7589,N_7286,N_7343);
nor U7590 (N_7590,N_7242,N_7219);
and U7591 (N_7591,N_7337,N_7356);
nand U7592 (N_7592,N_7284,N_7295);
or U7593 (N_7593,N_7267,N_7338);
nor U7594 (N_7594,N_7247,N_7393);
nor U7595 (N_7595,N_7283,N_7201);
and U7596 (N_7596,N_7282,N_7338);
nand U7597 (N_7597,N_7386,N_7210);
xnor U7598 (N_7598,N_7351,N_7311);
xnor U7599 (N_7599,N_7241,N_7218);
and U7600 (N_7600,N_7538,N_7509);
nand U7601 (N_7601,N_7476,N_7492);
nor U7602 (N_7602,N_7424,N_7419);
and U7603 (N_7603,N_7462,N_7529);
or U7604 (N_7604,N_7409,N_7523);
or U7605 (N_7605,N_7455,N_7483);
nor U7606 (N_7606,N_7494,N_7472);
nand U7607 (N_7607,N_7543,N_7408);
and U7608 (N_7608,N_7520,N_7429);
nand U7609 (N_7609,N_7593,N_7477);
nor U7610 (N_7610,N_7418,N_7478);
xnor U7611 (N_7611,N_7482,N_7566);
or U7612 (N_7612,N_7526,N_7510);
nand U7613 (N_7613,N_7578,N_7568);
xor U7614 (N_7614,N_7470,N_7406);
nand U7615 (N_7615,N_7515,N_7596);
or U7616 (N_7616,N_7546,N_7505);
and U7617 (N_7617,N_7503,N_7489);
and U7618 (N_7618,N_7496,N_7504);
and U7619 (N_7619,N_7458,N_7541);
or U7620 (N_7620,N_7443,N_7420);
or U7621 (N_7621,N_7464,N_7536);
nor U7622 (N_7622,N_7448,N_7539);
nor U7623 (N_7623,N_7513,N_7552);
or U7624 (N_7624,N_7548,N_7444);
or U7625 (N_7625,N_7577,N_7435);
xor U7626 (N_7626,N_7485,N_7498);
xor U7627 (N_7627,N_7574,N_7423);
or U7628 (N_7628,N_7595,N_7414);
nand U7629 (N_7629,N_7450,N_7521);
nand U7630 (N_7630,N_7572,N_7565);
nand U7631 (N_7631,N_7562,N_7517);
xor U7632 (N_7632,N_7570,N_7403);
nor U7633 (N_7633,N_7469,N_7530);
nor U7634 (N_7634,N_7533,N_7580);
nand U7635 (N_7635,N_7459,N_7584);
and U7636 (N_7636,N_7416,N_7586);
and U7637 (N_7637,N_7597,N_7415);
or U7638 (N_7638,N_7557,N_7466);
or U7639 (N_7639,N_7575,N_7528);
or U7640 (N_7640,N_7480,N_7491);
or U7641 (N_7641,N_7481,N_7413);
xor U7642 (N_7642,N_7412,N_7490);
and U7643 (N_7643,N_7454,N_7511);
xor U7644 (N_7644,N_7583,N_7425);
or U7645 (N_7645,N_7589,N_7417);
nand U7646 (N_7646,N_7407,N_7440);
and U7647 (N_7647,N_7564,N_7411);
nand U7648 (N_7648,N_7551,N_7559);
or U7649 (N_7649,N_7499,N_7463);
nor U7650 (N_7650,N_7453,N_7428);
nor U7651 (N_7651,N_7585,N_7554);
or U7652 (N_7652,N_7512,N_7486);
nand U7653 (N_7653,N_7442,N_7531);
or U7654 (N_7654,N_7433,N_7502);
nand U7655 (N_7655,N_7427,N_7446);
or U7656 (N_7656,N_7426,N_7506);
xnor U7657 (N_7657,N_7560,N_7422);
nand U7658 (N_7658,N_7519,N_7587);
xor U7659 (N_7659,N_7547,N_7474);
or U7660 (N_7660,N_7465,N_7467);
nor U7661 (N_7661,N_7598,N_7550);
or U7662 (N_7662,N_7582,N_7410);
nand U7663 (N_7663,N_7556,N_7449);
nor U7664 (N_7664,N_7500,N_7569);
or U7665 (N_7665,N_7592,N_7475);
and U7666 (N_7666,N_7430,N_7437);
nor U7667 (N_7667,N_7487,N_7402);
xnor U7668 (N_7668,N_7545,N_7447);
or U7669 (N_7669,N_7588,N_7544);
xnor U7670 (N_7670,N_7540,N_7573);
xor U7671 (N_7671,N_7488,N_7431);
nand U7672 (N_7672,N_7493,N_7525);
xor U7673 (N_7673,N_7599,N_7532);
xor U7674 (N_7674,N_7535,N_7558);
nand U7675 (N_7675,N_7468,N_7452);
or U7676 (N_7676,N_7542,N_7549);
and U7677 (N_7677,N_7518,N_7555);
nor U7678 (N_7678,N_7507,N_7457);
or U7679 (N_7679,N_7527,N_7501);
xnor U7680 (N_7680,N_7400,N_7524);
xor U7681 (N_7681,N_7436,N_7553);
nor U7682 (N_7682,N_7434,N_7590);
xor U7683 (N_7683,N_7497,N_7439);
or U7684 (N_7684,N_7460,N_7441);
and U7685 (N_7685,N_7576,N_7563);
xor U7686 (N_7686,N_7451,N_7594);
or U7687 (N_7687,N_7571,N_7461);
xnor U7688 (N_7688,N_7421,N_7404);
xor U7689 (N_7689,N_7484,N_7537);
nand U7690 (N_7690,N_7432,N_7534);
or U7691 (N_7691,N_7456,N_7591);
and U7692 (N_7692,N_7438,N_7471);
nand U7693 (N_7693,N_7579,N_7581);
nor U7694 (N_7694,N_7445,N_7405);
nor U7695 (N_7695,N_7473,N_7514);
or U7696 (N_7696,N_7516,N_7561);
xnor U7697 (N_7697,N_7522,N_7567);
nor U7698 (N_7698,N_7495,N_7508);
nand U7699 (N_7699,N_7479,N_7401);
nor U7700 (N_7700,N_7413,N_7498);
nand U7701 (N_7701,N_7590,N_7473);
and U7702 (N_7702,N_7520,N_7525);
xnor U7703 (N_7703,N_7456,N_7548);
xor U7704 (N_7704,N_7429,N_7537);
or U7705 (N_7705,N_7589,N_7517);
nand U7706 (N_7706,N_7551,N_7502);
xor U7707 (N_7707,N_7539,N_7433);
and U7708 (N_7708,N_7580,N_7541);
or U7709 (N_7709,N_7463,N_7527);
or U7710 (N_7710,N_7555,N_7556);
nor U7711 (N_7711,N_7556,N_7590);
or U7712 (N_7712,N_7495,N_7444);
nor U7713 (N_7713,N_7434,N_7493);
xnor U7714 (N_7714,N_7436,N_7589);
and U7715 (N_7715,N_7591,N_7502);
and U7716 (N_7716,N_7458,N_7482);
nand U7717 (N_7717,N_7424,N_7511);
nor U7718 (N_7718,N_7598,N_7594);
nand U7719 (N_7719,N_7588,N_7594);
or U7720 (N_7720,N_7408,N_7423);
nand U7721 (N_7721,N_7488,N_7503);
nor U7722 (N_7722,N_7512,N_7449);
nor U7723 (N_7723,N_7575,N_7422);
xnor U7724 (N_7724,N_7582,N_7561);
nand U7725 (N_7725,N_7536,N_7467);
nor U7726 (N_7726,N_7525,N_7403);
nor U7727 (N_7727,N_7430,N_7495);
xor U7728 (N_7728,N_7573,N_7408);
or U7729 (N_7729,N_7509,N_7546);
nor U7730 (N_7730,N_7450,N_7476);
or U7731 (N_7731,N_7464,N_7408);
nor U7732 (N_7732,N_7519,N_7491);
nand U7733 (N_7733,N_7447,N_7411);
nor U7734 (N_7734,N_7557,N_7548);
and U7735 (N_7735,N_7413,N_7432);
and U7736 (N_7736,N_7422,N_7496);
or U7737 (N_7737,N_7522,N_7544);
nand U7738 (N_7738,N_7591,N_7495);
xor U7739 (N_7739,N_7451,N_7558);
nor U7740 (N_7740,N_7509,N_7532);
or U7741 (N_7741,N_7512,N_7405);
nor U7742 (N_7742,N_7476,N_7493);
and U7743 (N_7743,N_7403,N_7488);
or U7744 (N_7744,N_7495,N_7553);
xnor U7745 (N_7745,N_7597,N_7417);
xnor U7746 (N_7746,N_7527,N_7477);
nand U7747 (N_7747,N_7514,N_7470);
nand U7748 (N_7748,N_7515,N_7436);
and U7749 (N_7749,N_7416,N_7455);
or U7750 (N_7750,N_7511,N_7421);
or U7751 (N_7751,N_7520,N_7576);
xor U7752 (N_7752,N_7433,N_7566);
nand U7753 (N_7753,N_7563,N_7583);
nor U7754 (N_7754,N_7496,N_7476);
nand U7755 (N_7755,N_7482,N_7516);
nand U7756 (N_7756,N_7492,N_7598);
or U7757 (N_7757,N_7590,N_7568);
nor U7758 (N_7758,N_7539,N_7560);
xor U7759 (N_7759,N_7437,N_7582);
or U7760 (N_7760,N_7412,N_7502);
or U7761 (N_7761,N_7578,N_7507);
or U7762 (N_7762,N_7599,N_7556);
nor U7763 (N_7763,N_7588,N_7438);
xnor U7764 (N_7764,N_7527,N_7511);
nor U7765 (N_7765,N_7572,N_7402);
nor U7766 (N_7766,N_7559,N_7555);
and U7767 (N_7767,N_7574,N_7571);
or U7768 (N_7768,N_7415,N_7577);
and U7769 (N_7769,N_7452,N_7416);
and U7770 (N_7770,N_7583,N_7411);
xnor U7771 (N_7771,N_7485,N_7568);
xor U7772 (N_7772,N_7411,N_7403);
or U7773 (N_7773,N_7574,N_7442);
nor U7774 (N_7774,N_7577,N_7526);
nand U7775 (N_7775,N_7448,N_7599);
nor U7776 (N_7776,N_7471,N_7507);
or U7777 (N_7777,N_7596,N_7548);
and U7778 (N_7778,N_7526,N_7547);
xnor U7779 (N_7779,N_7542,N_7503);
nand U7780 (N_7780,N_7509,N_7550);
nand U7781 (N_7781,N_7539,N_7420);
xnor U7782 (N_7782,N_7598,N_7485);
or U7783 (N_7783,N_7437,N_7468);
nor U7784 (N_7784,N_7448,N_7571);
or U7785 (N_7785,N_7583,N_7541);
and U7786 (N_7786,N_7538,N_7587);
and U7787 (N_7787,N_7436,N_7426);
xor U7788 (N_7788,N_7416,N_7449);
and U7789 (N_7789,N_7447,N_7502);
nor U7790 (N_7790,N_7547,N_7592);
nor U7791 (N_7791,N_7508,N_7491);
or U7792 (N_7792,N_7458,N_7539);
nand U7793 (N_7793,N_7597,N_7517);
xnor U7794 (N_7794,N_7500,N_7528);
nor U7795 (N_7795,N_7540,N_7574);
nor U7796 (N_7796,N_7518,N_7443);
nor U7797 (N_7797,N_7497,N_7477);
nor U7798 (N_7798,N_7546,N_7545);
xor U7799 (N_7799,N_7566,N_7511);
nand U7800 (N_7800,N_7721,N_7616);
and U7801 (N_7801,N_7768,N_7731);
nand U7802 (N_7802,N_7719,N_7686);
nor U7803 (N_7803,N_7669,N_7779);
and U7804 (N_7804,N_7663,N_7683);
or U7805 (N_7805,N_7693,N_7720);
or U7806 (N_7806,N_7724,N_7734);
nor U7807 (N_7807,N_7703,N_7667);
nor U7808 (N_7808,N_7676,N_7612);
xnor U7809 (N_7809,N_7690,N_7670);
and U7810 (N_7810,N_7786,N_7778);
xnor U7811 (N_7811,N_7775,N_7636);
nand U7812 (N_7812,N_7627,N_7696);
or U7813 (N_7813,N_7726,N_7613);
xnor U7814 (N_7814,N_7649,N_7615);
nor U7815 (N_7815,N_7680,N_7708);
nor U7816 (N_7816,N_7732,N_7665);
nor U7817 (N_7817,N_7664,N_7638);
or U7818 (N_7818,N_7785,N_7748);
nor U7819 (N_7819,N_7681,N_7780);
nor U7820 (N_7820,N_7620,N_7763);
xor U7821 (N_7821,N_7647,N_7611);
or U7822 (N_7822,N_7635,N_7675);
nand U7823 (N_7823,N_7655,N_7630);
nor U7824 (N_7824,N_7758,N_7709);
xor U7825 (N_7825,N_7767,N_7757);
xor U7826 (N_7826,N_7737,N_7714);
nand U7827 (N_7827,N_7705,N_7662);
or U7828 (N_7828,N_7741,N_7783);
nand U7829 (N_7829,N_7723,N_7771);
nand U7830 (N_7830,N_7601,N_7701);
and U7831 (N_7831,N_7622,N_7752);
nand U7832 (N_7832,N_7668,N_7756);
or U7833 (N_7833,N_7776,N_7782);
nor U7834 (N_7834,N_7722,N_7672);
nor U7835 (N_7835,N_7628,N_7742);
and U7836 (N_7836,N_7717,N_7608);
xnor U7837 (N_7837,N_7699,N_7702);
xor U7838 (N_7838,N_7711,N_7759);
xor U7839 (N_7839,N_7624,N_7792);
or U7840 (N_7840,N_7684,N_7787);
xnor U7841 (N_7841,N_7682,N_7637);
or U7842 (N_7842,N_7710,N_7730);
xnor U7843 (N_7843,N_7656,N_7614);
nor U7844 (N_7844,N_7642,N_7695);
and U7845 (N_7845,N_7650,N_7789);
or U7846 (N_7846,N_7619,N_7766);
nand U7847 (N_7847,N_7679,N_7729);
nor U7848 (N_7848,N_7755,N_7761);
nor U7849 (N_7849,N_7760,N_7799);
nand U7850 (N_7850,N_7725,N_7707);
and U7851 (N_7851,N_7745,N_7653);
xor U7852 (N_7852,N_7712,N_7618);
nor U7853 (N_7853,N_7629,N_7606);
xnor U7854 (N_7854,N_7600,N_7713);
xor U7855 (N_7855,N_7654,N_7743);
and U7856 (N_7856,N_7633,N_7793);
and U7857 (N_7857,N_7605,N_7735);
nor U7858 (N_7858,N_7651,N_7698);
and U7859 (N_7859,N_7639,N_7738);
nor U7860 (N_7860,N_7749,N_7727);
nand U7861 (N_7861,N_7677,N_7604);
or U7862 (N_7862,N_7674,N_7632);
nand U7863 (N_7863,N_7643,N_7772);
nor U7864 (N_7864,N_7704,N_7798);
and U7865 (N_7865,N_7795,N_7641);
nor U7866 (N_7866,N_7607,N_7784);
xor U7867 (N_7867,N_7716,N_7689);
xnor U7868 (N_7868,N_7739,N_7791);
and U7869 (N_7869,N_7781,N_7685);
or U7870 (N_7870,N_7706,N_7631);
nand U7871 (N_7871,N_7610,N_7744);
nand U7872 (N_7872,N_7626,N_7666);
nor U7873 (N_7873,N_7697,N_7671);
or U7874 (N_7874,N_7617,N_7621);
or U7875 (N_7875,N_7652,N_7797);
nand U7876 (N_7876,N_7746,N_7774);
xor U7877 (N_7877,N_7659,N_7796);
or U7878 (N_7878,N_7753,N_7692);
and U7879 (N_7879,N_7788,N_7609);
nand U7880 (N_7880,N_7694,N_7603);
nand U7881 (N_7881,N_7661,N_7687);
and U7882 (N_7882,N_7794,N_7715);
nor U7883 (N_7883,N_7747,N_7733);
nor U7884 (N_7884,N_7648,N_7740);
xor U7885 (N_7885,N_7700,N_7736);
or U7886 (N_7886,N_7770,N_7790);
or U7887 (N_7887,N_7657,N_7602);
or U7888 (N_7888,N_7678,N_7634);
nor U7889 (N_7889,N_7762,N_7754);
xor U7890 (N_7890,N_7688,N_7773);
nand U7891 (N_7891,N_7777,N_7625);
and U7892 (N_7892,N_7644,N_7673);
xnor U7893 (N_7893,N_7691,N_7645);
or U7894 (N_7894,N_7728,N_7658);
nor U7895 (N_7895,N_7765,N_7646);
nand U7896 (N_7896,N_7764,N_7718);
and U7897 (N_7897,N_7750,N_7769);
and U7898 (N_7898,N_7623,N_7751);
xor U7899 (N_7899,N_7660,N_7640);
nor U7900 (N_7900,N_7753,N_7777);
or U7901 (N_7901,N_7699,N_7786);
or U7902 (N_7902,N_7737,N_7602);
and U7903 (N_7903,N_7635,N_7717);
or U7904 (N_7904,N_7644,N_7751);
nor U7905 (N_7905,N_7630,N_7758);
or U7906 (N_7906,N_7632,N_7633);
and U7907 (N_7907,N_7655,N_7730);
and U7908 (N_7908,N_7768,N_7737);
or U7909 (N_7909,N_7767,N_7675);
or U7910 (N_7910,N_7751,N_7678);
nor U7911 (N_7911,N_7755,N_7772);
xor U7912 (N_7912,N_7733,N_7667);
nand U7913 (N_7913,N_7704,N_7700);
and U7914 (N_7914,N_7638,N_7698);
nand U7915 (N_7915,N_7708,N_7621);
xor U7916 (N_7916,N_7786,N_7664);
or U7917 (N_7917,N_7692,N_7778);
nand U7918 (N_7918,N_7617,N_7793);
or U7919 (N_7919,N_7652,N_7790);
and U7920 (N_7920,N_7714,N_7716);
nand U7921 (N_7921,N_7725,N_7600);
xnor U7922 (N_7922,N_7661,N_7655);
nand U7923 (N_7923,N_7642,N_7722);
or U7924 (N_7924,N_7602,N_7706);
xnor U7925 (N_7925,N_7667,N_7699);
and U7926 (N_7926,N_7679,N_7711);
nand U7927 (N_7927,N_7681,N_7605);
xor U7928 (N_7928,N_7658,N_7609);
nor U7929 (N_7929,N_7704,N_7739);
or U7930 (N_7930,N_7707,N_7611);
xor U7931 (N_7931,N_7665,N_7632);
nor U7932 (N_7932,N_7697,N_7647);
xnor U7933 (N_7933,N_7709,N_7769);
nand U7934 (N_7934,N_7649,N_7618);
and U7935 (N_7935,N_7696,N_7798);
and U7936 (N_7936,N_7640,N_7625);
nand U7937 (N_7937,N_7636,N_7756);
nand U7938 (N_7938,N_7647,N_7782);
nor U7939 (N_7939,N_7705,N_7788);
nor U7940 (N_7940,N_7636,N_7712);
nand U7941 (N_7941,N_7717,N_7737);
xnor U7942 (N_7942,N_7625,N_7712);
nand U7943 (N_7943,N_7618,N_7704);
and U7944 (N_7944,N_7624,N_7681);
or U7945 (N_7945,N_7712,N_7645);
xnor U7946 (N_7946,N_7664,N_7784);
and U7947 (N_7947,N_7709,N_7687);
nand U7948 (N_7948,N_7636,N_7799);
and U7949 (N_7949,N_7766,N_7698);
nand U7950 (N_7950,N_7740,N_7614);
xnor U7951 (N_7951,N_7707,N_7739);
or U7952 (N_7952,N_7714,N_7630);
or U7953 (N_7953,N_7742,N_7677);
nand U7954 (N_7954,N_7692,N_7740);
nand U7955 (N_7955,N_7796,N_7716);
nor U7956 (N_7956,N_7613,N_7733);
xor U7957 (N_7957,N_7782,N_7797);
xor U7958 (N_7958,N_7711,N_7609);
nand U7959 (N_7959,N_7609,N_7650);
nor U7960 (N_7960,N_7676,N_7759);
nor U7961 (N_7961,N_7692,N_7762);
or U7962 (N_7962,N_7787,N_7730);
or U7963 (N_7963,N_7669,N_7772);
xnor U7964 (N_7964,N_7708,N_7702);
and U7965 (N_7965,N_7689,N_7636);
or U7966 (N_7966,N_7742,N_7720);
xor U7967 (N_7967,N_7726,N_7743);
nor U7968 (N_7968,N_7642,N_7632);
xor U7969 (N_7969,N_7766,N_7773);
and U7970 (N_7970,N_7792,N_7681);
xnor U7971 (N_7971,N_7646,N_7738);
nand U7972 (N_7972,N_7670,N_7720);
nand U7973 (N_7973,N_7690,N_7688);
or U7974 (N_7974,N_7667,N_7630);
nor U7975 (N_7975,N_7742,N_7669);
and U7976 (N_7976,N_7700,N_7620);
nor U7977 (N_7977,N_7699,N_7692);
and U7978 (N_7978,N_7788,N_7797);
xor U7979 (N_7979,N_7665,N_7794);
nand U7980 (N_7980,N_7755,N_7615);
nand U7981 (N_7981,N_7672,N_7715);
xnor U7982 (N_7982,N_7613,N_7739);
or U7983 (N_7983,N_7660,N_7734);
and U7984 (N_7984,N_7603,N_7701);
xor U7985 (N_7985,N_7649,N_7678);
nand U7986 (N_7986,N_7602,N_7736);
xnor U7987 (N_7987,N_7692,N_7644);
nand U7988 (N_7988,N_7728,N_7619);
nand U7989 (N_7989,N_7795,N_7646);
xnor U7990 (N_7990,N_7610,N_7759);
and U7991 (N_7991,N_7722,N_7680);
nand U7992 (N_7992,N_7738,N_7655);
or U7993 (N_7993,N_7771,N_7658);
xnor U7994 (N_7994,N_7651,N_7681);
xor U7995 (N_7995,N_7660,N_7678);
xnor U7996 (N_7996,N_7699,N_7643);
and U7997 (N_7997,N_7743,N_7640);
nand U7998 (N_7998,N_7621,N_7603);
and U7999 (N_7999,N_7721,N_7789);
or U8000 (N_8000,N_7803,N_7801);
xnor U8001 (N_8001,N_7939,N_7808);
and U8002 (N_8002,N_7881,N_7841);
nor U8003 (N_8003,N_7832,N_7821);
or U8004 (N_8004,N_7872,N_7870);
or U8005 (N_8005,N_7885,N_7883);
nand U8006 (N_8006,N_7969,N_7974);
or U8007 (N_8007,N_7972,N_7968);
xor U8008 (N_8008,N_7865,N_7963);
nand U8009 (N_8009,N_7927,N_7847);
nor U8010 (N_8010,N_7863,N_7912);
and U8011 (N_8011,N_7941,N_7836);
xnor U8012 (N_8012,N_7923,N_7811);
and U8013 (N_8013,N_7917,N_7947);
xor U8014 (N_8014,N_7850,N_7879);
or U8015 (N_8015,N_7860,N_7871);
and U8016 (N_8016,N_7980,N_7815);
and U8017 (N_8017,N_7843,N_7986);
and U8018 (N_8018,N_7818,N_7862);
nand U8019 (N_8019,N_7902,N_7987);
nor U8020 (N_8020,N_7844,N_7944);
nor U8021 (N_8021,N_7971,N_7924);
nand U8022 (N_8022,N_7840,N_7960);
nand U8023 (N_8023,N_7846,N_7851);
xnor U8024 (N_8024,N_7956,N_7907);
or U8025 (N_8025,N_7904,N_7874);
nand U8026 (N_8026,N_7882,N_7985);
or U8027 (N_8027,N_7900,N_7855);
nor U8028 (N_8028,N_7994,N_7989);
nand U8029 (N_8029,N_7961,N_7978);
or U8030 (N_8030,N_7937,N_7829);
and U8031 (N_8031,N_7898,N_7822);
nand U8032 (N_8032,N_7861,N_7951);
and U8033 (N_8033,N_7970,N_7906);
nor U8034 (N_8034,N_7943,N_7830);
or U8035 (N_8035,N_7887,N_7893);
nand U8036 (N_8036,N_7929,N_7858);
xor U8037 (N_8037,N_7807,N_7992);
xor U8038 (N_8038,N_7935,N_7982);
xnor U8039 (N_8039,N_7814,N_7996);
or U8040 (N_8040,N_7838,N_7945);
nor U8041 (N_8041,N_7990,N_7848);
nand U8042 (N_8042,N_7856,N_7852);
nor U8043 (N_8043,N_7998,N_7901);
nor U8044 (N_8044,N_7888,N_7827);
xor U8045 (N_8045,N_7920,N_7853);
nor U8046 (N_8046,N_7905,N_7849);
nor U8047 (N_8047,N_7934,N_7991);
and U8048 (N_8048,N_7857,N_7875);
nand U8049 (N_8049,N_7819,N_7884);
nand U8050 (N_8050,N_7938,N_7936);
nand U8051 (N_8051,N_7957,N_7926);
or U8052 (N_8052,N_7979,N_7975);
nand U8053 (N_8053,N_7826,N_7959);
nand U8054 (N_8054,N_7997,N_7949);
and U8055 (N_8055,N_7984,N_7839);
nand U8056 (N_8056,N_7981,N_7824);
xor U8057 (N_8057,N_7834,N_7877);
xnor U8058 (N_8058,N_7810,N_7812);
xor U8059 (N_8059,N_7932,N_7876);
or U8060 (N_8060,N_7955,N_7962);
and U8061 (N_8061,N_7916,N_7805);
and U8062 (N_8062,N_7933,N_7817);
nand U8063 (N_8063,N_7813,N_7897);
nand U8064 (N_8064,N_7828,N_7894);
xor U8065 (N_8065,N_7940,N_7919);
nor U8066 (N_8066,N_7892,N_7953);
nand U8067 (N_8067,N_7964,N_7895);
nor U8068 (N_8068,N_7958,N_7845);
nand U8069 (N_8069,N_7899,N_7977);
nand U8070 (N_8070,N_7995,N_7809);
nor U8071 (N_8071,N_7952,N_7820);
xnor U8072 (N_8072,N_7993,N_7983);
and U8073 (N_8073,N_7867,N_7878);
nor U8074 (N_8074,N_7825,N_7948);
nand U8075 (N_8075,N_7823,N_7869);
and U8076 (N_8076,N_7890,N_7931);
and U8077 (N_8077,N_7833,N_7908);
and U8078 (N_8078,N_7928,N_7914);
and U8079 (N_8079,N_7854,N_7816);
nand U8080 (N_8080,N_7922,N_7913);
and U8081 (N_8081,N_7889,N_7800);
and U8082 (N_8082,N_7918,N_7950);
and U8083 (N_8083,N_7954,N_7831);
xnor U8084 (N_8084,N_7967,N_7925);
or U8085 (N_8085,N_7896,N_7886);
and U8086 (N_8086,N_7930,N_7911);
nand U8087 (N_8087,N_7842,N_7880);
and U8088 (N_8088,N_7942,N_7988);
xnor U8089 (N_8089,N_7891,N_7946);
xnor U8090 (N_8090,N_7866,N_7915);
or U8091 (N_8091,N_7868,N_7837);
and U8092 (N_8092,N_7806,N_7802);
xor U8093 (N_8093,N_7804,N_7909);
or U8094 (N_8094,N_7903,N_7859);
xnor U8095 (N_8095,N_7921,N_7966);
xnor U8096 (N_8096,N_7999,N_7835);
nand U8097 (N_8097,N_7973,N_7976);
or U8098 (N_8098,N_7910,N_7864);
and U8099 (N_8099,N_7873,N_7965);
and U8100 (N_8100,N_7801,N_7975);
nor U8101 (N_8101,N_7845,N_7818);
xor U8102 (N_8102,N_7918,N_7801);
or U8103 (N_8103,N_7966,N_7836);
and U8104 (N_8104,N_7835,N_7871);
or U8105 (N_8105,N_7940,N_7822);
or U8106 (N_8106,N_7828,N_7915);
or U8107 (N_8107,N_7852,N_7828);
nand U8108 (N_8108,N_7919,N_7874);
and U8109 (N_8109,N_7915,N_7831);
nand U8110 (N_8110,N_7856,N_7959);
nand U8111 (N_8111,N_7886,N_7835);
nand U8112 (N_8112,N_7918,N_7803);
and U8113 (N_8113,N_7830,N_7809);
xor U8114 (N_8114,N_7950,N_7829);
nand U8115 (N_8115,N_7915,N_7824);
or U8116 (N_8116,N_7910,N_7862);
or U8117 (N_8117,N_7946,N_7980);
and U8118 (N_8118,N_7888,N_7894);
nand U8119 (N_8119,N_7838,N_7894);
and U8120 (N_8120,N_7988,N_7944);
xnor U8121 (N_8121,N_7888,N_7957);
and U8122 (N_8122,N_7972,N_7917);
nand U8123 (N_8123,N_7890,N_7969);
or U8124 (N_8124,N_7929,N_7869);
nand U8125 (N_8125,N_7879,N_7964);
nor U8126 (N_8126,N_7859,N_7815);
nand U8127 (N_8127,N_7927,N_7917);
or U8128 (N_8128,N_7948,N_7902);
and U8129 (N_8129,N_7911,N_7998);
or U8130 (N_8130,N_7860,N_7870);
nand U8131 (N_8131,N_7835,N_7917);
or U8132 (N_8132,N_7993,N_7823);
nand U8133 (N_8133,N_7934,N_7831);
xor U8134 (N_8134,N_7881,N_7908);
nor U8135 (N_8135,N_7989,N_7949);
nand U8136 (N_8136,N_7976,N_7915);
xnor U8137 (N_8137,N_7917,N_7961);
nand U8138 (N_8138,N_7853,N_7854);
xor U8139 (N_8139,N_7858,N_7864);
or U8140 (N_8140,N_7996,N_7961);
and U8141 (N_8141,N_7800,N_7918);
and U8142 (N_8142,N_7826,N_7840);
xor U8143 (N_8143,N_7837,N_7934);
nor U8144 (N_8144,N_7995,N_7964);
and U8145 (N_8145,N_7947,N_7808);
and U8146 (N_8146,N_7963,N_7978);
nand U8147 (N_8147,N_7950,N_7933);
or U8148 (N_8148,N_7858,N_7807);
nand U8149 (N_8149,N_7859,N_7895);
nand U8150 (N_8150,N_7821,N_7998);
nand U8151 (N_8151,N_7964,N_7914);
nor U8152 (N_8152,N_7865,N_7863);
xnor U8153 (N_8153,N_7849,N_7863);
nor U8154 (N_8154,N_7955,N_7982);
nor U8155 (N_8155,N_7880,N_7939);
nor U8156 (N_8156,N_7889,N_7996);
or U8157 (N_8157,N_7879,N_7843);
nor U8158 (N_8158,N_7921,N_7973);
nor U8159 (N_8159,N_7975,N_7871);
nand U8160 (N_8160,N_7829,N_7935);
nand U8161 (N_8161,N_7896,N_7974);
or U8162 (N_8162,N_7861,N_7979);
nor U8163 (N_8163,N_7802,N_7817);
nand U8164 (N_8164,N_7861,N_7876);
or U8165 (N_8165,N_7965,N_7859);
or U8166 (N_8166,N_7977,N_7988);
nand U8167 (N_8167,N_7809,N_7914);
nor U8168 (N_8168,N_7906,N_7905);
and U8169 (N_8169,N_7966,N_7841);
and U8170 (N_8170,N_7960,N_7824);
xor U8171 (N_8171,N_7992,N_7900);
nand U8172 (N_8172,N_7845,N_7993);
nand U8173 (N_8173,N_7995,N_7985);
or U8174 (N_8174,N_7822,N_7862);
nor U8175 (N_8175,N_7927,N_7892);
nor U8176 (N_8176,N_7884,N_7992);
and U8177 (N_8177,N_7856,N_7995);
nor U8178 (N_8178,N_7917,N_7859);
or U8179 (N_8179,N_7896,N_7951);
xnor U8180 (N_8180,N_7808,N_7972);
and U8181 (N_8181,N_7981,N_7883);
or U8182 (N_8182,N_7816,N_7972);
or U8183 (N_8183,N_7857,N_7931);
and U8184 (N_8184,N_7903,N_7959);
xor U8185 (N_8185,N_7893,N_7831);
nand U8186 (N_8186,N_7981,N_7878);
nand U8187 (N_8187,N_7872,N_7933);
or U8188 (N_8188,N_7850,N_7978);
nor U8189 (N_8189,N_7936,N_7964);
xor U8190 (N_8190,N_7863,N_7885);
nor U8191 (N_8191,N_7834,N_7843);
or U8192 (N_8192,N_7901,N_7938);
nand U8193 (N_8193,N_7967,N_7968);
xor U8194 (N_8194,N_7848,N_7865);
nor U8195 (N_8195,N_7947,N_7923);
xnor U8196 (N_8196,N_7911,N_7865);
and U8197 (N_8197,N_7853,N_7868);
and U8198 (N_8198,N_7988,N_7843);
or U8199 (N_8199,N_7804,N_7806);
nor U8200 (N_8200,N_8166,N_8107);
and U8201 (N_8201,N_8087,N_8079);
xnor U8202 (N_8202,N_8122,N_8011);
and U8203 (N_8203,N_8168,N_8161);
or U8204 (N_8204,N_8041,N_8088);
or U8205 (N_8205,N_8045,N_8024);
nand U8206 (N_8206,N_8004,N_8185);
nand U8207 (N_8207,N_8021,N_8186);
and U8208 (N_8208,N_8006,N_8182);
or U8209 (N_8209,N_8148,N_8172);
xnor U8210 (N_8210,N_8129,N_8039);
xor U8211 (N_8211,N_8135,N_8068);
and U8212 (N_8212,N_8043,N_8030);
nor U8213 (N_8213,N_8173,N_8170);
xor U8214 (N_8214,N_8109,N_8092);
and U8215 (N_8215,N_8188,N_8123);
xnor U8216 (N_8216,N_8133,N_8037);
xnor U8217 (N_8217,N_8017,N_8091);
nor U8218 (N_8218,N_8199,N_8197);
or U8219 (N_8219,N_8141,N_8143);
or U8220 (N_8220,N_8074,N_8086);
nor U8221 (N_8221,N_8049,N_8183);
or U8222 (N_8222,N_8125,N_8142);
or U8223 (N_8223,N_8187,N_8016);
nor U8224 (N_8224,N_8127,N_8175);
and U8225 (N_8225,N_8014,N_8060);
xor U8226 (N_8226,N_8189,N_8002);
xor U8227 (N_8227,N_8146,N_8077);
or U8228 (N_8228,N_8075,N_8154);
nand U8229 (N_8229,N_8155,N_8126);
nand U8230 (N_8230,N_8137,N_8191);
nor U8231 (N_8231,N_8111,N_8108);
nor U8232 (N_8232,N_8029,N_8000);
xor U8233 (N_8233,N_8059,N_8181);
nor U8234 (N_8234,N_8012,N_8157);
nand U8235 (N_8235,N_8195,N_8140);
and U8236 (N_8236,N_8034,N_8040);
nor U8237 (N_8237,N_8171,N_8053);
and U8238 (N_8238,N_8019,N_8160);
and U8239 (N_8239,N_8009,N_8136);
xor U8240 (N_8240,N_8115,N_8196);
xor U8241 (N_8241,N_8102,N_8046);
and U8242 (N_8242,N_8116,N_8094);
nand U8243 (N_8243,N_8081,N_8067);
nor U8244 (N_8244,N_8112,N_8184);
xor U8245 (N_8245,N_8089,N_8058);
xnor U8246 (N_8246,N_8177,N_8159);
xnor U8247 (N_8247,N_8051,N_8130);
nor U8248 (N_8248,N_8179,N_8152);
or U8249 (N_8249,N_8038,N_8078);
nor U8250 (N_8250,N_8194,N_8026);
nand U8251 (N_8251,N_8072,N_8042);
and U8252 (N_8252,N_8165,N_8150);
or U8253 (N_8253,N_8156,N_8153);
and U8254 (N_8254,N_8158,N_8082);
and U8255 (N_8255,N_8015,N_8064);
or U8256 (N_8256,N_8139,N_8061);
nand U8257 (N_8257,N_8062,N_8114);
nand U8258 (N_8258,N_8027,N_8076);
nor U8259 (N_8259,N_8198,N_8063);
nor U8260 (N_8260,N_8022,N_8144);
xor U8261 (N_8261,N_8044,N_8098);
xor U8262 (N_8262,N_8120,N_8138);
nand U8263 (N_8263,N_8084,N_8128);
xor U8264 (N_8264,N_8023,N_8131);
or U8265 (N_8265,N_8080,N_8162);
or U8266 (N_8266,N_8121,N_8065);
and U8267 (N_8267,N_8178,N_8100);
nor U8268 (N_8268,N_8008,N_8105);
nor U8269 (N_8269,N_8192,N_8132);
xnor U8270 (N_8270,N_8007,N_8052);
xnor U8271 (N_8271,N_8118,N_8013);
xor U8272 (N_8272,N_8124,N_8145);
nand U8273 (N_8273,N_8180,N_8025);
or U8274 (N_8274,N_8099,N_8069);
xor U8275 (N_8275,N_8003,N_8070);
nor U8276 (N_8276,N_8164,N_8193);
nand U8277 (N_8277,N_8050,N_8055);
xor U8278 (N_8278,N_8095,N_8090);
or U8279 (N_8279,N_8169,N_8151);
nor U8280 (N_8280,N_8101,N_8020);
nand U8281 (N_8281,N_8028,N_8190);
nand U8282 (N_8282,N_8047,N_8032);
xor U8283 (N_8283,N_8066,N_8071);
xor U8284 (N_8284,N_8119,N_8048);
nor U8285 (N_8285,N_8097,N_8163);
nand U8286 (N_8286,N_8134,N_8005);
or U8287 (N_8287,N_8104,N_8035);
xor U8288 (N_8288,N_8036,N_8176);
nor U8289 (N_8289,N_8018,N_8110);
xnor U8290 (N_8290,N_8054,N_8117);
and U8291 (N_8291,N_8106,N_8174);
nor U8292 (N_8292,N_8096,N_8113);
nand U8293 (N_8293,N_8010,N_8167);
xnor U8294 (N_8294,N_8083,N_8147);
nand U8295 (N_8295,N_8001,N_8056);
and U8296 (N_8296,N_8093,N_8057);
or U8297 (N_8297,N_8103,N_8149);
nand U8298 (N_8298,N_8073,N_8033);
xor U8299 (N_8299,N_8031,N_8085);
nand U8300 (N_8300,N_8095,N_8195);
or U8301 (N_8301,N_8126,N_8143);
and U8302 (N_8302,N_8035,N_8173);
nand U8303 (N_8303,N_8074,N_8150);
nand U8304 (N_8304,N_8155,N_8034);
nand U8305 (N_8305,N_8046,N_8062);
and U8306 (N_8306,N_8123,N_8018);
nand U8307 (N_8307,N_8179,N_8175);
and U8308 (N_8308,N_8158,N_8194);
xnor U8309 (N_8309,N_8150,N_8054);
and U8310 (N_8310,N_8148,N_8126);
xor U8311 (N_8311,N_8108,N_8166);
nor U8312 (N_8312,N_8147,N_8115);
nor U8313 (N_8313,N_8197,N_8072);
and U8314 (N_8314,N_8066,N_8003);
or U8315 (N_8315,N_8074,N_8165);
nor U8316 (N_8316,N_8152,N_8016);
xor U8317 (N_8317,N_8137,N_8144);
and U8318 (N_8318,N_8022,N_8183);
nand U8319 (N_8319,N_8153,N_8117);
and U8320 (N_8320,N_8173,N_8054);
and U8321 (N_8321,N_8005,N_8113);
nor U8322 (N_8322,N_8028,N_8138);
xnor U8323 (N_8323,N_8100,N_8014);
or U8324 (N_8324,N_8164,N_8015);
xor U8325 (N_8325,N_8062,N_8146);
or U8326 (N_8326,N_8006,N_8038);
nand U8327 (N_8327,N_8059,N_8032);
or U8328 (N_8328,N_8164,N_8191);
and U8329 (N_8329,N_8169,N_8115);
xnor U8330 (N_8330,N_8136,N_8095);
nand U8331 (N_8331,N_8132,N_8194);
nor U8332 (N_8332,N_8163,N_8008);
nand U8333 (N_8333,N_8076,N_8063);
and U8334 (N_8334,N_8125,N_8133);
or U8335 (N_8335,N_8172,N_8089);
and U8336 (N_8336,N_8154,N_8024);
nor U8337 (N_8337,N_8000,N_8023);
nand U8338 (N_8338,N_8034,N_8140);
nand U8339 (N_8339,N_8099,N_8046);
xor U8340 (N_8340,N_8034,N_8160);
nor U8341 (N_8341,N_8042,N_8015);
or U8342 (N_8342,N_8048,N_8136);
xor U8343 (N_8343,N_8083,N_8106);
or U8344 (N_8344,N_8126,N_8046);
nand U8345 (N_8345,N_8119,N_8179);
nor U8346 (N_8346,N_8125,N_8176);
or U8347 (N_8347,N_8182,N_8031);
xor U8348 (N_8348,N_8057,N_8195);
nor U8349 (N_8349,N_8084,N_8139);
nor U8350 (N_8350,N_8150,N_8134);
xor U8351 (N_8351,N_8123,N_8063);
and U8352 (N_8352,N_8099,N_8127);
or U8353 (N_8353,N_8046,N_8115);
nand U8354 (N_8354,N_8176,N_8149);
xor U8355 (N_8355,N_8088,N_8012);
xor U8356 (N_8356,N_8085,N_8062);
or U8357 (N_8357,N_8161,N_8065);
nor U8358 (N_8358,N_8006,N_8026);
and U8359 (N_8359,N_8083,N_8100);
or U8360 (N_8360,N_8020,N_8147);
nor U8361 (N_8361,N_8163,N_8113);
or U8362 (N_8362,N_8134,N_8082);
nand U8363 (N_8363,N_8077,N_8121);
xor U8364 (N_8364,N_8021,N_8003);
or U8365 (N_8365,N_8034,N_8135);
and U8366 (N_8366,N_8028,N_8101);
nand U8367 (N_8367,N_8058,N_8195);
or U8368 (N_8368,N_8103,N_8080);
nor U8369 (N_8369,N_8101,N_8024);
xor U8370 (N_8370,N_8037,N_8190);
nor U8371 (N_8371,N_8032,N_8031);
and U8372 (N_8372,N_8022,N_8187);
and U8373 (N_8373,N_8013,N_8109);
or U8374 (N_8374,N_8124,N_8018);
xnor U8375 (N_8375,N_8059,N_8106);
nand U8376 (N_8376,N_8114,N_8021);
or U8377 (N_8377,N_8085,N_8077);
nand U8378 (N_8378,N_8185,N_8045);
and U8379 (N_8379,N_8132,N_8121);
xor U8380 (N_8380,N_8166,N_8114);
xnor U8381 (N_8381,N_8137,N_8099);
xor U8382 (N_8382,N_8139,N_8171);
nand U8383 (N_8383,N_8031,N_8034);
nor U8384 (N_8384,N_8191,N_8044);
xor U8385 (N_8385,N_8164,N_8087);
xnor U8386 (N_8386,N_8038,N_8036);
and U8387 (N_8387,N_8174,N_8155);
nand U8388 (N_8388,N_8100,N_8116);
or U8389 (N_8389,N_8091,N_8029);
xnor U8390 (N_8390,N_8052,N_8016);
xor U8391 (N_8391,N_8084,N_8099);
nor U8392 (N_8392,N_8022,N_8028);
nand U8393 (N_8393,N_8190,N_8104);
nand U8394 (N_8394,N_8091,N_8013);
nor U8395 (N_8395,N_8115,N_8019);
xor U8396 (N_8396,N_8142,N_8030);
nand U8397 (N_8397,N_8146,N_8098);
nor U8398 (N_8398,N_8097,N_8148);
xnor U8399 (N_8399,N_8197,N_8088);
or U8400 (N_8400,N_8392,N_8384);
xor U8401 (N_8401,N_8375,N_8258);
xnor U8402 (N_8402,N_8214,N_8382);
xor U8403 (N_8403,N_8268,N_8305);
nand U8404 (N_8404,N_8236,N_8373);
nor U8405 (N_8405,N_8307,N_8342);
or U8406 (N_8406,N_8275,N_8229);
and U8407 (N_8407,N_8388,N_8339);
or U8408 (N_8408,N_8309,N_8205);
or U8409 (N_8409,N_8243,N_8386);
nor U8410 (N_8410,N_8245,N_8274);
nor U8411 (N_8411,N_8237,N_8244);
nor U8412 (N_8412,N_8296,N_8312);
nand U8413 (N_8413,N_8304,N_8217);
nor U8414 (N_8414,N_8231,N_8396);
nor U8415 (N_8415,N_8207,N_8367);
nand U8416 (N_8416,N_8288,N_8201);
nor U8417 (N_8417,N_8356,N_8355);
or U8418 (N_8418,N_8262,N_8329);
nor U8419 (N_8419,N_8224,N_8393);
nor U8420 (N_8420,N_8354,N_8221);
nor U8421 (N_8421,N_8283,N_8265);
nor U8422 (N_8422,N_8253,N_8297);
xor U8423 (N_8423,N_8286,N_8238);
nor U8424 (N_8424,N_8223,N_8212);
nand U8425 (N_8425,N_8261,N_8206);
nand U8426 (N_8426,N_8289,N_8232);
nor U8427 (N_8427,N_8240,N_8226);
nor U8428 (N_8428,N_8324,N_8233);
and U8429 (N_8429,N_8228,N_8270);
xnor U8430 (N_8430,N_8280,N_8247);
or U8431 (N_8431,N_8284,N_8269);
nand U8432 (N_8432,N_8371,N_8241);
xnor U8433 (N_8433,N_8395,N_8372);
nor U8434 (N_8434,N_8316,N_8368);
xor U8435 (N_8435,N_8377,N_8353);
xnor U8436 (N_8436,N_8365,N_8204);
nand U8437 (N_8437,N_8248,N_8255);
xnor U8438 (N_8438,N_8336,N_8234);
xor U8439 (N_8439,N_8389,N_8338);
xor U8440 (N_8440,N_8218,N_8378);
nand U8441 (N_8441,N_8203,N_8318);
nor U8442 (N_8442,N_8293,N_8321);
and U8443 (N_8443,N_8374,N_8285);
nor U8444 (N_8444,N_8209,N_8310);
or U8445 (N_8445,N_8295,N_8350);
nor U8446 (N_8446,N_8302,N_8264);
nor U8447 (N_8447,N_8235,N_8225);
nand U8448 (N_8448,N_8366,N_8246);
nor U8449 (N_8449,N_8251,N_8202);
and U8450 (N_8450,N_8337,N_8344);
or U8451 (N_8451,N_8369,N_8271);
nand U8452 (N_8452,N_8357,N_8249);
or U8453 (N_8453,N_8299,N_8323);
and U8454 (N_8454,N_8327,N_8343);
nand U8455 (N_8455,N_8391,N_8325);
xor U8456 (N_8456,N_8379,N_8290);
and U8457 (N_8457,N_8326,N_8266);
nand U8458 (N_8458,N_8311,N_8359);
xnor U8459 (N_8459,N_8383,N_8213);
nand U8460 (N_8460,N_8227,N_8317);
nand U8461 (N_8461,N_8394,N_8260);
xor U8462 (N_8462,N_8294,N_8331);
nor U8463 (N_8463,N_8361,N_8282);
and U8464 (N_8464,N_8360,N_8298);
nand U8465 (N_8465,N_8276,N_8239);
or U8466 (N_8466,N_8281,N_8259);
and U8467 (N_8467,N_8222,N_8279);
nand U8468 (N_8468,N_8332,N_8345);
xnor U8469 (N_8469,N_8381,N_8363);
or U8470 (N_8470,N_8349,N_8267);
and U8471 (N_8471,N_8376,N_8328);
nor U8472 (N_8472,N_8320,N_8292);
nor U8473 (N_8473,N_8200,N_8230);
nand U8474 (N_8474,N_8273,N_8303);
or U8475 (N_8475,N_8347,N_8341);
nor U8476 (N_8476,N_8351,N_8256);
and U8477 (N_8477,N_8319,N_8219);
nand U8478 (N_8478,N_8335,N_8398);
and U8479 (N_8479,N_8210,N_8220);
nor U8480 (N_8480,N_8300,N_8370);
and U8481 (N_8481,N_8330,N_8352);
xnor U8482 (N_8482,N_8287,N_8291);
nor U8483 (N_8483,N_8257,N_8380);
and U8484 (N_8484,N_8301,N_8348);
or U8485 (N_8485,N_8277,N_8313);
and U8486 (N_8486,N_8358,N_8263);
or U8487 (N_8487,N_8387,N_8314);
xnor U8488 (N_8488,N_8346,N_8272);
or U8489 (N_8489,N_8399,N_8315);
nand U8490 (N_8490,N_8333,N_8322);
and U8491 (N_8491,N_8216,N_8390);
xor U8492 (N_8492,N_8362,N_8208);
nand U8493 (N_8493,N_8242,N_8254);
xor U8494 (N_8494,N_8278,N_8252);
nor U8495 (N_8495,N_8211,N_8308);
and U8496 (N_8496,N_8306,N_8340);
and U8497 (N_8497,N_8250,N_8215);
or U8498 (N_8498,N_8385,N_8334);
xnor U8499 (N_8499,N_8364,N_8397);
nor U8500 (N_8500,N_8352,N_8314);
nand U8501 (N_8501,N_8279,N_8333);
or U8502 (N_8502,N_8205,N_8259);
nand U8503 (N_8503,N_8350,N_8320);
nand U8504 (N_8504,N_8241,N_8321);
nor U8505 (N_8505,N_8231,N_8390);
or U8506 (N_8506,N_8386,N_8314);
nand U8507 (N_8507,N_8387,N_8362);
nand U8508 (N_8508,N_8276,N_8231);
xnor U8509 (N_8509,N_8349,N_8233);
nor U8510 (N_8510,N_8224,N_8332);
nand U8511 (N_8511,N_8345,N_8240);
and U8512 (N_8512,N_8265,N_8291);
nor U8513 (N_8513,N_8349,N_8346);
and U8514 (N_8514,N_8254,N_8211);
nor U8515 (N_8515,N_8286,N_8332);
and U8516 (N_8516,N_8397,N_8356);
or U8517 (N_8517,N_8288,N_8224);
or U8518 (N_8518,N_8226,N_8264);
and U8519 (N_8519,N_8212,N_8356);
xnor U8520 (N_8520,N_8353,N_8317);
nand U8521 (N_8521,N_8335,N_8200);
or U8522 (N_8522,N_8395,N_8381);
nor U8523 (N_8523,N_8355,N_8308);
nor U8524 (N_8524,N_8294,N_8350);
nand U8525 (N_8525,N_8214,N_8344);
and U8526 (N_8526,N_8354,N_8359);
xnor U8527 (N_8527,N_8316,N_8288);
nand U8528 (N_8528,N_8374,N_8325);
and U8529 (N_8529,N_8307,N_8287);
and U8530 (N_8530,N_8321,N_8332);
xor U8531 (N_8531,N_8397,N_8282);
or U8532 (N_8532,N_8312,N_8239);
nor U8533 (N_8533,N_8264,N_8379);
xnor U8534 (N_8534,N_8264,N_8358);
nor U8535 (N_8535,N_8313,N_8357);
nor U8536 (N_8536,N_8351,N_8324);
nor U8537 (N_8537,N_8229,N_8268);
nand U8538 (N_8538,N_8255,N_8333);
xor U8539 (N_8539,N_8205,N_8268);
or U8540 (N_8540,N_8243,N_8320);
nor U8541 (N_8541,N_8358,N_8337);
nand U8542 (N_8542,N_8345,N_8371);
xor U8543 (N_8543,N_8310,N_8372);
or U8544 (N_8544,N_8336,N_8387);
or U8545 (N_8545,N_8213,N_8262);
xor U8546 (N_8546,N_8350,N_8298);
xor U8547 (N_8547,N_8297,N_8227);
and U8548 (N_8548,N_8201,N_8222);
or U8549 (N_8549,N_8388,N_8381);
xnor U8550 (N_8550,N_8311,N_8257);
nand U8551 (N_8551,N_8284,N_8305);
and U8552 (N_8552,N_8365,N_8329);
xnor U8553 (N_8553,N_8342,N_8260);
nand U8554 (N_8554,N_8316,N_8242);
nor U8555 (N_8555,N_8291,N_8289);
and U8556 (N_8556,N_8207,N_8302);
nand U8557 (N_8557,N_8232,N_8257);
or U8558 (N_8558,N_8262,N_8318);
and U8559 (N_8559,N_8363,N_8273);
nor U8560 (N_8560,N_8252,N_8265);
and U8561 (N_8561,N_8324,N_8326);
or U8562 (N_8562,N_8288,N_8302);
or U8563 (N_8563,N_8288,N_8208);
and U8564 (N_8564,N_8387,N_8339);
xnor U8565 (N_8565,N_8348,N_8323);
nand U8566 (N_8566,N_8362,N_8349);
or U8567 (N_8567,N_8292,N_8243);
and U8568 (N_8568,N_8257,N_8244);
xnor U8569 (N_8569,N_8354,N_8226);
nand U8570 (N_8570,N_8385,N_8348);
and U8571 (N_8571,N_8311,N_8324);
xnor U8572 (N_8572,N_8230,N_8350);
nand U8573 (N_8573,N_8210,N_8268);
and U8574 (N_8574,N_8232,N_8207);
nor U8575 (N_8575,N_8369,N_8311);
nand U8576 (N_8576,N_8337,N_8348);
and U8577 (N_8577,N_8300,N_8255);
and U8578 (N_8578,N_8296,N_8244);
nor U8579 (N_8579,N_8238,N_8357);
nand U8580 (N_8580,N_8219,N_8243);
xnor U8581 (N_8581,N_8313,N_8256);
nor U8582 (N_8582,N_8275,N_8266);
and U8583 (N_8583,N_8336,N_8372);
xnor U8584 (N_8584,N_8280,N_8224);
and U8585 (N_8585,N_8276,N_8354);
nor U8586 (N_8586,N_8360,N_8277);
nor U8587 (N_8587,N_8205,N_8316);
xnor U8588 (N_8588,N_8272,N_8302);
or U8589 (N_8589,N_8372,N_8244);
nand U8590 (N_8590,N_8299,N_8287);
and U8591 (N_8591,N_8369,N_8381);
or U8592 (N_8592,N_8281,N_8363);
nand U8593 (N_8593,N_8263,N_8384);
and U8594 (N_8594,N_8385,N_8204);
or U8595 (N_8595,N_8277,N_8350);
nor U8596 (N_8596,N_8246,N_8385);
nand U8597 (N_8597,N_8284,N_8346);
nand U8598 (N_8598,N_8273,N_8351);
nor U8599 (N_8599,N_8354,N_8391);
or U8600 (N_8600,N_8518,N_8464);
or U8601 (N_8601,N_8594,N_8559);
and U8602 (N_8602,N_8436,N_8419);
nor U8603 (N_8603,N_8582,N_8598);
nand U8604 (N_8604,N_8413,N_8416);
or U8605 (N_8605,N_8405,N_8584);
nor U8606 (N_8606,N_8540,N_8472);
and U8607 (N_8607,N_8514,N_8430);
and U8608 (N_8608,N_8519,N_8505);
nor U8609 (N_8609,N_8572,N_8593);
nor U8610 (N_8610,N_8500,N_8415);
or U8611 (N_8611,N_8573,N_8507);
or U8612 (N_8612,N_8541,N_8468);
nand U8613 (N_8613,N_8467,N_8524);
nand U8614 (N_8614,N_8567,N_8482);
and U8615 (N_8615,N_8438,N_8520);
xnor U8616 (N_8616,N_8435,N_8565);
nand U8617 (N_8617,N_8485,N_8450);
nor U8618 (N_8618,N_8401,N_8599);
nor U8619 (N_8619,N_8466,N_8506);
nor U8620 (N_8620,N_8433,N_8568);
nand U8621 (N_8621,N_8560,N_8508);
and U8622 (N_8622,N_8510,N_8595);
xor U8623 (N_8623,N_8539,N_8421);
and U8624 (N_8624,N_8422,N_8457);
xor U8625 (N_8625,N_8471,N_8414);
and U8626 (N_8626,N_8420,N_8583);
and U8627 (N_8627,N_8554,N_8486);
xnor U8628 (N_8628,N_8418,N_8527);
nor U8629 (N_8629,N_8447,N_8571);
and U8630 (N_8630,N_8570,N_8417);
nand U8631 (N_8631,N_8569,N_8470);
xnor U8632 (N_8632,N_8452,N_8523);
nor U8633 (N_8633,N_8442,N_8548);
or U8634 (N_8634,N_8410,N_8478);
xor U8635 (N_8635,N_8460,N_8484);
nor U8636 (N_8636,N_8531,N_8516);
nor U8637 (N_8637,N_8495,N_8562);
or U8638 (N_8638,N_8443,N_8504);
xnor U8639 (N_8639,N_8465,N_8469);
and U8640 (N_8640,N_8425,N_8588);
or U8641 (N_8641,N_8532,N_8463);
nor U8642 (N_8642,N_8444,N_8493);
nand U8643 (N_8643,N_8563,N_8591);
nor U8644 (N_8644,N_8592,N_8546);
and U8645 (N_8645,N_8578,N_8581);
and U8646 (N_8646,N_8474,N_8530);
or U8647 (N_8647,N_8432,N_8533);
or U8648 (N_8648,N_8446,N_8441);
and U8649 (N_8649,N_8454,N_8542);
and U8650 (N_8650,N_8449,N_8407);
or U8651 (N_8651,N_8475,N_8445);
nand U8652 (N_8652,N_8458,N_8521);
nor U8653 (N_8653,N_8538,N_8587);
or U8654 (N_8654,N_8590,N_8488);
xnor U8655 (N_8655,N_8512,N_8580);
nor U8656 (N_8656,N_8491,N_8402);
and U8657 (N_8657,N_8575,N_8476);
nor U8658 (N_8658,N_8459,N_8544);
nand U8659 (N_8659,N_8456,N_8497);
nand U8660 (N_8660,N_8537,N_8503);
or U8661 (N_8661,N_8552,N_8564);
xor U8662 (N_8662,N_8557,N_8412);
and U8663 (N_8663,N_8492,N_8439);
nor U8664 (N_8664,N_8461,N_8424);
and U8665 (N_8665,N_8498,N_8525);
or U8666 (N_8666,N_8501,N_8403);
xor U8667 (N_8667,N_8423,N_8522);
nor U8668 (N_8668,N_8499,N_8409);
nand U8669 (N_8669,N_8487,N_8534);
xor U8670 (N_8670,N_8509,N_8547);
and U8671 (N_8671,N_8517,N_8528);
nand U8672 (N_8672,N_8427,N_8543);
nor U8673 (N_8673,N_8428,N_8490);
and U8674 (N_8674,N_8586,N_8545);
nor U8675 (N_8675,N_8555,N_8462);
nor U8676 (N_8676,N_8406,N_8479);
nor U8677 (N_8677,N_8536,N_8434);
nand U8678 (N_8678,N_8579,N_8513);
nand U8679 (N_8679,N_8526,N_8529);
nor U8680 (N_8680,N_8400,N_8496);
or U8681 (N_8681,N_8550,N_8426);
or U8682 (N_8682,N_8551,N_8483);
or U8683 (N_8683,N_8453,N_8549);
xnor U8684 (N_8684,N_8494,N_8440);
nand U8685 (N_8685,N_8566,N_8429);
nand U8686 (N_8686,N_8574,N_8561);
or U8687 (N_8687,N_8558,N_8553);
nand U8688 (N_8688,N_8585,N_8577);
nor U8689 (N_8689,N_8473,N_8515);
nor U8690 (N_8690,N_8448,N_8451);
nand U8691 (N_8691,N_8408,N_8477);
xnor U8692 (N_8692,N_8480,N_8597);
or U8693 (N_8693,N_8589,N_8502);
nand U8694 (N_8694,N_8481,N_8437);
nand U8695 (N_8695,N_8556,N_8489);
nor U8696 (N_8696,N_8411,N_8404);
and U8697 (N_8697,N_8455,N_8431);
xnor U8698 (N_8698,N_8535,N_8511);
nand U8699 (N_8699,N_8596,N_8576);
nand U8700 (N_8700,N_8406,N_8552);
or U8701 (N_8701,N_8517,N_8434);
nor U8702 (N_8702,N_8486,N_8523);
and U8703 (N_8703,N_8520,N_8592);
and U8704 (N_8704,N_8503,N_8432);
nor U8705 (N_8705,N_8430,N_8434);
nand U8706 (N_8706,N_8461,N_8534);
nor U8707 (N_8707,N_8540,N_8591);
xnor U8708 (N_8708,N_8455,N_8506);
and U8709 (N_8709,N_8525,N_8574);
nor U8710 (N_8710,N_8425,N_8470);
and U8711 (N_8711,N_8487,N_8450);
xnor U8712 (N_8712,N_8469,N_8490);
nand U8713 (N_8713,N_8545,N_8485);
or U8714 (N_8714,N_8492,N_8445);
or U8715 (N_8715,N_8544,N_8583);
xor U8716 (N_8716,N_8516,N_8437);
nor U8717 (N_8717,N_8541,N_8564);
xor U8718 (N_8718,N_8556,N_8536);
and U8719 (N_8719,N_8428,N_8557);
and U8720 (N_8720,N_8433,N_8591);
and U8721 (N_8721,N_8461,N_8445);
xor U8722 (N_8722,N_8563,N_8488);
nand U8723 (N_8723,N_8503,N_8456);
or U8724 (N_8724,N_8432,N_8471);
xnor U8725 (N_8725,N_8478,N_8471);
nand U8726 (N_8726,N_8466,N_8527);
xor U8727 (N_8727,N_8449,N_8493);
nand U8728 (N_8728,N_8494,N_8480);
nand U8729 (N_8729,N_8443,N_8425);
or U8730 (N_8730,N_8489,N_8582);
and U8731 (N_8731,N_8408,N_8428);
and U8732 (N_8732,N_8514,N_8551);
nand U8733 (N_8733,N_8530,N_8533);
and U8734 (N_8734,N_8531,N_8464);
and U8735 (N_8735,N_8559,N_8420);
and U8736 (N_8736,N_8484,N_8480);
and U8737 (N_8737,N_8430,N_8515);
or U8738 (N_8738,N_8597,N_8415);
nor U8739 (N_8739,N_8404,N_8516);
xnor U8740 (N_8740,N_8435,N_8534);
xnor U8741 (N_8741,N_8579,N_8470);
nand U8742 (N_8742,N_8572,N_8470);
or U8743 (N_8743,N_8496,N_8589);
xor U8744 (N_8744,N_8476,N_8534);
and U8745 (N_8745,N_8539,N_8437);
nand U8746 (N_8746,N_8447,N_8588);
nand U8747 (N_8747,N_8421,N_8498);
nor U8748 (N_8748,N_8480,N_8434);
nor U8749 (N_8749,N_8407,N_8547);
and U8750 (N_8750,N_8521,N_8539);
xnor U8751 (N_8751,N_8570,N_8402);
xor U8752 (N_8752,N_8584,N_8599);
nor U8753 (N_8753,N_8413,N_8434);
nand U8754 (N_8754,N_8512,N_8400);
xor U8755 (N_8755,N_8475,N_8490);
nor U8756 (N_8756,N_8405,N_8574);
xnor U8757 (N_8757,N_8468,N_8401);
and U8758 (N_8758,N_8466,N_8450);
or U8759 (N_8759,N_8591,N_8547);
xor U8760 (N_8760,N_8413,N_8484);
xor U8761 (N_8761,N_8406,N_8446);
nand U8762 (N_8762,N_8422,N_8561);
xnor U8763 (N_8763,N_8589,N_8430);
and U8764 (N_8764,N_8556,N_8557);
and U8765 (N_8765,N_8420,N_8438);
nand U8766 (N_8766,N_8402,N_8458);
and U8767 (N_8767,N_8492,N_8453);
and U8768 (N_8768,N_8438,N_8526);
or U8769 (N_8769,N_8573,N_8516);
nand U8770 (N_8770,N_8561,N_8479);
and U8771 (N_8771,N_8587,N_8542);
nand U8772 (N_8772,N_8460,N_8519);
or U8773 (N_8773,N_8519,N_8473);
or U8774 (N_8774,N_8407,N_8508);
nor U8775 (N_8775,N_8440,N_8454);
nor U8776 (N_8776,N_8431,N_8496);
nand U8777 (N_8777,N_8514,N_8464);
and U8778 (N_8778,N_8553,N_8422);
xor U8779 (N_8779,N_8482,N_8457);
and U8780 (N_8780,N_8554,N_8403);
or U8781 (N_8781,N_8475,N_8531);
nand U8782 (N_8782,N_8492,N_8454);
xor U8783 (N_8783,N_8497,N_8565);
xnor U8784 (N_8784,N_8493,N_8504);
xnor U8785 (N_8785,N_8494,N_8484);
nor U8786 (N_8786,N_8444,N_8485);
xnor U8787 (N_8787,N_8433,N_8415);
or U8788 (N_8788,N_8564,N_8463);
and U8789 (N_8789,N_8466,N_8509);
or U8790 (N_8790,N_8504,N_8401);
xnor U8791 (N_8791,N_8581,N_8592);
nand U8792 (N_8792,N_8448,N_8547);
nand U8793 (N_8793,N_8575,N_8543);
nand U8794 (N_8794,N_8434,N_8502);
nand U8795 (N_8795,N_8484,N_8595);
or U8796 (N_8796,N_8429,N_8435);
or U8797 (N_8797,N_8415,N_8430);
xor U8798 (N_8798,N_8575,N_8443);
nand U8799 (N_8799,N_8506,N_8551);
nand U8800 (N_8800,N_8797,N_8738);
and U8801 (N_8801,N_8725,N_8761);
nand U8802 (N_8802,N_8643,N_8607);
and U8803 (N_8803,N_8749,N_8685);
nor U8804 (N_8804,N_8731,N_8666);
and U8805 (N_8805,N_8795,N_8732);
nand U8806 (N_8806,N_8648,N_8694);
nand U8807 (N_8807,N_8611,N_8602);
nor U8808 (N_8808,N_8695,N_8659);
or U8809 (N_8809,N_8723,N_8672);
or U8810 (N_8810,N_8651,N_8728);
nor U8811 (N_8811,N_8698,N_8783);
and U8812 (N_8812,N_8702,N_8781);
xnor U8813 (N_8813,N_8724,N_8771);
and U8814 (N_8814,N_8791,N_8677);
or U8815 (N_8815,N_8600,N_8630);
or U8816 (N_8816,N_8641,N_8755);
and U8817 (N_8817,N_8645,N_8650);
nand U8818 (N_8818,N_8633,N_8774);
or U8819 (N_8819,N_8626,N_8625);
and U8820 (N_8820,N_8740,N_8624);
and U8821 (N_8821,N_8713,N_8644);
and U8822 (N_8822,N_8693,N_8606);
and U8823 (N_8823,N_8608,N_8766);
xnor U8824 (N_8824,N_8734,N_8722);
and U8825 (N_8825,N_8619,N_8726);
nor U8826 (N_8826,N_8690,N_8746);
and U8827 (N_8827,N_8748,N_8753);
and U8828 (N_8828,N_8776,N_8711);
xor U8829 (N_8829,N_8668,N_8744);
and U8830 (N_8830,N_8796,N_8664);
nand U8831 (N_8831,N_8681,N_8620);
and U8832 (N_8832,N_8629,N_8621);
nor U8833 (N_8833,N_8727,N_8770);
or U8834 (N_8834,N_8736,N_8660);
nor U8835 (N_8835,N_8788,N_8710);
or U8836 (N_8836,N_8762,N_8640);
or U8837 (N_8837,N_8730,N_8721);
or U8838 (N_8838,N_8707,N_8669);
or U8839 (N_8839,N_8705,N_8635);
and U8840 (N_8840,N_8623,N_8793);
and U8841 (N_8841,N_8604,N_8657);
nand U8842 (N_8842,N_8637,N_8649);
and U8843 (N_8843,N_8778,N_8691);
nand U8844 (N_8844,N_8696,N_8786);
nor U8845 (N_8845,N_8618,N_8703);
nand U8846 (N_8846,N_8794,N_8772);
xnor U8847 (N_8847,N_8706,N_8658);
nor U8848 (N_8848,N_8751,N_8739);
xnor U8849 (N_8849,N_8647,N_8759);
xor U8850 (N_8850,N_8743,N_8716);
or U8851 (N_8851,N_8775,N_8714);
or U8852 (N_8852,N_8735,N_8675);
nor U8853 (N_8853,N_8684,N_8639);
and U8854 (N_8854,N_8653,N_8792);
xor U8855 (N_8855,N_8697,N_8613);
and U8856 (N_8856,N_8718,N_8634);
and U8857 (N_8857,N_8603,N_8757);
xor U8858 (N_8858,N_8642,N_8656);
and U8859 (N_8859,N_8686,N_8687);
xnor U8860 (N_8860,N_8747,N_8756);
nor U8861 (N_8861,N_8750,N_8679);
nor U8862 (N_8862,N_8689,N_8622);
or U8863 (N_8863,N_8717,N_8671);
or U8864 (N_8864,N_8674,N_8767);
nor U8865 (N_8865,N_8737,N_8708);
nand U8866 (N_8866,N_8779,N_8760);
nor U8867 (N_8867,N_8652,N_8601);
nor U8868 (N_8868,N_8646,N_8758);
and U8869 (N_8869,N_8662,N_8719);
and U8870 (N_8870,N_8628,N_8754);
or U8871 (N_8871,N_8673,N_8667);
and U8872 (N_8872,N_8614,N_8638);
and U8873 (N_8873,N_8665,N_8789);
and U8874 (N_8874,N_8798,N_8780);
nand U8875 (N_8875,N_8785,N_8654);
nand U8876 (N_8876,N_8773,N_8699);
and U8877 (N_8877,N_8605,N_8741);
and U8878 (N_8878,N_8670,N_8701);
xor U8879 (N_8879,N_8733,N_8612);
nand U8880 (N_8880,N_8700,N_8631);
nand U8881 (N_8881,N_8636,N_8715);
or U8882 (N_8882,N_8765,N_8678);
xor U8883 (N_8883,N_8676,N_8627);
nand U8884 (N_8884,N_8720,N_8769);
nor U8885 (N_8885,N_8777,N_8768);
and U8886 (N_8886,N_8682,N_8729);
nand U8887 (N_8887,N_8712,N_8661);
xnor U8888 (N_8888,N_8799,N_8763);
and U8889 (N_8889,N_8683,N_8709);
or U8890 (N_8890,N_8704,N_8655);
and U8891 (N_8891,N_8745,N_8617);
or U8892 (N_8892,N_8680,N_8782);
nor U8893 (N_8893,N_8784,N_8688);
and U8894 (N_8894,N_8610,N_8787);
or U8895 (N_8895,N_8790,N_8752);
xnor U8896 (N_8896,N_8764,N_8616);
nand U8897 (N_8897,N_8615,N_8632);
xnor U8898 (N_8898,N_8742,N_8609);
xnor U8899 (N_8899,N_8663,N_8692);
and U8900 (N_8900,N_8624,N_8692);
and U8901 (N_8901,N_8732,N_8790);
nor U8902 (N_8902,N_8686,N_8771);
nand U8903 (N_8903,N_8672,N_8601);
nand U8904 (N_8904,N_8655,N_8618);
and U8905 (N_8905,N_8655,N_8673);
nor U8906 (N_8906,N_8716,N_8740);
xor U8907 (N_8907,N_8618,N_8632);
xor U8908 (N_8908,N_8763,N_8790);
or U8909 (N_8909,N_8706,N_8700);
nand U8910 (N_8910,N_8652,N_8634);
xnor U8911 (N_8911,N_8757,N_8698);
or U8912 (N_8912,N_8663,N_8622);
and U8913 (N_8913,N_8798,N_8769);
xor U8914 (N_8914,N_8749,N_8648);
xor U8915 (N_8915,N_8601,N_8732);
and U8916 (N_8916,N_8785,N_8675);
or U8917 (N_8917,N_8752,N_8751);
and U8918 (N_8918,N_8670,N_8698);
nand U8919 (N_8919,N_8767,N_8666);
xor U8920 (N_8920,N_8786,N_8721);
nand U8921 (N_8921,N_8727,N_8621);
xnor U8922 (N_8922,N_8652,N_8698);
or U8923 (N_8923,N_8740,N_8706);
or U8924 (N_8924,N_8748,N_8789);
xnor U8925 (N_8925,N_8613,N_8666);
and U8926 (N_8926,N_8760,N_8666);
xnor U8927 (N_8927,N_8622,N_8629);
nand U8928 (N_8928,N_8661,N_8631);
xor U8929 (N_8929,N_8730,N_8784);
nor U8930 (N_8930,N_8735,N_8681);
or U8931 (N_8931,N_8726,N_8751);
and U8932 (N_8932,N_8649,N_8642);
nand U8933 (N_8933,N_8633,N_8779);
and U8934 (N_8934,N_8683,N_8634);
nor U8935 (N_8935,N_8767,N_8684);
or U8936 (N_8936,N_8763,N_8689);
nand U8937 (N_8937,N_8789,N_8765);
or U8938 (N_8938,N_8610,N_8601);
and U8939 (N_8939,N_8695,N_8614);
nor U8940 (N_8940,N_8720,N_8657);
nand U8941 (N_8941,N_8647,N_8605);
nor U8942 (N_8942,N_8713,N_8692);
nor U8943 (N_8943,N_8643,N_8692);
or U8944 (N_8944,N_8612,N_8646);
and U8945 (N_8945,N_8684,N_8678);
or U8946 (N_8946,N_8602,N_8747);
nand U8947 (N_8947,N_8605,N_8624);
xor U8948 (N_8948,N_8754,N_8686);
nor U8949 (N_8949,N_8755,N_8691);
nand U8950 (N_8950,N_8704,N_8681);
nand U8951 (N_8951,N_8786,N_8668);
xor U8952 (N_8952,N_8685,N_8741);
xor U8953 (N_8953,N_8704,N_8731);
or U8954 (N_8954,N_8756,N_8739);
nor U8955 (N_8955,N_8786,N_8763);
nor U8956 (N_8956,N_8779,N_8753);
xnor U8957 (N_8957,N_8701,N_8726);
nor U8958 (N_8958,N_8757,N_8618);
nand U8959 (N_8959,N_8659,N_8613);
nor U8960 (N_8960,N_8687,N_8651);
nand U8961 (N_8961,N_8702,N_8722);
nor U8962 (N_8962,N_8696,N_8727);
and U8963 (N_8963,N_8612,N_8698);
and U8964 (N_8964,N_8605,N_8622);
nand U8965 (N_8965,N_8736,N_8667);
xor U8966 (N_8966,N_8722,N_8657);
or U8967 (N_8967,N_8764,N_8762);
nor U8968 (N_8968,N_8745,N_8646);
nor U8969 (N_8969,N_8610,N_8732);
nor U8970 (N_8970,N_8707,N_8643);
or U8971 (N_8971,N_8779,N_8656);
xnor U8972 (N_8972,N_8749,N_8763);
nor U8973 (N_8973,N_8657,N_8735);
xnor U8974 (N_8974,N_8677,N_8766);
xnor U8975 (N_8975,N_8645,N_8755);
or U8976 (N_8976,N_8727,N_8793);
and U8977 (N_8977,N_8644,N_8743);
or U8978 (N_8978,N_8749,N_8641);
nand U8979 (N_8979,N_8710,N_8761);
nand U8980 (N_8980,N_8679,N_8663);
nor U8981 (N_8981,N_8624,N_8736);
nand U8982 (N_8982,N_8666,N_8668);
or U8983 (N_8983,N_8734,N_8620);
xnor U8984 (N_8984,N_8615,N_8641);
or U8985 (N_8985,N_8781,N_8744);
or U8986 (N_8986,N_8785,N_8793);
nand U8987 (N_8987,N_8605,N_8731);
nand U8988 (N_8988,N_8703,N_8732);
xnor U8989 (N_8989,N_8738,N_8637);
and U8990 (N_8990,N_8642,N_8623);
and U8991 (N_8991,N_8751,N_8657);
nor U8992 (N_8992,N_8763,N_8683);
nand U8993 (N_8993,N_8638,N_8787);
and U8994 (N_8994,N_8799,N_8738);
nand U8995 (N_8995,N_8768,N_8675);
and U8996 (N_8996,N_8743,N_8751);
xor U8997 (N_8997,N_8664,N_8637);
nor U8998 (N_8998,N_8725,N_8626);
or U8999 (N_8999,N_8717,N_8664);
and U9000 (N_9000,N_8950,N_8881);
or U9001 (N_9001,N_8988,N_8948);
nor U9002 (N_9002,N_8982,N_8840);
nand U9003 (N_9003,N_8888,N_8921);
xor U9004 (N_9004,N_8857,N_8917);
or U9005 (N_9005,N_8860,N_8871);
nor U9006 (N_9006,N_8933,N_8838);
nand U9007 (N_9007,N_8851,N_8943);
nand U9008 (N_9008,N_8910,N_8971);
nand U9009 (N_9009,N_8949,N_8855);
and U9010 (N_9010,N_8873,N_8832);
nand U9011 (N_9011,N_8807,N_8898);
xnor U9012 (N_9012,N_8986,N_8821);
xnor U9013 (N_9013,N_8876,N_8895);
nand U9014 (N_9014,N_8992,N_8997);
nand U9015 (N_9015,N_8893,N_8908);
xor U9016 (N_9016,N_8830,N_8822);
or U9017 (N_9017,N_8818,N_8810);
and U9018 (N_9018,N_8934,N_8942);
nand U9019 (N_9019,N_8843,N_8935);
xor U9020 (N_9020,N_8983,N_8841);
and U9021 (N_9021,N_8834,N_8975);
xnor U9022 (N_9022,N_8804,N_8813);
and U9023 (N_9023,N_8977,N_8823);
nand U9024 (N_9024,N_8985,N_8845);
or U9025 (N_9025,N_8809,N_8803);
nor U9026 (N_9026,N_8800,N_8815);
or U9027 (N_9027,N_8909,N_8850);
or U9028 (N_9028,N_8839,N_8964);
nor U9029 (N_9029,N_8951,N_8966);
or U9030 (N_9030,N_8945,N_8849);
or U9031 (N_9031,N_8907,N_8998);
xor U9032 (N_9032,N_8848,N_8884);
nor U9033 (N_9033,N_8903,N_8938);
or U9034 (N_9034,N_8928,N_8811);
nor U9035 (N_9035,N_8906,N_8872);
and U9036 (N_9036,N_8926,N_8931);
nand U9037 (N_9037,N_8896,N_8930);
xnor U9038 (N_9038,N_8885,N_8980);
and U9039 (N_9039,N_8987,N_8847);
or U9040 (N_9040,N_8905,N_8874);
or U9041 (N_9041,N_8941,N_8958);
nand U9042 (N_9042,N_8814,N_8877);
or U9043 (N_9043,N_8904,N_8954);
and U9044 (N_9044,N_8918,N_8853);
nand U9045 (N_9045,N_8865,N_8861);
xnor U9046 (N_9046,N_8858,N_8944);
and U9047 (N_9047,N_8835,N_8867);
or U9048 (N_9048,N_8925,N_8869);
nand U9049 (N_9049,N_8891,N_8916);
xnor U9050 (N_9050,N_8828,N_8882);
xnor U9051 (N_9051,N_8863,N_8956);
or U9052 (N_9052,N_8939,N_8940);
nor U9053 (N_9053,N_8808,N_8991);
and U9054 (N_9054,N_8864,N_8883);
nand U9055 (N_9055,N_8880,N_8802);
nand U9056 (N_9056,N_8923,N_8886);
or U9057 (N_9057,N_8947,N_8955);
or U9058 (N_9058,N_8854,N_8967);
nand U9059 (N_9059,N_8961,N_8932);
xnor U9060 (N_9060,N_8833,N_8959);
nand U9061 (N_9061,N_8870,N_8929);
nand U9062 (N_9062,N_8887,N_8826);
nor U9063 (N_9063,N_8825,N_8989);
or U9064 (N_9064,N_8969,N_8936);
and U9065 (N_9065,N_8911,N_8900);
and U9066 (N_9066,N_8819,N_8820);
nor U9067 (N_9067,N_8914,N_8862);
or U9068 (N_9068,N_8852,N_8879);
xnor U9069 (N_9069,N_8801,N_8920);
xor U9070 (N_9070,N_8994,N_8972);
xnor U9071 (N_9071,N_8999,N_8846);
or U9072 (N_9072,N_8868,N_8993);
and U9073 (N_9073,N_8995,N_8806);
nand U9074 (N_9074,N_8842,N_8957);
xnor U9075 (N_9075,N_8829,N_8902);
or U9076 (N_9076,N_8831,N_8875);
or U9077 (N_9077,N_8976,N_8952);
or U9078 (N_9078,N_8897,N_8894);
nor U9079 (N_9079,N_8979,N_8922);
nor U9080 (N_9080,N_8946,N_8970);
or U9081 (N_9081,N_8973,N_8984);
nand U9082 (N_9082,N_8913,N_8963);
xnor U9083 (N_9083,N_8892,N_8901);
and U9084 (N_9084,N_8990,N_8981);
and U9085 (N_9085,N_8924,N_8899);
nand U9086 (N_9086,N_8859,N_8965);
nor U9087 (N_9087,N_8844,N_8974);
xor U9088 (N_9088,N_8827,N_8915);
nor U9089 (N_9089,N_8836,N_8978);
or U9090 (N_9090,N_8837,N_8962);
and U9091 (N_9091,N_8805,N_8866);
and U9092 (N_9092,N_8889,N_8927);
nor U9093 (N_9093,N_8812,N_8816);
or U9094 (N_9094,N_8824,N_8817);
xnor U9095 (N_9095,N_8890,N_8878);
nand U9096 (N_9096,N_8968,N_8919);
xor U9097 (N_9097,N_8960,N_8856);
nor U9098 (N_9098,N_8953,N_8937);
and U9099 (N_9099,N_8912,N_8996);
nand U9100 (N_9100,N_8812,N_8828);
and U9101 (N_9101,N_8805,N_8918);
nand U9102 (N_9102,N_8956,N_8895);
and U9103 (N_9103,N_8930,N_8915);
nand U9104 (N_9104,N_8893,N_8964);
and U9105 (N_9105,N_8833,N_8956);
or U9106 (N_9106,N_8995,N_8881);
nand U9107 (N_9107,N_8929,N_8820);
nand U9108 (N_9108,N_8981,N_8999);
or U9109 (N_9109,N_8931,N_8851);
nor U9110 (N_9110,N_8923,N_8882);
or U9111 (N_9111,N_8872,N_8845);
and U9112 (N_9112,N_8997,N_8949);
nand U9113 (N_9113,N_8832,N_8868);
nor U9114 (N_9114,N_8878,N_8951);
xnor U9115 (N_9115,N_8866,N_8902);
nand U9116 (N_9116,N_8838,N_8810);
nor U9117 (N_9117,N_8988,N_8908);
and U9118 (N_9118,N_8807,N_8958);
nand U9119 (N_9119,N_8905,N_8839);
and U9120 (N_9120,N_8961,N_8942);
nand U9121 (N_9121,N_8876,N_8875);
xnor U9122 (N_9122,N_8926,N_8999);
and U9123 (N_9123,N_8899,N_8922);
or U9124 (N_9124,N_8965,N_8842);
or U9125 (N_9125,N_8963,N_8998);
nand U9126 (N_9126,N_8919,N_8870);
and U9127 (N_9127,N_8873,N_8860);
and U9128 (N_9128,N_8970,N_8923);
or U9129 (N_9129,N_8925,N_8868);
and U9130 (N_9130,N_8837,N_8970);
and U9131 (N_9131,N_8936,N_8853);
or U9132 (N_9132,N_8830,N_8920);
xor U9133 (N_9133,N_8831,N_8977);
nor U9134 (N_9134,N_8853,N_8897);
or U9135 (N_9135,N_8952,N_8838);
or U9136 (N_9136,N_8991,N_8984);
and U9137 (N_9137,N_8821,N_8839);
and U9138 (N_9138,N_8975,N_8844);
xor U9139 (N_9139,N_8939,N_8805);
and U9140 (N_9140,N_8951,N_8834);
nand U9141 (N_9141,N_8915,N_8923);
nand U9142 (N_9142,N_8990,N_8987);
and U9143 (N_9143,N_8879,N_8951);
nand U9144 (N_9144,N_8869,N_8927);
xor U9145 (N_9145,N_8819,N_8865);
nand U9146 (N_9146,N_8947,N_8905);
and U9147 (N_9147,N_8934,N_8881);
xor U9148 (N_9148,N_8861,N_8973);
and U9149 (N_9149,N_8923,N_8995);
nand U9150 (N_9150,N_8926,N_8904);
nand U9151 (N_9151,N_8996,N_8884);
or U9152 (N_9152,N_8841,N_8953);
or U9153 (N_9153,N_8860,N_8964);
xor U9154 (N_9154,N_8991,N_8850);
or U9155 (N_9155,N_8974,N_8996);
and U9156 (N_9156,N_8817,N_8985);
or U9157 (N_9157,N_8986,N_8872);
xnor U9158 (N_9158,N_8858,N_8947);
or U9159 (N_9159,N_8968,N_8913);
or U9160 (N_9160,N_8992,N_8891);
nor U9161 (N_9161,N_8883,N_8983);
or U9162 (N_9162,N_8807,N_8976);
xnor U9163 (N_9163,N_8984,N_8912);
or U9164 (N_9164,N_8837,N_8866);
and U9165 (N_9165,N_8905,N_8934);
and U9166 (N_9166,N_8985,N_8968);
or U9167 (N_9167,N_8919,N_8924);
or U9168 (N_9168,N_8804,N_8901);
xor U9169 (N_9169,N_8801,N_8906);
nand U9170 (N_9170,N_8935,N_8944);
nand U9171 (N_9171,N_8967,N_8886);
xnor U9172 (N_9172,N_8949,N_8871);
xnor U9173 (N_9173,N_8904,N_8836);
xor U9174 (N_9174,N_8842,N_8900);
nand U9175 (N_9175,N_8913,N_8817);
or U9176 (N_9176,N_8950,N_8947);
nor U9177 (N_9177,N_8921,N_8990);
and U9178 (N_9178,N_8893,N_8825);
xor U9179 (N_9179,N_8879,N_8950);
xnor U9180 (N_9180,N_8903,N_8902);
nor U9181 (N_9181,N_8978,N_8821);
nor U9182 (N_9182,N_8851,N_8925);
and U9183 (N_9183,N_8842,N_8929);
nand U9184 (N_9184,N_8879,N_8960);
or U9185 (N_9185,N_8936,N_8907);
nand U9186 (N_9186,N_8898,N_8887);
and U9187 (N_9187,N_8937,N_8805);
or U9188 (N_9188,N_8924,N_8857);
xor U9189 (N_9189,N_8872,N_8978);
or U9190 (N_9190,N_8902,N_8865);
nor U9191 (N_9191,N_8979,N_8958);
xor U9192 (N_9192,N_8968,N_8833);
xnor U9193 (N_9193,N_8839,N_8871);
xnor U9194 (N_9194,N_8914,N_8996);
or U9195 (N_9195,N_8873,N_8941);
and U9196 (N_9196,N_8968,N_8974);
nor U9197 (N_9197,N_8994,N_8870);
and U9198 (N_9198,N_8904,N_8860);
nor U9199 (N_9199,N_8835,N_8876);
and U9200 (N_9200,N_9188,N_9093);
xnor U9201 (N_9201,N_9033,N_9105);
nor U9202 (N_9202,N_9059,N_9176);
and U9203 (N_9203,N_9127,N_9139);
or U9204 (N_9204,N_9118,N_9027);
nand U9205 (N_9205,N_9116,N_9121);
xor U9206 (N_9206,N_9091,N_9166);
xor U9207 (N_9207,N_9154,N_9014);
or U9208 (N_9208,N_9173,N_9081);
nand U9209 (N_9209,N_9045,N_9064);
or U9210 (N_9210,N_9049,N_9142);
or U9211 (N_9211,N_9025,N_9022);
and U9212 (N_9212,N_9174,N_9066);
xor U9213 (N_9213,N_9072,N_9075);
xnor U9214 (N_9214,N_9197,N_9067);
nand U9215 (N_9215,N_9042,N_9169);
or U9216 (N_9216,N_9103,N_9119);
and U9217 (N_9217,N_9088,N_9069);
xor U9218 (N_9218,N_9035,N_9147);
xnor U9219 (N_9219,N_9010,N_9018);
nand U9220 (N_9220,N_9160,N_9183);
nand U9221 (N_9221,N_9054,N_9082);
or U9222 (N_9222,N_9001,N_9086);
and U9223 (N_9223,N_9175,N_9016);
or U9224 (N_9224,N_9165,N_9040);
or U9225 (N_9225,N_9132,N_9194);
and U9226 (N_9226,N_9019,N_9151);
nor U9227 (N_9227,N_9052,N_9095);
nand U9228 (N_9228,N_9138,N_9156);
nand U9229 (N_9229,N_9078,N_9159);
and U9230 (N_9230,N_9092,N_9180);
nand U9231 (N_9231,N_9106,N_9074);
xnor U9232 (N_9232,N_9195,N_9006);
nand U9233 (N_9233,N_9189,N_9157);
and U9234 (N_9234,N_9123,N_9136);
or U9235 (N_9235,N_9161,N_9062);
nor U9236 (N_9236,N_9198,N_9083);
nand U9237 (N_9237,N_9050,N_9191);
nor U9238 (N_9238,N_9079,N_9131);
or U9239 (N_9239,N_9051,N_9094);
or U9240 (N_9240,N_9167,N_9104);
nand U9241 (N_9241,N_9005,N_9087);
nand U9242 (N_9242,N_9065,N_9076);
or U9243 (N_9243,N_9039,N_9000);
or U9244 (N_9244,N_9084,N_9110);
nor U9245 (N_9245,N_9008,N_9182);
and U9246 (N_9246,N_9057,N_9192);
nand U9247 (N_9247,N_9199,N_9044);
or U9248 (N_9248,N_9141,N_9061);
nor U9249 (N_9249,N_9117,N_9007);
or U9250 (N_9250,N_9185,N_9015);
nor U9251 (N_9251,N_9190,N_9187);
and U9252 (N_9252,N_9055,N_9150);
and U9253 (N_9253,N_9068,N_9026);
nand U9254 (N_9254,N_9135,N_9120);
xnor U9255 (N_9255,N_9171,N_9140);
xnor U9256 (N_9256,N_9113,N_9073);
xor U9257 (N_9257,N_9046,N_9090);
or U9258 (N_9258,N_9098,N_9181);
or U9259 (N_9259,N_9029,N_9060);
nand U9260 (N_9260,N_9089,N_9012);
and U9261 (N_9261,N_9178,N_9080);
xnor U9262 (N_9262,N_9137,N_9126);
xor U9263 (N_9263,N_9097,N_9168);
and U9264 (N_9264,N_9047,N_9164);
nand U9265 (N_9265,N_9145,N_9053);
and U9266 (N_9266,N_9036,N_9108);
or U9267 (N_9267,N_9063,N_9107);
nand U9268 (N_9268,N_9133,N_9096);
or U9269 (N_9269,N_9041,N_9085);
nand U9270 (N_9270,N_9038,N_9101);
or U9271 (N_9271,N_9149,N_9122);
xor U9272 (N_9272,N_9153,N_9077);
nand U9273 (N_9273,N_9009,N_9186);
or U9274 (N_9274,N_9170,N_9048);
nand U9275 (N_9275,N_9172,N_9011);
or U9276 (N_9276,N_9111,N_9056);
and U9277 (N_9277,N_9158,N_9058);
nor U9278 (N_9278,N_9163,N_9020);
xor U9279 (N_9279,N_9143,N_9179);
nor U9280 (N_9280,N_9144,N_9102);
and U9281 (N_9281,N_9128,N_9037);
xnor U9282 (N_9282,N_9124,N_9146);
or U9283 (N_9283,N_9099,N_9024);
nand U9284 (N_9284,N_9115,N_9109);
and U9285 (N_9285,N_9134,N_9031);
nand U9286 (N_9286,N_9193,N_9032);
nor U9287 (N_9287,N_9129,N_9023);
xor U9288 (N_9288,N_9021,N_9013);
or U9289 (N_9289,N_9152,N_9184);
nor U9290 (N_9290,N_9148,N_9003);
nor U9291 (N_9291,N_9155,N_9002);
and U9292 (N_9292,N_9112,N_9114);
and U9293 (N_9293,N_9043,N_9004);
and U9294 (N_9294,N_9196,N_9030);
and U9295 (N_9295,N_9034,N_9130);
nand U9296 (N_9296,N_9071,N_9017);
nand U9297 (N_9297,N_9162,N_9177);
or U9298 (N_9298,N_9070,N_9028);
and U9299 (N_9299,N_9125,N_9100);
xor U9300 (N_9300,N_9050,N_9064);
nor U9301 (N_9301,N_9065,N_9058);
xnor U9302 (N_9302,N_9116,N_9093);
nor U9303 (N_9303,N_9003,N_9066);
nand U9304 (N_9304,N_9088,N_9006);
xor U9305 (N_9305,N_9056,N_9121);
nor U9306 (N_9306,N_9050,N_9134);
nand U9307 (N_9307,N_9130,N_9103);
nor U9308 (N_9308,N_9005,N_9177);
and U9309 (N_9309,N_9113,N_9099);
xnor U9310 (N_9310,N_9068,N_9067);
nor U9311 (N_9311,N_9198,N_9192);
nand U9312 (N_9312,N_9197,N_9050);
nand U9313 (N_9313,N_9019,N_9102);
xor U9314 (N_9314,N_9041,N_9182);
xnor U9315 (N_9315,N_9040,N_9113);
nor U9316 (N_9316,N_9170,N_9008);
or U9317 (N_9317,N_9042,N_9117);
or U9318 (N_9318,N_9015,N_9158);
nor U9319 (N_9319,N_9164,N_9163);
nor U9320 (N_9320,N_9166,N_9082);
nand U9321 (N_9321,N_9098,N_9076);
xor U9322 (N_9322,N_9185,N_9151);
nor U9323 (N_9323,N_9180,N_9045);
nand U9324 (N_9324,N_9045,N_9179);
nand U9325 (N_9325,N_9059,N_9013);
and U9326 (N_9326,N_9114,N_9142);
nand U9327 (N_9327,N_9165,N_9115);
nand U9328 (N_9328,N_9073,N_9008);
and U9329 (N_9329,N_9122,N_9080);
nand U9330 (N_9330,N_9099,N_9180);
nand U9331 (N_9331,N_9075,N_9173);
xnor U9332 (N_9332,N_9197,N_9107);
and U9333 (N_9333,N_9078,N_9147);
or U9334 (N_9334,N_9176,N_9084);
nand U9335 (N_9335,N_9156,N_9199);
xnor U9336 (N_9336,N_9039,N_9121);
or U9337 (N_9337,N_9040,N_9184);
nand U9338 (N_9338,N_9172,N_9040);
nor U9339 (N_9339,N_9055,N_9094);
or U9340 (N_9340,N_9168,N_9068);
nand U9341 (N_9341,N_9040,N_9094);
nand U9342 (N_9342,N_9193,N_9173);
and U9343 (N_9343,N_9016,N_9020);
or U9344 (N_9344,N_9008,N_9101);
nor U9345 (N_9345,N_9047,N_9186);
nand U9346 (N_9346,N_9118,N_9062);
nor U9347 (N_9347,N_9135,N_9128);
nand U9348 (N_9348,N_9010,N_9077);
nor U9349 (N_9349,N_9173,N_9037);
nand U9350 (N_9350,N_9181,N_9184);
or U9351 (N_9351,N_9167,N_9159);
or U9352 (N_9352,N_9119,N_9180);
nor U9353 (N_9353,N_9121,N_9066);
nor U9354 (N_9354,N_9051,N_9181);
or U9355 (N_9355,N_9021,N_9157);
or U9356 (N_9356,N_9096,N_9197);
or U9357 (N_9357,N_9141,N_9148);
nor U9358 (N_9358,N_9153,N_9101);
nor U9359 (N_9359,N_9157,N_9089);
or U9360 (N_9360,N_9091,N_9107);
xor U9361 (N_9361,N_9031,N_9099);
nor U9362 (N_9362,N_9104,N_9091);
or U9363 (N_9363,N_9086,N_9182);
and U9364 (N_9364,N_9145,N_9161);
or U9365 (N_9365,N_9128,N_9166);
or U9366 (N_9366,N_9172,N_9003);
xnor U9367 (N_9367,N_9152,N_9044);
nor U9368 (N_9368,N_9190,N_9063);
nor U9369 (N_9369,N_9149,N_9100);
nor U9370 (N_9370,N_9184,N_9176);
and U9371 (N_9371,N_9071,N_9070);
nor U9372 (N_9372,N_9118,N_9022);
nand U9373 (N_9373,N_9009,N_9129);
nand U9374 (N_9374,N_9056,N_9152);
or U9375 (N_9375,N_9113,N_9162);
nor U9376 (N_9376,N_9129,N_9180);
xnor U9377 (N_9377,N_9025,N_9002);
or U9378 (N_9378,N_9172,N_9197);
xor U9379 (N_9379,N_9064,N_9122);
nand U9380 (N_9380,N_9179,N_9165);
nor U9381 (N_9381,N_9024,N_9124);
nor U9382 (N_9382,N_9060,N_9043);
and U9383 (N_9383,N_9145,N_9118);
nand U9384 (N_9384,N_9186,N_9054);
nand U9385 (N_9385,N_9124,N_9131);
nand U9386 (N_9386,N_9080,N_9184);
nor U9387 (N_9387,N_9067,N_9102);
xor U9388 (N_9388,N_9131,N_9012);
nand U9389 (N_9389,N_9031,N_9019);
xor U9390 (N_9390,N_9192,N_9137);
and U9391 (N_9391,N_9160,N_9042);
xnor U9392 (N_9392,N_9036,N_9035);
and U9393 (N_9393,N_9198,N_9143);
and U9394 (N_9394,N_9077,N_9125);
and U9395 (N_9395,N_9058,N_9061);
nor U9396 (N_9396,N_9189,N_9017);
nor U9397 (N_9397,N_9117,N_9124);
nand U9398 (N_9398,N_9079,N_9152);
and U9399 (N_9399,N_9172,N_9069);
nand U9400 (N_9400,N_9393,N_9255);
xor U9401 (N_9401,N_9341,N_9366);
nand U9402 (N_9402,N_9285,N_9391);
nor U9403 (N_9403,N_9307,N_9305);
or U9404 (N_9404,N_9370,N_9266);
nor U9405 (N_9405,N_9247,N_9236);
xor U9406 (N_9406,N_9258,N_9245);
and U9407 (N_9407,N_9298,N_9371);
nor U9408 (N_9408,N_9268,N_9326);
xor U9409 (N_9409,N_9383,N_9214);
nand U9410 (N_9410,N_9224,N_9287);
xor U9411 (N_9411,N_9382,N_9299);
nand U9412 (N_9412,N_9396,N_9257);
and U9413 (N_9413,N_9328,N_9385);
nand U9414 (N_9414,N_9377,N_9292);
nand U9415 (N_9415,N_9252,N_9388);
and U9416 (N_9416,N_9319,N_9329);
nand U9417 (N_9417,N_9246,N_9306);
xor U9418 (N_9418,N_9264,N_9358);
or U9419 (N_9419,N_9290,N_9270);
or U9420 (N_9420,N_9230,N_9351);
nand U9421 (N_9421,N_9202,N_9233);
xnor U9422 (N_9422,N_9372,N_9229);
or U9423 (N_9423,N_9347,N_9205);
and U9424 (N_9424,N_9283,N_9390);
or U9425 (N_9425,N_9316,N_9309);
and U9426 (N_9426,N_9310,N_9280);
nor U9427 (N_9427,N_9339,N_9267);
or U9428 (N_9428,N_9384,N_9336);
or U9429 (N_9429,N_9303,N_9218);
nand U9430 (N_9430,N_9361,N_9277);
xnor U9431 (N_9431,N_9363,N_9200);
and U9432 (N_9432,N_9362,N_9313);
and U9433 (N_9433,N_9203,N_9220);
nand U9434 (N_9434,N_9387,N_9279);
nand U9435 (N_9435,N_9232,N_9227);
nand U9436 (N_9436,N_9338,N_9308);
nand U9437 (N_9437,N_9201,N_9321);
and U9438 (N_9438,N_9212,N_9373);
and U9439 (N_9439,N_9323,N_9209);
nor U9440 (N_9440,N_9335,N_9248);
or U9441 (N_9441,N_9318,N_9211);
and U9442 (N_9442,N_9282,N_9369);
xor U9443 (N_9443,N_9325,N_9225);
nand U9444 (N_9444,N_9350,N_9356);
and U9445 (N_9445,N_9260,N_9295);
or U9446 (N_9446,N_9273,N_9238);
or U9447 (N_9447,N_9375,N_9251);
or U9448 (N_9448,N_9348,N_9380);
nand U9449 (N_9449,N_9256,N_9253);
xor U9450 (N_9450,N_9226,N_9311);
or U9451 (N_9451,N_9315,N_9330);
or U9452 (N_9452,N_9234,N_9345);
xnor U9453 (N_9453,N_9265,N_9217);
xor U9454 (N_9454,N_9223,N_9337);
and U9455 (N_9455,N_9320,N_9346);
and U9456 (N_9456,N_9300,N_9243);
and U9457 (N_9457,N_9365,N_9357);
nor U9458 (N_9458,N_9322,N_9378);
nand U9459 (N_9459,N_9215,N_9389);
xnor U9460 (N_9460,N_9242,N_9376);
and U9461 (N_9461,N_9239,N_9333);
and U9462 (N_9462,N_9304,N_9340);
and U9463 (N_9463,N_9301,N_9360);
or U9464 (N_9464,N_9219,N_9204);
and U9465 (N_9465,N_9314,N_9222);
and U9466 (N_9466,N_9259,N_9221);
and U9467 (N_9467,N_9284,N_9349);
xnor U9468 (N_9468,N_9216,N_9367);
nand U9469 (N_9469,N_9342,N_9286);
xnor U9470 (N_9470,N_9237,N_9276);
nor U9471 (N_9471,N_9274,N_9208);
and U9472 (N_9472,N_9288,N_9293);
or U9473 (N_9473,N_9381,N_9364);
or U9474 (N_9474,N_9206,N_9359);
nand U9475 (N_9475,N_9317,N_9250);
or U9476 (N_9476,N_9394,N_9291);
xor U9477 (N_9477,N_9261,N_9281);
or U9478 (N_9478,N_9235,N_9302);
xnor U9479 (N_9479,N_9228,N_9324);
nor U9480 (N_9480,N_9353,N_9397);
or U9481 (N_9481,N_9263,N_9374);
xor U9482 (N_9482,N_9240,N_9344);
and U9483 (N_9483,N_9231,N_9278);
nand U9484 (N_9484,N_9210,N_9213);
or U9485 (N_9485,N_9395,N_9352);
nor U9486 (N_9486,N_9354,N_9275);
xor U9487 (N_9487,N_9392,N_9398);
nand U9488 (N_9488,N_9296,N_9262);
and U9489 (N_9489,N_9272,N_9254);
or U9490 (N_9490,N_9334,N_9312);
nand U9491 (N_9491,N_9343,N_9327);
xor U9492 (N_9492,N_9241,N_9271);
nor U9493 (N_9493,N_9294,N_9207);
xnor U9494 (N_9494,N_9297,N_9379);
nor U9495 (N_9495,N_9368,N_9289);
nand U9496 (N_9496,N_9331,N_9269);
nand U9497 (N_9497,N_9399,N_9244);
nand U9498 (N_9498,N_9332,N_9355);
xor U9499 (N_9499,N_9386,N_9249);
or U9500 (N_9500,N_9326,N_9368);
nor U9501 (N_9501,N_9398,N_9240);
and U9502 (N_9502,N_9327,N_9265);
or U9503 (N_9503,N_9313,N_9344);
or U9504 (N_9504,N_9355,N_9242);
or U9505 (N_9505,N_9249,N_9347);
or U9506 (N_9506,N_9302,N_9211);
or U9507 (N_9507,N_9294,N_9203);
xor U9508 (N_9508,N_9321,N_9323);
xnor U9509 (N_9509,N_9385,N_9314);
nor U9510 (N_9510,N_9336,N_9214);
or U9511 (N_9511,N_9258,N_9342);
nor U9512 (N_9512,N_9229,N_9337);
and U9513 (N_9513,N_9203,N_9215);
or U9514 (N_9514,N_9383,N_9236);
and U9515 (N_9515,N_9360,N_9346);
nor U9516 (N_9516,N_9372,N_9358);
nand U9517 (N_9517,N_9327,N_9315);
and U9518 (N_9518,N_9234,N_9383);
nor U9519 (N_9519,N_9385,N_9208);
xnor U9520 (N_9520,N_9385,N_9370);
and U9521 (N_9521,N_9277,N_9264);
xnor U9522 (N_9522,N_9362,N_9331);
nor U9523 (N_9523,N_9265,N_9307);
nand U9524 (N_9524,N_9284,N_9325);
nand U9525 (N_9525,N_9370,N_9357);
or U9526 (N_9526,N_9388,N_9276);
nor U9527 (N_9527,N_9310,N_9350);
nor U9528 (N_9528,N_9249,N_9353);
nand U9529 (N_9529,N_9299,N_9296);
and U9530 (N_9530,N_9211,N_9258);
and U9531 (N_9531,N_9328,N_9361);
xor U9532 (N_9532,N_9309,N_9332);
xor U9533 (N_9533,N_9305,N_9366);
or U9534 (N_9534,N_9287,N_9278);
nand U9535 (N_9535,N_9318,N_9376);
xor U9536 (N_9536,N_9316,N_9260);
nand U9537 (N_9537,N_9397,N_9243);
and U9538 (N_9538,N_9356,N_9217);
xnor U9539 (N_9539,N_9278,N_9318);
or U9540 (N_9540,N_9316,N_9399);
nand U9541 (N_9541,N_9273,N_9224);
nor U9542 (N_9542,N_9286,N_9259);
xor U9543 (N_9543,N_9387,N_9243);
nor U9544 (N_9544,N_9235,N_9389);
and U9545 (N_9545,N_9297,N_9211);
nand U9546 (N_9546,N_9230,N_9228);
xnor U9547 (N_9547,N_9220,N_9235);
nor U9548 (N_9548,N_9219,N_9269);
nand U9549 (N_9549,N_9398,N_9243);
nor U9550 (N_9550,N_9313,N_9293);
nand U9551 (N_9551,N_9268,N_9329);
or U9552 (N_9552,N_9262,N_9280);
xnor U9553 (N_9553,N_9324,N_9251);
nor U9554 (N_9554,N_9343,N_9288);
or U9555 (N_9555,N_9305,N_9219);
nor U9556 (N_9556,N_9396,N_9383);
nor U9557 (N_9557,N_9240,N_9337);
and U9558 (N_9558,N_9282,N_9233);
and U9559 (N_9559,N_9271,N_9322);
xor U9560 (N_9560,N_9340,N_9338);
xnor U9561 (N_9561,N_9397,N_9272);
nor U9562 (N_9562,N_9358,N_9346);
and U9563 (N_9563,N_9263,N_9341);
and U9564 (N_9564,N_9264,N_9374);
or U9565 (N_9565,N_9376,N_9295);
nand U9566 (N_9566,N_9205,N_9344);
nand U9567 (N_9567,N_9289,N_9297);
and U9568 (N_9568,N_9229,N_9309);
xor U9569 (N_9569,N_9371,N_9287);
nand U9570 (N_9570,N_9351,N_9355);
and U9571 (N_9571,N_9386,N_9381);
and U9572 (N_9572,N_9269,N_9234);
nand U9573 (N_9573,N_9399,N_9257);
or U9574 (N_9574,N_9356,N_9337);
nand U9575 (N_9575,N_9371,N_9324);
nor U9576 (N_9576,N_9289,N_9274);
and U9577 (N_9577,N_9326,N_9353);
xnor U9578 (N_9578,N_9306,N_9238);
and U9579 (N_9579,N_9244,N_9236);
nand U9580 (N_9580,N_9245,N_9203);
xnor U9581 (N_9581,N_9381,N_9377);
and U9582 (N_9582,N_9356,N_9341);
nand U9583 (N_9583,N_9268,N_9352);
nand U9584 (N_9584,N_9237,N_9323);
xor U9585 (N_9585,N_9241,N_9212);
nor U9586 (N_9586,N_9353,N_9388);
and U9587 (N_9587,N_9304,N_9336);
nand U9588 (N_9588,N_9257,N_9263);
and U9589 (N_9589,N_9340,N_9380);
nand U9590 (N_9590,N_9232,N_9332);
nor U9591 (N_9591,N_9252,N_9323);
or U9592 (N_9592,N_9398,N_9280);
or U9593 (N_9593,N_9344,N_9280);
nand U9594 (N_9594,N_9357,N_9267);
nand U9595 (N_9595,N_9336,N_9367);
and U9596 (N_9596,N_9344,N_9356);
xnor U9597 (N_9597,N_9314,N_9211);
xor U9598 (N_9598,N_9239,N_9288);
nor U9599 (N_9599,N_9242,N_9297);
nand U9600 (N_9600,N_9518,N_9537);
nor U9601 (N_9601,N_9573,N_9580);
or U9602 (N_9602,N_9487,N_9429);
and U9603 (N_9603,N_9508,N_9426);
or U9604 (N_9604,N_9574,N_9484);
xnor U9605 (N_9605,N_9445,N_9486);
nor U9606 (N_9606,N_9504,N_9497);
or U9607 (N_9607,N_9461,N_9506);
and U9608 (N_9608,N_9581,N_9453);
xnor U9609 (N_9609,N_9400,N_9452);
or U9610 (N_9610,N_9407,N_9565);
nand U9611 (N_9611,N_9469,N_9468);
xnor U9612 (N_9612,N_9414,N_9410);
xor U9613 (N_9613,N_9440,N_9511);
xor U9614 (N_9614,N_9417,N_9491);
xor U9615 (N_9615,N_9462,N_9542);
nand U9616 (N_9616,N_9431,N_9442);
xor U9617 (N_9617,N_9424,N_9454);
nor U9618 (N_9618,N_9599,N_9411);
nor U9619 (N_9619,N_9568,N_9570);
and U9620 (N_9620,N_9524,N_9436);
nor U9621 (N_9621,N_9510,N_9513);
nand U9622 (N_9622,N_9408,N_9529);
nor U9623 (N_9623,N_9561,N_9433);
nand U9624 (N_9624,N_9585,N_9463);
nand U9625 (N_9625,N_9413,N_9479);
xnor U9626 (N_9626,N_9582,N_9578);
xnor U9627 (N_9627,N_9488,N_9465);
and U9628 (N_9628,N_9552,N_9548);
nor U9629 (N_9629,N_9447,N_9525);
and U9630 (N_9630,N_9430,N_9406);
and U9631 (N_9631,N_9512,N_9412);
or U9632 (N_9632,N_9450,N_9477);
nor U9633 (N_9633,N_9594,N_9528);
xnor U9634 (N_9634,N_9534,N_9519);
nand U9635 (N_9635,N_9522,N_9490);
or U9636 (N_9636,N_9423,N_9457);
and U9637 (N_9637,N_9416,N_9472);
and U9638 (N_9638,N_9434,N_9421);
nor U9639 (N_9639,N_9405,N_9509);
nand U9640 (N_9640,N_9569,N_9559);
and U9641 (N_9641,N_9485,N_9443);
xnor U9642 (N_9642,N_9562,N_9418);
and U9643 (N_9643,N_9514,N_9590);
xor U9644 (N_9644,N_9535,N_9517);
nand U9645 (N_9645,N_9481,N_9455);
and U9646 (N_9646,N_9547,N_9532);
xor U9647 (N_9647,N_9571,N_9500);
nand U9648 (N_9648,N_9476,N_9498);
nand U9649 (N_9649,N_9464,N_9543);
nor U9650 (N_9650,N_9438,N_9567);
or U9651 (N_9651,N_9576,N_9493);
and U9652 (N_9652,N_9446,N_9495);
or U9653 (N_9653,N_9483,N_9587);
xnor U9654 (N_9654,N_9432,N_9520);
xnor U9655 (N_9655,N_9589,N_9536);
or U9656 (N_9656,N_9415,N_9557);
or U9657 (N_9657,N_9563,N_9460);
nand U9658 (N_9658,N_9550,N_9456);
xor U9659 (N_9659,N_9502,N_9404);
or U9660 (N_9660,N_9556,N_9503);
nor U9661 (N_9661,N_9546,N_9471);
xor U9662 (N_9662,N_9419,N_9592);
or U9663 (N_9663,N_9523,N_9551);
nand U9664 (N_9664,N_9521,N_9588);
nand U9665 (N_9665,N_9494,N_9409);
nor U9666 (N_9666,N_9473,N_9449);
nor U9667 (N_9667,N_9475,N_9467);
and U9668 (N_9668,N_9597,N_9584);
xnor U9669 (N_9669,N_9577,N_9437);
and U9670 (N_9670,N_9402,N_9501);
xnor U9671 (N_9671,N_9526,N_9586);
nor U9672 (N_9672,N_9593,N_9598);
nand U9673 (N_9673,N_9505,N_9527);
nand U9674 (N_9674,N_9480,N_9572);
xor U9675 (N_9675,N_9444,N_9596);
nor U9676 (N_9676,N_9507,N_9544);
nand U9677 (N_9677,N_9427,N_9553);
xor U9678 (N_9678,N_9470,N_9541);
xnor U9679 (N_9679,N_9558,N_9560);
or U9680 (N_9680,N_9591,N_9458);
and U9681 (N_9681,N_9439,N_9420);
xor U9682 (N_9682,N_9545,N_9482);
xnor U9683 (N_9683,N_9435,N_9401);
nand U9684 (N_9684,N_9533,N_9549);
and U9685 (N_9685,N_9539,N_9489);
nor U9686 (N_9686,N_9466,N_9575);
and U9687 (N_9687,N_9441,N_9451);
xor U9688 (N_9688,N_9492,N_9531);
nand U9689 (N_9689,N_9425,N_9538);
xnor U9690 (N_9690,N_9595,N_9403);
xnor U9691 (N_9691,N_9474,N_9540);
or U9692 (N_9692,N_9530,N_9459);
or U9693 (N_9693,N_9516,N_9579);
nor U9694 (N_9694,N_9554,N_9566);
xnor U9695 (N_9695,N_9496,N_9515);
and U9696 (N_9696,N_9555,N_9583);
or U9697 (N_9697,N_9428,N_9448);
nor U9698 (N_9698,N_9564,N_9478);
nand U9699 (N_9699,N_9422,N_9499);
or U9700 (N_9700,N_9507,N_9417);
and U9701 (N_9701,N_9560,N_9413);
or U9702 (N_9702,N_9492,N_9541);
nand U9703 (N_9703,N_9431,N_9596);
nor U9704 (N_9704,N_9419,N_9586);
nor U9705 (N_9705,N_9583,N_9528);
nand U9706 (N_9706,N_9411,N_9452);
nand U9707 (N_9707,N_9476,N_9489);
nand U9708 (N_9708,N_9493,N_9442);
or U9709 (N_9709,N_9537,N_9506);
nand U9710 (N_9710,N_9553,N_9505);
or U9711 (N_9711,N_9421,N_9570);
nor U9712 (N_9712,N_9521,N_9443);
or U9713 (N_9713,N_9461,N_9537);
nor U9714 (N_9714,N_9553,N_9484);
xor U9715 (N_9715,N_9448,N_9528);
and U9716 (N_9716,N_9493,N_9591);
nand U9717 (N_9717,N_9577,N_9488);
nor U9718 (N_9718,N_9559,N_9552);
nand U9719 (N_9719,N_9412,N_9555);
or U9720 (N_9720,N_9470,N_9423);
or U9721 (N_9721,N_9435,N_9433);
or U9722 (N_9722,N_9437,N_9435);
nand U9723 (N_9723,N_9417,N_9497);
nor U9724 (N_9724,N_9429,N_9505);
xnor U9725 (N_9725,N_9549,N_9544);
nand U9726 (N_9726,N_9457,N_9500);
nor U9727 (N_9727,N_9465,N_9420);
or U9728 (N_9728,N_9488,N_9517);
nor U9729 (N_9729,N_9529,N_9511);
nand U9730 (N_9730,N_9580,N_9429);
nand U9731 (N_9731,N_9449,N_9500);
and U9732 (N_9732,N_9538,N_9594);
and U9733 (N_9733,N_9564,N_9524);
nand U9734 (N_9734,N_9510,N_9590);
nand U9735 (N_9735,N_9548,N_9512);
and U9736 (N_9736,N_9551,N_9512);
xor U9737 (N_9737,N_9508,N_9558);
nand U9738 (N_9738,N_9593,N_9445);
or U9739 (N_9739,N_9576,N_9444);
nand U9740 (N_9740,N_9475,N_9599);
nor U9741 (N_9741,N_9482,N_9581);
nor U9742 (N_9742,N_9551,N_9479);
xor U9743 (N_9743,N_9557,N_9594);
or U9744 (N_9744,N_9569,N_9557);
or U9745 (N_9745,N_9445,N_9583);
and U9746 (N_9746,N_9448,N_9450);
nand U9747 (N_9747,N_9582,N_9412);
xnor U9748 (N_9748,N_9515,N_9509);
nor U9749 (N_9749,N_9413,N_9570);
xor U9750 (N_9750,N_9428,N_9558);
nand U9751 (N_9751,N_9436,N_9414);
nand U9752 (N_9752,N_9561,N_9402);
nor U9753 (N_9753,N_9539,N_9403);
nand U9754 (N_9754,N_9595,N_9520);
or U9755 (N_9755,N_9515,N_9517);
nor U9756 (N_9756,N_9416,N_9584);
nand U9757 (N_9757,N_9526,N_9536);
and U9758 (N_9758,N_9531,N_9498);
xor U9759 (N_9759,N_9590,N_9490);
nand U9760 (N_9760,N_9591,N_9544);
and U9761 (N_9761,N_9417,N_9582);
xor U9762 (N_9762,N_9492,N_9475);
or U9763 (N_9763,N_9407,N_9451);
or U9764 (N_9764,N_9482,N_9532);
and U9765 (N_9765,N_9586,N_9444);
and U9766 (N_9766,N_9594,N_9404);
xor U9767 (N_9767,N_9564,N_9578);
nand U9768 (N_9768,N_9435,N_9467);
nand U9769 (N_9769,N_9420,N_9534);
nor U9770 (N_9770,N_9445,N_9476);
nand U9771 (N_9771,N_9412,N_9428);
xnor U9772 (N_9772,N_9446,N_9482);
nand U9773 (N_9773,N_9416,N_9506);
nand U9774 (N_9774,N_9496,N_9512);
nor U9775 (N_9775,N_9456,N_9544);
or U9776 (N_9776,N_9457,N_9519);
nand U9777 (N_9777,N_9429,N_9436);
and U9778 (N_9778,N_9504,N_9540);
xnor U9779 (N_9779,N_9488,N_9400);
xnor U9780 (N_9780,N_9513,N_9562);
nor U9781 (N_9781,N_9447,N_9411);
nand U9782 (N_9782,N_9466,N_9598);
nand U9783 (N_9783,N_9416,N_9460);
nand U9784 (N_9784,N_9444,N_9565);
xor U9785 (N_9785,N_9580,N_9507);
nor U9786 (N_9786,N_9561,N_9596);
nand U9787 (N_9787,N_9545,N_9500);
or U9788 (N_9788,N_9521,N_9519);
nor U9789 (N_9789,N_9546,N_9508);
xnor U9790 (N_9790,N_9528,N_9582);
and U9791 (N_9791,N_9510,N_9538);
nand U9792 (N_9792,N_9473,N_9569);
or U9793 (N_9793,N_9499,N_9458);
or U9794 (N_9794,N_9460,N_9516);
or U9795 (N_9795,N_9541,N_9447);
xor U9796 (N_9796,N_9533,N_9467);
xor U9797 (N_9797,N_9426,N_9592);
nor U9798 (N_9798,N_9545,N_9478);
and U9799 (N_9799,N_9452,N_9587);
xor U9800 (N_9800,N_9650,N_9628);
xnor U9801 (N_9801,N_9648,N_9743);
nand U9802 (N_9802,N_9621,N_9731);
and U9803 (N_9803,N_9709,N_9687);
nor U9804 (N_9804,N_9735,N_9613);
or U9805 (N_9805,N_9758,N_9614);
and U9806 (N_9806,N_9636,N_9702);
or U9807 (N_9807,N_9633,N_9671);
or U9808 (N_9808,N_9639,N_9718);
and U9809 (N_9809,N_9798,N_9646);
nor U9810 (N_9810,N_9723,N_9658);
or U9811 (N_9811,N_9789,N_9770);
and U9812 (N_9812,N_9739,N_9727);
or U9813 (N_9813,N_9662,N_9710);
and U9814 (N_9814,N_9726,N_9750);
nand U9815 (N_9815,N_9787,N_9734);
nand U9816 (N_9816,N_9752,N_9763);
nor U9817 (N_9817,N_9657,N_9655);
or U9818 (N_9818,N_9607,N_9696);
and U9819 (N_9819,N_9707,N_9720);
nand U9820 (N_9820,N_9721,N_9701);
and U9821 (N_9821,N_9651,N_9623);
or U9822 (N_9822,N_9654,N_9790);
xnor U9823 (N_9823,N_9774,N_9794);
nor U9824 (N_9824,N_9793,N_9730);
nor U9825 (N_9825,N_9716,N_9757);
nor U9826 (N_9826,N_9737,N_9796);
and U9827 (N_9827,N_9729,N_9640);
nor U9828 (N_9828,N_9698,N_9629);
nand U9829 (N_9829,N_9622,N_9783);
xnor U9830 (N_9830,N_9781,N_9767);
nand U9831 (N_9831,N_9602,N_9732);
and U9832 (N_9832,N_9736,N_9711);
nor U9833 (N_9833,N_9765,N_9616);
xor U9834 (N_9834,N_9766,N_9667);
and U9835 (N_9835,N_9652,N_9680);
and U9836 (N_9836,N_9620,N_9756);
or U9837 (N_9837,N_9780,N_9626);
nand U9838 (N_9838,N_9769,N_9631);
and U9839 (N_9839,N_9638,N_9659);
nor U9840 (N_9840,N_9773,N_9666);
or U9841 (N_9841,N_9605,N_9738);
or U9842 (N_9842,N_9786,N_9691);
nor U9843 (N_9843,N_9797,N_9719);
nand U9844 (N_9844,N_9768,N_9660);
and U9845 (N_9845,N_9603,N_9608);
nand U9846 (N_9846,N_9784,N_9697);
and U9847 (N_9847,N_9664,N_9725);
or U9848 (N_9848,N_9647,N_9625);
xor U9849 (N_9849,N_9703,N_9741);
or U9850 (N_9850,N_9776,N_9692);
nor U9851 (N_9851,N_9779,N_9717);
or U9852 (N_9852,N_9627,N_9791);
nand U9853 (N_9853,N_9751,N_9624);
and U9854 (N_9854,N_9744,N_9615);
nand U9855 (N_9855,N_9740,N_9759);
nand U9856 (N_9856,N_9618,N_9782);
nor U9857 (N_9857,N_9683,N_9665);
xor U9858 (N_9858,N_9699,N_9641);
nand U9859 (N_9859,N_9749,N_9611);
xnor U9860 (N_9860,N_9748,N_9601);
nand U9861 (N_9861,N_9661,N_9728);
nand U9862 (N_9862,N_9674,N_9742);
and U9863 (N_9863,N_9637,N_9753);
nand U9864 (N_9864,N_9775,N_9693);
and U9865 (N_9865,N_9619,N_9676);
nor U9866 (N_9866,N_9681,N_9672);
nand U9867 (N_9867,N_9649,N_9713);
and U9868 (N_9868,N_9706,N_9788);
nor U9869 (N_9869,N_9606,N_9760);
nand U9870 (N_9870,N_9670,N_9690);
and U9871 (N_9871,N_9771,N_9792);
xnor U9872 (N_9872,N_9630,N_9678);
nand U9873 (N_9873,N_9610,N_9604);
xor U9874 (N_9874,N_9634,N_9612);
or U9875 (N_9875,N_9686,N_9632);
nor U9876 (N_9876,N_9609,N_9673);
nor U9877 (N_9877,N_9745,N_9764);
nand U9878 (N_9878,N_9677,N_9714);
and U9879 (N_9879,N_9715,N_9635);
nand U9880 (N_9880,N_9695,N_9675);
nor U9881 (N_9881,N_9704,N_9755);
nor U9882 (N_9882,N_9795,N_9722);
nand U9883 (N_9883,N_9747,N_9600);
xor U9884 (N_9884,N_9679,N_9724);
nor U9885 (N_9885,N_9668,N_9645);
and U9886 (N_9886,N_9746,N_9669);
nand U9887 (N_9887,N_9785,N_9733);
nand U9888 (N_9888,N_9682,N_9689);
or U9889 (N_9889,N_9772,N_9663);
and U9890 (N_9890,N_9777,N_9656);
and U9891 (N_9891,N_9653,N_9700);
nand U9892 (N_9892,N_9684,N_9644);
xnor U9893 (N_9893,N_9762,N_9685);
nor U9894 (N_9894,N_9643,N_9708);
and U9895 (N_9895,N_9761,N_9799);
nand U9896 (N_9896,N_9712,N_9705);
or U9897 (N_9897,N_9642,N_9688);
nand U9898 (N_9898,N_9754,N_9778);
and U9899 (N_9899,N_9617,N_9694);
nor U9900 (N_9900,N_9678,N_9638);
and U9901 (N_9901,N_9785,N_9723);
or U9902 (N_9902,N_9684,N_9756);
and U9903 (N_9903,N_9797,N_9753);
xor U9904 (N_9904,N_9797,N_9609);
nand U9905 (N_9905,N_9728,N_9609);
or U9906 (N_9906,N_9763,N_9772);
nand U9907 (N_9907,N_9611,N_9753);
xor U9908 (N_9908,N_9750,N_9754);
and U9909 (N_9909,N_9692,N_9637);
and U9910 (N_9910,N_9657,N_9632);
or U9911 (N_9911,N_9648,N_9697);
xnor U9912 (N_9912,N_9675,N_9736);
and U9913 (N_9913,N_9650,N_9793);
and U9914 (N_9914,N_9641,N_9763);
nand U9915 (N_9915,N_9718,N_9618);
and U9916 (N_9916,N_9691,N_9695);
and U9917 (N_9917,N_9744,N_9645);
and U9918 (N_9918,N_9765,N_9775);
nor U9919 (N_9919,N_9789,N_9643);
or U9920 (N_9920,N_9784,N_9610);
xor U9921 (N_9921,N_9684,N_9610);
nand U9922 (N_9922,N_9725,N_9603);
and U9923 (N_9923,N_9608,N_9604);
nor U9924 (N_9924,N_9614,N_9772);
and U9925 (N_9925,N_9795,N_9656);
nand U9926 (N_9926,N_9793,N_9797);
xnor U9927 (N_9927,N_9698,N_9644);
and U9928 (N_9928,N_9754,N_9664);
xnor U9929 (N_9929,N_9635,N_9662);
or U9930 (N_9930,N_9679,N_9760);
nand U9931 (N_9931,N_9789,N_9727);
xor U9932 (N_9932,N_9750,N_9707);
nor U9933 (N_9933,N_9778,N_9737);
nand U9934 (N_9934,N_9667,N_9754);
nor U9935 (N_9935,N_9619,N_9785);
or U9936 (N_9936,N_9630,N_9717);
xor U9937 (N_9937,N_9790,N_9763);
and U9938 (N_9938,N_9750,N_9609);
and U9939 (N_9939,N_9722,N_9785);
xor U9940 (N_9940,N_9787,N_9795);
and U9941 (N_9941,N_9620,N_9678);
or U9942 (N_9942,N_9793,N_9739);
or U9943 (N_9943,N_9605,N_9706);
nor U9944 (N_9944,N_9709,N_9650);
and U9945 (N_9945,N_9711,N_9653);
nand U9946 (N_9946,N_9780,N_9749);
or U9947 (N_9947,N_9736,N_9790);
and U9948 (N_9948,N_9717,N_9751);
xor U9949 (N_9949,N_9641,N_9785);
or U9950 (N_9950,N_9792,N_9791);
and U9951 (N_9951,N_9697,N_9702);
nand U9952 (N_9952,N_9668,N_9692);
nor U9953 (N_9953,N_9652,N_9783);
and U9954 (N_9954,N_9755,N_9753);
nor U9955 (N_9955,N_9675,N_9708);
nor U9956 (N_9956,N_9763,N_9610);
xnor U9957 (N_9957,N_9677,N_9704);
nand U9958 (N_9958,N_9663,N_9764);
or U9959 (N_9959,N_9636,N_9706);
or U9960 (N_9960,N_9734,N_9683);
nand U9961 (N_9961,N_9625,N_9612);
or U9962 (N_9962,N_9652,N_9653);
nand U9963 (N_9963,N_9761,N_9650);
nand U9964 (N_9964,N_9638,N_9669);
xor U9965 (N_9965,N_9646,N_9635);
nor U9966 (N_9966,N_9679,N_9628);
or U9967 (N_9967,N_9641,N_9646);
or U9968 (N_9968,N_9751,N_9696);
or U9969 (N_9969,N_9685,N_9654);
or U9970 (N_9970,N_9776,N_9777);
and U9971 (N_9971,N_9637,N_9786);
nor U9972 (N_9972,N_9798,N_9768);
xor U9973 (N_9973,N_9790,N_9626);
xnor U9974 (N_9974,N_9737,N_9791);
xnor U9975 (N_9975,N_9751,N_9745);
and U9976 (N_9976,N_9672,N_9666);
xor U9977 (N_9977,N_9723,N_9746);
nand U9978 (N_9978,N_9628,N_9617);
nand U9979 (N_9979,N_9616,N_9702);
and U9980 (N_9980,N_9742,N_9605);
xnor U9981 (N_9981,N_9792,N_9674);
nand U9982 (N_9982,N_9641,N_9634);
xor U9983 (N_9983,N_9626,N_9676);
and U9984 (N_9984,N_9783,N_9757);
nor U9985 (N_9985,N_9608,N_9622);
nand U9986 (N_9986,N_9663,N_9767);
and U9987 (N_9987,N_9746,N_9674);
and U9988 (N_9988,N_9699,N_9647);
nand U9989 (N_9989,N_9710,N_9672);
xnor U9990 (N_9990,N_9712,N_9645);
or U9991 (N_9991,N_9784,N_9667);
or U9992 (N_9992,N_9780,N_9714);
nor U9993 (N_9993,N_9707,N_9613);
nor U9994 (N_9994,N_9788,N_9643);
xnor U9995 (N_9995,N_9766,N_9797);
xnor U9996 (N_9996,N_9660,N_9624);
and U9997 (N_9997,N_9733,N_9741);
nand U9998 (N_9998,N_9729,N_9750);
nand U9999 (N_9999,N_9781,N_9736);
xor U10000 (N_10000,N_9943,N_9886);
and U10001 (N_10001,N_9990,N_9849);
and U10002 (N_10002,N_9970,N_9958);
or U10003 (N_10003,N_9848,N_9927);
or U10004 (N_10004,N_9835,N_9864);
nor U10005 (N_10005,N_9800,N_9862);
nor U10006 (N_10006,N_9861,N_9998);
xnor U10007 (N_10007,N_9865,N_9814);
xnor U10008 (N_10008,N_9857,N_9962);
nand U10009 (N_10009,N_9887,N_9807);
xor U10010 (N_10010,N_9893,N_9982);
xnor U10011 (N_10011,N_9965,N_9853);
and U10012 (N_10012,N_9838,N_9996);
nor U10013 (N_10013,N_9922,N_9926);
or U10014 (N_10014,N_9819,N_9892);
or U10015 (N_10015,N_9846,N_9878);
and U10016 (N_10016,N_9916,N_9841);
and U10017 (N_10017,N_9812,N_9872);
and U10018 (N_10018,N_9948,N_9946);
or U10019 (N_10019,N_9815,N_9899);
nand U10020 (N_10020,N_9909,N_9975);
nor U10021 (N_10021,N_9842,N_9830);
or U10022 (N_10022,N_9947,N_9906);
nor U10023 (N_10023,N_9908,N_9900);
and U10024 (N_10024,N_9968,N_9960);
and U10025 (N_10025,N_9974,N_9873);
nand U10026 (N_10026,N_9839,N_9804);
nor U10027 (N_10027,N_9999,N_9959);
xnor U10028 (N_10028,N_9997,N_9805);
xor U10029 (N_10029,N_9869,N_9847);
nand U10030 (N_10030,N_9833,N_9858);
nor U10031 (N_10031,N_9986,N_9897);
nor U10032 (N_10032,N_9816,N_9994);
and U10033 (N_10033,N_9874,N_9939);
nand U10034 (N_10034,N_9931,N_9910);
and U10035 (N_10035,N_9980,N_9844);
nand U10036 (N_10036,N_9942,N_9941);
nand U10037 (N_10037,N_9920,N_9914);
nand U10038 (N_10038,N_9981,N_9876);
xnor U10039 (N_10039,N_9905,N_9966);
nand U10040 (N_10040,N_9810,N_9852);
or U10041 (N_10041,N_9924,N_9850);
nand U10042 (N_10042,N_9978,N_9933);
nor U10043 (N_10043,N_9930,N_9915);
or U10044 (N_10044,N_9949,N_9825);
and U10045 (N_10045,N_9851,N_9928);
and U10046 (N_10046,N_9832,N_9936);
and U10047 (N_10047,N_9976,N_9856);
xor U10048 (N_10048,N_9984,N_9871);
xor U10049 (N_10049,N_9964,N_9836);
or U10050 (N_10050,N_9956,N_9827);
xor U10051 (N_10051,N_9803,N_9967);
nand U10052 (N_10052,N_9884,N_9891);
and U10053 (N_10053,N_9988,N_9813);
or U10054 (N_10054,N_9954,N_9888);
nor U10055 (N_10055,N_9937,N_9961);
and U10056 (N_10056,N_9957,N_9823);
xor U10057 (N_10057,N_9889,N_9902);
or U10058 (N_10058,N_9896,N_9829);
nor U10059 (N_10059,N_9863,N_9929);
nand U10060 (N_10060,N_9995,N_9843);
nand U10061 (N_10061,N_9867,N_9881);
xnor U10062 (N_10062,N_9882,N_9987);
nand U10063 (N_10063,N_9808,N_9894);
or U10064 (N_10064,N_9854,N_9880);
and U10065 (N_10065,N_9925,N_9883);
or U10066 (N_10066,N_9870,N_9877);
or U10067 (N_10067,N_9875,N_9879);
xor U10068 (N_10068,N_9971,N_9821);
nand U10069 (N_10069,N_9932,N_9903);
and U10070 (N_10070,N_9945,N_9921);
xor U10071 (N_10071,N_9963,N_9989);
and U10072 (N_10072,N_9972,N_9952);
nor U10073 (N_10073,N_9923,N_9826);
nand U10074 (N_10074,N_9919,N_9901);
and U10075 (N_10075,N_9944,N_9811);
nand U10076 (N_10076,N_9969,N_9890);
nor U10077 (N_10077,N_9904,N_9831);
xor U10078 (N_10078,N_9860,N_9845);
and U10079 (N_10079,N_9912,N_9977);
and U10080 (N_10080,N_9820,N_9824);
nor U10081 (N_10081,N_9985,N_9951);
nand U10082 (N_10082,N_9898,N_9822);
nand U10083 (N_10083,N_9868,N_9991);
nor U10084 (N_10084,N_9913,N_9802);
nor U10085 (N_10085,N_9953,N_9828);
xor U10086 (N_10086,N_9934,N_9917);
or U10087 (N_10087,N_9973,N_9950);
and U10088 (N_10088,N_9818,N_9938);
nor U10089 (N_10089,N_9955,N_9840);
nand U10090 (N_10090,N_9801,N_9979);
nor U10091 (N_10091,N_9993,N_9983);
and U10092 (N_10092,N_9935,N_9809);
or U10093 (N_10093,N_9834,N_9817);
nand U10094 (N_10094,N_9911,N_9866);
and U10095 (N_10095,N_9895,N_9907);
xnor U10096 (N_10096,N_9940,N_9855);
and U10097 (N_10097,N_9992,N_9918);
and U10098 (N_10098,N_9885,N_9859);
and U10099 (N_10099,N_9806,N_9837);
and U10100 (N_10100,N_9944,N_9852);
xnor U10101 (N_10101,N_9805,N_9941);
nor U10102 (N_10102,N_9933,N_9848);
nand U10103 (N_10103,N_9862,N_9972);
xor U10104 (N_10104,N_9842,N_9888);
xor U10105 (N_10105,N_9895,N_9801);
nand U10106 (N_10106,N_9915,N_9985);
nand U10107 (N_10107,N_9918,N_9964);
or U10108 (N_10108,N_9867,N_9981);
xnor U10109 (N_10109,N_9931,N_9875);
nor U10110 (N_10110,N_9975,N_9927);
or U10111 (N_10111,N_9865,N_9988);
nand U10112 (N_10112,N_9995,N_9879);
and U10113 (N_10113,N_9880,N_9877);
nor U10114 (N_10114,N_9903,N_9823);
or U10115 (N_10115,N_9863,N_9989);
nand U10116 (N_10116,N_9913,N_9806);
nand U10117 (N_10117,N_9957,N_9971);
nor U10118 (N_10118,N_9958,N_9903);
and U10119 (N_10119,N_9803,N_9801);
and U10120 (N_10120,N_9846,N_9997);
xnor U10121 (N_10121,N_9858,N_9874);
and U10122 (N_10122,N_9938,N_9808);
or U10123 (N_10123,N_9910,N_9995);
xor U10124 (N_10124,N_9978,N_9875);
and U10125 (N_10125,N_9964,N_9986);
nor U10126 (N_10126,N_9817,N_9811);
xor U10127 (N_10127,N_9989,N_9810);
nor U10128 (N_10128,N_9841,N_9839);
nand U10129 (N_10129,N_9884,N_9951);
or U10130 (N_10130,N_9916,N_9970);
and U10131 (N_10131,N_9850,N_9883);
and U10132 (N_10132,N_9957,N_9937);
xnor U10133 (N_10133,N_9952,N_9881);
nand U10134 (N_10134,N_9902,N_9850);
nand U10135 (N_10135,N_9817,N_9846);
and U10136 (N_10136,N_9954,N_9846);
nand U10137 (N_10137,N_9850,N_9939);
nand U10138 (N_10138,N_9874,N_9918);
nand U10139 (N_10139,N_9845,N_9984);
nand U10140 (N_10140,N_9979,N_9915);
nand U10141 (N_10141,N_9843,N_9885);
or U10142 (N_10142,N_9933,N_9814);
xnor U10143 (N_10143,N_9917,N_9806);
or U10144 (N_10144,N_9848,N_9891);
nand U10145 (N_10145,N_9898,N_9805);
xnor U10146 (N_10146,N_9802,N_9878);
nor U10147 (N_10147,N_9871,N_9811);
and U10148 (N_10148,N_9929,N_9838);
nor U10149 (N_10149,N_9983,N_9973);
or U10150 (N_10150,N_9911,N_9920);
xor U10151 (N_10151,N_9932,N_9832);
nand U10152 (N_10152,N_9935,N_9993);
nand U10153 (N_10153,N_9886,N_9912);
nor U10154 (N_10154,N_9800,N_9866);
nand U10155 (N_10155,N_9920,N_9957);
xnor U10156 (N_10156,N_9970,N_9866);
or U10157 (N_10157,N_9808,N_9941);
or U10158 (N_10158,N_9898,N_9836);
nor U10159 (N_10159,N_9816,N_9895);
nor U10160 (N_10160,N_9810,N_9861);
and U10161 (N_10161,N_9806,N_9984);
nand U10162 (N_10162,N_9865,N_9931);
xor U10163 (N_10163,N_9969,N_9841);
nor U10164 (N_10164,N_9811,N_9837);
nand U10165 (N_10165,N_9981,N_9995);
or U10166 (N_10166,N_9878,N_9831);
or U10167 (N_10167,N_9969,N_9891);
nand U10168 (N_10168,N_9962,N_9921);
and U10169 (N_10169,N_9855,N_9886);
nand U10170 (N_10170,N_9974,N_9864);
nand U10171 (N_10171,N_9904,N_9956);
or U10172 (N_10172,N_9844,N_9862);
xnor U10173 (N_10173,N_9907,N_9847);
nand U10174 (N_10174,N_9921,N_9865);
nor U10175 (N_10175,N_9928,N_9907);
nor U10176 (N_10176,N_9894,N_9835);
or U10177 (N_10177,N_9973,N_9991);
and U10178 (N_10178,N_9901,N_9979);
nor U10179 (N_10179,N_9938,N_9804);
or U10180 (N_10180,N_9862,N_9880);
nor U10181 (N_10181,N_9937,N_9878);
nand U10182 (N_10182,N_9884,N_9995);
or U10183 (N_10183,N_9857,N_9854);
xnor U10184 (N_10184,N_9962,N_9805);
nor U10185 (N_10185,N_9925,N_9860);
and U10186 (N_10186,N_9806,N_9980);
or U10187 (N_10187,N_9884,N_9868);
nor U10188 (N_10188,N_9929,N_9818);
nor U10189 (N_10189,N_9881,N_9962);
nand U10190 (N_10190,N_9809,N_9814);
nand U10191 (N_10191,N_9914,N_9991);
and U10192 (N_10192,N_9974,N_9983);
or U10193 (N_10193,N_9814,N_9800);
nand U10194 (N_10194,N_9838,N_9915);
and U10195 (N_10195,N_9992,N_9882);
and U10196 (N_10196,N_9935,N_9874);
xnor U10197 (N_10197,N_9952,N_9838);
nand U10198 (N_10198,N_9809,N_9854);
xor U10199 (N_10199,N_9991,N_9906);
nand U10200 (N_10200,N_10090,N_10085);
and U10201 (N_10201,N_10067,N_10106);
nand U10202 (N_10202,N_10129,N_10154);
xor U10203 (N_10203,N_10033,N_10005);
xor U10204 (N_10204,N_10160,N_10004);
and U10205 (N_10205,N_10130,N_10092);
or U10206 (N_10206,N_10177,N_10042);
or U10207 (N_10207,N_10128,N_10073);
or U10208 (N_10208,N_10168,N_10032);
and U10209 (N_10209,N_10058,N_10124);
and U10210 (N_10210,N_10146,N_10010);
and U10211 (N_10211,N_10025,N_10165);
nand U10212 (N_10212,N_10122,N_10104);
and U10213 (N_10213,N_10054,N_10173);
or U10214 (N_10214,N_10096,N_10055);
nor U10215 (N_10215,N_10011,N_10115);
nor U10216 (N_10216,N_10070,N_10187);
xor U10217 (N_10217,N_10072,N_10143);
nor U10218 (N_10218,N_10188,N_10066);
or U10219 (N_10219,N_10041,N_10174);
and U10220 (N_10220,N_10121,N_10053);
or U10221 (N_10221,N_10193,N_10157);
nand U10222 (N_10222,N_10197,N_10148);
nand U10223 (N_10223,N_10110,N_10134);
or U10224 (N_10224,N_10030,N_10133);
xor U10225 (N_10225,N_10152,N_10138);
and U10226 (N_10226,N_10035,N_10182);
nor U10227 (N_10227,N_10175,N_10196);
xor U10228 (N_10228,N_10161,N_10063);
and U10229 (N_10229,N_10060,N_10028);
xor U10230 (N_10230,N_10084,N_10052);
xnor U10231 (N_10231,N_10051,N_10099);
and U10232 (N_10232,N_10023,N_10153);
nand U10233 (N_10233,N_10167,N_10108);
or U10234 (N_10234,N_10094,N_10150);
and U10235 (N_10235,N_10001,N_10093);
nor U10236 (N_10236,N_10008,N_10185);
or U10237 (N_10237,N_10132,N_10095);
xnor U10238 (N_10238,N_10044,N_10176);
nor U10239 (N_10239,N_10075,N_10027);
xor U10240 (N_10240,N_10172,N_10199);
nor U10241 (N_10241,N_10117,N_10105);
and U10242 (N_10242,N_10020,N_10000);
nor U10243 (N_10243,N_10147,N_10198);
nor U10244 (N_10244,N_10109,N_10149);
nor U10245 (N_10245,N_10181,N_10040);
nor U10246 (N_10246,N_10123,N_10111);
or U10247 (N_10247,N_10114,N_10191);
nand U10248 (N_10248,N_10194,N_10192);
nand U10249 (N_10249,N_10140,N_10116);
xor U10250 (N_10250,N_10048,N_10136);
and U10251 (N_10251,N_10195,N_10034);
or U10252 (N_10252,N_10159,N_10078);
and U10253 (N_10253,N_10098,N_10164);
and U10254 (N_10254,N_10036,N_10170);
nor U10255 (N_10255,N_10118,N_10037);
nand U10256 (N_10256,N_10069,N_10135);
nand U10257 (N_10257,N_10065,N_10127);
xnor U10258 (N_10258,N_10026,N_10071);
nand U10259 (N_10259,N_10144,N_10077);
nor U10260 (N_10260,N_10083,N_10076);
and U10261 (N_10261,N_10113,N_10183);
or U10262 (N_10262,N_10029,N_10080);
and U10263 (N_10263,N_10101,N_10017);
or U10264 (N_10264,N_10009,N_10125);
and U10265 (N_10265,N_10006,N_10137);
nor U10266 (N_10266,N_10081,N_10163);
or U10267 (N_10267,N_10142,N_10186);
or U10268 (N_10268,N_10003,N_10031);
and U10269 (N_10269,N_10171,N_10086);
xnor U10270 (N_10270,N_10180,N_10156);
xnor U10271 (N_10271,N_10139,N_10014);
and U10272 (N_10272,N_10126,N_10047);
nor U10273 (N_10273,N_10064,N_10131);
xnor U10274 (N_10274,N_10087,N_10059);
and U10275 (N_10275,N_10184,N_10019);
and U10276 (N_10276,N_10151,N_10162);
and U10277 (N_10277,N_10145,N_10107);
or U10278 (N_10278,N_10103,N_10021);
nand U10279 (N_10279,N_10112,N_10082);
and U10280 (N_10280,N_10120,N_10024);
and U10281 (N_10281,N_10119,N_10013);
and U10282 (N_10282,N_10061,N_10155);
or U10283 (N_10283,N_10062,N_10015);
nor U10284 (N_10284,N_10079,N_10097);
nor U10285 (N_10285,N_10049,N_10141);
and U10286 (N_10286,N_10089,N_10158);
nor U10287 (N_10287,N_10169,N_10022);
xor U10288 (N_10288,N_10088,N_10007);
nor U10289 (N_10289,N_10045,N_10050);
xor U10290 (N_10290,N_10100,N_10043);
xor U10291 (N_10291,N_10016,N_10102);
and U10292 (N_10292,N_10018,N_10074);
xnor U10293 (N_10293,N_10056,N_10012);
nand U10294 (N_10294,N_10190,N_10178);
or U10295 (N_10295,N_10189,N_10179);
xnor U10296 (N_10296,N_10046,N_10057);
nor U10297 (N_10297,N_10038,N_10002);
or U10298 (N_10298,N_10039,N_10166);
nor U10299 (N_10299,N_10068,N_10091);
nor U10300 (N_10300,N_10099,N_10158);
nand U10301 (N_10301,N_10046,N_10047);
xor U10302 (N_10302,N_10082,N_10100);
xnor U10303 (N_10303,N_10169,N_10011);
nor U10304 (N_10304,N_10126,N_10039);
nor U10305 (N_10305,N_10149,N_10119);
xor U10306 (N_10306,N_10012,N_10001);
nand U10307 (N_10307,N_10181,N_10012);
nor U10308 (N_10308,N_10056,N_10122);
or U10309 (N_10309,N_10046,N_10170);
and U10310 (N_10310,N_10064,N_10078);
nor U10311 (N_10311,N_10094,N_10142);
nand U10312 (N_10312,N_10157,N_10075);
xnor U10313 (N_10313,N_10100,N_10003);
nand U10314 (N_10314,N_10081,N_10129);
xor U10315 (N_10315,N_10157,N_10108);
nor U10316 (N_10316,N_10090,N_10123);
and U10317 (N_10317,N_10160,N_10144);
nand U10318 (N_10318,N_10063,N_10000);
nand U10319 (N_10319,N_10077,N_10072);
and U10320 (N_10320,N_10103,N_10094);
and U10321 (N_10321,N_10159,N_10151);
nand U10322 (N_10322,N_10070,N_10007);
nor U10323 (N_10323,N_10053,N_10025);
nor U10324 (N_10324,N_10175,N_10030);
xnor U10325 (N_10325,N_10157,N_10015);
or U10326 (N_10326,N_10159,N_10190);
nor U10327 (N_10327,N_10087,N_10174);
xor U10328 (N_10328,N_10104,N_10127);
nand U10329 (N_10329,N_10005,N_10181);
xor U10330 (N_10330,N_10038,N_10106);
nor U10331 (N_10331,N_10151,N_10085);
nor U10332 (N_10332,N_10005,N_10198);
nand U10333 (N_10333,N_10036,N_10153);
nor U10334 (N_10334,N_10130,N_10121);
nand U10335 (N_10335,N_10025,N_10047);
or U10336 (N_10336,N_10029,N_10104);
xnor U10337 (N_10337,N_10144,N_10028);
xnor U10338 (N_10338,N_10141,N_10187);
or U10339 (N_10339,N_10062,N_10175);
nand U10340 (N_10340,N_10037,N_10079);
nand U10341 (N_10341,N_10046,N_10099);
nor U10342 (N_10342,N_10043,N_10106);
nand U10343 (N_10343,N_10097,N_10199);
xor U10344 (N_10344,N_10185,N_10091);
and U10345 (N_10345,N_10068,N_10088);
and U10346 (N_10346,N_10193,N_10131);
or U10347 (N_10347,N_10116,N_10064);
or U10348 (N_10348,N_10129,N_10023);
nor U10349 (N_10349,N_10067,N_10190);
or U10350 (N_10350,N_10096,N_10066);
nor U10351 (N_10351,N_10198,N_10119);
or U10352 (N_10352,N_10099,N_10031);
and U10353 (N_10353,N_10124,N_10089);
nand U10354 (N_10354,N_10013,N_10087);
or U10355 (N_10355,N_10107,N_10115);
and U10356 (N_10356,N_10065,N_10087);
xnor U10357 (N_10357,N_10132,N_10120);
nand U10358 (N_10358,N_10006,N_10075);
nor U10359 (N_10359,N_10022,N_10012);
nor U10360 (N_10360,N_10120,N_10016);
nand U10361 (N_10361,N_10155,N_10100);
and U10362 (N_10362,N_10097,N_10013);
and U10363 (N_10363,N_10068,N_10161);
xor U10364 (N_10364,N_10020,N_10194);
nor U10365 (N_10365,N_10007,N_10091);
or U10366 (N_10366,N_10030,N_10107);
and U10367 (N_10367,N_10036,N_10017);
and U10368 (N_10368,N_10031,N_10127);
nand U10369 (N_10369,N_10046,N_10105);
xor U10370 (N_10370,N_10083,N_10193);
and U10371 (N_10371,N_10052,N_10186);
or U10372 (N_10372,N_10128,N_10151);
nor U10373 (N_10373,N_10085,N_10054);
or U10374 (N_10374,N_10195,N_10139);
nor U10375 (N_10375,N_10167,N_10120);
and U10376 (N_10376,N_10039,N_10040);
xnor U10377 (N_10377,N_10102,N_10140);
xor U10378 (N_10378,N_10042,N_10139);
nand U10379 (N_10379,N_10077,N_10069);
and U10380 (N_10380,N_10047,N_10103);
and U10381 (N_10381,N_10080,N_10049);
and U10382 (N_10382,N_10151,N_10197);
xor U10383 (N_10383,N_10085,N_10196);
and U10384 (N_10384,N_10006,N_10090);
and U10385 (N_10385,N_10007,N_10120);
xor U10386 (N_10386,N_10044,N_10093);
nand U10387 (N_10387,N_10080,N_10038);
or U10388 (N_10388,N_10042,N_10017);
xnor U10389 (N_10389,N_10141,N_10064);
or U10390 (N_10390,N_10068,N_10013);
nor U10391 (N_10391,N_10051,N_10080);
xor U10392 (N_10392,N_10104,N_10037);
nand U10393 (N_10393,N_10074,N_10051);
xor U10394 (N_10394,N_10138,N_10110);
or U10395 (N_10395,N_10054,N_10043);
nor U10396 (N_10396,N_10123,N_10094);
or U10397 (N_10397,N_10001,N_10106);
or U10398 (N_10398,N_10179,N_10130);
or U10399 (N_10399,N_10022,N_10008);
nor U10400 (N_10400,N_10201,N_10341);
and U10401 (N_10401,N_10300,N_10374);
and U10402 (N_10402,N_10386,N_10213);
xor U10403 (N_10403,N_10265,N_10384);
and U10404 (N_10404,N_10259,N_10226);
nor U10405 (N_10405,N_10223,N_10367);
or U10406 (N_10406,N_10372,N_10364);
nand U10407 (N_10407,N_10375,N_10254);
or U10408 (N_10408,N_10320,N_10214);
nor U10409 (N_10409,N_10250,N_10277);
nand U10410 (N_10410,N_10286,N_10340);
and U10411 (N_10411,N_10337,N_10228);
nor U10412 (N_10412,N_10326,N_10330);
nor U10413 (N_10413,N_10304,N_10356);
or U10414 (N_10414,N_10302,N_10296);
nor U10415 (N_10415,N_10362,N_10258);
xnor U10416 (N_10416,N_10343,N_10331);
nor U10417 (N_10417,N_10390,N_10352);
xor U10418 (N_10418,N_10312,N_10270);
or U10419 (N_10419,N_10212,N_10204);
nand U10420 (N_10420,N_10260,N_10227);
nor U10421 (N_10421,N_10385,N_10393);
xor U10422 (N_10422,N_10378,N_10282);
and U10423 (N_10423,N_10342,N_10392);
or U10424 (N_10424,N_10285,N_10338);
or U10425 (N_10425,N_10377,N_10244);
nand U10426 (N_10426,N_10269,N_10247);
and U10427 (N_10427,N_10321,N_10242);
xnor U10428 (N_10428,N_10280,N_10200);
or U10429 (N_10429,N_10287,N_10257);
and U10430 (N_10430,N_10301,N_10249);
xnor U10431 (N_10431,N_10314,N_10294);
and U10432 (N_10432,N_10366,N_10264);
and U10433 (N_10433,N_10293,N_10399);
xnor U10434 (N_10434,N_10335,N_10297);
nand U10435 (N_10435,N_10311,N_10334);
nor U10436 (N_10436,N_10327,N_10336);
xor U10437 (N_10437,N_10291,N_10281);
or U10438 (N_10438,N_10389,N_10373);
nand U10439 (N_10439,N_10332,N_10325);
nor U10440 (N_10440,N_10348,N_10288);
nand U10441 (N_10441,N_10262,N_10350);
xor U10442 (N_10442,N_10395,N_10205);
xor U10443 (N_10443,N_10383,N_10253);
nand U10444 (N_10444,N_10307,N_10239);
or U10445 (N_10445,N_10363,N_10278);
xor U10446 (N_10446,N_10353,N_10359);
or U10447 (N_10447,N_10209,N_10308);
or U10448 (N_10448,N_10273,N_10231);
and U10449 (N_10449,N_10255,N_10360);
or U10450 (N_10450,N_10243,N_10319);
nor U10451 (N_10451,N_10382,N_10279);
or U10452 (N_10452,N_10391,N_10222);
and U10453 (N_10453,N_10346,N_10230);
nand U10454 (N_10454,N_10380,N_10345);
or U10455 (N_10455,N_10216,N_10206);
nor U10456 (N_10456,N_10272,N_10397);
or U10457 (N_10457,N_10323,N_10203);
and U10458 (N_10458,N_10354,N_10349);
or U10459 (N_10459,N_10256,N_10238);
nor U10460 (N_10460,N_10347,N_10322);
or U10461 (N_10461,N_10351,N_10284);
nand U10462 (N_10462,N_10370,N_10202);
nand U10463 (N_10463,N_10365,N_10251);
xor U10464 (N_10464,N_10224,N_10219);
or U10465 (N_10465,N_10207,N_10261);
and U10466 (N_10466,N_10233,N_10339);
and U10467 (N_10467,N_10317,N_10266);
xor U10468 (N_10468,N_10358,N_10248);
or U10469 (N_10469,N_10394,N_10225);
nand U10470 (N_10470,N_10376,N_10234);
nor U10471 (N_10471,N_10274,N_10271);
and U10472 (N_10472,N_10221,N_10276);
nor U10473 (N_10473,N_10240,N_10298);
nand U10474 (N_10474,N_10299,N_10211);
xnor U10475 (N_10475,N_10267,N_10220);
or U10476 (N_10476,N_10357,N_10381);
xnor U10477 (N_10477,N_10268,N_10292);
nor U10478 (N_10478,N_10355,N_10313);
xnor U10479 (N_10479,N_10218,N_10246);
nor U10480 (N_10480,N_10263,N_10329);
nor U10481 (N_10481,N_10369,N_10368);
xor U10482 (N_10482,N_10318,N_10245);
and U10483 (N_10483,N_10210,N_10232);
xnor U10484 (N_10484,N_10316,N_10333);
nor U10485 (N_10485,N_10387,N_10241);
or U10486 (N_10486,N_10324,N_10295);
nor U10487 (N_10487,N_10235,N_10361);
and U10488 (N_10488,N_10283,N_10306);
and U10489 (N_10489,N_10236,N_10305);
nor U10490 (N_10490,N_10309,N_10229);
xnor U10491 (N_10491,N_10208,N_10388);
or U10492 (N_10492,N_10315,N_10398);
or U10493 (N_10493,N_10396,N_10303);
xor U10494 (N_10494,N_10252,N_10237);
or U10495 (N_10495,N_10310,N_10371);
xor U10496 (N_10496,N_10275,N_10290);
xor U10497 (N_10497,N_10328,N_10344);
nor U10498 (N_10498,N_10215,N_10379);
nor U10499 (N_10499,N_10289,N_10217);
nand U10500 (N_10500,N_10298,N_10223);
nor U10501 (N_10501,N_10207,N_10221);
nand U10502 (N_10502,N_10383,N_10318);
xnor U10503 (N_10503,N_10295,N_10302);
nand U10504 (N_10504,N_10393,N_10236);
or U10505 (N_10505,N_10355,N_10365);
nand U10506 (N_10506,N_10210,N_10275);
and U10507 (N_10507,N_10293,N_10258);
nor U10508 (N_10508,N_10254,N_10387);
nor U10509 (N_10509,N_10327,N_10200);
xnor U10510 (N_10510,N_10365,N_10276);
xor U10511 (N_10511,N_10286,N_10232);
nand U10512 (N_10512,N_10280,N_10239);
nand U10513 (N_10513,N_10273,N_10226);
nand U10514 (N_10514,N_10387,N_10249);
nor U10515 (N_10515,N_10330,N_10362);
and U10516 (N_10516,N_10216,N_10260);
nand U10517 (N_10517,N_10310,N_10341);
and U10518 (N_10518,N_10352,N_10256);
nor U10519 (N_10519,N_10215,N_10234);
nand U10520 (N_10520,N_10378,N_10371);
or U10521 (N_10521,N_10339,N_10270);
and U10522 (N_10522,N_10211,N_10239);
xnor U10523 (N_10523,N_10232,N_10267);
nand U10524 (N_10524,N_10255,N_10297);
and U10525 (N_10525,N_10394,N_10359);
and U10526 (N_10526,N_10365,N_10366);
xor U10527 (N_10527,N_10330,N_10260);
and U10528 (N_10528,N_10379,N_10225);
and U10529 (N_10529,N_10354,N_10346);
nor U10530 (N_10530,N_10249,N_10271);
xor U10531 (N_10531,N_10203,N_10357);
or U10532 (N_10532,N_10272,N_10205);
xor U10533 (N_10533,N_10321,N_10250);
xnor U10534 (N_10534,N_10219,N_10318);
or U10535 (N_10535,N_10246,N_10222);
nor U10536 (N_10536,N_10228,N_10241);
and U10537 (N_10537,N_10281,N_10246);
xnor U10538 (N_10538,N_10358,N_10222);
nor U10539 (N_10539,N_10246,N_10357);
nand U10540 (N_10540,N_10394,N_10253);
and U10541 (N_10541,N_10274,N_10353);
and U10542 (N_10542,N_10338,N_10215);
nand U10543 (N_10543,N_10376,N_10369);
or U10544 (N_10544,N_10251,N_10287);
xnor U10545 (N_10545,N_10347,N_10381);
xor U10546 (N_10546,N_10354,N_10311);
or U10547 (N_10547,N_10370,N_10278);
or U10548 (N_10548,N_10331,N_10367);
or U10549 (N_10549,N_10229,N_10313);
xnor U10550 (N_10550,N_10239,N_10273);
or U10551 (N_10551,N_10206,N_10200);
and U10552 (N_10552,N_10246,N_10356);
and U10553 (N_10553,N_10263,N_10249);
and U10554 (N_10554,N_10254,N_10275);
or U10555 (N_10555,N_10238,N_10252);
nor U10556 (N_10556,N_10345,N_10292);
nor U10557 (N_10557,N_10333,N_10326);
or U10558 (N_10558,N_10250,N_10371);
xnor U10559 (N_10559,N_10260,N_10247);
nand U10560 (N_10560,N_10347,N_10388);
or U10561 (N_10561,N_10299,N_10336);
xnor U10562 (N_10562,N_10235,N_10320);
nand U10563 (N_10563,N_10346,N_10228);
nand U10564 (N_10564,N_10216,N_10291);
and U10565 (N_10565,N_10233,N_10368);
nor U10566 (N_10566,N_10383,N_10229);
or U10567 (N_10567,N_10368,N_10259);
nor U10568 (N_10568,N_10289,N_10324);
nand U10569 (N_10569,N_10333,N_10222);
or U10570 (N_10570,N_10350,N_10369);
xor U10571 (N_10571,N_10224,N_10273);
xnor U10572 (N_10572,N_10258,N_10369);
or U10573 (N_10573,N_10241,N_10208);
or U10574 (N_10574,N_10278,N_10386);
nand U10575 (N_10575,N_10344,N_10250);
nor U10576 (N_10576,N_10338,N_10281);
nor U10577 (N_10577,N_10214,N_10240);
or U10578 (N_10578,N_10228,N_10382);
and U10579 (N_10579,N_10325,N_10242);
xnor U10580 (N_10580,N_10232,N_10229);
and U10581 (N_10581,N_10297,N_10202);
nor U10582 (N_10582,N_10346,N_10349);
or U10583 (N_10583,N_10311,N_10355);
and U10584 (N_10584,N_10265,N_10364);
and U10585 (N_10585,N_10323,N_10366);
nand U10586 (N_10586,N_10278,N_10365);
nand U10587 (N_10587,N_10389,N_10237);
nor U10588 (N_10588,N_10262,N_10268);
xnor U10589 (N_10589,N_10308,N_10273);
nor U10590 (N_10590,N_10329,N_10214);
xor U10591 (N_10591,N_10310,N_10225);
or U10592 (N_10592,N_10311,N_10253);
nor U10593 (N_10593,N_10295,N_10381);
xnor U10594 (N_10594,N_10205,N_10206);
nor U10595 (N_10595,N_10210,N_10261);
nor U10596 (N_10596,N_10224,N_10296);
nor U10597 (N_10597,N_10390,N_10361);
and U10598 (N_10598,N_10332,N_10355);
nand U10599 (N_10599,N_10301,N_10373);
nand U10600 (N_10600,N_10470,N_10599);
or U10601 (N_10601,N_10443,N_10469);
nor U10602 (N_10602,N_10447,N_10451);
xor U10603 (N_10603,N_10406,N_10492);
or U10604 (N_10604,N_10577,N_10506);
nand U10605 (N_10605,N_10432,N_10485);
or U10606 (N_10606,N_10550,N_10593);
xnor U10607 (N_10607,N_10412,N_10415);
nand U10608 (N_10608,N_10572,N_10414);
and U10609 (N_10609,N_10422,N_10528);
and U10610 (N_10610,N_10501,N_10571);
xnor U10611 (N_10611,N_10520,N_10454);
nor U10612 (N_10612,N_10574,N_10585);
nand U10613 (N_10613,N_10569,N_10487);
and U10614 (N_10614,N_10507,N_10486);
nor U10615 (N_10615,N_10563,N_10423);
and U10616 (N_10616,N_10519,N_10595);
nor U10617 (N_10617,N_10436,N_10512);
xor U10618 (N_10618,N_10483,N_10578);
or U10619 (N_10619,N_10541,N_10554);
nor U10620 (N_10620,N_10521,N_10437);
nor U10621 (N_10621,N_10476,N_10544);
xnor U10622 (N_10622,N_10568,N_10559);
nand U10623 (N_10623,N_10474,N_10530);
and U10624 (N_10624,N_10460,N_10409);
nor U10625 (N_10625,N_10404,N_10416);
xnor U10626 (N_10626,N_10418,N_10427);
nand U10627 (N_10627,N_10534,N_10518);
or U10628 (N_10628,N_10539,N_10430);
nand U10629 (N_10629,N_10558,N_10537);
nand U10630 (N_10630,N_10576,N_10400);
or U10631 (N_10631,N_10450,N_10497);
and U10632 (N_10632,N_10459,N_10582);
xor U10633 (N_10633,N_10489,N_10555);
or U10634 (N_10634,N_10535,N_10581);
nor U10635 (N_10635,N_10560,N_10548);
and U10636 (N_10636,N_10570,N_10442);
nand U10637 (N_10637,N_10538,N_10439);
and U10638 (N_10638,N_10529,N_10573);
and U10639 (N_10639,N_10495,N_10549);
or U10640 (N_10640,N_10401,N_10435);
xor U10641 (N_10641,N_10477,N_10511);
nor U10642 (N_10642,N_10446,N_10444);
nand U10643 (N_10643,N_10562,N_10480);
and U10644 (N_10644,N_10588,N_10473);
nand U10645 (N_10645,N_10407,N_10502);
or U10646 (N_10646,N_10566,N_10543);
xor U10647 (N_10647,N_10499,N_10546);
xor U10648 (N_10648,N_10516,N_10405);
nand U10649 (N_10649,N_10510,N_10457);
nand U10650 (N_10650,N_10551,N_10448);
xnor U10651 (N_10651,N_10488,N_10475);
xor U10652 (N_10652,N_10458,N_10493);
and U10653 (N_10653,N_10567,N_10453);
or U10654 (N_10654,N_10471,N_10402);
nor U10655 (N_10655,N_10526,N_10425);
or U10656 (N_10656,N_10408,N_10592);
nand U10657 (N_10657,N_10490,N_10597);
nand U10658 (N_10658,N_10417,N_10517);
nand U10659 (N_10659,N_10433,N_10533);
nor U10660 (N_10660,N_10419,N_10461);
nand U10661 (N_10661,N_10403,N_10557);
nand U10662 (N_10662,N_10410,N_10500);
and U10663 (N_10663,N_10428,N_10411);
xnor U10664 (N_10664,N_10484,N_10579);
or U10665 (N_10665,N_10564,N_10455);
nor U10666 (N_10666,N_10561,N_10532);
and U10667 (N_10667,N_10431,N_10525);
nand U10668 (N_10668,N_10509,N_10547);
and U10669 (N_10669,N_10494,N_10498);
or U10670 (N_10670,N_10527,N_10496);
nand U10671 (N_10671,N_10424,N_10591);
nor U10672 (N_10672,N_10514,N_10463);
or U10673 (N_10673,N_10465,N_10552);
nor U10674 (N_10674,N_10504,N_10429);
nor U10675 (N_10675,N_10590,N_10464);
xor U10676 (N_10676,N_10438,N_10522);
or U10677 (N_10677,N_10505,N_10553);
xnor U10678 (N_10678,N_10575,N_10580);
xor U10679 (N_10679,N_10508,N_10478);
xnor U10680 (N_10680,N_10440,N_10524);
or U10681 (N_10681,N_10531,N_10540);
nor U10682 (N_10682,N_10466,N_10583);
xor U10683 (N_10683,N_10542,N_10556);
or U10684 (N_10684,N_10598,N_10545);
and U10685 (N_10685,N_10479,N_10434);
or U10686 (N_10686,N_10565,N_10467);
and U10687 (N_10687,N_10462,N_10536);
and U10688 (N_10688,N_10426,N_10452);
or U10689 (N_10689,N_10523,N_10456);
xnor U10690 (N_10690,N_10413,N_10421);
xnor U10691 (N_10691,N_10441,N_10491);
xor U10692 (N_10692,N_10596,N_10515);
xnor U10693 (N_10693,N_10584,N_10587);
and U10694 (N_10694,N_10449,N_10481);
xor U10695 (N_10695,N_10445,N_10468);
or U10696 (N_10696,N_10586,N_10513);
or U10697 (N_10697,N_10472,N_10503);
nand U10698 (N_10698,N_10594,N_10482);
nor U10699 (N_10699,N_10589,N_10420);
or U10700 (N_10700,N_10495,N_10461);
xor U10701 (N_10701,N_10451,N_10496);
or U10702 (N_10702,N_10431,N_10409);
or U10703 (N_10703,N_10531,N_10425);
and U10704 (N_10704,N_10448,N_10468);
and U10705 (N_10705,N_10458,N_10496);
and U10706 (N_10706,N_10400,N_10461);
nor U10707 (N_10707,N_10529,N_10566);
nor U10708 (N_10708,N_10591,N_10506);
nand U10709 (N_10709,N_10504,N_10592);
or U10710 (N_10710,N_10586,N_10439);
nand U10711 (N_10711,N_10474,N_10522);
and U10712 (N_10712,N_10555,N_10504);
nand U10713 (N_10713,N_10485,N_10537);
and U10714 (N_10714,N_10514,N_10543);
and U10715 (N_10715,N_10421,N_10492);
xnor U10716 (N_10716,N_10430,N_10495);
nor U10717 (N_10717,N_10476,N_10431);
nor U10718 (N_10718,N_10573,N_10407);
and U10719 (N_10719,N_10490,N_10441);
and U10720 (N_10720,N_10496,N_10459);
xnor U10721 (N_10721,N_10483,N_10555);
xor U10722 (N_10722,N_10550,N_10548);
and U10723 (N_10723,N_10503,N_10475);
nor U10724 (N_10724,N_10413,N_10574);
or U10725 (N_10725,N_10420,N_10580);
or U10726 (N_10726,N_10416,N_10493);
or U10727 (N_10727,N_10413,N_10486);
nor U10728 (N_10728,N_10558,N_10526);
nand U10729 (N_10729,N_10464,N_10543);
nand U10730 (N_10730,N_10496,N_10516);
or U10731 (N_10731,N_10574,N_10422);
nor U10732 (N_10732,N_10498,N_10512);
nand U10733 (N_10733,N_10565,N_10571);
nand U10734 (N_10734,N_10502,N_10442);
and U10735 (N_10735,N_10473,N_10596);
and U10736 (N_10736,N_10588,N_10563);
xor U10737 (N_10737,N_10524,N_10584);
or U10738 (N_10738,N_10496,N_10429);
and U10739 (N_10739,N_10401,N_10553);
and U10740 (N_10740,N_10533,N_10431);
xor U10741 (N_10741,N_10581,N_10502);
nor U10742 (N_10742,N_10457,N_10569);
nor U10743 (N_10743,N_10488,N_10505);
nand U10744 (N_10744,N_10510,N_10539);
nor U10745 (N_10745,N_10545,N_10430);
xnor U10746 (N_10746,N_10401,N_10476);
or U10747 (N_10747,N_10580,N_10516);
or U10748 (N_10748,N_10581,N_10490);
and U10749 (N_10749,N_10492,N_10465);
xnor U10750 (N_10750,N_10492,N_10581);
xnor U10751 (N_10751,N_10443,N_10402);
or U10752 (N_10752,N_10408,N_10576);
and U10753 (N_10753,N_10500,N_10434);
or U10754 (N_10754,N_10437,N_10458);
or U10755 (N_10755,N_10561,N_10490);
and U10756 (N_10756,N_10534,N_10455);
nand U10757 (N_10757,N_10521,N_10400);
nor U10758 (N_10758,N_10483,N_10493);
nand U10759 (N_10759,N_10464,N_10572);
nand U10760 (N_10760,N_10506,N_10558);
nor U10761 (N_10761,N_10510,N_10578);
nand U10762 (N_10762,N_10537,N_10411);
and U10763 (N_10763,N_10514,N_10524);
and U10764 (N_10764,N_10544,N_10461);
nand U10765 (N_10765,N_10431,N_10420);
and U10766 (N_10766,N_10550,N_10436);
nand U10767 (N_10767,N_10414,N_10470);
or U10768 (N_10768,N_10571,N_10570);
and U10769 (N_10769,N_10593,N_10401);
nor U10770 (N_10770,N_10510,N_10460);
nor U10771 (N_10771,N_10475,N_10422);
or U10772 (N_10772,N_10550,N_10473);
and U10773 (N_10773,N_10423,N_10428);
nor U10774 (N_10774,N_10452,N_10506);
nor U10775 (N_10775,N_10597,N_10581);
nand U10776 (N_10776,N_10422,N_10588);
nor U10777 (N_10777,N_10448,N_10455);
xnor U10778 (N_10778,N_10562,N_10582);
nor U10779 (N_10779,N_10531,N_10406);
nand U10780 (N_10780,N_10591,N_10445);
nand U10781 (N_10781,N_10469,N_10467);
and U10782 (N_10782,N_10524,N_10408);
nand U10783 (N_10783,N_10514,N_10562);
and U10784 (N_10784,N_10453,N_10410);
nor U10785 (N_10785,N_10402,N_10484);
nand U10786 (N_10786,N_10571,N_10521);
or U10787 (N_10787,N_10465,N_10512);
nand U10788 (N_10788,N_10429,N_10483);
xnor U10789 (N_10789,N_10477,N_10537);
nor U10790 (N_10790,N_10410,N_10485);
or U10791 (N_10791,N_10597,N_10562);
nor U10792 (N_10792,N_10492,N_10546);
nand U10793 (N_10793,N_10493,N_10445);
and U10794 (N_10794,N_10550,N_10597);
or U10795 (N_10795,N_10520,N_10577);
and U10796 (N_10796,N_10412,N_10544);
xnor U10797 (N_10797,N_10588,N_10553);
nand U10798 (N_10798,N_10411,N_10541);
nand U10799 (N_10799,N_10412,N_10515);
and U10800 (N_10800,N_10719,N_10749);
nand U10801 (N_10801,N_10732,N_10603);
xor U10802 (N_10802,N_10616,N_10614);
or U10803 (N_10803,N_10629,N_10692);
and U10804 (N_10804,N_10631,N_10745);
or U10805 (N_10805,N_10799,N_10764);
and U10806 (N_10806,N_10766,N_10604);
and U10807 (N_10807,N_10789,N_10755);
xnor U10808 (N_10808,N_10610,N_10717);
xnor U10809 (N_10809,N_10793,N_10611);
and U10810 (N_10810,N_10770,N_10765);
xnor U10811 (N_10811,N_10754,N_10763);
and U10812 (N_10812,N_10675,N_10605);
nor U10813 (N_10813,N_10659,N_10637);
nand U10814 (N_10814,N_10679,N_10787);
xor U10815 (N_10815,N_10761,N_10662);
nand U10816 (N_10816,N_10711,N_10698);
nand U10817 (N_10817,N_10690,N_10669);
xor U10818 (N_10818,N_10791,N_10652);
nor U10819 (N_10819,N_10686,N_10664);
nor U10820 (N_10820,N_10758,N_10790);
or U10821 (N_10821,N_10621,N_10784);
nand U10822 (N_10822,N_10794,N_10792);
and U10823 (N_10823,N_10641,N_10709);
nor U10824 (N_10824,N_10747,N_10798);
xnor U10825 (N_10825,N_10665,N_10620);
xor U10826 (N_10826,N_10632,N_10689);
xor U10827 (N_10827,N_10617,N_10696);
or U10828 (N_10828,N_10772,N_10744);
xor U10829 (N_10829,N_10738,N_10721);
nand U10830 (N_10830,N_10716,N_10618);
and U10831 (N_10831,N_10737,N_10724);
or U10832 (N_10832,N_10708,N_10673);
and U10833 (N_10833,N_10704,N_10683);
nand U10834 (N_10834,N_10691,N_10672);
or U10835 (N_10835,N_10756,N_10615);
xor U10836 (N_10836,N_10788,N_10796);
nand U10837 (N_10837,N_10642,N_10701);
or U10838 (N_10838,N_10778,N_10657);
nor U10839 (N_10839,N_10760,N_10619);
nor U10840 (N_10840,N_10718,N_10702);
xor U10841 (N_10841,N_10668,N_10627);
and U10842 (N_10842,N_10650,N_10694);
or U10843 (N_10843,N_10685,N_10630);
and U10844 (N_10844,N_10628,N_10644);
and U10845 (N_10845,N_10748,N_10636);
or U10846 (N_10846,N_10783,N_10722);
or U10847 (N_10847,N_10622,N_10648);
nor U10848 (N_10848,N_10661,N_10751);
nor U10849 (N_10849,N_10731,N_10601);
nor U10850 (N_10850,N_10678,N_10705);
and U10851 (N_10851,N_10695,N_10735);
nor U10852 (N_10852,N_10707,N_10762);
or U10853 (N_10853,N_10774,N_10728);
xor U10854 (N_10854,N_10640,N_10688);
xor U10855 (N_10855,N_10660,N_10676);
or U10856 (N_10856,N_10634,N_10753);
and U10857 (N_10857,N_10677,N_10656);
nand U10858 (N_10858,N_10693,N_10713);
and U10859 (N_10859,N_10706,N_10782);
or U10860 (N_10860,N_10723,N_10714);
nor U10861 (N_10861,N_10666,N_10667);
or U10862 (N_10862,N_10730,N_10626);
xnor U10863 (N_10863,N_10703,N_10670);
xnor U10864 (N_10864,N_10795,N_10727);
nand U10865 (N_10865,N_10752,N_10699);
or U10866 (N_10866,N_10741,N_10743);
or U10867 (N_10867,N_10658,N_10746);
nor U10868 (N_10868,N_10715,N_10725);
nor U10869 (N_10869,N_10797,N_10647);
and U10870 (N_10870,N_10623,N_10645);
or U10871 (N_10871,N_10775,N_10740);
and U10872 (N_10872,N_10776,N_10742);
or U10873 (N_10873,N_10733,N_10684);
xnor U10874 (N_10874,N_10773,N_10633);
nand U10875 (N_10875,N_10779,N_10734);
or U10876 (N_10876,N_10712,N_10769);
nand U10877 (N_10877,N_10608,N_10607);
nor U10878 (N_10878,N_10674,N_10757);
and U10879 (N_10879,N_10682,N_10655);
and U10880 (N_10880,N_10643,N_10710);
and U10881 (N_10881,N_10663,N_10600);
nand U10882 (N_10882,N_10671,N_10609);
nor U10883 (N_10883,N_10750,N_10771);
nand U10884 (N_10884,N_10639,N_10638);
or U10885 (N_10885,N_10781,N_10651);
nor U10886 (N_10886,N_10625,N_10700);
nor U10887 (N_10887,N_10720,N_10606);
xor U10888 (N_10888,N_10624,N_10697);
and U10889 (N_10889,N_10759,N_10680);
or U10890 (N_10890,N_10777,N_10649);
nor U10891 (N_10891,N_10768,N_10736);
nor U10892 (N_10892,N_10613,N_10681);
or U10893 (N_10893,N_10739,N_10767);
xnor U10894 (N_10894,N_10726,N_10687);
nand U10895 (N_10895,N_10602,N_10786);
or U10896 (N_10896,N_10612,N_10780);
xnor U10897 (N_10897,N_10653,N_10729);
nor U10898 (N_10898,N_10785,N_10646);
and U10899 (N_10899,N_10635,N_10654);
or U10900 (N_10900,N_10690,N_10706);
xnor U10901 (N_10901,N_10710,N_10730);
and U10902 (N_10902,N_10788,N_10705);
and U10903 (N_10903,N_10767,N_10645);
nand U10904 (N_10904,N_10676,N_10707);
nand U10905 (N_10905,N_10790,N_10638);
nand U10906 (N_10906,N_10701,N_10681);
and U10907 (N_10907,N_10600,N_10732);
nand U10908 (N_10908,N_10618,N_10604);
or U10909 (N_10909,N_10753,N_10605);
xor U10910 (N_10910,N_10725,N_10787);
xor U10911 (N_10911,N_10689,N_10622);
and U10912 (N_10912,N_10600,N_10700);
nand U10913 (N_10913,N_10669,N_10697);
nor U10914 (N_10914,N_10682,N_10702);
and U10915 (N_10915,N_10638,N_10774);
nand U10916 (N_10916,N_10731,N_10756);
nand U10917 (N_10917,N_10665,N_10742);
xnor U10918 (N_10918,N_10642,N_10754);
nor U10919 (N_10919,N_10734,N_10778);
nor U10920 (N_10920,N_10777,N_10639);
xor U10921 (N_10921,N_10780,N_10614);
or U10922 (N_10922,N_10794,N_10746);
or U10923 (N_10923,N_10715,N_10789);
nand U10924 (N_10924,N_10785,N_10649);
nor U10925 (N_10925,N_10658,N_10737);
nand U10926 (N_10926,N_10757,N_10799);
or U10927 (N_10927,N_10622,N_10703);
nand U10928 (N_10928,N_10697,N_10783);
xor U10929 (N_10929,N_10778,N_10742);
and U10930 (N_10930,N_10624,N_10637);
nor U10931 (N_10931,N_10607,N_10666);
nand U10932 (N_10932,N_10767,N_10638);
and U10933 (N_10933,N_10753,N_10638);
nand U10934 (N_10934,N_10720,N_10626);
nor U10935 (N_10935,N_10783,N_10719);
and U10936 (N_10936,N_10601,N_10678);
nor U10937 (N_10937,N_10728,N_10609);
nor U10938 (N_10938,N_10658,N_10648);
xor U10939 (N_10939,N_10788,N_10642);
nand U10940 (N_10940,N_10750,N_10709);
nand U10941 (N_10941,N_10736,N_10627);
nand U10942 (N_10942,N_10601,N_10609);
nor U10943 (N_10943,N_10735,N_10782);
xor U10944 (N_10944,N_10657,N_10686);
xor U10945 (N_10945,N_10708,N_10627);
xnor U10946 (N_10946,N_10715,N_10726);
xor U10947 (N_10947,N_10716,N_10623);
nor U10948 (N_10948,N_10745,N_10675);
nor U10949 (N_10949,N_10661,N_10691);
nor U10950 (N_10950,N_10707,N_10610);
nand U10951 (N_10951,N_10630,N_10735);
nor U10952 (N_10952,N_10785,N_10717);
nand U10953 (N_10953,N_10787,N_10631);
xor U10954 (N_10954,N_10657,N_10652);
xnor U10955 (N_10955,N_10794,N_10713);
xnor U10956 (N_10956,N_10696,N_10764);
xnor U10957 (N_10957,N_10648,N_10705);
or U10958 (N_10958,N_10710,N_10732);
nand U10959 (N_10959,N_10652,N_10631);
and U10960 (N_10960,N_10717,N_10747);
and U10961 (N_10961,N_10621,N_10652);
nor U10962 (N_10962,N_10744,N_10782);
nor U10963 (N_10963,N_10764,N_10784);
or U10964 (N_10964,N_10602,N_10768);
nor U10965 (N_10965,N_10602,N_10617);
nor U10966 (N_10966,N_10753,N_10725);
or U10967 (N_10967,N_10730,N_10772);
or U10968 (N_10968,N_10695,N_10741);
nand U10969 (N_10969,N_10647,N_10737);
and U10970 (N_10970,N_10602,N_10736);
and U10971 (N_10971,N_10772,N_10725);
and U10972 (N_10972,N_10639,N_10667);
xnor U10973 (N_10973,N_10724,N_10666);
and U10974 (N_10974,N_10643,N_10764);
nand U10975 (N_10975,N_10693,N_10744);
or U10976 (N_10976,N_10732,N_10696);
xor U10977 (N_10977,N_10755,N_10798);
and U10978 (N_10978,N_10719,N_10686);
xor U10979 (N_10979,N_10681,N_10669);
or U10980 (N_10980,N_10662,N_10728);
and U10981 (N_10981,N_10798,N_10794);
nand U10982 (N_10982,N_10725,N_10672);
xor U10983 (N_10983,N_10612,N_10681);
and U10984 (N_10984,N_10790,N_10624);
xnor U10985 (N_10985,N_10619,N_10651);
nand U10986 (N_10986,N_10605,N_10742);
nand U10987 (N_10987,N_10654,N_10722);
xnor U10988 (N_10988,N_10767,N_10649);
and U10989 (N_10989,N_10646,N_10703);
or U10990 (N_10990,N_10777,N_10644);
nor U10991 (N_10991,N_10631,N_10683);
nor U10992 (N_10992,N_10718,N_10624);
nand U10993 (N_10993,N_10622,N_10669);
xnor U10994 (N_10994,N_10783,N_10621);
and U10995 (N_10995,N_10691,N_10716);
or U10996 (N_10996,N_10614,N_10685);
xnor U10997 (N_10997,N_10613,N_10761);
nor U10998 (N_10998,N_10735,N_10698);
or U10999 (N_10999,N_10729,N_10784);
nand U11000 (N_11000,N_10920,N_10864);
nor U11001 (N_11001,N_10947,N_10809);
or U11002 (N_11002,N_10904,N_10818);
nor U11003 (N_11003,N_10926,N_10982);
and U11004 (N_11004,N_10832,N_10951);
or U11005 (N_11005,N_10981,N_10999);
nor U11006 (N_11006,N_10942,N_10934);
xnor U11007 (N_11007,N_10849,N_10836);
and U11008 (N_11008,N_10929,N_10997);
xnor U11009 (N_11009,N_10949,N_10819);
nand U11010 (N_11010,N_10924,N_10862);
or U11011 (N_11011,N_10917,N_10941);
and U11012 (N_11012,N_10800,N_10987);
and U11013 (N_11013,N_10954,N_10980);
nand U11014 (N_11014,N_10815,N_10892);
nor U11015 (N_11015,N_10974,N_10966);
nor U11016 (N_11016,N_10936,N_10884);
nor U11017 (N_11017,N_10841,N_10945);
nor U11018 (N_11018,N_10810,N_10910);
xor U11019 (N_11019,N_10906,N_10994);
nor U11020 (N_11020,N_10975,N_10890);
or U11021 (N_11021,N_10842,N_10971);
nor U11022 (N_11022,N_10881,N_10855);
and U11023 (N_11023,N_10877,N_10880);
and U11024 (N_11024,N_10883,N_10958);
or U11025 (N_11025,N_10955,N_10932);
nand U11026 (N_11026,N_10854,N_10911);
nand U11027 (N_11027,N_10889,N_10878);
xnor U11028 (N_11028,N_10960,N_10825);
and U11029 (N_11029,N_10843,N_10953);
and U11030 (N_11030,N_10938,N_10845);
or U11031 (N_11031,N_10978,N_10868);
or U11032 (N_11032,N_10871,N_10894);
nor U11033 (N_11033,N_10990,N_10872);
and U11034 (N_11034,N_10963,N_10950);
and U11035 (N_11035,N_10882,N_10914);
and U11036 (N_11036,N_10930,N_10909);
nor U11037 (N_11037,N_10946,N_10863);
and U11038 (N_11038,N_10927,N_10874);
nand U11039 (N_11039,N_10984,N_10879);
nor U11040 (N_11040,N_10834,N_10859);
or U11041 (N_11041,N_10875,N_10952);
and U11042 (N_11042,N_10940,N_10967);
and U11043 (N_11043,N_10891,N_10885);
or U11044 (N_11044,N_10916,N_10820);
or U11045 (N_11045,N_10933,N_10833);
nand U11046 (N_11046,N_10886,N_10801);
xnor U11047 (N_11047,N_10893,N_10812);
and U11048 (N_11048,N_10931,N_10873);
nor U11049 (N_11049,N_10957,N_10811);
nand U11050 (N_11050,N_10976,N_10817);
or U11051 (N_11051,N_10847,N_10956);
nand U11052 (N_11052,N_10935,N_10870);
and U11053 (N_11053,N_10851,N_10876);
xnor U11054 (N_11054,N_10857,N_10995);
and U11055 (N_11055,N_10991,N_10977);
nand U11056 (N_11056,N_10943,N_10866);
nand U11057 (N_11057,N_10838,N_10858);
or U11058 (N_11058,N_10830,N_10805);
xor U11059 (N_11059,N_10816,N_10804);
and U11060 (N_11060,N_10973,N_10867);
and U11061 (N_11061,N_10813,N_10856);
and U11062 (N_11062,N_10802,N_10828);
nor U11063 (N_11063,N_10839,N_10923);
nand U11064 (N_11064,N_10860,N_10852);
nor U11065 (N_11065,N_10964,N_10992);
or U11066 (N_11066,N_10988,N_10996);
or U11067 (N_11067,N_10918,N_10896);
or U11068 (N_11068,N_10835,N_10948);
and U11069 (N_11069,N_10837,N_10962);
or U11070 (N_11070,N_10822,N_10848);
and U11071 (N_11071,N_10827,N_10865);
nand U11072 (N_11072,N_10826,N_10823);
xor U11073 (N_11073,N_10998,N_10900);
and U11074 (N_11074,N_10831,N_10993);
and U11075 (N_11075,N_10869,N_10821);
and U11076 (N_11076,N_10928,N_10983);
xnor U11077 (N_11077,N_10985,N_10902);
xor U11078 (N_11078,N_10829,N_10807);
nor U11079 (N_11079,N_10915,N_10925);
or U11080 (N_11080,N_10846,N_10895);
nor U11081 (N_11081,N_10903,N_10961);
xnor U11082 (N_11082,N_10887,N_10907);
nor U11083 (N_11083,N_10972,N_10965);
nor U11084 (N_11084,N_10808,N_10969);
nor U11085 (N_11085,N_10970,N_10840);
xnor U11086 (N_11086,N_10908,N_10888);
and U11087 (N_11087,N_10939,N_10986);
and U11088 (N_11088,N_10944,N_10921);
nand U11089 (N_11089,N_10861,N_10937);
xnor U11090 (N_11090,N_10853,N_10844);
and U11091 (N_11091,N_10824,N_10850);
xnor U11092 (N_11092,N_10968,N_10814);
and U11093 (N_11093,N_10979,N_10959);
or U11094 (N_11094,N_10913,N_10912);
and U11095 (N_11095,N_10897,N_10898);
nor U11096 (N_11096,N_10922,N_10806);
and U11097 (N_11097,N_10803,N_10905);
nand U11098 (N_11098,N_10901,N_10989);
nand U11099 (N_11099,N_10899,N_10919);
or U11100 (N_11100,N_10861,N_10983);
nor U11101 (N_11101,N_10860,N_10917);
nor U11102 (N_11102,N_10864,N_10939);
or U11103 (N_11103,N_10996,N_10992);
xnor U11104 (N_11104,N_10808,N_10814);
and U11105 (N_11105,N_10851,N_10916);
and U11106 (N_11106,N_10824,N_10994);
nand U11107 (N_11107,N_10928,N_10933);
and U11108 (N_11108,N_10998,N_10928);
and U11109 (N_11109,N_10987,N_10819);
or U11110 (N_11110,N_10823,N_10838);
nand U11111 (N_11111,N_10880,N_10870);
or U11112 (N_11112,N_10856,N_10997);
nand U11113 (N_11113,N_10910,N_10942);
xnor U11114 (N_11114,N_10937,N_10943);
xor U11115 (N_11115,N_10997,N_10833);
nor U11116 (N_11116,N_10869,N_10948);
xnor U11117 (N_11117,N_10952,N_10868);
nor U11118 (N_11118,N_10823,N_10812);
nand U11119 (N_11119,N_10880,N_10957);
nor U11120 (N_11120,N_10874,N_10966);
or U11121 (N_11121,N_10996,N_10870);
and U11122 (N_11122,N_10900,N_10879);
nor U11123 (N_11123,N_10899,N_10809);
nor U11124 (N_11124,N_10967,N_10812);
nor U11125 (N_11125,N_10988,N_10898);
and U11126 (N_11126,N_10839,N_10858);
or U11127 (N_11127,N_10830,N_10843);
xor U11128 (N_11128,N_10840,N_10983);
or U11129 (N_11129,N_10966,N_10813);
and U11130 (N_11130,N_10908,N_10830);
nand U11131 (N_11131,N_10970,N_10937);
and U11132 (N_11132,N_10930,N_10896);
and U11133 (N_11133,N_10922,N_10864);
and U11134 (N_11134,N_10909,N_10810);
nor U11135 (N_11135,N_10879,N_10807);
nor U11136 (N_11136,N_10808,N_10805);
nor U11137 (N_11137,N_10943,N_10898);
nand U11138 (N_11138,N_10919,N_10825);
xnor U11139 (N_11139,N_10916,N_10830);
nor U11140 (N_11140,N_10992,N_10898);
nand U11141 (N_11141,N_10865,N_10876);
nand U11142 (N_11142,N_10851,N_10841);
and U11143 (N_11143,N_10912,N_10953);
nor U11144 (N_11144,N_10937,N_10907);
nand U11145 (N_11145,N_10858,N_10810);
and U11146 (N_11146,N_10887,N_10846);
and U11147 (N_11147,N_10992,N_10852);
nor U11148 (N_11148,N_10970,N_10947);
and U11149 (N_11149,N_10908,N_10954);
and U11150 (N_11150,N_10838,N_10926);
or U11151 (N_11151,N_10959,N_10878);
nor U11152 (N_11152,N_10847,N_10865);
xor U11153 (N_11153,N_10824,N_10856);
nand U11154 (N_11154,N_10845,N_10847);
nor U11155 (N_11155,N_10978,N_10930);
or U11156 (N_11156,N_10949,N_10931);
or U11157 (N_11157,N_10854,N_10862);
xor U11158 (N_11158,N_10978,N_10835);
nor U11159 (N_11159,N_10822,N_10915);
and U11160 (N_11160,N_10831,N_10858);
or U11161 (N_11161,N_10886,N_10940);
xor U11162 (N_11162,N_10841,N_10804);
nand U11163 (N_11163,N_10837,N_10992);
and U11164 (N_11164,N_10843,N_10946);
nor U11165 (N_11165,N_10986,N_10890);
nor U11166 (N_11166,N_10897,N_10991);
nor U11167 (N_11167,N_10843,N_10966);
and U11168 (N_11168,N_10889,N_10886);
nand U11169 (N_11169,N_10965,N_10914);
or U11170 (N_11170,N_10873,N_10817);
or U11171 (N_11171,N_10881,N_10872);
nor U11172 (N_11172,N_10926,N_10867);
nor U11173 (N_11173,N_10963,N_10922);
nor U11174 (N_11174,N_10942,N_10874);
nand U11175 (N_11175,N_10896,N_10856);
nand U11176 (N_11176,N_10910,N_10959);
nand U11177 (N_11177,N_10908,N_10934);
xnor U11178 (N_11178,N_10995,N_10938);
and U11179 (N_11179,N_10937,N_10837);
or U11180 (N_11180,N_10924,N_10814);
xnor U11181 (N_11181,N_10862,N_10930);
nor U11182 (N_11182,N_10926,N_10974);
and U11183 (N_11183,N_10926,N_10886);
nand U11184 (N_11184,N_10857,N_10943);
or U11185 (N_11185,N_10966,N_10980);
nand U11186 (N_11186,N_10887,N_10952);
and U11187 (N_11187,N_10832,N_10826);
xor U11188 (N_11188,N_10838,N_10805);
and U11189 (N_11189,N_10977,N_10849);
xnor U11190 (N_11190,N_10890,N_10966);
and U11191 (N_11191,N_10987,N_10940);
and U11192 (N_11192,N_10992,N_10841);
xor U11193 (N_11193,N_10922,N_10877);
nand U11194 (N_11194,N_10813,N_10986);
or U11195 (N_11195,N_10830,N_10941);
xor U11196 (N_11196,N_10809,N_10982);
xor U11197 (N_11197,N_10966,N_10932);
xor U11198 (N_11198,N_10835,N_10808);
xor U11199 (N_11199,N_10912,N_10921);
nand U11200 (N_11200,N_11098,N_11060);
nor U11201 (N_11201,N_11036,N_11044);
and U11202 (N_11202,N_11080,N_11008);
nand U11203 (N_11203,N_11181,N_11110);
or U11204 (N_11204,N_11111,N_11195);
or U11205 (N_11205,N_11091,N_11024);
nor U11206 (N_11206,N_11174,N_11007);
nor U11207 (N_11207,N_11131,N_11179);
nor U11208 (N_11208,N_11094,N_11010);
xnor U11209 (N_11209,N_11009,N_11081);
nor U11210 (N_11210,N_11021,N_11020);
or U11211 (N_11211,N_11082,N_11148);
nor U11212 (N_11212,N_11023,N_11054);
nand U11213 (N_11213,N_11086,N_11027);
nor U11214 (N_11214,N_11083,N_11193);
or U11215 (N_11215,N_11022,N_11116);
and U11216 (N_11216,N_11068,N_11052);
nor U11217 (N_11217,N_11173,N_11093);
nand U11218 (N_11218,N_11159,N_11078);
or U11219 (N_11219,N_11030,N_11154);
nand U11220 (N_11220,N_11047,N_11090);
xor U11221 (N_11221,N_11186,N_11095);
and U11222 (N_11222,N_11139,N_11037);
xor U11223 (N_11223,N_11124,N_11133);
or U11224 (N_11224,N_11045,N_11017);
and U11225 (N_11225,N_11121,N_11178);
xor U11226 (N_11226,N_11145,N_11029);
nor U11227 (N_11227,N_11185,N_11016);
nand U11228 (N_11228,N_11171,N_11142);
nor U11229 (N_11229,N_11168,N_11119);
nor U11230 (N_11230,N_11109,N_11135);
and U11231 (N_11231,N_11101,N_11042);
nor U11232 (N_11232,N_11088,N_11143);
and U11233 (N_11233,N_11025,N_11084);
or U11234 (N_11234,N_11126,N_11040);
or U11235 (N_11235,N_11153,N_11170);
xnor U11236 (N_11236,N_11163,N_11097);
or U11237 (N_11237,N_11117,N_11100);
xnor U11238 (N_11238,N_11072,N_11151);
nand U11239 (N_11239,N_11141,N_11166);
and U11240 (N_11240,N_11187,N_11031);
nor U11241 (N_11241,N_11191,N_11180);
or U11242 (N_11242,N_11028,N_11085);
xnor U11243 (N_11243,N_11129,N_11053);
nand U11244 (N_11244,N_11011,N_11184);
or U11245 (N_11245,N_11099,N_11177);
or U11246 (N_11246,N_11120,N_11070);
or U11247 (N_11247,N_11164,N_11074);
nor U11248 (N_11248,N_11102,N_11150);
or U11249 (N_11249,N_11076,N_11089);
xor U11250 (N_11250,N_11136,N_11061);
and U11251 (N_11251,N_11073,N_11169);
or U11252 (N_11252,N_11161,N_11063);
nor U11253 (N_11253,N_11146,N_11162);
and U11254 (N_11254,N_11048,N_11188);
nor U11255 (N_11255,N_11182,N_11050);
nand U11256 (N_11256,N_11152,N_11033);
or U11257 (N_11257,N_11147,N_11134);
or U11258 (N_11258,N_11155,N_11003);
nand U11259 (N_11259,N_11183,N_11104);
nand U11260 (N_11260,N_11114,N_11189);
nor U11261 (N_11261,N_11115,N_11103);
or U11262 (N_11262,N_11056,N_11199);
xnor U11263 (N_11263,N_11140,N_11156);
nor U11264 (N_11264,N_11012,N_11165);
nand U11265 (N_11265,N_11127,N_11041);
or U11266 (N_11266,N_11032,N_11071);
xnor U11267 (N_11267,N_11014,N_11034);
or U11268 (N_11268,N_11130,N_11049);
xnor U11269 (N_11269,N_11075,N_11176);
nand U11270 (N_11270,N_11038,N_11160);
nor U11271 (N_11271,N_11077,N_11144);
xor U11272 (N_11272,N_11055,N_11051);
and U11273 (N_11273,N_11128,N_11105);
and U11274 (N_11274,N_11059,N_11096);
nor U11275 (N_11275,N_11112,N_11057);
or U11276 (N_11276,N_11197,N_11196);
and U11277 (N_11277,N_11158,N_11026);
nand U11278 (N_11278,N_11107,N_11125);
or U11279 (N_11279,N_11079,N_11043);
nor U11280 (N_11280,N_11190,N_11018);
and U11281 (N_11281,N_11013,N_11064);
nand U11282 (N_11282,N_11118,N_11194);
nor U11283 (N_11283,N_11035,N_11001);
xnor U11284 (N_11284,N_11066,N_11019);
and U11285 (N_11285,N_11065,N_11108);
xor U11286 (N_11286,N_11092,N_11087);
or U11287 (N_11287,N_11172,N_11137);
nand U11288 (N_11288,N_11149,N_11058);
or U11289 (N_11289,N_11004,N_11113);
or U11290 (N_11290,N_11015,N_11062);
and U11291 (N_11291,N_11039,N_11106);
xor U11292 (N_11292,N_11002,N_11157);
nor U11293 (N_11293,N_11069,N_11175);
nor U11294 (N_11294,N_11046,N_11123);
nor U11295 (N_11295,N_11132,N_11122);
nor U11296 (N_11296,N_11198,N_11192);
nand U11297 (N_11297,N_11005,N_11167);
xnor U11298 (N_11298,N_11006,N_11067);
and U11299 (N_11299,N_11000,N_11138);
xnor U11300 (N_11300,N_11113,N_11053);
or U11301 (N_11301,N_11053,N_11080);
xor U11302 (N_11302,N_11123,N_11087);
xnor U11303 (N_11303,N_11118,N_11090);
xnor U11304 (N_11304,N_11007,N_11011);
and U11305 (N_11305,N_11109,N_11190);
nand U11306 (N_11306,N_11085,N_11093);
or U11307 (N_11307,N_11058,N_11196);
nor U11308 (N_11308,N_11101,N_11010);
nand U11309 (N_11309,N_11107,N_11024);
nor U11310 (N_11310,N_11171,N_11182);
nand U11311 (N_11311,N_11088,N_11062);
nor U11312 (N_11312,N_11006,N_11196);
xor U11313 (N_11313,N_11135,N_11022);
xnor U11314 (N_11314,N_11042,N_11017);
and U11315 (N_11315,N_11076,N_11013);
nor U11316 (N_11316,N_11199,N_11124);
xnor U11317 (N_11317,N_11182,N_11159);
nor U11318 (N_11318,N_11179,N_11077);
xnor U11319 (N_11319,N_11087,N_11183);
and U11320 (N_11320,N_11018,N_11161);
nor U11321 (N_11321,N_11081,N_11058);
xor U11322 (N_11322,N_11085,N_11099);
nand U11323 (N_11323,N_11089,N_11166);
or U11324 (N_11324,N_11133,N_11130);
and U11325 (N_11325,N_11010,N_11114);
or U11326 (N_11326,N_11149,N_11007);
nor U11327 (N_11327,N_11097,N_11188);
nor U11328 (N_11328,N_11015,N_11074);
xor U11329 (N_11329,N_11065,N_11059);
or U11330 (N_11330,N_11186,N_11170);
nor U11331 (N_11331,N_11124,N_11198);
nand U11332 (N_11332,N_11048,N_11183);
xnor U11333 (N_11333,N_11153,N_11144);
nand U11334 (N_11334,N_11069,N_11130);
or U11335 (N_11335,N_11046,N_11111);
or U11336 (N_11336,N_11162,N_11140);
nor U11337 (N_11337,N_11006,N_11097);
xor U11338 (N_11338,N_11063,N_11108);
xnor U11339 (N_11339,N_11021,N_11015);
nand U11340 (N_11340,N_11195,N_11155);
or U11341 (N_11341,N_11078,N_11022);
and U11342 (N_11342,N_11103,N_11038);
nand U11343 (N_11343,N_11147,N_11013);
or U11344 (N_11344,N_11158,N_11109);
and U11345 (N_11345,N_11130,N_11151);
nor U11346 (N_11346,N_11111,N_11044);
or U11347 (N_11347,N_11018,N_11046);
or U11348 (N_11348,N_11105,N_11059);
and U11349 (N_11349,N_11110,N_11140);
nor U11350 (N_11350,N_11117,N_11193);
xnor U11351 (N_11351,N_11172,N_11167);
nand U11352 (N_11352,N_11137,N_11040);
and U11353 (N_11353,N_11018,N_11052);
xor U11354 (N_11354,N_11123,N_11122);
nand U11355 (N_11355,N_11092,N_11043);
nand U11356 (N_11356,N_11012,N_11013);
xnor U11357 (N_11357,N_11147,N_11170);
nor U11358 (N_11358,N_11058,N_11028);
nand U11359 (N_11359,N_11099,N_11115);
nor U11360 (N_11360,N_11034,N_11122);
and U11361 (N_11361,N_11023,N_11183);
and U11362 (N_11362,N_11042,N_11065);
nor U11363 (N_11363,N_11010,N_11048);
nand U11364 (N_11364,N_11075,N_11159);
xor U11365 (N_11365,N_11054,N_11019);
nor U11366 (N_11366,N_11113,N_11068);
xor U11367 (N_11367,N_11018,N_11199);
or U11368 (N_11368,N_11002,N_11013);
or U11369 (N_11369,N_11075,N_11062);
and U11370 (N_11370,N_11000,N_11183);
nor U11371 (N_11371,N_11055,N_11135);
nand U11372 (N_11372,N_11027,N_11002);
and U11373 (N_11373,N_11054,N_11020);
nand U11374 (N_11374,N_11046,N_11114);
nand U11375 (N_11375,N_11179,N_11142);
nor U11376 (N_11376,N_11121,N_11070);
and U11377 (N_11377,N_11035,N_11130);
and U11378 (N_11378,N_11049,N_11023);
or U11379 (N_11379,N_11096,N_11068);
or U11380 (N_11380,N_11060,N_11077);
or U11381 (N_11381,N_11139,N_11073);
xnor U11382 (N_11382,N_11074,N_11063);
nand U11383 (N_11383,N_11137,N_11111);
or U11384 (N_11384,N_11113,N_11161);
or U11385 (N_11385,N_11179,N_11035);
and U11386 (N_11386,N_11002,N_11145);
xor U11387 (N_11387,N_11144,N_11195);
nand U11388 (N_11388,N_11064,N_11071);
nor U11389 (N_11389,N_11185,N_11143);
nor U11390 (N_11390,N_11108,N_11148);
nand U11391 (N_11391,N_11038,N_11096);
and U11392 (N_11392,N_11176,N_11072);
nand U11393 (N_11393,N_11112,N_11151);
or U11394 (N_11394,N_11007,N_11181);
and U11395 (N_11395,N_11162,N_11028);
or U11396 (N_11396,N_11037,N_11076);
and U11397 (N_11397,N_11060,N_11124);
or U11398 (N_11398,N_11108,N_11062);
nor U11399 (N_11399,N_11129,N_11044);
xor U11400 (N_11400,N_11319,N_11271);
xor U11401 (N_11401,N_11299,N_11244);
and U11402 (N_11402,N_11283,N_11200);
nand U11403 (N_11403,N_11296,N_11362);
xor U11404 (N_11404,N_11209,N_11327);
nor U11405 (N_11405,N_11225,N_11398);
nor U11406 (N_11406,N_11323,N_11353);
nor U11407 (N_11407,N_11245,N_11379);
xor U11408 (N_11408,N_11221,N_11263);
xor U11409 (N_11409,N_11330,N_11346);
nor U11410 (N_11410,N_11358,N_11295);
or U11411 (N_11411,N_11356,N_11257);
nand U11412 (N_11412,N_11291,N_11348);
or U11413 (N_11413,N_11278,N_11369);
nand U11414 (N_11414,N_11277,N_11314);
nand U11415 (N_11415,N_11297,N_11241);
xor U11416 (N_11416,N_11266,N_11212);
nor U11417 (N_11417,N_11370,N_11325);
or U11418 (N_11418,N_11338,N_11233);
xor U11419 (N_11419,N_11280,N_11268);
nand U11420 (N_11420,N_11363,N_11269);
nor U11421 (N_11421,N_11276,N_11290);
or U11422 (N_11422,N_11343,N_11286);
or U11423 (N_11423,N_11273,N_11380);
and U11424 (N_11424,N_11249,N_11218);
or U11425 (N_11425,N_11267,N_11237);
or U11426 (N_11426,N_11252,N_11315);
nor U11427 (N_11427,N_11395,N_11216);
nand U11428 (N_11428,N_11377,N_11240);
or U11429 (N_11429,N_11376,N_11224);
xnor U11430 (N_11430,N_11384,N_11328);
or U11431 (N_11431,N_11382,N_11366);
xor U11432 (N_11432,N_11331,N_11208);
nor U11433 (N_11433,N_11349,N_11258);
xnor U11434 (N_11434,N_11372,N_11205);
xor U11435 (N_11435,N_11220,N_11235);
or U11436 (N_11436,N_11303,N_11270);
or U11437 (N_11437,N_11206,N_11204);
or U11438 (N_11438,N_11333,N_11246);
nand U11439 (N_11439,N_11207,N_11311);
nor U11440 (N_11440,N_11238,N_11371);
or U11441 (N_11441,N_11393,N_11318);
nor U11442 (N_11442,N_11236,N_11234);
nand U11443 (N_11443,N_11394,N_11306);
nand U11444 (N_11444,N_11274,N_11389);
nand U11445 (N_11445,N_11298,N_11375);
nor U11446 (N_11446,N_11254,N_11354);
nand U11447 (N_11447,N_11396,N_11392);
nand U11448 (N_11448,N_11391,N_11322);
and U11449 (N_11449,N_11340,N_11373);
and U11450 (N_11450,N_11344,N_11272);
nor U11451 (N_11451,N_11211,N_11347);
nor U11452 (N_11452,N_11386,N_11302);
or U11453 (N_11453,N_11201,N_11399);
and U11454 (N_11454,N_11219,N_11239);
nand U11455 (N_11455,N_11251,N_11329);
nor U11456 (N_11456,N_11289,N_11351);
nand U11457 (N_11457,N_11294,N_11214);
nand U11458 (N_11458,N_11223,N_11210);
xnor U11459 (N_11459,N_11364,N_11281);
nor U11460 (N_11460,N_11230,N_11305);
and U11461 (N_11461,N_11320,N_11222);
or U11462 (N_11462,N_11255,N_11374);
xnor U11463 (N_11463,N_11317,N_11350);
nand U11464 (N_11464,N_11253,N_11335);
nor U11465 (N_11465,N_11321,N_11326);
and U11466 (N_11466,N_11287,N_11313);
or U11467 (N_11467,N_11309,N_11361);
and U11468 (N_11468,N_11231,N_11334);
or U11469 (N_11469,N_11229,N_11381);
xor U11470 (N_11470,N_11316,N_11345);
xor U11471 (N_11471,N_11203,N_11378);
xor U11472 (N_11472,N_11310,N_11259);
nor U11473 (N_11473,N_11390,N_11284);
nand U11474 (N_11474,N_11265,N_11293);
and U11475 (N_11475,N_11262,N_11243);
nand U11476 (N_11476,N_11217,N_11368);
and U11477 (N_11477,N_11285,N_11388);
and U11478 (N_11478,N_11248,N_11359);
and U11479 (N_11479,N_11292,N_11275);
xnor U11480 (N_11480,N_11228,N_11339);
nor U11481 (N_11481,N_11301,N_11324);
xor U11482 (N_11482,N_11242,N_11387);
nand U11483 (N_11483,N_11227,N_11304);
nor U11484 (N_11484,N_11247,N_11308);
or U11485 (N_11485,N_11232,N_11385);
xor U11486 (N_11486,N_11337,N_11260);
nand U11487 (N_11487,N_11355,N_11215);
and U11488 (N_11488,N_11226,N_11365);
and U11489 (N_11489,N_11397,N_11312);
xnor U11490 (N_11490,N_11383,N_11264);
or U11491 (N_11491,N_11357,N_11341);
nand U11492 (N_11492,N_11202,N_11261);
nor U11493 (N_11493,N_11352,N_11342);
nand U11494 (N_11494,N_11213,N_11307);
or U11495 (N_11495,N_11336,N_11360);
xor U11496 (N_11496,N_11367,N_11256);
nand U11497 (N_11497,N_11300,N_11279);
and U11498 (N_11498,N_11288,N_11332);
xor U11499 (N_11499,N_11250,N_11282);
or U11500 (N_11500,N_11280,N_11219);
nand U11501 (N_11501,N_11314,N_11348);
nor U11502 (N_11502,N_11249,N_11358);
nand U11503 (N_11503,N_11386,N_11384);
nand U11504 (N_11504,N_11375,N_11309);
or U11505 (N_11505,N_11306,N_11305);
nor U11506 (N_11506,N_11215,N_11300);
nor U11507 (N_11507,N_11310,N_11277);
or U11508 (N_11508,N_11350,N_11383);
nand U11509 (N_11509,N_11394,N_11327);
or U11510 (N_11510,N_11395,N_11241);
nor U11511 (N_11511,N_11381,N_11208);
nand U11512 (N_11512,N_11381,N_11341);
nand U11513 (N_11513,N_11327,N_11343);
and U11514 (N_11514,N_11384,N_11217);
or U11515 (N_11515,N_11306,N_11261);
nor U11516 (N_11516,N_11363,N_11247);
nor U11517 (N_11517,N_11204,N_11200);
nor U11518 (N_11518,N_11335,N_11263);
xor U11519 (N_11519,N_11255,N_11257);
nor U11520 (N_11520,N_11295,N_11312);
and U11521 (N_11521,N_11323,N_11251);
or U11522 (N_11522,N_11204,N_11309);
nor U11523 (N_11523,N_11230,N_11285);
nand U11524 (N_11524,N_11254,N_11242);
nand U11525 (N_11525,N_11353,N_11237);
nor U11526 (N_11526,N_11236,N_11365);
nor U11527 (N_11527,N_11390,N_11294);
and U11528 (N_11528,N_11241,N_11330);
nand U11529 (N_11529,N_11228,N_11200);
nand U11530 (N_11530,N_11282,N_11244);
and U11531 (N_11531,N_11231,N_11378);
xnor U11532 (N_11532,N_11296,N_11220);
or U11533 (N_11533,N_11394,N_11248);
nand U11534 (N_11534,N_11213,N_11336);
nor U11535 (N_11535,N_11227,N_11220);
and U11536 (N_11536,N_11380,N_11392);
xor U11537 (N_11537,N_11269,N_11253);
nor U11538 (N_11538,N_11245,N_11275);
xnor U11539 (N_11539,N_11262,N_11329);
xor U11540 (N_11540,N_11208,N_11313);
xor U11541 (N_11541,N_11256,N_11318);
or U11542 (N_11542,N_11262,N_11363);
or U11543 (N_11543,N_11273,N_11220);
or U11544 (N_11544,N_11216,N_11253);
nor U11545 (N_11545,N_11363,N_11357);
nand U11546 (N_11546,N_11251,N_11306);
nor U11547 (N_11547,N_11231,N_11262);
xor U11548 (N_11548,N_11371,N_11203);
xor U11549 (N_11549,N_11220,N_11367);
and U11550 (N_11550,N_11277,N_11250);
nor U11551 (N_11551,N_11389,N_11287);
nand U11552 (N_11552,N_11365,N_11275);
nor U11553 (N_11553,N_11383,N_11217);
or U11554 (N_11554,N_11318,N_11374);
or U11555 (N_11555,N_11254,N_11370);
xnor U11556 (N_11556,N_11203,N_11369);
nor U11557 (N_11557,N_11372,N_11304);
nor U11558 (N_11558,N_11236,N_11256);
nor U11559 (N_11559,N_11249,N_11294);
and U11560 (N_11560,N_11250,N_11210);
nor U11561 (N_11561,N_11322,N_11365);
or U11562 (N_11562,N_11336,N_11343);
nor U11563 (N_11563,N_11287,N_11211);
nand U11564 (N_11564,N_11377,N_11367);
nand U11565 (N_11565,N_11202,N_11216);
xor U11566 (N_11566,N_11293,N_11304);
or U11567 (N_11567,N_11394,N_11226);
nor U11568 (N_11568,N_11209,N_11238);
xnor U11569 (N_11569,N_11253,N_11285);
xnor U11570 (N_11570,N_11225,N_11257);
nor U11571 (N_11571,N_11268,N_11214);
and U11572 (N_11572,N_11331,N_11308);
nand U11573 (N_11573,N_11318,N_11214);
and U11574 (N_11574,N_11348,N_11322);
or U11575 (N_11575,N_11346,N_11360);
or U11576 (N_11576,N_11278,N_11334);
xnor U11577 (N_11577,N_11201,N_11343);
and U11578 (N_11578,N_11268,N_11369);
and U11579 (N_11579,N_11363,N_11353);
and U11580 (N_11580,N_11306,N_11218);
xor U11581 (N_11581,N_11207,N_11261);
nor U11582 (N_11582,N_11285,N_11393);
nand U11583 (N_11583,N_11209,N_11232);
or U11584 (N_11584,N_11355,N_11358);
xnor U11585 (N_11585,N_11265,N_11260);
nand U11586 (N_11586,N_11318,N_11326);
or U11587 (N_11587,N_11238,N_11366);
or U11588 (N_11588,N_11349,N_11238);
xnor U11589 (N_11589,N_11309,N_11304);
and U11590 (N_11590,N_11391,N_11218);
and U11591 (N_11591,N_11286,N_11339);
xor U11592 (N_11592,N_11353,N_11367);
xor U11593 (N_11593,N_11316,N_11331);
and U11594 (N_11594,N_11304,N_11354);
and U11595 (N_11595,N_11346,N_11251);
or U11596 (N_11596,N_11348,N_11357);
or U11597 (N_11597,N_11331,N_11209);
and U11598 (N_11598,N_11299,N_11342);
nor U11599 (N_11599,N_11262,N_11210);
or U11600 (N_11600,N_11593,N_11441);
xnor U11601 (N_11601,N_11486,N_11404);
nand U11602 (N_11602,N_11500,N_11439);
nor U11603 (N_11603,N_11480,N_11401);
xnor U11604 (N_11604,N_11574,N_11564);
nand U11605 (N_11605,N_11563,N_11493);
and U11606 (N_11606,N_11478,N_11422);
nand U11607 (N_11607,N_11408,N_11565);
and U11608 (N_11608,N_11538,N_11470);
nand U11609 (N_11609,N_11561,N_11528);
nand U11610 (N_11610,N_11529,N_11590);
or U11611 (N_11611,N_11572,N_11598);
nand U11612 (N_11612,N_11535,N_11537);
nand U11613 (N_11613,N_11578,N_11418);
and U11614 (N_11614,N_11502,N_11458);
or U11615 (N_11615,N_11508,N_11497);
nand U11616 (N_11616,N_11550,N_11540);
nand U11617 (N_11617,N_11446,N_11510);
nor U11618 (N_11618,N_11543,N_11507);
and U11619 (N_11619,N_11440,N_11549);
nand U11620 (N_11620,N_11423,N_11551);
nand U11621 (N_11621,N_11424,N_11432);
xnor U11622 (N_11622,N_11585,N_11447);
nor U11623 (N_11623,N_11419,N_11456);
xnor U11624 (N_11624,N_11589,N_11442);
and U11625 (N_11625,N_11469,N_11496);
nor U11626 (N_11626,N_11444,N_11568);
xnor U11627 (N_11627,N_11426,N_11473);
nor U11628 (N_11628,N_11571,N_11438);
or U11629 (N_11629,N_11526,N_11567);
or U11630 (N_11630,N_11457,N_11466);
or U11631 (N_11631,N_11584,N_11521);
nand U11632 (N_11632,N_11556,N_11461);
or U11633 (N_11633,N_11481,N_11501);
xnor U11634 (N_11634,N_11494,N_11415);
xnor U11635 (N_11635,N_11489,N_11479);
nor U11636 (N_11636,N_11580,N_11450);
nor U11637 (N_11637,N_11587,N_11455);
and U11638 (N_11638,N_11428,N_11558);
and U11639 (N_11639,N_11517,N_11490);
nand U11640 (N_11640,N_11531,N_11525);
or U11641 (N_11641,N_11506,N_11512);
xor U11642 (N_11642,N_11462,N_11474);
or U11643 (N_11643,N_11464,N_11454);
xor U11644 (N_11644,N_11575,N_11583);
and U11645 (N_11645,N_11421,N_11449);
xnor U11646 (N_11646,N_11505,N_11542);
xor U11647 (N_11647,N_11483,N_11523);
xor U11648 (N_11648,N_11416,N_11488);
xnor U11649 (N_11649,N_11557,N_11579);
xor U11650 (N_11650,N_11524,N_11569);
and U11651 (N_11651,N_11541,N_11536);
and U11652 (N_11652,N_11471,N_11453);
nand U11653 (N_11653,N_11425,N_11554);
or U11654 (N_11654,N_11485,N_11520);
nand U11655 (N_11655,N_11463,N_11492);
and U11656 (N_11656,N_11576,N_11553);
nor U11657 (N_11657,N_11592,N_11532);
nor U11658 (N_11658,N_11559,N_11511);
xnor U11659 (N_11659,N_11433,N_11588);
or U11660 (N_11660,N_11434,N_11599);
nand U11661 (N_11661,N_11594,N_11468);
or U11662 (N_11662,N_11465,N_11487);
nand U11663 (N_11663,N_11555,N_11431);
nor U11664 (N_11664,N_11445,N_11499);
nand U11665 (N_11665,N_11527,N_11548);
or U11666 (N_11666,N_11427,N_11443);
nand U11667 (N_11667,N_11591,N_11566);
nand U11668 (N_11668,N_11546,N_11400);
nor U11669 (N_11669,N_11503,N_11515);
nor U11670 (N_11670,N_11484,N_11477);
nor U11671 (N_11671,N_11498,N_11534);
xnor U11672 (N_11672,N_11452,N_11430);
or U11673 (N_11673,N_11435,N_11417);
xor U11674 (N_11674,N_11544,N_11516);
or U11675 (N_11675,N_11406,N_11581);
and U11676 (N_11676,N_11519,N_11402);
xnor U11677 (N_11677,N_11411,N_11562);
and U11678 (N_11678,N_11595,N_11573);
xnor U11679 (N_11679,N_11533,N_11405);
or U11680 (N_11680,N_11475,N_11545);
nor U11681 (N_11681,N_11577,N_11403);
nand U11682 (N_11682,N_11491,N_11570);
xor U11683 (N_11683,N_11539,N_11459);
and U11684 (N_11684,N_11509,N_11460);
and U11685 (N_11685,N_11504,N_11451);
xnor U11686 (N_11686,N_11518,N_11552);
xor U11687 (N_11687,N_11414,N_11597);
and U11688 (N_11688,N_11530,N_11413);
nor U11689 (N_11689,N_11522,N_11436);
xor U11690 (N_11690,N_11472,N_11410);
xor U11691 (N_11691,N_11513,N_11547);
nor U11692 (N_11692,N_11448,N_11596);
xnor U11693 (N_11693,N_11495,N_11582);
nor U11694 (N_11694,N_11476,N_11514);
nor U11695 (N_11695,N_11586,N_11429);
xor U11696 (N_11696,N_11437,N_11409);
xor U11697 (N_11697,N_11412,N_11420);
and U11698 (N_11698,N_11482,N_11467);
xor U11699 (N_11699,N_11407,N_11560);
or U11700 (N_11700,N_11488,N_11486);
and U11701 (N_11701,N_11516,N_11565);
xor U11702 (N_11702,N_11463,N_11579);
nand U11703 (N_11703,N_11485,N_11400);
and U11704 (N_11704,N_11585,N_11519);
and U11705 (N_11705,N_11523,N_11465);
nand U11706 (N_11706,N_11470,N_11483);
or U11707 (N_11707,N_11586,N_11451);
nand U11708 (N_11708,N_11547,N_11552);
and U11709 (N_11709,N_11550,N_11463);
nand U11710 (N_11710,N_11499,N_11500);
or U11711 (N_11711,N_11536,N_11498);
xor U11712 (N_11712,N_11495,N_11574);
nor U11713 (N_11713,N_11557,N_11444);
nor U11714 (N_11714,N_11498,N_11508);
nor U11715 (N_11715,N_11410,N_11581);
nor U11716 (N_11716,N_11541,N_11595);
and U11717 (N_11717,N_11407,N_11541);
nor U11718 (N_11718,N_11438,N_11514);
or U11719 (N_11719,N_11554,N_11447);
xnor U11720 (N_11720,N_11465,N_11504);
xor U11721 (N_11721,N_11568,N_11555);
nand U11722 (N_11722,N_11481,N_11411);
nand U11723 (N_11723,N_11568,N_11508);
and U11724 (N_11724,N_11538,N_11477);
or U11725 (N_11725,N_11457,N_11482);
or U11726 (N_11726,N_11431,N_11548);
or U11727 (N_11727,N_11542,N_11478);
and U11728 (N_11728,N_11581,N_11451);
xor U11729 (N_11729,N_11512,N_11521);
nand U11730 (N_11730,N_11462,N_11583);
nor U11731 (N_11731,N_11530,N_11500);
and U11732 (N_11732,N_11410,N_11437);
nor U11733 (N_11733,N_11547,N_11489);
nor U11734 (N_11734,N_11552,N_11409);
nand U11735 (N_11735,N_11570,N_11468);
nand U11736 (N_11736,N_11566,N_11479);
xor U11737 (N_11737,N_11471,N_11489);
xnor U11738 (N_11738,N_11574,N_11593);
or U11739 (N_11739,N_11597,N_11581);
or U11740 (N_11740,N_11551,N_11495);
or U11741 (N_11741,N_11427,N_11563);
nor U11742 (N_11742,N_11472,N_11560);
xnor U11743 (N_11743,N_11423,N_11549);
or U11744 (N_11744,N_11493,N_11430);
nor U11745 (N_11745,N_11450,N_11406);
or U11746 (N_11746,N_11483,N_11404);
nor U11747 (N_11747,N_11431,N_11572);
nor U11748 (N_11748,N_11403,N_11561);
nand U11749 (N_11749,N_11548,N_11475);
or U11750 (N_11750,N_11587,N_11450);
xnor U11751 (N_11751,N_11430,N_11492);
nor U11752 (N_11752,N_11590,N_11585);
nand U11753 (N_11753,N_11577,N_11528);
and U11754 (N_11754,N_11568,N_11573);
or U11755 (N_11755,N_11512,N_11421);
nor U11756 (N_11756,N_11502,N_11571);
nand U11757 (N_11757,N_11580,N_11590);
nand U11758 (N_11758,N_11524,N_11537);
nor U11759 (N_11759,N_11575,N_11489);
nand U11760 (N_11760,N_11493,N_11485);
and U11761 (N_11761,N_11526,N_11472);
or U11762 (N_11762,N_11570,N_11523);
xnor U11763 (N_11763,N_11552,N_11473);
and U11764 (N_11764,N_11450,N_11418);
or U11765 (N_11765,N_11429,N_11545);
and U11766 (N_11766,N_11473,N_11490);
nand U11767 (N_11767,N_11486,N_11541);
nor U11768 (N_11768,N_11438,N_11401);
nand U11769 (N_11769,N_11454,N_11582);
nand U11770 (N_11770,N_11434,N_11563);
nand U11771 (N_11771,N_11400,N_11596);
nand U11772 (N_11772,N_11470,N_11443);
nor U11773 (N_11773,N_11456,N_11565);
nor U11774 (N_11774,N_11450,N_11428);
nor U11775 (N_11775,N_11460,N_11504);
xor U11776 (N_11776,N_11524,N_11525);
nor U11777 (N_11777,N_11546,N_11450);
nand U11778 (N_11778,N_11502,N_11544);
xnor U11779 (N_11779,N_11551,N_11414);
nand U11780 (N_11780,N_11517,N_11454);
and U11781 (N_11781,N_11427,N_11502);
and U11782 (N_11782,N_11514,N_11491);
and U11783 (N_11783,N_11447,N_11495);
and U11784 (N_11784,N_11552,N_11416);
nor U11785 (N_11785,N_11552,N_11415);
xor U11786 (N_11786,N_11532,N_11527);
and U11787 (N_11787,N_11447,N_11469);
nor U11788 (N_11788,N_11504,N_11475);
xor U11789 (N_11789,N_11435,N_11406);
and U11790 (N_11790,N_11448,N_11409);
nand U11791 (N_11791,N_11537,N_11428);
and U11792 (N_11792,N_11462,N_11421);
nor U11793 (N_11793,N_11475,N_11473);
nand U11794 (N_11794,N_11429,N_11597);
nand U11795 (N_11795,N_11586,N_11532);
nor U11796 (N_11796,N_11521,N_11502);
and U11797 (N_11797,N_11553,N_11428);
xnor U11798 (N_11798,N_11582,N_11598);
xor U11799 (N_11799,N_11564,N_11494);
and U11800 (N_11800,N_11751,N_11663);
and U11801 (N_11801,N_11610,N_11728);
nand U11802 (N_11802,N_11770,N_11780);
nand U11803 (N_11803,N_11744,N_11771);
or U11804 (N_11804,N_11692,N_11773);
nand U11805 (N_11805,N_11726,N_11667);
nand U11806 (N_11806,N_11603,N_11644);
or U11807 (N_11807,N_11746,N_11627);
and U11808 (N_11808,N_11750,N_11641);
xnor U11809 (N_11809,N_11697,N_11732);
and U11810 (N_11810,N_11614,N_11607);
nor U11811 (N_11811,N_11690,N_11688);
nand U11812 (N_11812,N_11649,N_11685);
nand U11813 (N_11813,N_11789,N_11735);
xnor U11814 (N_11814,N_11643,N_11619);
or U11815 (N_11815,N_11752,N_11717);
nor U11816 (N_11816,N_11673,N_11689);
nand U11817 (N_11817,N_11777,N_11768);
or U11818 (N_11818,N_11714,N_11748);
xor U11819 (N_11819,N_11753,N_11708);
or U11820 (N_11820,N_11631,N_11754);
and U11821 (N_11821,N_11675,N_11785);
or U11822 (N_11822,N_11760,N_11799);
or U11823 (N_11823,N_11624,N_11656);
or U11824 (N_11824,N_11794,N_11783);
xor U11825 (N_11825,N_11615,N_11602);
xnor U11826 (N_11826,N_11634,N_11694);
xor U11827 (N_11827,N_11740,N_11775);
and U11828 (N_11828,N_11761,N_11616);
nand U11829 (N_11829,N_11787,N_11764);
and U11830 (N_11830,N_11719,N_11763);
nor U11831 (N_11831,N_11716,N_11796);
nand U11832 (N_11832,N_11755,N_11696);
nor U11833 (N_11833,N_11622,N_11629);
nor U11834 (N_11834,N_11762,N_11670);
nor U11835 (N_11835,N_11691,N_11757);
or U11836 (N_11836,N_11782,N_11654);
and U11837 (N_11837,N_11666,N_11661);
nand U11838 (N_11838,N_11650,N_11605);
nor U11839 (N_11839,N_11766,N_11680);
nor U11840 (N_11840,N_11684,N_11682);
or U11841 (N_11841,N_11635,N_11638);
or U11842 (N_11842,N_11679,N_11671);
and U11843 (N_11843,N_11628,N_11729);
or U11844 (N_11844,N_11797,N_11738);
and U11845 (N_11845,N_11640,N_11779);
nor U11846 (N_11846,N_11723,N_11788);
xnor U11847 (N_11847,N_11672,N_11645);
nand U11848 (N_11848,N_11778,N_11711);
and U11849 (N_11849,N_11699,N_11608);
nand U11850 (N_11850,N_11646,N_11706);
xnor U11851 (N_11851,N_11659,N_11625);
nor U11852 (N_11852,N_11657,N_11677);
nand U11853 (N_11853,N_11705,N_11664);
xnor U11854 (N_11854,N_11665,N_11623);
nor U11855 (N_11855,N_11745,N_11715);
and U11856 (N_11856,N_11700,N_11759);
and U11857 (N_11857,N_11724,N_11687);
xor U11858 (N_11858,N_11639,N_11718);
nand U11859 (N_11859,N_11713,N_11731);
xnor U11860 (N_11860,N_11648,N_11668);
nand U11861 (N_11861,N_11736,N_11791);
and U11862 (N_11862,N_11756,N_11707);
and U11863 (N_11863,N_11693,N_11606);
and U11864 (N_11864,N_11795,N_11765);
and U11865 (N_11865,N_11734,N_11793);
nor U11866 (N_11866,N_11747,N_11655);
and U11867 (N_11867,N_11609,N_11686);
or U11868 (N_11868,N_11636,N_11758);
or U11869 (N_11869,N_11651,N_11702);
nand U11870 (N_11870,N_11642,N_11601);
xnor U11871 (N_11871,N_11722,N_11769);
xnor U11872 (N_11872,N_11767,N_11683);
or U11873 (N_11873,N_11709,N_11674);
and U11874 (N_11874,N_11660,N_11612);
and U11875 (N_11875,N_11786,N_11698);
xnor U11876 (N_11876,N_11617,N_11781);
xor U11877 (N_11877,N_11695,N_11703);
or U11878 (N_11878,N_11630,N_11743);
and U11879 (N_11879,N_11637,N_11681);
xnor U11880 (N_11880,N_11749,N_11613);
xnor U11881 (N_11881,N_11647,N_11669);
nand U11882 (N_11882,N_11712,N_11725);
xnor U11883 (N_11883,N_11658,N_11704);
xnor U11884 (N_11884,N_11772,N_11633);
nor U11885 (N_11885,N_11737,N_11632);
and U11886 (N_11886,N_11792,N_11600);
and U11887 (N_11887,N_11733,N_11730);
xnor U11888 (N_11888,N_11626,N_11678);
nand U11889 (N_11889,N_11720,N_11662);
or U11890 (N_11890,N_11790,N_11784);
nand U11891 (N_11891,N_11727,N_11721);
xor U11892 (N_11892,N_11621,N_11653);
nand U11893 (N_11893,N_11739,N_11776);
nor U11894 (N_11894,N_11701,N_11676);
and U11895 (N_11895,N_11652,N_11742);
xor U11896 (N_11896,N_11741,N_11620);
or U11897 (N_11897,N_11774,N_11798);
nand U11898 (N_11898,N_11611,N_11618);
and U11899 (N_11899,N_11604,N_11710);
nand U11900 (N_11900,N_11636,N_11799);
xor U11901 (N_11901,N_11777,N_11749);
or U11902 (N_11902,N_11726,N_11643);
nor U11903 (N_11903,N_11639,N_11787);
xor U11904 (N_11904,N_11603,N_11661);
nand U11905 (N_11905,N_11702,N_11664);
nand U11906 (N_11906,N_11647,N_11637);
and U11907 (N_11907,N_11709,N_11731);
nand U11908 (N_11908,N_11719,N_11681);
or U11909 (N_11909,N_11703,N_11655);
xnor U11910 (N_11910,N_11710,N_11672);
xnor U11911 (N_11911,N_11658,N_11789);
and U11912 (N_11912,N_11631,N_11630);
or U11913 (N_11913,N_11762,N_11721);
or U11914 (N_11914,N_11700,N_11685);
or U11915 (N_11915,N_11654,N_11632);
and U11916 (N_11916,N_11735,N_11682);
and U11917 (N_11917,N_11638,N_11741);
or U11918 (N_11918,N_11667,N_11635);
xor U11919 (N_11919,N_11675,N_11797);
and U11920 (N_11920,N_11790,N_11676);
nor U11921 (N_11921,N_11752,N_11720);
xnor U11922 (N_11922,N_11768,N_11606);
and U11923 (N_11923,N_11691,N_11741);
and U11924 (N_11924,N_11765,N_11611);
or U11925 (N_11925,N_11654,N_11614);
nor U11926 (N_11926,N_11715,N_11769);
or U11927 (N_11927,N_11710,N_11722);
nor U11928 (N_11928,N_11706,N_11688);
nor U11929 (N_11929,N_11686,N_11782);
xor U11930 (N_11930,N_11607,N_11798);
xnor U11931 (N_11931,N_11745,N_11743);
nor U11932 (N_11932,N_11730,N_11640);
nand U11933 (N_11933,N_11793,N_11681);
nor U11934 (N_11934,N_11701,N_11799);
nor U11935 (N_11935,N_11671,N_11648);
nor U11936 (N_11936,N_11677,N_11751);
and U11937 (N_11937,N_11727,N_11632);
nor U11938 (N_11938,N_11636,N_11714);
xor U11939 (N_11939,N_11656,N_11654);
nand U11940 (N_11940,N_11798,N_11696);
or U11941 (N_11941,N_11702,N_11649);
nor U11942 (N_11942,N_11758,N_11743);
nand U11943 (N_11943,N_11728,N_11640);
xor U11944 (N_11944,N_11715,N_11604);
nor U11945 (N_11945,N_11759,N_11679);
nand U11946 (N_11946,N_11765,N_11655);
xor U11947 (N_11947,N_11667,N_11742);
and U11948 (N_11948,N_11643,N_11671);
nand U11949 (N_11949,N_11709,N_11644);
and U11950 (N_11950,N_11699,N_11775);
xnor U11951 (N_11951,N_11626,N_11637);
nand U11952 (N_11952,N_11741,N_11742);
or U11953 (N_11953,N_11671,N_11799);
or U11954 (N_11954,N_11777,N_11612);
nand U11955 (N_11955,N_11761,N_11794);
nand U11956 (N_11956,N_11644,N_11624);
nor U11957 (N_11957,N_11701,N_11689);
and U11958 (N_11958,N_11648,N_11714);
xor U11959 (N_11959,N_11641,N_11638);
and U11960 (N_11960,N_11692,N_11619);
nor U11961 (N_11961,N_11755,N_11621);
or U11962 (N_11962,N_11641,N_11663);
and U11963 (N_11963,N_11724,N_11612);
nor U11964 (N_11964,N_11625,N_11620);
and U11965 (N_11965,N_11724,N_11646);
nand U11966 (N_11966,N_11689,N_11627);
nor U11967 (N_11967,N_11769,N_11613);
nand U11968 (N_11968,N_11714,N_11780);
nor U11969 (N_11969,N_11717,N_11604);
nand U11970 (N_11970,N_11647,N_11656);
or U11971 (N_11971,N_11713,N_11792);
and U11972 (N_11972,N_11719,N_11674);
or U11973 (N_11973,N_11718,N_11770);
or U11974 (N_11974,N_11644,N_11745);
or U11975 (N_11975,N_11747,N_11658);
and U11976 (N_11976,N_11771,N_11644);
nand U11977 (N_11977,N_11752,N_11710);
xnor U11978 (N_11978,N_11625,N_11640);
nor U11979 (N_11979,N_11722,N_11641);
nor U11980 (N_11980,N_11697,N_11730);
nand U11981 (N_11981,N_11628,N_11604);
nor U11982 (N_11982,N_11620,N_11733);
and U11983 (N_11983,N_11719,N_11706);
and U11984 (N_11984,N_11702,N_11797);
and U11985 (N_11985,N_11622,N_11776);
or U11986 (N_11986,N_11791,N_11787);
and U11987 (N_11987,N_11716,N_11600);
nand U11988 (N_11988,N_11717,N_11636);
nor U11989 (N_11989,N_11733,N_11657);
xnor U11990 (N_11990,N_11654,N_11641);
xor U11991 (N_11991,N_11711,N_11771);
nand U11992 (N_11992,N_11747,N_11682);
or U11993 (N_11993,N_11779,N_11613);
nor U11994 (N_11994,N_11627,N_11657);
xnor U11995 (N_11995,N_11713,N_11680);
or U11996 (N_11996,N_11785,N_11609);
or U11997 (N_11997,N_11719,N_11729);
nand U11998 (N_11998,N_11601,N_11644);
or U11999 (N_11999,N_11791,N_11667);
nor U12000 (N_12000,N_11987,N_11988);
xnor U12001 (N_12001,N_11927,N_11800);
xnor U12002 (N_12002,N_11959,N_11999);
nand U12003 (N_12003,N_11836,N_11841);
xor U12004 (N_12004,N_11881,N_11819);
or U12005 (N_12005,N_11886,N_11972);
and U12006 (N_12006,N_11816,N_11901);
and U12007 (N_12007,N_11880,N_11813);
and U12008 (N_12008,N_11818,N_11829);
nor U12009 (N_12009,N_11846,N_11820);
nor U12010 (N_12010,N_11909,N_11843);
nor U12011 (N_12011,N_11848,N_11957);
xor U12012 (N_12012,N_11981,N_11810);
nand U12013 (N_12013,N_11899,N_11921);
xnor U12014 (N_12014,N_11929,N_11907);
xor U12015 (N_12015,N_11885,N_11941);
or U12016 (N_12016,N_11996,N_11809);
and U12017 (N_12017,N_11857,N_11939);
nor U12018 (N_12018,N_11815,N_11905);
xor U12019 (N_12019,N_11982,N_11855);
nand U12020 (N_12020,N_11943,N_11863);
and U12021 (N_12021,N_11891,N_11940);
or U12022 (N_12022,N_11969,N_11938);
nor U12023 (N_12023,N_11887,N_11835);
nand U12024 (N_12024,N_11871,N_11903);
nor U12025 (N_12025,N_11971,N_11961);
or U12026 (N_12026,N_11849,N_11878);
nand U12027 (N_12027,N_11873,N_11944);
nor U12028 (N_12028,N_11934,N_11928);
nand U12029 (N_12029,N_11931,N_11882);
nor U12030 (N_12030,N_11974,N_11898);
nor U12031 (N_12031,N_11842,N_11875);
nand U12032 (N_12032,N_11935,N_11990);
nor U12033 (N_12033,N_11801,N_11922);
xnor U12034 (N_12034,N_11869,N_11844);
and U12035 (N_12035,N_11883,N_11989);
or U12036 (N_12036,N_11992,N_11917);
or U12037 (N_12037,N_11879,N_11906);
or U12038 (N_12038,N_11876,N_11805);
nor U12039 (N_12039,N_11954,N_11868);
xor U12040 (N_12040,N_11867,N_11978);
or U12041 (N_12041,N_11908,N_11824);
and U12042 (N_12042,N_11806,N_11980);
or U12043 (N_12043,N_11986,N_11822);
and U12044 (N_12044,N_11919,N_11930);
and U12045 (N_12045,N_11968,N_11918);
nor U12046 (N_12046,N_11893,N_11832);
and U12047 (N_12047,N_11812,N_11942);
nor U12048 (N_12048,N_11933,N_11964);
or U12049 (N_12049,N_11834,N_11993);
or U12050 (N_12050,N_11897,N_11946);
nor U12051 (N_12051,N_11896,N_11932);
or U12052 (N_12052,N_11977,N_11924);
nand U12053 (N_12053,N_11960,N_11970);
or U12054 (N_12054,N_11973,N_11851);
nand U12055 (N_12055,N_11870,N_11975);
or U12056 (N_12056,N_11866,N_11865);
xnor U12057 (N_12057,N_11902,N_11884);
xor U12058 (N_12058,N_11953,N_11847);
xor U12059 (N_12059,N_11952,N_11831);
nand U12060 (N_12060,N_11825,N_11966);
or U12061 (N_12061,N_11998,N_11888);
xor U12062 (N_12062,N_11874,N_11923);
nand U12063 (N_12063,N_11828,N_11913);
and U12064 (N_12064,N_11861,N_11955);
or U12065 (N_12065,N_11900,N_11925);
xnor U12066 (N_12066,N_11949,N_11811);
nor U12067 (N_12067,N_11951,N_11963);
nor U12068 (N_12068,N_11991,N_11948);
nor U12069 (N_12069,N_11804,N_11823);
or U12070 (N_12070,N_11833,N_11864);
nor U12071 (N_12071,N_11856,N_11950);
xnor U12072 (N_12072,N_11912,N_11814);
or U12073 (N_12073,N_11817,N_11936);
xor U12074 (N_12074,N_11956,N_11854);
or U12075 (N_12075,N_11872,N_11808);
xor U12076 (N_12076,N_11997,N_11937);
and U12077 (N_12077,N_11916,N_11904);
xnor U12078 (N_12078,N_11807,N_11994);
nor U12079 (N_12079,N_11895,N_11860);
xor U12080 (N_12080,N_11889,N_11850);
nand U12081 (N_12081,N_11985,N_11839);
nor U12082 (N_12082,N_11984,N_11976);
nand U12083 (N_12083,N_11995,N_11920);
or U12084 (N_12084,N_11945,N_11853);
xnor U12085 (N_12085,N_11858,N_11827);
and U12086 (N_12086,N_11830,N_11862);
nand U12087 (N_12087,N_11859,N_11821);
or U12088 (N_12088,N_11915,N_11845);
nand U12089 (N_12089,N_11983,N_11838);
or U12090 (N_12090,N_11826,N_11967);
xor U12091 (N_12091,N_11803,N_11802);
nand U12092 (N_12092,N_11911,N_11837);
xnor U12093 (N_12093,N_11926,N_11877);
or U12094 (N_12094,N_11852,N_11962);
nor U12095 (N_12095,N_11890,N_11958);
nor U12096 (N_12096,N_11910,N_11840);
nor U12097 (N_12097,N_11965,N_11914);
nor U12098 (N_12098,N_11979,N_11892);
and U12099 (N_12099,N_11947,N_11894);
nand U12100 (N_12100,N_11854,N_11868);
nor U12101 (N_12101,N_11981,N_11851);
nor U12102 (N_12102,N_11893,N_11884);
xnor U12103 (N_12103,N_11886,N_11802);
and U12104 (N_12104,N_11965,N_11853);
or U12105 (N_12105,N_11916,N_11997);
or U12106 (N_12106,N_11858,N_11811);
xor U12107 (N_12107,N_11908,N_11809);
xnor U12108 (N_12108,N_11937,N_11994);
or U12109 (N_12109,N_11941,N_11894);
and U12110 (N_12110,N_11964,N_11852);
nor U12111 (N_12111,N_11945,N_11824);
nor U12112 (N_12112,N_11815,N_11910);
and U12113 (N_12113,N_11818,N_11802);
xnor U12114 (N_12114,N_11978,N_11887);
xnor U12115 (N_12115,N_11812,N_11840);
nand U12116 (N_12116,N_11899,N_11983);
nor U12117 (N_12117,N_11808,N_11853);
xnor U12118 (N_12118,N_11869,N_11971);
and U12119 (N_12119,N_11881,N_11942);
or U12120 (N_12120,N_11838,N_11988);
nand U12121 (N_12121,N_11849,N_11980);
or U12122 (N_12122,N_11869,N_11961);
or U12123 (N_12123,N_11804,N_11882);
or U12124 (N_12124,N_11930,N_11814);
xor U12125 (N_12125,N_11952,N_11933);
nand U12126 (N_12126,N_11990,N_11932);
xnor U12127 (N_12127,N_11808,N_11848);
or U12128 (N_12128,N_11931,N_11871);
and U12129 (N_12129,N_11853,N_11949);
nand U12130 (N_12130,N_11901,N_11995);
nor U12131 (N_12131,N_11938,N_11856);
nand U12132 (N_12132,N_11820,N_11879);
xor U12133 (N_12133,N_11922,N_11837);
and U12134 (N_12134,N_11966,N_11885);
nand U12135 (N_12135,N_11998,N_11807);
nand U12136 (N_12136,N_11953,N_11921);
and U12137 (N_12137,N_11913,N_11888);
nand U12138 (N_12138,N_11953,N_11845);
and U12139 (N_12139,N_11833,N_11924);
and U12140 (N_12140,N_11950,N_11854);
nor U12141 (N_12141,N_11837,N_11944);
nand U12142 (N_12142,N_11906,N_11987);
xor U12143 (N_12143,N_11932,N_11924);
and U12144 (N_12144,N_11802,N_11817);
and U12145 (N_12145,N_11848,N_11831);
nand U12146 (N_12146,N_11867,N_11847);
and U12147 (N_12147,N_11889,N_11986);
and U12148 (N_12148,N_11862,N_11803);
xnor U12149 (N_12149,N_11898,N_11806);
or U12150 (N_12150,N_11872,N_11820);
and U12151 (N_12151,N_11888,N_11926);
xor U12152 (N_12152,N_11977,N_11917);
and U12153 (N_12153,N_11860,N_11901);
xnor U12154 (N_12154,N_11885,N_11827);
xnor U12155 (N_12155,N_11839,N_11908);
xor U12156 (N_12156,N_11995,N_11935);
xor U12157 (N_12157,N_11905,N_11964);
nand U12158 (N_12158,N_11990,N_11969);
nor U12159 (N_12159,N_11985,N_11918);
nor U12160 (N_12160,N_11800,N_11834);
and U12161 (N_12161,N_11936,N_11802);
nor U12162 (N_12162,N_11947,N_11935);
or U12163 (N_12163,N_11850,N_11897);
xnor U12164 (N_12164,N_11921,N_11950);
and U12165 (N_12165,N_11926,N_11825);
nor U12166 (N_12166,N_11830,N_11802);
or U12167 (N_12167,N_11975,N_11873);
nor U12168 (N_12168,N_11988,N_11966);
or U12169 (N_12169,N_11825,N_11981);
nand U12170 (N_12170,N_11929,N_11996);
and U12171 (N_12171,N_11891,N_11992);
and U12172 (N_12172,N_11996,N_11964);
and U12173 (N_12173,N_11873,N_11801);
nand U12174 (N_12174,N_11825,N_11828);
and U12175 (N_12175,N_11927,N_11882);
nor U12176 (N_12176,N_11952,N_11873);
nor U12177 (N_12177,N_11862,N_11956);
nand U12178 (N_12178,N_11957,N_11821);
nor U12179 (N_12179,N_11841,N_11831);
xor U12180 (N_12180,N_11986,N_11933);
nand U12181 (N_12181,N_11818,N_11925);
nand U12182 (N_12182,N_11851,N_11814);
nor U12183 (N_12183,N_11879,N_11985);
nor U12184 (N_12184,N_11984,N_11931);
or U12185 (N_12185,N_11854,N_11968);
nand U12186 (N_12186,N_11874,N_11975);
xor U12187 (N_12187,N_11978,N_11876);
nand U12188 (N_12188,N_11983,N_11941);
xor U12189 (N_12189,N_11818,N_11861);
and U12190 (N_12190,N_11952,N_11983);
xor U12191 (N_12191,N_11979,N_11888);
or U12192 (N_12192,N_11806,N_11997);
and U12193 (N_12193,N_11802,N_11898);
nor U12194 (N_12194,N_11942,N_11955);
nand U12195 (N_12195,N_11949,N_11987);
nand U12196 (N_12196,N_11936,N_11937);
and U12197 (N_12197,N_11897,N_11912);
and U12198 (N_12198,N_11811,N_11845);
and U12199 (N_12199,N_11914,N_11969);
or U12200 (N_12200,N_12056,N_12032);
and U12201 (N_12201,N_12130,N_12080);
or U12202 (N_12202,N_12180,N_12091);
nor U12203 (N_12203,N_12093,N_12144);
xnor U12204 (N_12204,N_12078,N_12189);
xor U12205 (N_12205,N_12148,N_12063);
nand U12206 (N_12206,N_12003,N_12147);
nor U12207 (N_12207,N_12060,N_12145);
xnor U12208 (N_12208,N_12140,N_12134);
and U12209 (N_12209,N_12036,N_12132);
nand U12210 (N_12210,N_12109,N_12046);
xor U12211 (N_12211,N_12156,N_12016);
nor U12212 (N_12212,N_12164,N_12153);
xnor U12213 (N_12213,N_12123,N_12191);
nand U12214 (N_12214,N_12054,N_12021);
nand U12215 (N_12215,N_12157,N_12069);
xnor U12216 (N_12216,N_12150,N_12182);
nand U12217 (N_12217,N_12135,N_12065);
xnor U12218 (N_12218,N_12126,N_12187);
nor U12219 (N_12219,N_12117,N_12040);
nand U12220 (N_12220,N_12152,N_12105);
nand U12221 (N_12221,N_12181,N_12029);
xnor U12222 (N_12222,N_12172,N_12097);
nand U12223 (N_12223,N_12088,N_12111);
or U12224 (N_12224,N_12095,N_12124);
or U12225 (N_12225,N_12163,N_12002);
nand U12226 (N_12226,N_12106,N_12050);
xnor U12227 (N_12227,N_12007,N_12179);
and U12228 (N_12228,N_12121,N_12118);
xnor U12229 (N_12229,N_12012,N_12011);
or U12230 (N_12230,N_12115,N_12096);
and U12231 (N_12231,N_12155,N_12197);
xnor U12232 (N_12232,N_12188,N_12034);
nand U12233 (N_12233,N_12185,N_12039);
and U12234 (N_12234,N_12049,N_12186);
and U12235 (N_12235,N_12005,N_12042);
nor U12236 (N_12236,N_12061,N_12072);
xnor U12237 (N_12237,N_12128,N_12085);
and U12238 (N_12238,N_12077,N_12141);
nor U12239 (N_12239,N_12161,N_12070);
nor U12240 (N_12240,N_12138,N_12024);
or U12241 (N_12241,N_12103,N_12000);
nor U12242 (N_12242,N_12110,N_12025);
nor U12243 (N_12243,N_12166,N_12139);
and U12244 (N_12244,N_12009,N_12019);
or U12245 (N_12245,N_12073,N_12099);
nor U12246 (N_12246,N_12041,N_12053);
nand U12247 (N_12247,N_12031,N_12127);
and U12248 (N_12248,N_12030,N_12165);
or U12249 (N_12249,N_12014,N_12146);
or U12250 (N_12250,N_12159,N_12055);
nand U12251 (N_12251,N_12028,N_12169);
and U12252 (N_12252,N_12116,N_12154);
xor U12253 (N_12253,N_12047,N_12120);
or U12254 (N_12254,N_12066,N_12190);
nand U12255 (N_12255,N_12195,N_12086);
nor U12256 (N_12256,N_12044,N_12052);
nand U12257 (N_12257,N_12058,N_12089);
nor U12258 (N_12258,N_12175,N_12017);
xnor U12259 (N_12259,N_12081,N_12125);
xnor U12260 (N_12260,N_12136,N_12162);
nand U12261 (N_12261,N_12168,N_12033);
xor U12262 (N_12262,N_12177,N_12022);
nand U12263 (N_12263,N_12059,N_12026);
and U12264 (N_12264,N_12149,N_12020);
and U12265 (N_12265,N_12129,N_12083);
nand U12266 (N_12266,N_12075,N_12027);
and U12267 (N_12267,N_12067,N_12004);
and U12268 (N_12268,N_12107,N_12018);
or U12269 (N_12269,N_12114,N_12074);
or U12270 (N_12270,N_12167,N_12001);
or U12271 (N_12271,N_12119,N_12023);
xnor U12272 (N_12272,N_12196,N_12015);
nor U12273 (N_12273,N_12006,N_12192);
nor U12274 (N_12274,N_12194,N_12198);
xor U12275 (N_12275,N_12170,N_12100);
and U12276 (N_12276,N_12184,N_12101);
nor U12277 (N_12277,N_12090,N_12158);
nor U12278 (N_12278,N_12104,N_12122);
or U12279 (N_12279,N_12176,N_12143);
nor U12280 (N_12280,N_12112,N_12057);
nor U12281 (N_12281,N_12102,N_12193);
or U12282 (N_12282,N_12171,N_12051);
and U12283 (N_12283,N_12048,N_12076);
xor U12284 (N_12284,N_12173,N_12113);
xnor U12285 (N_12285,N_12199,N_12013);
nand U12286 (N_12286,N_12108,N_12160);
nor U12287 (N_12287,N_12062,N_12098);
nor U12288 (N_12288,N_12037,N_12183);
nand U12289 (N_12289,N_12178,N_12092);
and U12290 (N_12290,N_12043,N_12038);
xnor U12291 (N_12291,N_12151,N_12094);
and U12292 (N_12292,N_12133,N_12084);
and U12293 (N_12293,N_12045,N_12079);
nor U12294 (N_12294,N_12035,N_12082);
and U12295 (N_12295,N_12064,N_12087);
nor U12296 (N_12296,N_12137,N_12071);
nor U12297 (N_12297,N_12142,N_12131);
nand U12298 (N_12298,N_12068,N_12008);
xor U12299 (N_12299,N_12010,N_12174);
nor U12300 (N_12300,N_12157,N_12013);
nor U12301 (N_12301,N_12027,N_12093);
nand U12302 (N_12302,N_12005,N_12105);
nor U12303 (N_12303,N_12085,N_12119);
nor U12304 (N_12304,N_12170,N_12188);
and U12305 (N_12305,N_12076,N_12082);
nand U12306 (N_12306,N_12193,N_12037);
xor U12307 (N_12307,N_12047,N_12048);
nor U12308 (N_12308,N_12103,N_12060);
nor U12309 (N_12309,N_12143,N_12154);
nand U12310 (N_12310,N_12076,N_12155);
nand U12311 (N_12311,N_12115,N_12003);
or U12312 (N_12312,N_12141,N_12178);
nand U12313 (N_12313,N_12154,N_12106);
xor U12314 (N_12314,N_12002,N_12064);
and U12315 (N_12315,N_12100,N_12002);
or U12316 (N_12316,N_12018,N_12083);
nor U12317 (N_12317,N_12115,N_12036);
nand U12318 (N_12318,N_12191,N_12082);
and U12319 (N_12319,N_12198,N_12001);
or U12320 (N_12320,N_12131,N_12083);
or U12321 (N_12321,N_12000,N_12100);
and U12322 (N_12322,N_12054,N_12166);
or U12323 (N_12323,N_12050,N_12150);
or U12324 (N_12324,N_12158,N_12055);
and U12325 (N_12325,N_12199,N_12054);
and U12326 (N_12326,N_12041,N_12086);
nor U12327 (N_12327,N_12029,N_12180);
xnor U12328 (N_12328,N_12144,N_12166);
or U12329 (N_12329,N_12167,N_12136);
nand U12330 (N_12330,N_12180,N_12163);
nand U12331 (N_12331,N_12021,N_12171);
xnor U12332 (N_12332,N_12030,N_12173);
or U12333 (N_12333,N_12075,N_12082);
nand U12334 (N_12334,N_12095,N_12049);
xnor U12335 (N_12335,N_12179,N_12189);
xor U12336 (N_12336,N_12162,N_12076);
or U12337 (N_12337,N_12169,N_12102);
xor U12338 (N_12338,N_12121,N_12137);
nor U12339 (N_12339,N_12104,N_12063);
and U12340 (N_12340,N_12045,N_12126);
nand U12341 (N_12341,N_12067,N_12185);
xor U12342 (N_12342,N_12026,N_12013);
nor U12343 (N_12343,N_12172,N_12094);
nor U12344 (N_12344,N_12113,N_12190);
nand U12345 (N_12345,N_12173,N_12151);
xnor U12346 (N_12346,N_12154,N_12178);
xnor U12347 (N_12347,N_12018,N_12126);
nor U12348 (N_12348,N_12017,N_12049);
nand U12349 (N_12349,N_12076,N_12161);
and U12350 (N_12350,N_12100,N_12198);
or U12351 (N_12351,N_12155,N_12095);
and U12352 (N_12352,N_12148,N_12152);
nand U12353 (N_12353,N_12086,N_12155);
and U12354 (N_12354,N_12196,N_12000);
xor U12355 (N_12355,N_12155,N_12032);
xor U12356 (N_12356,N_12076,N_12037);
nand U12357 (N_12357,N_12117,N_12093);
nand U12358 (N_12358,N_12073,N_12170);
and U12359 (N_12359,N_12074,N_12092);
and U12360 (N_12360,N_12179,N_12158);
nor U12361 (N_12361,N_12015,N_12169);
xnor U12362 (N_12362,N_12163,N_12084);
or U12363 (N_12363,N_12083,N_12191);
or U12364 (N_12364,N_12085,N_12140);
or U12365 (N_12365,N_12147,N_12062);
nor U12366 (N_12366,N_12004,N_12120);
or U12367 (N_12367,N_12024,N_12193);
and U12368 (N_12368,N_12061,N_12137);
nor U12369 (N_12369,N_12166,N_12176);
xor U12370 (N_12370,N_12061,N_12095);
or U12371 (N_12371,N_12114,N_12138);
nor U12372 (N_12372,N_12070,N_12051);
or U12373 (N_12373,N_12085,N_12172);
xnor U12374 (N_12374,N_12063,N_12049);
nand U12375 (N_12375,N_12033,N_12172);
xor U12376 (N_12376,N_12010,N_12179);
nor U12377 (N_12377,N_12016,N_12168);
nor U12378 (N_12378,N_12137,N_12191);
xor U12379 (N_12379,N_12028,N_12012);
nand U12380 (N_12380,N_12179,N_12075);
nor U12381 (N_12381,N_12133,N_12099);
xor U12382 (N_12382,N_12189,N_12155);
or U12383 (N_12383,N_12039,N_12196);
nand U12384 (N_12384,N_12064,N_12041);
or U12385 (N_12385,N_12107,N_12058);
or U12386 (N_12386,N_12126,N_12174);
and U12387 (N_12387,N_12069,N_12071);
and U12388 (N_12388,N_12047,N_12063);
or U12389 (N_12389,N_12069,N_12195);
nor U12390 (N_12390,N_12110,N_12001);
xor U12391 (N_12391,N_12066,N_12009);
xnor U12392 (N_12392,N_12110,N_12006);
and U12393 (N_12393,N_12160,N_12010);
nor U12394 (N_12394,N_12164,N_12141);
or U12395 (N_12395,N_12065,N_12139);
nor U12396 (N_12396,N_12172,N_12004);
nor U12397 (N_12397,N_12086,N_12016);
nor U12398 (N_12398,N_12170,N_12056);
or U12399 (N_12399,N_12087,N_12072);
nand U12400 (N_12400,N_12374,N_12230);
xor U12401 (N_12401,N_12347,N_12293);
nor U12402 (N_12402,N_12394,N_12270);
and U12403 (N_12403,N_12205,N_12327);
and U12404 (N_12404,N_12399,N_12256);
and U12405 (N_12405,N_12322,N_12378);
nor U12406 (N_12406,N_12294,N_12359);
xnor U12407 (N_12407,N_12283,N_12364);
nand U12408 (N_12408,N_12365,N_12231);
and U12409 (N_12409,N_12206,N_12325);
nor U12410 (N_12410,N_12393,N_12309);
and U12411 (N_12411,N_12334,N_12329);
and U12412 (N_12412,N_12244,N_12336);
nand U12413 (N_12413,N_12245,N_12261);
nor U12414 (N_12414,N_12284,N_12201);
nand U12415 (N_12415,N_12333,N_12302);
and U12416 (N_12416,N_12383,N_12389);
nand U12417 (N_12417,N_12298,N_12275);
or U12418 (N_12418,N_12377,N_12211);
xor U12419 (N_12419,N_12235,N_12266);
nor U12420 (N_12420,N_12306,N_12285);
and U12421 (N_12421,N_12220,N_12208);
or U12422 (N_12422,N_12318,N_12386);
or U12423 (N_12423,N_12369,N_12346);
nand U12424 (N_12424,N_12357,N_12355);
or U12425 (N_12425,N_12370,N_12305);
nand U12426 (N_12426,N_12350,N_12239);
nor U12427 (N_12427,N_12320,N_12288);
nand U12428 (N_12428,N_12332,N_12345);
and U12429 (N_12429,N_12277,N_12321);
or U12430 (N_12430,N_12311,N_12247);
nand U12431 (N_12431,N_12328,N_12280);
nand U12432 (N_12432,N_12248,N_12356);
or U12433 (N_12433,N_12213,N_12398);
or U12434 (N_12434,N_12272,N_12297);
nor U12435 (N_12435,N_12287,N_12217);
xnor U12436 (N_12436,N_12202,N_12268);
and U12437 (N_12437,N_12281,N_12250);
or U12438 (N_12438,N_12351,N_12241);
nand U12439 (N_12439,N_12278,N_12229);
nor U12440 (N_12440,N_12253,N_12246);
and U12441 (N_12441,N_12242,N_12344);
or U12442 (N_12442,N_12326,N_12228);
or U12443 (N_12443,N_12237,N_12214);
nand U12444 (N_12444,N_12341,N_12338);
nor U12445 (N_12445,N_12381,N_12296);
nand U12446 (N_12446,N_12225,N_12372);
nand U12447 (N_12447,N_12363,N_12279);
and U12448 (N_12448,N_12215,N_12240);
xnor U12449 (N_12449,N_12371,N_12373);
and U12450 (N_12450,N_12223,N_12203);
nor U12451 (N_12451,N_12312,N_12366);
or U12452 (N_12452,N_12360,N_12331);
nor U12453 (N_12453,N_12282,N_12330);
nor U12454 (N_12454,N_12361,N_12388);
or U12455 (N_12455,N_12339,N_12258);
xor U12456 (N_12456,N_12216,N_12204);
and U12457 (N_12457,N_12210,N_12348);
or U12458 (N_12458,N_12264,N_12238);
nor U12459 (N_12459,N_12286,N_12385);
nor U12460 (N_12460,N_12335,N_12362);
nand U12461 (N_12461,N_12352,N_12295);
nor U12462 (N_12462,N_12317,N_12269);
nand U12463 (N_12463,N_12340,N_12207);
xnor U12464 (N_12464,N_12218,N_12380);
and U12465 (N_12465,N_12232,N_12234);
nand U12466 (N_12466,N_12392,N_12379);
and U12467 (N_12467,N_12274,N_12376);
nor U12468 (N_12468,N_12243,N_12252);
nand U12469 (N_12469,N_12349,N_12358);
nor U12470 (N_12470,N_12368,N_12276);
and U12471 (N_12471,N_12273,N_12224);
and U12472 (N_12472,N_12375,N_12308);
nor U12473 (N_12473,N_12384,N_12263);
nand U12474 (N_12474,N_12292,N_12315);
or U12475 (N_12475,N_12249,N_12313);
and U12476 (N_12476,N_12353,N_12291);
nand U12477 (N_12477,N_12271,N_12260);
or U12478 (N_12478,N_12342,N_12227);
and U12479 (N_12479,N_12254,N_12212);
nand U12480 (N_12480,N_12299,N_12391);
nor U12481 (N_12481,N_12221,N_12301);
nor U12482 (N_12482,N_12395,N_12303);
or U12483 (N_12483,N_12262,N_12337);
and U12484 (N_12484,N_12259,N_12265);
or U12485 (N_12485,N_12367,N_12387);
or U12486 (N_12486,N_12343,N_12397);
xnor U12487 (N_12487,N_12354,N_12255);
nand U12488 (N_12488,N_12324,N_12290);
xnor U12489 (N_12489,N_12236,N_12304);
or U12490 (N_12490,N_12323,N_12257);
nor U12491 (N_12491,N_12251,N_12390);
or U12492 (N_12492,N_12300,N_12219);
or U12493 (N_12493,N_12319,N_12310);
or U12494 (N_12494,N_12209,N_12314);
nor U12495 (N_12495,N_12267,N_12200);
xnor U12496 (N_12496,N_12222,N_12316);
xor U12497 (N_12497,N_12307,N_12226);
and U12498 (N_12498,N_12382,N_12233);
or U12499 (N_12499,N_12289,N_12396);
and U12500 (N_12500,N_12344,N_12226);
and U12501 (N_12501,N_12369,N_12238);
and U12502 (N_12502,N_12247,N_12333);
nor U12503 (N_12503,N_12261,N_12259);
and U12504 (N_12504,N_12316,N_12377);
or U12505 (N_12505,N_12354,N_12391);
nor U12506 (N_12506,N_12205,N_12330);
and U12507 (N_12507,N_12335,N_12333);
nor U12508 (N_12508,N_12387,N_12306);
and U12509 (N_12509,N_12267,N_12270);
or U12510 (N_12510,N_12243,N_12310);
xor U12511 (N_12511,N_12249,N_12206);
and U12512 (N_12512,N_12224,N_12341);
nand U12513 (N_12513,N_12387,N_12348);
or U12514 (N_12514,N_12263,N_12365);
or U12515 (N_12515,N_12313,N_12360);
nand U12516 (N_12516,N_12338,N_12384);
xor U12517 (N_12517,N_12350,N_12347);
or U12518 (N_12518,N_12211,N_12365);
xnor U12519 (N_12519,N_12289,N_12374);
xnor U12520 (N_12520,N_12378,N_12201);
xor U12521 (N_12521,N_12263,N_12251);
nor U12522 (N_12522,N_12254,N_12240);
nor U12523 (N_12523,N_12295,N_12372);
and U12524 (N_12524,N_12338,N_12364);
nor U12525 (N_12525,N_12309,N_12211);
or U12526 (N_12526,N_12219,N_12228);
xor U12527 (N_12527,N_12363,N_12367);
nor U12528 (N_12528,N_12233,N_12285);
xnor U12529 (N_12529,N_12359,N_12210);
and U12530 (N_12530,N_12390,N_12304);
xnor U12531 (N_12531,N_12384,N_12283);
nor U12532 (N_12532,N_12331,N_12308);
nand U12533 (N_12533,N_12243,N_12362);
or U12534 (N_12534,N_12328,N_12245);
xnor U12535 (N_12535,N_12313,N_12244);
nand U12536 (N_12536,N_12397,N_12260);
or U12537 (N_12537,N_12363,N_12264);
xnor U12538 (N_12538,N_12267,N_12266);
and U12539 (N_12539,N_12276,N_12299);
and U12540 (N_12540,N_12273,N_12362);
nor U12541 (N_12541,N_12316,N_12337);
or U12542 (N_12542,N_12267,N_12215);
xnor U12543 (N_12543,N_12247,N_12358);
or U12544 (N_12544,N_12331,N_12219);
xnor U12545 (N_12545,N_12302,N_12327);
xnor U12546 (N_12546,N_12216,N_12393);
nor U12547 (N_12547,N_12382,N_12279);
nand U12548 (N_12548,N_12218,N_12214);
nand U12549 (N_12549,N_12304,N_12391);
nor U12550 (N_12550,N_12398,N_12263);
nand U12551 (N_12551,N_12391,N_12360);
nor U12552 (N_12552,N_12217,N_12253);
nand U12553 (N_12553,N_12283,N_12337);
nor U12554 (N_12554,N_12208,N_12235);
nor U12555 (N_12555,N_12219,N_12294);
nor U12556 (N_12556,N_12361,N_12375);
nand U12557 (N_12557,N_12302,N_12305);
or U12558 (N_12558,N_12300,N_12306);
and U12559 (N_12559,N_12220,N_12236);
and U12560 (N_12560,N_12276,N_12280);
nor U12561 (N_12561,N_12365,N_12266);
or U12562 (N_12562,N_12239,N_12319);
or U12563 (N_12563,N_12369,N_12298);
nand U12564 (N_12564,N_12282,N_12304);
or U12565 (N_12565,N_12390,N_12252);
and U12566 (N_12566,N_12212,N_12228);
xnor U12567 (N_12567,N_12318,N_12230);
nor U12568 (N_12568,N_12375,N_12228);
nor U12569 (N_12569,N_12397,N_12210);
nand U12570 (N_12570,N_12218,N_12390);
xnor U12571 (N_12571,N_12381,N_12232);
or U12572 (N_12572,N_12238,N_12210);
xor U12573 (N_12573,N_12262,N_12369);
nor U12574 (N_12574,N_12368,N_12244);
or U12575 (N_12575,N_12380,N_12207);
or U12576 (N_12576,N_12329,N_12296);
and U12577 (N_12577,N_12256,N_12236);
or U12578 (N_12578,N_12286,N_12352);
nand U12579 (N_12579,N_12323,N_12271);
and U12580 (N_12580,N_12278,N_12363);
xor U12581 (N_12581,N_12204,N_12276);
and U12582 (N_12582,N_12205,N_12298);
xnor U12583 (N_12583,N_12367,N_12300);
nor U12584 (N_12584,N_12216,N_12314);
or U12585 (N_12585,N_12310,N_12395);
xnor U12586 (N_12586,N_12236,N_12281);
nor U12587 (N_12587,N_12233,N_12328);
and U12588 (N_12588,N_12359,N_12295);
nor U12589 (N_12589,N_12382,N_12362);
nor U12590 (N_12590,N_12235,N_12399);
xor U12591 (N_12591,N_12336,N_12327);
or U12592 (N_12592,N_12348,N_12211);
nand U12593 (N_12593,N_12344,N_12394);
nor U12594 (N_12594,N_12299,N_12281);
or U12595 (N_12595,N_12349,N_12235);
nor U12596 (N_12596,N_12316,N_12256);
and U12597 (N_12597,N_12276,N_12374);
nand U12598 (N_12598,N_12240,N_12323);
xnor U12599 (N_12599,N_12309,N_12299);
xnor U12600 (N_12600,N_12472,N_12504);
and U12601 (N_12601,N_12452,N_12581);
nand U12602 (N_12602,N_12422,N_12443);
and U12603 (N_12603,N_12575,N_12435);
xnor U12604 (N_12604,N_12417,N_12448);
nor U12605 (N_12605,N_12523,N_12552);
and U12606 (N_12606,N_12468,N_12496);
or U12607 (N_12607,N_12545,N_12474);
or U12608 (N_12608,N_12550,N_12480);
or U12609 (N_12609,N_12503,N_12521);
nor U12610 (N_12610,N_12506,N_12459);
or U12611 (N_12611,N_12533,N_12495);
xnor U12612 (N_12612,N_12419,N_12527);
and U12613 (N_12613,N_12481,N_12439);
nand U12614 (N_12614,N_12593,N_12408);
nor U12615 (N_12615,N_12436,N_12410);
nor U12616 (N_12616,N_12470,N_12402);
nand U12617 (N_12617,N_12591,N_12528);
and U12618 (N_12618,N_12401,N_12429);
xor U12619 (N_12619,N_12413,N_12457);
or U12620 (N_12620,N_12421,N_12493);
and U12621 (N_12621,N_12458,N_12515);
nor U12622 (N_12622,N_12573,N_12534);
and U12623 (N_12623,N_12592,N_12513);
or U12624 (N_12624,N_12540,N_12478);
nand U12625 (N_12625,N_12547,N_12529);
or U12626 (N_12626,N_12490,N_12416);
nor U12627 (N_12627,N_12568,N_12596);
xnor U12628 (N_12628,N_12412,N_12444);
or U12629 (N_12629,N_12432,N_12510);
or U12630 (N_12630,N_12505,N_12426);
nor U12631 (N_12631,N_12438,N_12524);
nand U12632 (N_12632,N_12464,N_12462);
nor U12633 (N_12633,N_12576,N_12442);
and U12634 (N_12634,N_12569,N_12473);
and U12635 (N_12635,N_12548,N_12491);
and U12636 (N_12636,N_12562,N_12456);
and U12637 (N_12637,N_12570,N_12558);
xnor U12638 (N_12638,N_12530,N_12508);
nor U12639 (N_12639,N_12501,N_12498);
nand U12640 (N_12640,N_12433,N_12580);
xnor U12641 (N_12641,N_12541,N_12567);
or U12642 (N_12642,N_12411,N_12579);
and U12643 (N_12643,N_12526,N_12409);
and U12644 (N_12644,N_12400,N_12586);
xor U12645 (N_12645,N_12598,N_12477);
or U12646 (N_12646,N_12549,N_12475);
nor U12647 (N_12647,N_12538,N_12406);
and U12648 (N_12648,N_12465,N_12451);
xnor U12649 (N_12649,N_12423,N_12499);
or U12650 (N_12650,N_12425,N_12407);
and U12651 (N_12651,N_12471,N_12561);
nor U12652 (N_12652,N_12560,N_12430);
nor U12653 (N_12653,N_12588,N_12445);
nor U12654 (N_12654,N_12553,N_12518);
or U12655 (N_12655,N_12492,N_12418);
and U12656 (N_12656,N_12420,N_12449);
or U12657 (N_12657,N_12557,N_12546);
xor U12658 (N_12658,N_12502,N_12454);
or U12659 (N_12659,N_12469,N_12428);
nor U12660 (N_12660,N_12486,N_12440);
or U12661 (N_12661,N_12494,N_12565);
nand U12662 (N_12662,N_12554,N_12590);
or U12663 (N_12663,N_12595,N_12564);
and U12664 (N_12664,N_12453,N_12587);
nor U12665 (N_12665,N_12461,N_12582);
and U12666 (N_12666,N_12597,N_12447);
nand U12667 (N_12667,N_12522,N_12427);
xor U12668 (N_12668,N_12446,N_12460);
and U12669 (N_12669,N_12497,N_12466);
nor U12670 (N_12670,N_12536,N_12509);
nor U12671 (N_12671,N_12559,N_12441);
nor U12672 (N_12672,N_12537,N_12563);
xnor U12673 (N_12673,N_12424,N_12437);
and U12674 (N_12674,N_12405,N_12532);
or U12675 (N_12675,N_12566,N_12450);
and U12676 (N_12676,N_12543,N_12484);
xor U12677 (N_12677,N_12488,N_12479);
nor U12678 (N_12678,N_12467,N_12489);
and U12679 (N_12679,N_12583,N_12507);
or U12680 (N_12680,N_12525,N_12415);
or U12681 (N_12681,N_12574,N_12577);
and U12682 (N_12682,N_12404,N_12542);
nand U12683 (N_12683,N_12511,N_12585);
nor U12684 (N_12684,N_12517,N_12463);
and U12685 (N_12685,N_12500,N_12539);
and U12686 (N_12686,N_12544,N_12584);
nor U12687 (N_12687,N_12535,N_12594);
or U12688 (N_12688,N_12482,N_12556);
nor U12689 (N_12689,N_12431,N_12531);
nand U12690 (N_12690,N_12551,N_12571);
or U12691 (N_12691,N_12589,N_12520);
xor U12692 (N_12692,N_12434,N_12414);
and U12693 (N_12693,N_12483,N_12403);
xnor U12694 (N_12694,N_12514,N_12516);
or U12695 (N_12695,N_12519,N_12555);
or U12696 (N_12696,N_12485,N_12476);
xnor U12697 (N_12697,N_12578,N_12487);
or U12698 (N_12698,N_12599,N_12455);
and U12699 (N_12699,N_12572,N_12512);
nor U12700 (N_12700,N_12513,N_12515);
or U12701 (N_12701,N_12570,N_12547);
or U12702 (N_12702,N_12547,N_12528);
and U12703 (N_12703,N_12474,N_12508);
or U12704 (N_12704,N_12468,N_12560);
or U12705 (N_12705,N_12517,N_12486);
nor U12706 (N_12706,N_12566,N_12432);
and U12707 (N_12707,N_12531,N_12403);
xor U12708 (N_12708,N_12565,N_12422);
nand U12709 (N_12709,N_12561,N_12551);
nor U12710 (N_12710,N_12447,N_12515);
xnor U12711 (N_12711,N_12448,N_12492);
xor U12712 (N_12712,N_12402,N_12531);
and U12713 (N_12713,N_12458,N_12566);
and U12714 (N_12714,N_12475,N_12497);
nor U12715 (N_12715,N_12585,N_12506);
or U12716 (N_12716,N_12540,N_12569);
and U12717 (N_12717,N_12512,N_12534);
xnor U12718 (N_12718,N_12561,N_12447);
and U12719 (N_12719,N_12495,N_12586);
or U12720 (N_12720,N_12529,N_12599);
xor U12721 (N_12721,N_12408,N_12505);
nor U12722 (N_12722,N_12437,N_12412);
nand U12723 (N_12723,N_12590,N_12465);
nor U12724 (N_12724,N_12426,N_12475);
or U12725 (N_12725,N_12584,N_12598);
or U12726 (N_12726,N_12403,N_12481);
or U12727 (N_12727,N_12453,N_12438);
nand U12728 (N_12728,N_12516,N_12511);
and U12729 (N_12729,N_12555,N_12457);
xnor U12730 (N_12730,N_12404,N_12592);
or U12731 (N_12731,N_12440,N_12589);
or U12732 (N_12732,N_12405,N_12408);
nand U12733 (N_12733,N_12596,N_12557);
xnor U12734 (N_12734,N_12587,N_12521);
and U12735 (N_12735,N_12510,N_12502);
xor U12736 (N_12736,N_12593,N_12482);
or U12737 (N_12737,N_12588,N_12570);
nand U12738 (N_12738,N_12412,N_12525);
and U12739 (N_12739,N_12445,N_12427);
xor U12740 (N_12740,N_12535,N_12407);
nor U12741 (N_12741,N_12437,N_12525);
nand U12742 (N_12742,N_12585,N_12513);
or U12743 (N_12743,N_12549,N_12521);
nor U12744 (N_12744,N_12579,N_12526);
and U12745 (N_12745,N_12454,N_12442);
xor U12746 (N_12746,N_12495,N_12599);
and U12747 (N_12747,N_12508,N_12427);
xor U12748 (N_12748,N_12417,N_12577);
nand U12749 (N_12749,N_12569,N_12465);
nand U12750 (N_12750,N_12461,N_12426);
xor U12751 (N_12751,N_12447,N_12523);
nand U12752 (N_12752,N_12579,N_12578);
xnor U12753 (N_12753,N_12535,N_12452);
xnor U12754 (N_12754,N_12429,N_12428);
nand U12755 (N_12755,N_12585,N_12503);
nor U12756 (N_12756,N_12525,N_12523);
and U12757 (N_12757,N_12527,N_12480);
nand U12758 (N_12758,N_12528,N_12531);
xnor U12759 (N_12759,N_12590,N_12441);
nor U12760 (N_12760,N_12506,N_12407);
nand U12761 (N_12761,N_12465,N_12454);
nor U12762 (N_12762,N_12478,N_12547);
and U12763 (N_12763,N_12472,N_12405);
nor U12764 (N_12764,N_12450,N_12520);
and U12765 (N_12765,N_12433,N_12567);
or U12766 (N_12766,N_12596,N_12591);
nor U12767 (N_12767,N_12413,N_12441);
nor U12768 (N_12768,N_12555,N_12549);
nand U12769 (N_12769,N_12402,N_12599);
xnor U12770 (N_12770,N_12551,N_12568);
and U12771 (N_12771,N_12438,N_12510);
or U12772 (N_12772,N_12591,N_12512);
and U12773 (N_12773,N_12477,N_12420);
and U12774 (N_12774,N_12405,N_12516);
xor U12775 (N_12775,N_12439,N_12467);
nor U12776 (N_12776,N_12514,N_12582);
and U12777 (N_12777,N_12525,N_12521);
nand U12778 (N_12778,N_12437,N_12470);
nand U12779 (N_12779,N_12411,N_12597);
nor U12780 (N_12780,N_12499,N_12506);
nand U12781 (N_12781,N_12590,N_12503);
nor U12782 (N_12782,N_12593,N_12427);
nand U12783 (N_12783,N_12569,N_12533);
nor U12784 (N_12784,N_12531,N_12440);
nor U12785 (N_12785,N_12539,N_12515);
nor U12786 (N_12786,N_12482,N_12473);
xor U12787 (N_12787,N_12450,N_12581);
xnor U12788 (N_12788,N_12572,N_12545);
and U12789 (N_12789,N_12457,N_12426);
xnor U12790 (N_12790,N_12583,N_12587);
and U12791 (N_12791,N_12482,N_12528);
nor U12792 (N_12792,N_12552,N_12463);
and U12793 (N_12793,N_12407,N_12536);
nor U12794 (N_12794,N_12462,N_12495);
xor U12795 (N_12795,N_12524,N_12457);
and U12796 (N_12796,N_12583,N_12485);
or U12797 (N_12797,N_12535,N_12577);
or U12798 (N_12798,N_12478,N_12433);
or U12799 (N_12799,N_12473,N_12472);
nor U12800 (N_12800,N_12617,N_12713);
xnor U12801 (N_12801,N_12664,N_12601);
xor U12802 (N_12802,N_12734,N_12740);
xnor U12803 (N_12803,N_12790,N_12789);
nand U12804 (N_12804,N_12652,N_12649);
xnor U12805 (N_12805,N_12756,N_12741);
and U12806 (N_12806,N_12607,N_12742);
and U12807 (N_12807,N_12752,N_12715);
nor U12808 (N_12808,N_12766,N_12714);
and U12809 (N_12809,N_12787,N_12773);
xnor U12810 (N_12810,N_12744,N_12748);
nand U12811 (N_12811,N_12696,N_12783);
xnor U12812 (N_12812,N_12768,N_12663);
nor U12813 (N_12813,N_12602,N_12637);
nor U12814 (N_12814,N_12717,N_12699);
nor U12815 (N_12815,N_12743,N_12606);
or U12816 (N_12816,N_12733,N_12710);
nand U12817 (N_12817,N_12634,N_12684);
nor U12818 (N_12818,N_12661,N_12700);
xor U12819 (N_12819,N_12686,N_12749);
nand U12820 (N_12820,N_12764,N_12648);
nand U12821 (N_12821,N_12640,N_12757);
nand U12822 (N_12822,N_12687,N_12711);
or U12823 (N_12823,N_12679,N_12737);
nor U12824 (N_12824,N_12646,N_12695);
or U12825 (N_12825,N_12799,N_12656);
nand U12826 (N_12826,N_12777,N_12784);
and U12827 (N_12827,N_12765,N_12726);
nor U12828 (N_12828,N_12635,N_12724);
or U12829 (N_12829,N_12680,N_12792);
nor U12830 (N_12830,N_12643,N_12767);
nor U12831 (N_12831,N_12780,N_12628);
nand U12832 (N_12832,N_12745,N_12716);
nor U12833 (N_12833,N_12609,N_12677);
nand U12834 (N_12834,N_12697,N_12639);
nand U12835 (N_12835,N_12755,N_12683);
nor U12836 (N_12836,N_12675,N_12753);
nand U12837 (N_12837,N_12691,N_12709);
and U12838 (N_12838,N_12624,N_12786);
and U12839 (N_12839,N_12702,N_12622);
or U12840 (N_12840,N_12754,N_12795);
xnor U12841 (N_12841,N_12681,N_12625);
nor U12842 (N_12842,N_12738,N_12612);
or U12843 (N_12843,N_12781,N_12688);
or U12844 (N_12844,N_12721,N_12621);
or U12845 (N_12845,N_12651,N_12707);
xnor U12846 (N_12846,N_12660,N_12673);
xnor U12847 (N_12847,N_12794,N_12618);
and U12848 (N_12848,N_12650,N_12730);
xnor U12849 (N_12849,N_12670,N_12759);
and U12850 (N_12850,N_12775,N_12620);
nor U12851 (N_12851,N_12778,N_12729);
xnor U12852 (N_12852,N_12623,N_12782);
xor U12853 (N_12853,N_12615,N_12662);
xnor U12854 (N_12854,N_12626,N_12632);
xor U12855 (N_12855,N_12659,N_12665);
xnor U12856 (N_12856,N_12608,N_12629);
or U12857 (N_12857,N_12692,N_12614);
nor U12858 (N_12858,N_12703,N_12678);
nand U12859 (N_12859,N_12772,N_12701);
xnor U12860 (N_12860,N_12739,N_12676);
xnor U12861 (N_12861,N_12732,N_12666);
or U12862 (N_12862,N_12785,N_12758);
or U12863 (N_12863,N_12712,N_12630);
and U12864 (N_12864,N_12723,N_12727);
nand U12865 (N_12865,N_12672,N_12698);
nor U12866 (N_12866,N_12644,N_12728);
or U12867 (N_12867,N_12796,N_12667);
xnor U12868 (N_12868,N_12627,N_12731);
or U12869 (N_12869,N_12771,N_12605);
nand U12870 (N_12870,N_12638,N_12763);
xor U12871 (N_12871,N_12671,N_12633);
xor U12872 (N_12872,N_12776,N_12631);
nor U12873 (N_12873,N_12722,N_12706);
nor U12874 (N_12874,N_12600,N_12705);
xnor U12875 (N_12875,N_12658,N_12655);
or U12876 (N_12876,N_12769,N_12797);
or U12877 (N_12877,N_12760,N_12657);
and U12878 (N_12878,N_12791,N_12690);
nor U12879 (N_12879,N_12653,N_12693);
or U12880 (N_12880,N_12770,N_12761);
nand U12881 (N_12881,N_12708,N_12603);
or U12882 (N_12882,N_12694,N_12685);
nor U12883 (N_12883,N_12718,N_12798);
nand U12884 (N_12884,N_12645,N_12611);
and U12885 (N_12885,N_12735,N_12750);
and U12886 (N_12886,N_12689,N_12793);
nor U12887 (N_12887,N_12610,N_12779);
nor U12888 (N_12888,N_12788,N_12746);
or U12889 (N_12889,N_12751,N_12762);
nor U12890 (N_12890,N_12642,N_12674);
nor U12891 (N_12891,N_12647,N_12704);
or U12892 (N_12892,N_12641,N_12774);
or U12893 (N_12893,N_12636,N_12719);
and U12894 (N_12894,N_12616,N_12654);
nor U12895 (N_12895,N_12736,N_12725);
or U12896 (N_12896,N_12682,N_12619);
and U12897 (N_12897,N_12668,N_12747);
xor U12898 (N_12898,N_12613,N_12669);
or U12899 (N_12899,N_12604,N_12720);
and U12900 (N_12900,N_12656,N_12717);
or U12901 (N_12901,N_12625,N_12747);
or U12902 (N_12902,N_12712,N_12768);
and U12903 (N_12903,N_12619,N_12613);
xor U12904 (N_12904,N_12710,N_12626);
nor U12905 (N_12905,N_12603,N_12674);
and U12906 (N_12906,N_12667,N_12750);
and U12907 (N_12907,N_12785,N_12653);
or U12908 (N_12908,N_12723,N_12755);
nor U12909 (N_12909,N_12798,N_12675);
or U12910 (N_12910,N_12673,N_12696);
and U12911 (N_12911,N_12668,N_12768);
nor U12912 (N_12912,N_12766,N_12747);
or U12913 (N_12913,N_12708,N_12761);
nand U12914 (N_12914,N_12707,N_12793);
xor U12915 (N_12915,N_12684,N_12796);
nand U12916 (N_12916,N_12773,N_12713);
nor U12917 (N_12917,N_12622,N_12761);
and U12918 (N_12918,N_12777,N_12790);
xnor U12919 (N_12919,N_12774,N_12743);
nor U12920 (N_12920,N_12615,N_12718);
and U12921 (N_12921,N_12731,N_12698);
or U12922 (N_12922,N_12753,N_12694);
and U12923 (N_12923,N_12609,N_12737);
and U12924 (N_12924,N_12780,N_12626);
xnor U12925 (N_12925,N_12669,N_12605);
nor U12926 (N_12926,N_12603,N_12727);
and U12927 (N_12927,N_12767,N_12610);
or U12928 (N_12928,N_12629,N_12743);
or U12929 (N_12929,N_12731,N_12795);
xnor U12930 (N_12930,N_12665,N_12658);
and U12931 (N_12931,N_12695,N_12748);
nand U12932 (N_12932,N_12798,N_12606);
and U12933 (N_12933,N_12782,N_12787);
and U12934 (N_12934,N_12720,N_12759);
and U12935 (N_12935,N_12645,N_12732);
or U12936 (N_12936,N_12760,N_12683);
nand U12937 (N_12937,N_12785,N_12692);
xnor U12938 (N_12938,N_12682,N_12705);
nor U12939 (N_12939,N_12622,N_12668);
and U12940 (N_12940,N_12627,N_12701);
xor U12941 (N_12941,N_12776,N_12789);
nor U12942 (N_12942,N_12621,N_12663);
and U12943 (N_12943,N_12737,N_12666);
and U12944 (N_12944,N_12646,N_12742);
and U12945 (N_12945,N_12617,N_12695);
nor U12946 (N_12946,N_12659,N_12673);
and U12947 (N_12947,N_12626,N_12697);
nand U12948 (N_12948,N_12664,N_12781);
xor U12949 (N_12949,N_12757,N_12615);
nor U12950 (N_12950,N_12695,N_12762);
nor U12951 (N_12951,N_12746,N_12677);
nor U12952 (N_12952,N_12641,N_12737);
nand U12953 (N_12953,N_12677,N_12637);
and U12954 (N_12954,N_12663,N_12697);
nor U12955 (N_12955,N_12656,N_12680);
and U12956 (N_12956,N_12699,N_12782);
xnor U12957 (N_12957,N_12783,N_12731);
or U12958 (N_12958,N_12790,N_12780);
xor U12959 (N_12959,N_12611,N_12738);
xor U12960 (N_12960,N_12619,N_12661);
and U12961 (N_12961,N_12756,N_12727);
and U12962 (N_12962,N_12776,N_12768);
or U12963 (N_12963,N_12628,N_12633);
nor U12964 (N_12964,N_12652,N_12701);
nand U12965 (N_12965,N_12791,N_12686);
and U12966 (N_12966,N_12677,N_12671);
and U12967 (N_12967,N_12779,N_12762);
or U12968 (N_12968,N_12628,N_12674);
nor U12969 (N_12969,N_12623,N_12624);
or U12970 (N_12970,N_12732,N_12639);
or U12971 (N_12971,N_12789,N_12649);
and U12972 (N_12972,N_12747,N_12786);
or U12973 (N_12973,N_12699,N_12713);
nor U12974 (N_12974,N_12614,N_12659);
or U12975 (N_12975,N_12680,N_12643);
nand U12976 (N_12976,N_12648,N_12622);
nor U12977 (N_12977,N_12656,N_12719);
nand U12978 (N_12978,N_12642,N_12761);
nor U12979 (N_12979,N_12657,N_12626);
nor U12980 (N_12980,N_12645,N_12722);
and U12981 (N_12981,N_12664,N_12712);
nor U12982 (N_12982,N_12794,N_12713);
and U12983 (N_12983,N_12642,N_12746);
xnor U12984 (N_12984,N_12671,N_12724);
and U12985 (N_12985,N_12734,N_12795);
nor U12986 (N_12986,N_12755,N_12634);
nor U12987 (N_12987,N_12644,N_12720);
nand U12988 (N_12988,N_12655,N_12679);
nor U12989 (N_12989,N_12695,N_12722);
xnor U12990 (N_12990,N_12661,N_12626);
or U12991 (N_12991,N_12618,N_12691);
or U12992 (N_12992,N_12753,N_12775);
or U12993 (N_12993,N_12685,N_12761);
or U12994 (N_12994,N_12629,N_12658);
xnor U12995 (N_12995,N_12715,N_12619);
or U12996 (N_12996,N_12688,N_12619);
and U12997 (N_12997,N_12634,N_12632);
and U12998 (N_12998,N_12732,N_12753);
or U12999 (N_12999,N_12724,N_12739);
nand U13000 (N_13000,N_12946,N_12800);
or U13001 (N_13001,N_12807,N_12868);
and U13002 (N_13002,N_12937,N_12955);
or U13003 (N_13003,N_12926,N_12836);
or U13004 (N_13004,N_12921,N_12907);
or U13005 (N_13005,N_12848,N_12932);
and U13006 (N_13006,N_12948,N_12902);
xor U13007 (N_13007,N_12985,N_12867);
xnor U13008 (N_13008,N_12850,N_12942);
nor U13009 (N_13009,N_12855,N_12898);
nand U13010 (N_13010,N_12826,N_12925);
xor U13011 (N_13011,N_12882,N_12810);
nand U13012 (N_13012,N_12831,N_12938);
or U13013 (N_13013,N_12920,N_12928);
xnor U13014 (N_13014,N_12896,N_12816);
and U13015 (N_13015,N_12947,N_12889);
or U13016 (N_13016,N_12841,N_12853);
or U13017 (N_13017,N_12990,N_12832);
or U13018 (N_13018,N_12805,N_12852);
xnor U13019 (N_13019,N_12954,N_12843);
or U13020 (N_13020,N_12977,N_12981);
nand U13021 (N_13021,N_12872,N_12865);
xnor U13022 (N_13022,N_12908,N_12941);
nand U13023 (N_13023,N_12887,N_12900);
and U13024 (N_13024,N_12924,N_12812);
and U13025 (N_13025,N_12824,N_12993);
and U13026 (N_13026,N_12809,N_12875);
and U13027 (N_13027,N_12840,N_12984);
or U13028 (N_13028,N_12933,N_12846);
or U13029 (N_13029,N_12811,N_12974);
and U13030 (N_13030,N_12881,N_12817);
or U13031 (N_13031,N_12992,N_12964);
or U13032 (N_13032,N_12821,N_12895);
nand U13033 (N_13033,N_12897,N_12891);
nand U13034 (N_13034,N_12986,N_12962);
and U13035 (N_13035,N_12972,N_12913);
xor U13036 (N_13036,N_12859,N_12927);
and U13037 (N_13037,N_12862,N_12929);
and U13038 (N_13038,N_12940,N_12967);
nand U13039 (N_13039,N_12910,N_12911);
xor U13040 (N_13040,N_12995,N_12828);
nand U13041 (N_13041,N_12866,N_12915);
and U13042 (N_13042,N_12830,N_12982);
or U13043 (N_13043,N_12936,N_12975);
xor U13044 (N_13044,N_12970,N_12863);
and U13045 (N_13045,N_12973,N_12833);
xnor U13046 (N_13046,N_12971,N_12991);
and U13047 (N_13047,N_12871,N_12901);
and U13048 (N_13048,N_12903,N_12904);
xnor U13049 (N_13049,N_12861,N_12879);
xnor U13050 (N_13050,N_12820,N_12958);
nor U13051 (N_13051,N_12998,N_12969);
nor U13052 (N_13052,N_12997,N_12884);
nor U13053 (N_13053,N_12952,N_12883);
and U13054 (N_13054,N_12894,N_12944);
or U13055 (N_13055,N_12804,N_12876);
nand U13056 (N_13056,N_12999,N_12918);
or U13057 (N_13057,N_12827,N_12945);
xnor U13058 (N_13058,N_12893,N_12834);
nor U13059 (N_13059,N_12983,N_12890);
nor U13060 (N_13060,N_12813,N_12814);
nand U13061 (N_13061,N_12856,N_12950);
or U13062 (N_13062,N_12905,N_12909);
and U13063 (N_13063,N_12842,N_12851);
nand U13064 (N_13064,N_12818,N_12892);
xor U13065 (N_13065,N_12886,N_12829);
and U13066 (N_13066,N_12939,N_12860);
nor U13067 (N_13067,N_12870,N_12877);
or U13068 (N_13068,N_12980,N_12953);
and U13069 (N_13069,N_12930,N_12965);
and U13070 (N_13070,N_12916,N_12873);
and U13071 (N_13071,N_12854,N_12822);
nand U13072 (N_13072,N_12899,N_12923);
xor U13073 (N_13073,N_12988,N_12943);
xnor U13074 (N_13074,N_12906,N_12857);
or U13075 (N_13075,N_12815,N_12847);
xnor U13076 (N_13076,N_12931,N_12858);
xor U13077 (N_13077,N_12935,N_12922);
or U13078 (N_13078,N_12869,N_12888);
or U13079 (N_13079,N_12874,N_12885);
xor U13080 (N_13080,N_12949,N_12803);
nand U13081 (N_13081,N_12837,N_12960);
and U13082 (N_13082,N_12801,N_12808);
nand U13083 (N_13083,N_12994,N_12912);
or U13084 (N_13084,N_12864,N_12963);
or U13085 (N_13085,N_12844,N_12823);
nor U13086 (N_13086,N_12979,N_12917);
nor U13087 (N_13087,N_12839,N_12819);
xor U13088 (N_13088,N_12966,N_12835);
and U13089 (N_13089,N_12806,N_12838);
xnor U13090 (N_13090,N_12959,N_12961);
and U13091 (N_13091,N_12968,N_12919);
nand U13092 (N_13092,N_12934,N_12996);
xnor U13093 (N_13093,N_12802,N_12914);
nand U13094 (N_13094,N_12989,N_12849);
nand U13095 (N_13095,N_12880,N_12987);
xor U13096 (N_13096,N_12825,N_12845);
or U13097 (N_13097,N_12956,N_12978);
or U13098 (N_13098,N_12957,N_12878);
or U13099 (N_13099,N_12976,N_12951);
nor U13100 (N_13100,N_12981,N_12936);
and U13101 (N_13101,N_12903,N_12913);
nor U13102 (N_13102,N_12947,N_12842);
xor U13103 (N_13103,N_12908,N_12895);
or U13104 (N_13104,N_12865,N_12977);
nor U13105 (N_13105,N_12869,N_12885);
and U13106 (N_13106,N_12939,N_12947);
xnor U13107 (N_13107,N_12911,N_12831);
and U13108 (N_13108,N_12974,N_12803);
xor U13109 (N_13109,N_12808,N_12844);
xor U13110 (N_13110,N_12814,N_12906);
xnor U13111 (N_13111,N_12863,N_12817);
and U13112 (N_13112,N_12837,N_12985);
nand U13113 (N_13113,N_12871,N_12843);
xnor U13114 (N_13114,N_12935,N_12999);
nor U13115 (N_13115,N_12973,N_12938);
nor U13116 (N_13116,N_12803,N_12858);
nor U13117 (N_13117,N_12840,N_12985);
xor U13118 (N_13118,N_12890,N_12817);
nand U13119 (N_13119,N_12989,N_12949);
xor U13120 (N_13120,N_12966,N_12915);
xor U13121 (N_13121,N_12918,N_12909);
xnor U13122 (N_13122,N_12902,N_12997);
xor U13123 (N_13123,N_12907,N_12937);
or U13124 (N_13124,N_12866,N_12920);
or U13125 (N_13125,N_12994,N_12997);
and U13126 (N_13126,N_12916,N_12844);
xor U13127 (N_13127,N_12918,N_12963);
and U13128 (N_13128,N_12800,N_12942);
nand U13129 (N_13129,N_12973,N_12871);
or U13130 (N_13130,N_12818,N_12922);
nor U13131 (N_13131,N_12837,N_12955);
or U13132 (N_13132,N_12898,N_12985);
nor U13133 (N_13133,N_12940,N_12871);
nor U13134 (N_13134,N_12920,N_12988);
nand U13135 (N_13135,N_12850,N_12882);
xnor U13136 (N_13136,N_12890,N_12842);
nand U13137 (N_13137,N_12926,N_12979);
and U13138 (N_13138,N_12812,N_12888);
nand U13139 (N_13139,N_12996,N_12920);
nand U13140 (N_13140,N_12998,N_12962);
xnor U13141 (N_13141,N_12823,N_12999);
and U13142 (N_13142,N_12891,N_12944);
nor U13143 (N_13143,N_12940,N_12853);
nand U13144 (N_13144,N_12919,N_12924);
nor U13145 (N_13145,N_12861,N_12803);
nand U13146 (N_13146,N_12941,N_12991);
or U13147 (N_13147,N_12855,N_12905);
or U13148 (N_13148,N_12804,N_12945);
or U13149 (N_13149,N_12947,N_12958);
and U13150 (N_13150,N_12836,N_12831);
nor U13151 (N_13151,N_12822,N_12808);
xnor U13152 (N_13152,N_12999,N_12841);
or U13153 (N_13153,N_12912,N_12976);
and U13154 (N_13154,N_12800,N_12982);
xnor U13155 (N_13155,N_12941,N_12911);
nor U13156 (N_13156,N_12848,N_12857);
and U13157 (N_13157,N_12820,N_12816);
nor U13158 (N_13158,N_12877,N_12889);
xor U13159 (N_13159,N_12924,N_12986);
or U13160 (N_13160,N_12839,N_12986);
xor U13161 (N_13161,N_12992,N_12967);
nand U13162 (N_13162,N_12976,N_12969);
and U13163 (N_13163,N_12880,N_12867);
xnor U13164 (N_13164,N_12849,N_12903);
nand U13165 (N_13165,N_12825,N_12900);
or U13166 (N_13166,N_12826,N_12942);
nand U13167 (N_13167,N_12808,N_12814);
and U13168 (N_13168,N_12803,N_12887);
nor U13169 (N_13169,N_12974,N_12816);
xnor U13170 (N_13170,N_12876,N_12921);
nand U13171 (N_13171,N_12860,N_12899);
and U13172 (N_13172,N_12938,N_12863);
or U13173 (N_13173,N_12998,N_12990);
nand U13174 (N_13174,N_12997,N_12809);
or U13175 (N_13175,N_12935,N_12956);
nor U13176 (N_13176,N_12828,N_12940);
or U13177 (N_13177,N_12818,N_12919);
or U13178 (N_13178,N_12857,N_12899);
and U13179 (N_13179,N_12815,N_12886);
nand U13180 (N_13180,N_12922,N_12813);
or U13181 (N_13181,N_12926,N_12852);
or U13182 (N_13182,N_12903,N_12905);
nand U13183 (N_13183,N_12941,N_12903);
and U13184 (N_13184,N_12964,N_12935);
and U13185 (N_13185,N_12937,N_12936);
nand U13186 (N_13186,N_12887,N_12910);
xor U13187 (N_13187,N_12832,N_12908);
xor U13188 (N_13188,N_12954,N_12933);
and U13189 (N_13189,N_12896,N_12911);
or U13190 (N_13190,N_12990,N_12822);
nor U13191 (N_13191,N_12845,N_12924);
xor U13192 (N_13192,N_12988,N_12808);
nor U13193 (N_13193,N_12958,N_12840);
and U13194 (N_13194,N_12947,N_12937);
and U13195 (N_13195,N_12883,N_12999);
and U13196 (N_13196,N_12810,N_12825);
and U13197 (N_13197,N_12859,N_12919);
or U13198 (N_13198,N_12916,N_12897);
xnor U13199 (N_13199,N_12940,N_12935);
or U13200 (N_13200,N_13191,N_13182);
and U13201 (N_13201,N_13096,N_13118);
xnor U13202 (N_13202,N_13113,N_13060);
nand U13203 (N_13203,N_13126,N_13095);
xor U13204 (N_13204,N_13196,N_13097);
xnor U13205 (N_13205,N_13039,N_13088);
nor U13206 (N_13206,N_13172,N_13124);
and U13207 (N_13207,N_13143,N_13035);
nand U13208 (N_13208,N_13160,N_13112);
nor U13209 (N_13209,N_13068,N_13041);
xor U13210 (N_13210,N_13059,N_13158);
and U13211 (N_13211,N_13043,N_13111);
nand U13212 (N_13212,N_13104,N_13188);
and U13213 (N_13213,N_13163,N_13026);
xor U13214 (N_13214,N_13110,N_13166);
nand U13215 (N_13215,N_13017,N_13168);
or U13216 (N_13216,N_13178,N_13194);
or U13217 (N_13217,N_13077,N_13164);
or U13218 (N_13218,N_13055,N_13010);
xnor U13219 (N_13219,N_13148,N_13065);
and U13220 (N_13220,N_13130,N_13103);
or U13221 (N_13221,N_13031,N_13181);
and U13222 (N_13222,N_13193,N_13081);
nand U13223 (N_13223,N_13140,N_13094);
nand U13224 (N_13224,N_13129,N_13195);
xnor U13225 (N_13225,N_13187,N_13177);
nand U13226 (N_13226,N_13133,N_13090);
nand U13227 (N_13227,N_13016,N_13098);
nor U13228 (N_13228,N_13179,N_13058);
nor U13229 (N_13229,N_13037,N_13052);
and U13230 (N_13230,N_13165,N_13075);
and U13231 (N_13231,N_13125,N_13076);
nand U13232 (N_13232,N_13069,N_13099);
or U13233 (N_13233,N_13120,N_13048);
and U13234 (N_13234,N_13171,N_13061);
nor U13235 (N_13235,N_13064,N_13024);
xnor U13236 (N_13236,N_13092,N_13114);
nor U13237 (N_13237,N_13149,N_13128);
xnor U13238 (N_13238,N_13006,N_13087);
xor U13239 (N_13239,N_13131,N_13074);
xor U13240 (N_13240,N_13009,N_13199);
nand U13241 (N_13241,N_13000,N_13038);
xor U13242 (N_13242,N_13091,N_13070);
nand U13243 (N_13243,N_13062,N_13086);
nor U13244 (N_13244,N_13011,N_13054);
nand U13245 (N_13245,N_13014,N_13145);
or U13246 (N_13246,N_13004,N_13132);
or U13247 (N_13247,N_13170,N_13071);
nor U13248 (N_13248,N_13190,N_13078);
nand U13249 (N_13249,N_13192,N_13073);
or U13250 (N_13250,N_13005,N_13159);
nor U13251 (N_13251,N_13046,N_13079);
nor U13252 (N_13252,N_13066,N_13063);
and U13253 (N_13253,N_13117,N_13044);
and U13254 (N_13254,N_13001,N_13056);
nand U13255 (N_13255,N_13007,N_13169);
or U13256 (N_13256,N_13013,N_13034);
nor U13257 (N_13257,N_13156,N_13072);
nand U13258 (N_13258,N_13085,N_13174);
nor U13259 (N_13259,N_13134,N_13189);
nand U13260 (N_13260,N_13157,N_13021);
xnor U13261 (N_13261,N_13008,N_13101);
xor U13262 (N_13262,N_13082,N_13153);
nor U13263 (N_13263,N_13151,N_13067);
and U13264 (N_13264,N_13049,N_13184);
xor U13265 (N_13265,N_13197,N_13050);
nor U13266 (N_13266,N_13146,N_13135);
or U13267 (N_13267,N_13180,N_13102);
and U13268 (N_13268,N_13127,N_13036);
or U13269 (N_13269,N_13183,N_13047);
or U13270 (N_13270,N_13139,N_13100);
nor U13271 (N_13271,N_13028,N_13122);
and U13272 (N_13272,N_13109,N_13175);
or U13273 (N_13273,N_13053,N_13161);
xnor U13274 (N_13274,N_13015,N_13147);
nand U13275 (N_13275,N_13123,N_13027);
nand U13276 (N_13276,N_13185,N_13012);
nand U13277 (N_13277,N_13167,N_13198);
xor U13278 (N_13278,N_13020,N_13119);
and U13279 (N_13279,N_13057,N_13042);
and U13280 (N_13280,N_13136,N_13138);
or U13281 (N_13281,N_13150,N_13023);
xor U13282 (N_13282,N_13142,N_13040);
xnor U13283 (N_13283,N_13108,N_13105);
and U13284 (N_13284,N_13033,N_13106);
and U13285 (N_13285,N_13144,N_13121);
and U13286 (N_13286,N_13002,N_13003);
and U13287 (N_13287,N_13116,N_13089);
nand U13288 (N_13288,N_13186,N_13162);
xnor U13289 (N_13289,N_13022,N_13154);
nand U13290 (N_13290,N_13083,N_13173);
nand U13291 (N_13291,N_13030,N_13032);
nand U13292 (N_13292,N_13045,N_13155);
nor U13293 (N_13293,N_13084,N_13115);
or U13294 (N_13294,N_13019,N_13176);
xnor U13295 (N_13295,N_13137,N_13029);
xor U13296 (N_13296,N_13152,N_13025);
xor U13297 (N_13297,N_13051,N_13080);
nand U13298 (N_13298,N_13018,N_13141);
nand U13299 (N_13299,N_13107,N_13093);
nand U13300 (N_13300,N_13115,N_13065);
xnor U13301 (N_13301,N_13087,N_13064);
or U13302 (N_13302,N_13077,N_13036);
nor U13303 (N_13303,N_13184,N_13178);
nand U13304 (N_13304,N_13002,N_13153);
nand U13305 (N_13305,N_13076,N_13011);
and U13306 (N_13306,N_13116,N_13074);
or U13307 (N_13307,N_13180,N_13168);
or U13308 (N_13308,N_13013,N_13123);
and U13309 (N_13309,N_13097,N_13061);
xor U13310 (N_13310,N_13039,N_13173);
nor U13311 (N_13311,N_13167,N_13029);
nor U13312 (N_13312,N_13056,N_13160);
nor U13313 (N_13313,N_13088,N_13115);
xor U13314 (N_13314,N_13102,N_13012);
nand U13315 (N_13315,N_13076,N_13072);
xnor U13316 (N_13316,N_13171,N_13063);
and U13317 (N_13317,N_13139,N_13107);
nand U13318 (N_13318,N_13104,N_13028);
and U13319 (N_13319,N_13152,N_13192);
xnor U13320 (N_13320,N_13099,N_13054);
or U13321 (N_13321,N_13162,N_13093);
nand U13322 (N_13322,N_13161,N_13187);
or U13323 (N_13323,N_13091,N_13182);
nor U13324 (N_13324,N_13183,N_13157);
nor U13325 (N_13325,N_13108,N_13070);
xnor U13326 (N_13326,N_13123,N_13088);
nor U13327 (N_13327,N_13132,N_13013);
and U13328 (N_13328,N_13105,N_13168);
xor U13329 (N_13329,N_13012,N_13114);
xnor U13330 (N_13330,N_13043,N_13054);
xnor U13331 (N_13331,N_13148,N_13195);
or U13332 (N_13332,N_13074,N_13154);
nor U13333 (N_13333,N_13004,N_13129);
nor U13334 (N_13334,N_13034,N_13020);
nand U13335 (N_13335,N_13058,N_13039);
and U13336 (N_13336,N_13002,N_13044);
xnor U13337 (N_13337,N_13041,N_13014);
and U13338 (N_13338,N_13117,N_13128);
nand U13339 (N_13339,N_13122,N_13050);
nand U13340 (N_13340,N_13124,N_13113);
nand U13341 (N_13341,N_13178,N_13197);
nor U13342 (N_13342,N_13092,N_13012);
and U13343 (N_13343,N_13001,N_13093);
or U13344 (N_13344,N_13020,N_13197);
xor U13345 (N_13345,N_13084,N_13121);
and U13346 (N_13346,N_13071,N_13197);
nor U13347 (N_13347,N_13129,N_13053);
xor U13348 (N_13348,N_13083,N_13148);
nor U13349 (N_13349,N_13123,N_13002);
nor U13350 (N_13350,N_13093,N_13054);
and U13351 (N_13351,N_13138,N_13189);
xor U13352 (N_13352,N_13130,N_13063);
nand U13353 (N_13353,N_13116,N_13121);
and U13354 (N_13354,N_13060,N_13176);
xnor U13355 (N_13355,N_13007,N_13177);
xor U13356 (N_13356,N_13062,N_13060);
xor U13357 (N_13357,N_13075,N_13122);
nor U13358 (N_13358,N_13034,N_13070);
nor U13359 (N_13359,N_13072,N_13003);
xor U13360 (N_13360,N_13049,N_13004);
xor U13361 (N_13361,N_13062,N_13047);
xor U13362 (N_13362,N_13084,N_13048);
or U13363 (N_13363,N_13112,N_13007);
nand U13364 (N_13364,N_13143,N_13089);
xor U13365 (N_13365,N_13084,N_13017);
or U13366 (N_13366,N_13000,N_13123);
xor U13367 (N_13367,N_13042,N_13077);
xor U13368 (N_13368,N_13029,N_13050);
nor U13369 (N_13369,N_13011,N_13110);
xor U13370 (N_13370,N_13062,N_13146);
nor U13371 (N_13371,N_13132,N_13197);
xnor U13372 (N_13372,N_13186,N_13100);
xnor U13373 (N_13373,N_13130,N_13139);
nor U13374 (N_13374,N_13034,N_13161);
nor U13375 (N_13375,N_13076,N_13043);
or U13376 (N_13376,N_13047,N_13128);
or U13377 (N_13377,N_13101,N_13003);
or U13378 (N_13378,N_13140,N_13144);
and U13379 (N_13379,N_13167,N_13130);
nor U13380 (N_13380,N_13046,N_13191);
and U13381 (N_13381,N_13031,N_13107);
nand U13382 (N_13382,N_13096,N_13114);
or U13383 (N_13383,N_13018,N_13059);
and U13384 (N_13384,N_13086,N_13060);
nor U13385 (N_13385,N_13178,N_13118);
xor U13386 (N_13386,N_13045,N_13089);
nand U13387 (N_13387,N_13122,N_13135);
or U13388 (N_13388,N_13048,N_13199);
nor U13389 (N_13389,N_13093,N_13174);
nor U13390 (N_13390,N_13044,N_13141);
or U13391 (N_13391,N_13096,N_13157);
nand U13392 (N_13392,N_13066,N_13023);
xor U13393 (N_13393,N_13022,N_13099);
nand U13394 (N_13394,N_13043,N_13050);
or U13395 (N_13395,N_13191,N_13014);
and U13396 (N_13396,N_13144,N_13128);
nand U13397 (N_13397,N_13112,N_13170);
or U13398 (N_13398,N_13080,N_13194);
and U13399 (N_13399,N_13136,N_13039);
or U13400 (N_13400,N_13399,N_13246);
nand U13401 (N_13401,N_13288,N_13219);
xor U13402 (N_13402,N_13229,N_13224);
nor U13403 (N_13403,N_13367,N_13317);
or U13404 (N_13404,N_13263,N_13221);
and U13405 (N_13405,N_13375,N_13311);
or U13406 (N_13406,N_13363,N_13328);
nand U13407 (N_13407,N_13379,N_13325);
and U13408 (N_13408,N_13248,N_13322);
nand U13409 (N_13409,N_13210,N_13298);
or U13410 (N_13410,N_13344,N_13257);
and U13411 (N_13411,N_13216,N_13289);
nor U13412 (N_13412,N_13241,N_13254);
nor U13413 (N_13413,N_13300,N_13266);
xnor U13414 (N_13414,N_13277,N_13228);
and U13415 (N_13415,N_13307,N_13268);
nor U13416 (N_13416,N_13334,N_13286);
and U13417 (N_13417,N_13275,N_13321);
or U13418 (N_13418,N_13330,N_13350);
nor U13419 (N_13419,N_13358,N_13270);
nor U13420 (N_13420,N_13214,N_13284);
and U13421 (N_13421,N_13377,N_13208);
or U13422 (N_13422,N_13226,N_13359);
xnor U13423 (N_13423,N_13372,N_13292);
nand U13424 (N_13424,N_13264,N_13369);
and U13425 (N_13425,N_13362,N_13249);
and U13426 (N_13426,N_13297,N_13240);
nor U13427 (N_13427,N_13366,N_13385);
and U13428 (N_13428,N_13343,N_13250);
xnor U13429 (N_13429,N_13395,N_13352);
xor U13430 (N_13430,N_13276,N_13294);
nand U13431 (N_13431,N_13361,N_13389);
or U13432 (N_13432,N_13376,N_13290);
and U13433 (N_13433,N_13243,N_13331);
xnor U13434 (N_13434,N_13244,N_13320);
nor U13435 (N_13435,N_13341,N_13368);
or U13436 (N_13436,N_13365,N_13213);
or U13437 (N_13437,N_13394,N_13205);
and U13438 (N_13438,N_13370,N_13283);
or U13439 (N_13439,N_13239,N_13312);
nor U13440 (N_13440,N_13282,N_13342);
or U13441 (N_13441,N_13347,N_13333);
or U13442 (N_13442,N_13353,N_13381);
and U13443 (N_13443,N_13204,N_13233);
or U13444 (N_13444,N_13260,N_13397);
and U13445 (N_13445,N_13371,N_13235);
or U13446 (N_13446,N_13220,N_13287);
nor U13447 (N_13447,N_13332,N_13346);
xor U13448 (N_13448,N_13339,N_13201);
and U13449 (N_13449,N_13354,N_13258);
and U13450 (N_13450,N_13313,N_13234);
xor U13451 (N_13451,N_13338,N_13384);
and U13452 (N_13452,N_13206,N_13203);
xnor U13453 (N_13453,N_13316,N_13261);
xnor U13454 (N_13454,N_13308,N_13273);
nand U13455 (N_13455,N_13253,N_13351);
nor U13456 (N_13456,N_13323,N_13374);
nor U13457 (N_13457,N_13310,N_13251);
nand U13458 (N_13458,N_13295,N_13274);
xor U13459 (N_13459,N_13390,N_13265);
xnor U13460 (N_13460,N_13373,N_13303);
xor U13461 (N_13461,N_13291,N_13315);
or U13462 (N_13462,N_13252,N_13259);
xor U13463 (N_13463,N_13256,N_13242);
nand U13464 (N_13464,N_13231,N_13225);
xor U13465 (N_13465,N_13336,N_13247);
and U13466 (N_13466,N_13230,N_13306);
and U13467 (N_13467,N_13380,N_13272);
nand U13468 (N_13468,N_13319,N_13262);
nor U13469 (N_13469,N_13398,N_13237);
xnor U13470 (N_13470,N_13255,N_13236);
nor U13471 (N_13471,N_13305,N_13393);
or U13472 (N_13472,N_13357,N_13269);
or U13473 (N_13473,N_13238,N_13337);
xor U13474 (N_13474,N_13378,N_13267);
or U13475 (N_13475,N_13209,N_13293);
xnor U13476 (N_13476,N_13324,N_13392);
or U13477 (N_13477,N_13207,N_13388);
and U13478 (N_13478,N_13329,N_13200);
or U13479 (N_13479,N_13218,N_13285);
and U13480 (N_13480,N_13304,N_13296);
and U13481 (N_13481,N_13211,N_13222);
xnor U13482 (N_13482,N_13245,N_13396);
xnor U13483 (N_13483,N_13279,N_13364);
and U13484 (N_13484,N_13348,N_13386);
nor U13485 (N_13485,N_13227,N_13281);
or U13486 (N_13486,N_13301,N_13340);
nor U13487 (N_13487,N_13314,N_13309);
and U13488 (N_13488,N_13271,N_13299);
xor U13489 (N_13489,N_13232,N_13360);
and U13490 (N_13490,N_13387,N_13302);
nor U13491 (N_13491,N_13326,N_13280);
and U13492 (N_13492,N_13391,N_13327);
and U13493 (N_13493,N_13335,N_13382);
or U13494 (N_13494,N_13202,N_13345);
xnor U13495 (N_13495,N_13355,N_13383);
nand U13496 (N_13496,N_13356,N_13215);
and U13497 (N_13497,N_13217,N_13349);
nor U13498 (N_13498,N_13318,N_13212);
and U13499 (N_13499,N_13278,N_13223);
nor U13500 (N_13500,N_13261,N_13315);
nand U13501 (N_13501,N_13316,N_13347);
and U13502 (N_13502,N_13318,N_13277);
and U13503 (N_13503,N_13295,N_13389);
nand U13504 (N_13504,N_13383,N_13362);
and U13505 (N_13505,N_13322,N_13321);
or U13506 (N_13506,N_13358,N_13242);
or U13507 (N_13507,N_13296,N_13226);
nor U13508 (N_13508,N_13204,N_13257);
and U13509 (N_13509,N_13222,N_13367);
nor U13510 (N_13510,N_13221,N_13268);
nand U13511 (N_13511,N_13318,N_13331);
or U13512 (N_13512,N_13361,N_13257);
and U13513 (N_13513,N_13296,N_13206);
xnor U13514 (N_13514,N_13366,N_13215);
and U13515 (N_13515,N_13306,N_13305);
nor U13516 (N_13516,N_13349,N_13321);
nand U13517 (N_13517,N_13248,N_13298);
and U13518 (N_13518,N_13368,N_13375);
and U13519 (N_13519,N_13283,N_13202);
nor U13520 (N_13520,N_13276,N_13203);
and U13521 (N_13521,N_13394,N_13312);
nand U13522 (N_13522,N_13265,N_13244);
xor U13523 (N_13523,N_13295,N_13203);
xor U13524 (N_13524,N_13318,N_13369);
and U13525 (N_13525,N_13350,N_13388);
and U13526 (N_13526,N_13227,N_13286);
or U13527 (N_13527,N_13206,N_13383);
xnor U13528 (N_13528,N_13368,N_13328);
and U13529 (N_13529,N_13345,N_13208);
xor U13530 (N_13530,N_13370,N_13223);
xnor U13531 (N_13531,N_13243,N_13323);
nand U13532 (N_13532,N_13319,N_13398);
and U13533 (N_13533,N_13276,N_13217);
nand U13534 (N_13534,N_13270,N_13361);
and U13535 (N_13535,N_13223,N_13307);
xnor U13536 (N_13536,N_13369,N_13281);
xor U13537 (N_13537,N_13200,N_13223);
and U13538 (N_13538,N_13274,N_13320);
nand U13539 (N_13539,N_13342,N_13332);
and U13540 (N_13540,N_13366,N_13319);
nor U13541 (N_13541,N_13235,N_13234);
and U13542 (N_13542,N_13393,N_13254);
xnor U13543 (N_13543,N_13294,N_13357);
and U13544 (N_13544,N_13211,N_13258);
nor U13545 (N_13545,N_13224,N_13284);
nor U13546 (N_13546,N_13222,N_13344);
xor U13547 (N_13547,N_13293,N_13266);
nand U13548 (N_13548,N_13364,N_13397);
or U13549 (N_13549,N_13255,N_13241);
and U13550 (N_13550,N_13342,N_13279);
nor U13551 (N_13551,N_13365,N_13218);
or U13552 (N_13552,N_13395,N_13387);
nor U13553 (N_13553,N_13302,N_13383);
and U13554 (N_13554,N_13377,N_13308);
and U13555 (N_13555,N_13367,N_13207);
nor U13556 (N_13556,N_13358,N_13201);
or U13557 (N_13557,N_13234,N_13381);
nor U13558 (N_13558,N_13301,N_13338);
nand U13559 (N_13559,N_13398,N_13315);
or U13560 (N_13560,N_13306,N_13363);
nor U13561 (N_13561,N_13374,N_13225);
xnor U13562 (N_13562,N_13344,N_13353);
xnor U13563 (N_13563,N_13311,N_13372);
nor U13564 (N_13564,N_13213,N_13386);
xnor U13565 (N_13565,N_13364,N_13251);
nand U13566 (N_13566,N_13335,N_13229);
xnor U13567 (N_13567,N_13237,N_13356);
xnor U13568 (N_13568,N_13313,N_13396);
and U13569 (N_13569,N_13233,N_13295);
nand U13570 (N_13570,N_13387,N_13329);
nor U13571 (N_13571,N_13317,N_13214);
nor U13572 (N_13572,N_13303,N_13307);
nand U13573 (N_13573,N_13353,N_13366);
xor U13574 (N_13574,N_13220,N_13222);
nand U13575 (N_13575,N_13262,N_13300);
and U13576 (N_13576,N_13383,N_13350);
and U13577 (N_13577,N_13325,N_13349);
nor U13578 (N_13578,N_13358,N_13217);
and U13579 (N_13579,N_13255,N_13221);
or U13580 (N_13580,N_13242,N_13387);
nor U13581 (N_13581,N_13356,N_13300);
nand U13582 (N_13582,N_13388,N_13291);
nor U13583 (N_13583,N_13315,N_13382);
or U13584 (N_13584,N_13353,N_13331);
or U13585 (N_13585,N_13250,N_13203);
or U13586 (N_13586,N_13381,N_13391);
or U13587 (N_13587,N_13342,N_13374);
nor U13588 (N_13588,N_13207,N_13353);
xor U13589 (N_13589,N_13328,N_13348);
xor U13590 (N_13590,N_13306,N_13392);
xnor U13591 (N_13591,N_13380,N_13257);
nand U13592 (N_13592,N_13328,N_13217);
or U13593 (N_13593,N_13280,N_13351);
or U13594 (N_13594,N_13281,N_13371);
nand U13595 (N_13595,N_13291,N_13318);
and U13596 (N_13596,N_13267,N_13200);
nand U13597 (N_13597,N_13360,N_13283);
nor U13598 (N_13598,N_13306,N_13212);
nand U13599 (N_13599,N_13389,N_13251);
nor U13600 (N_13600,N_13497,N_13510);
nor U13601 (N_13601,N_13402,N_13522);
or U13602 (N_13602,N_13489,N_13438);
nor U13603 (N_13603,N_13552,N_13463);
xnor U13604 (N_13604,N_13513,N_13565);
xor U13605 (N_13605,N_13423,N_13570);
xnor U13606 (N_13606,N_13585,N_13426);
nand U13607 (N_13607,N_13542,N_13411);
xnor U13608 (N_13608,N_13450,N_13469);
nand U13609 (N_13609,N_13443,N_13418);
and U13610 (N_13610,N_13459,N_13456);
and U13611 (N_13611,N_13533,N_13435);
xnor U13612 (N_13612,N_13512,N_13567);
nand U13613 (N_13613,N_13578,N_13442);
xor U13614 (N_13614,N_13517,N_13501);
and U13615 (N_13615,N_13587,N_13477);
or U13616 (N_13616,N_13491,N_13593);
or U13617 (N_13617,N_13597,N_13556);
or U13618 (N_13618,N_13466,N_13467);
and U13619 (N_13619,N_13461,N_13596);
nor U13620 (N_13620,N_13540,N_13483);
xnor U13621 (N_13621,N_13562,N_13505);
xnor U13622 (N_13622,N_13400,N_13462);
and U13623 (N_13623,N_13569,N_13584);
nor U13624 (N_13624,N_13481,N_13473);
and U13625 (N_13625,N_13504,N_13539);
xor U13626 (N_13626,N_13547,N_13493);
and U13627 (N_13627,N_13424,N_13433);
nand U13628 (N_13628,N_13437,N_13495);
and U13629 (N_13629,N_13520,N_13531);
nand U13630 (N_13630,N_13553,N_13465);
or U13631 (N_13631,N_13591,N_13416);
or U13632 (N_13632,N_13445,N_13586);
or U13633 (N_13633,N_13490,N_13480);
nand U13634 (N_13634,N_13516,N_13492);
xnor U13635 (N_13635,N_13428,N_13452);
and U13636 (N_13636,N_13551,N_13519);
nor U13637 (N_13637,N_13496,N_13472);
nand U13638 (N_13638,N_13538,N_13577);
xnor U13639 (N_13639,N_13448,N_13415);
and U13640 (N_13640,N_13545,N_13447);
and U13641 (N_13641,N_13508,N_13529);
or U13642 (N_13642,N_13590,N_13409);
and U13643 (N_13643,N_13527,N_13460);
nand U13644 (N_13644,N_13579,N_13580);
xor U13645 (N_13645,N_13588,N_13576);
nor U13646 (N_13646,N_13475,N_13482);
nor U13647 (N_13647,N_13509,N_13430);
xor U13648 (N_13648,N_13449,N_13468);
and U13649 (N_13649,N_13521,N_13589);
or U13650 (N_13650,N_13573,N_13454);
xnor U13651 (N_13651,N_13431,N_13524);
or U13652 (N_13652,N_13421,N_13559);
nand U13653 (N_13653,N_13534,N_13549);
or U13654 (N_13654,N_13500,N_13506);
xor U13655 (N_13655,N_13476,N_13582);
xor U13656 (N_13656,N_13439,N_13478);
xnor U13657 (N_13657,N_13571,N_13403);
nor U13658 (N_13658,N_13457,N_13494);
or U13659 (N_13659,N_13499,N_13432);
or U13660 (N_13660,N_13484,N_13436);
and U13661 (N_13661,N_13440,N_13548);
nand U13662 (N_13662,N_13557,N_13518);
and U13663 (N_13663,N_13404,N_13444);
nand U13664 (N_13664,N_13486,N_13572);
and U13665 (N_13665,N_13446,N_13474);
and U13666 (N_13666,N_13554,N_13406);
nand U13667 (N_13667,N_13498,N_13470);
or U13668 (N_13668,N_13544,N_13511);
nand U13669 (N_13669,N_13427,N_13414);
nand U13670 (N_13670,N_13417,N_13599);
and U13671 (N_13671,N_13455,N_13488);
or U13672 (N_13672,N_13575,N_13598);
xor U13673 (N_13673,N_13537,N_13407);
nor U13674 (N_13674,N_13425,N_13543);
or U13675 (N_13675,N_13583,N_13558);
and U13676 (N_13676,N_13479,N_13581);
or U13677 (N_13677,N_13507,N_13550);
xor U13678 (N_13678,N_13555,N_13530);
xnor U13679 (N_13679,N_13526,N_13405);
nor U13680 (N_13680,N_13528,N_13429);
nand U13681 (N_13681,N_13422,N_13453);
and U13682 (N_13682,N_13458,N_13546);
xnor U13683 (N_13683,N_13592,N_13523);
nand U13684 (N_13684,N_13568,N_13560);
and U13685 (N_13685,N_13564,N_13485);
or U13686 (N_13686,N_13420,N_13412);
and U13687 (N_13687,N_13561,N_13541);
nor U13688 (N_13688,N_13535,N_13408);
nor U13689 (N_13689,N_13595,N_13594);
xor U13690 (N_13690,N_13515,N_13464);
nand U13691 (N_13691,N_13410,N_13419);
or U13692 (N_13692,N_13503,N_13441);
and U13693 (N_13693,N_13536,N_13401);
nand U13694 (N_13694,N_13451,N_13574);
or U13695 (N_13695,N_13471,N_13413);
xnor U13696 (N_13696,N_13514,N_13502);
nand U13697 (N_13697,N_13563,N_13487);
nand U13698 (N_13698,N_13566,N_13532);
nand U13699 (N_13699,N_13525,N_13434);
and U13700 (N_13700,N_13445,N_13574);
or U13701 (N_13701,N_13599,N_13503);
nor U13702 (N_13702,N_13404,N_13439);
xnor U13703 (N_13703,N_13576,N_13552);
xor U13704 (N_13704,N_13435,N_13491);
xnor U13705 (N_13705,N_13428,N_13575);
xnor U13706 (N_13706,N_13402,N_13561);
nand U13707 (N_13707,N_13532,N_13429);
nand U13708 (N_13708,N_13514,N_13442);
nand U13709 (N_13709,N_13404,N_13453);
nor U13710 (N_13710,N_13496,N_13498);
nand U13711 (N_13711,N_13496,N_13500);
or U13712 (N_13712,N_13486,N_13456);
nand U13713 (N_13713,N_13583,N_13497);
nor U13714 (N_13714,N_13533,N_13550);
or U13715 (N_13715,N_13400,N_13423);
xnor U13716 (N_13716,N_13547,N_13401);
and U13717 (N_13717,N_13590,N_13556);
nor U13718 (N_13718,N_13462,N_13441);
xor U13719 (N_13719,N_13405,N_13414);
nor U13720 (N_13720,N_13527,N_13567);
xnor U13721 (N_13721,N_13447,N_13555);
nor U13722 (N_13722,N_13469,N_13594);
nor U13723 (N_13723,N_13574,N_13500);
nand U13724 (N_13724,N_13478,N_13492);
or U13725 (N_13725,N_13475,N_13519);
or U13726 (N_13726,N_13455,N_13535);
and U13727 (N_13727,N_13408,N_13481);
xor U13728 (N_13728,N_13599,N_13461);
nand U13729 (N_13729,N_13556,N_13554);
nand U13730 (N_13730,N_13521,N_13595);
or U13731 (N_13731,N_13588,N_13448);
or U13732 (N_13732,N_13586,N_13464);
nand U13733 (N_13733,N_13402,N_13578);
xor U13734 (N_13734,N_13455,N_13475);
and U13735 (N_13735,N_13513,N_13419);
or U13736 (N_13736,N_13572,N_13503);
nor U13737 (N_13737,N_13419,N_13453);
nand U13738 (N_13738,N_13535,N_13523);
or U13739 (N_13739,N_13406,N_13435);
and U13740 (N_13740,N_13401,N_13429);
or U13741 (N_13741,N_13507,N_13413);
xor U13742 (N_13742,N_13508,N_13540);
nand U13743 (N_13743,N_13417,N_13466);
nand U13744 (N_13744,N_13559,N_13501);
or U13745 (N_13745,N_13443,N_13434);
and U13746 (N_13746,N_13575,N_13466);
nand U13747 (N_13747,N_13552,N_13489);
nor U13748 (N_13748,N_13438,N_13466);
or U13749 (N_13749,N_13439,N_13412);
and U13750 (N_13750,N_13472,N_13540);
nor U13751 (N_13751,N_13432,N_13523);
nand U13752 (N_13752,N_13577,N_13435);
or U13753 (N_13753,N_13515,N_13540);
xor U13754 (N_13754,N_13444,N_13507);
xor U13755 (N_13755,N_13563,N_13503);
xor U13756 (N_13756,N_13536,N_13473);
nor U13757 (N_13757,N_13568,N_13445);
nor U13758 (N_13758,N_13489,N_13465);
and U13759 (N_13759,N_13511,N_13593);
nand U13760 (N_13760,N_13489,N_13594);
nor U13761 (N_13761,N_13468,N_13526);
xnor U13762 (N_13762,N_13465,N_13413);
or U13763 (N_13763,N_13417,N_13506);
nand U13764 (N_13764,N_13570,N_13528);
and U13765 (N_13765,N_13565,N_13557);
nor U13766 (N_13766,N_13419,N_13598);
nor U13767 (N_13767,N_13534,N_13579);
xor U13768 (N_13768,N_13424,N_13559);
xnor U13769 (N_13769,N_13484,N_13432);
nor U13770 (N_13770,N_13447,N_13540);
xor U13771 (N_13771,N_13589,N_13479);
or U13772 (N_13772,N_13400,N_13597);
xor U13773 (N_13773,N_13439,N_13549);
and U13774 (N_13774,N_13446,N_13494);
xnor U13775 (N_13775,N_13514,N_13415);
and U13776 (N_13776,N_13593,N_13530);
nor U13777 (N_13777,N_13435,N_13574);
nor U13778 (N_13778,N_13485,N_13503);
xnor U13779 (N_13779,N_13499,N_13522);
and U13780 (N_13780,N_13400,N_13538);
nand U13781 (N_13781,N_13507,N_13573);
or U13782 (N_13782,N_13406,N_13545);
nor U13783 (N_13783,N_13495,N_13401);
and U13784 (N_13784,N_13457,N_13554);
xor U13785 (N_13785,N_13441,N_13495);
nor U13786 (N_13786,N_13543,N_13583);
nor U13787 (N_13787,N_13556,N_13499);
xor U13788 (N_13788,N_13568,N_13420);
nand U13789 (N_13789,N_13549,N_13451);
and U13790 (N_13790,N_13458,N_13465);
or U13791 (N_13791,N_13530,N_13570);
nand U13792 (N_13792,N_13567,N_13448);
and U13793 (N_13793,N_13546,N_13568);
xor U13794 (N_13794,N_13554,N_13527);
xnor U13795 (N_13795,N_13494,N_13540);
xor U13796 (N_13796,N_13587,N_13565);
or U13797 (N_13797,N_13465,N_13503);
xor U13798 (N_13798,N_13454,N_13516);
xor U13799 (N_13799,N_13519,N_13450);
nor U13800 (N_13800,N_13696,N_13711);
nand U13801 (N_13801,N_13743,N_13716);
nor U13802 (N_13802,N_13732,N_13715);
or U13803 (N_13803,N_13608,N_13700);
xnor U13804 (N_13804,N_13778,N_13672);
nor U13805 (N_13805,N_13767,N_13657);
xnor U13806 (N_13806,N_13603,N_13652);
nand U13807 (N_13807,N_13607,N_13624);
nand U13808 (N_13808,N_13610,N_13787);
nor U13809 (N_13809,N_13773,N_13704);
and U13810 (N_13810,N_13761,N_13695);
xor U13811 (N_13811,N_13739,N_13661);
nor U13812 (N_13812,N_13643,N_13650);
nor U13813 (N_13813,N_13762,N_13648);
xnor U13814 (N_13814,N_13702,N_13782);
xnor U13815 (N_13815,N_13678,N_13633);
xnor U13816 (N_13816,N_13737,N_13632);
or U13817 (N_13817,N_13668,N_13793);
nand U13818 (N_13818,N_13682,N_13645);
or U13819 (N_13819,N_13790,N_13740);
nor U13820 (N_13820,N_13636,N_13799);
or U13821 (N_13821,N_13712,N_13600);
or U13822 (N_13822,N_13685,N_13694);
and U13823 (N_13823,N_13775,N_13691);
nor U13824 (N_13824,N_13714,N_13635);
and U13825 (N_13825,N_13768,N_13659);
xnor U13826 (N_13826,N_13677,N_13663);
and U13827 (N_13827,N_13614,N_13777);
xor U13828 (N_13828,N_13748,N_13660);
and U13829 (N_13829,N_13779,N_13744);
and U13830 (N_13830,N_13713,N_13618);
xor U13831 (N_13831,N_13728,N_13670);
xor U13832 (N_13832,N_13613,N_13602);
nor U13833 (N_13833,N_13766,N_13674);
nor U13834 (N_13834,N_13604,N_13753);
nor U13835 (N_13835,N_13738,N_13725);
nor U13836 (N_13836,N_13797,N_13693);
and U13837 (N_13837,N_13798,N_13644);
and U13838 (N_13838,N_13749,N_13680);
and U13839 (N_13839,N_13745,N_13656);
nand U13840 (N_13840,N_13615,N_13789);
xnor U13841 (N_13841,N_13783,N_13795);
or U13842 (N_13842,N_13623,N_13676);
and U13843 (N_13843,N_13786,N_13770);
nand U13844 (N_13844,N_13673,N_13675);
nor U13845 (N_13845,N_13664,N_13781);
or U13846 (N_13846,N_13763,N_13637);
and U13847 (N_13847,N_13697,N_13785);
and U13848 (N_13848,N_13669,N_13751);
nor U13849 (N_13849,N_13601,N_13667);
nand U13850 (N_13850,N_13634,N_13662);
or U13851 (N_13851,N_13747,N_13752);
xnor U13852 (N_13852,N_13729,N_13654);
nand U13853 (N_13853,N_13709,N_13612);
nand U13854 (N_13854,N_13619,N_13622);
xnor U13855 (N_13855,N_13630,N_13647);
nor U13856 (N_13856,N_13687,N_13684);
nor U13857 (N_13857,N_13765,N_13791);
nand U13858 (N_13858,N_13774,N_13658);
nand U13859 (N_13859,N_13651,N_13719);
or U13860 (N_13860,N_13776,N_13616);
nand U13861 (N_13861,N_13655,N_13772);
nor U13862 (N_13862,N_13796,N_13758);
and U13863 (N_13863,N_13692,N_13681);
or U13864 (N_13864,N_13671,N_13717);
or U13865 (N_13865,N_13617,N_13609);
and U13866 (N_13866,N_13769,N_13741);
xor U13867 (N_13867,N_13706,N_13683);
nand U13868 (N_13868,N_13605,N_13625);
or U13869 (N_13869,N_13780,N_13720);
xor U13870 (N_13870,N_13649,N_13629);
nand U13871 (N_13871,N_13638,N_13699);
or U13872 (N_13872,N_13665,N_13701);
xor U13873 (N_13873,N_13756,N_13707);
nand U13874 (N_13874,N_13639,N_13771);
nor U13875 (N_13875,N_13759,N_13679);
xnor U13876 (N_13876,N_13606,N_13628);
and U13877 (N_13877,N_13631,N_13710);
nor U13878 (N_13878,N_13727,N_13627);
nor U13879 (N_13879,N_13734,N_13621);
nor U13880 (N_13880,N_13640,N_13689);
or U13881 (N_13881,N_13723,N_13750);
or U13882 (N_13882,N_13626,N_13754);
nand U13883 (N_13883,N_13722,N_13792);
and U13884 (N_13884,N_13794,N_13703);
and U13885 (N_13885,N_13736,N_13705);
and U13886 (N_13886,N_13666,N_13611);
xor U13887 (N_13887,N_13764,N_13698);
nor U13888 (N_13888,N_13788,N_13686);
xor U13889 (N_13889,N_13731,N_13784);
or U13890 (N_13890,N_13726,N_13620);
nand U13891 (N_13891,N_13653,N_13721);
nor U13892 (N_13892,N_13733,N_13760);
nor U13893 (N_13893,N_13646,N_13718);
xnor U13894 (N_13894,N_13735,N_13730);
nor U13895 (N_13895,N_13724,N_13708);
xnor U13896 (N_13896,N_13690,N_13742);
xnor U13897 (N_13897,N_13642,N_13688);
nor U13898 (N_13898,N_13757,N_13641);
xor U13899 (N_13899,N_13755,N_13746);
nand U13900 (N_13900,N_13623,N_13697);
xnor U13901 (N_13901,N_13621,N_13620);
and U13902 (N_13902,N_13666,N_13604);
xor U13903 (N_13903,N_13725,N_13658);
nand U13904 (N_13904,N_13734,N_13737);
nor U13905 (N_13905,N_13633,N_13709);
and U13906 (N_13906,N_13754,N_13661);
or U13907 (N_13907,N_13624,N_13625);
nand U13908 (N_13908,N_13757,N_13795);
nand U13909 (N_13909,N_13686,N_13630);
nor U13910 (N_13910,N_13796,N_13743);
nand U13911 (N_13911,N_13736,N_13726);
nand U13912 (N_13912,N_13718,N_13773);
nor U13913 (N_13913,N_13601,N_13627);
nor U13914 (N_13914,N_13637,N_13618);
or U13915 (N_13915,N_13770,N_13672);
or U13916 (N_13916,N_13723,N_13727);
and U13917 (N_13917,N_13655,N_13612);
nand U13918 (N_13918,N_13607,N_13792);
xnor U13919 (N_13919,N_13784,N_13765);
or U13920 (N_13920,N_13707,N_13709);
nor U13921 (N_13921,N_13718,N_13711);
or U13922 (N_13922,N_13617,N_13743);
or U13923 (N_13923,N_13773,N_13658);
nand U13924 (N_13924,N_13606,N_13799);
xnor U13925 (N_13925,N_13741,N_13787);
nor U13926 (N_13926,N_13646,N_13747);
or U13927 (N_13927,N_13763,N_13731);
or U13928 (N_13928,N_13752,N_13706);
xor U13929 (N_13929,N_13658,N_13637);
and U13930 (N_13930,N_13653,N_13748);
nand U13931 (N_13931,N_13721,N_13677);
xor U13932 (N_13932,N_13602,N_13645);
nor U13933 (N_13933,N_13620,N_13762);
nor U13934 (N_13934,N_13703,N_13764);
nand U13935 (N_13935,N_13679,N_13752);
or U13936 (N_13936,N_13792,N_13669);
and U13937 (N_13937,N_13648,N_13732);
or U13938 (N_13938,N_13611,N_13741);
or U13939 (N_13939,N_13768,N_13667);
and U13940 (N_13940,N_13622,N_13675);
nand U13941 (N_13941,N_13788,N_13670);
or U13942 (N_13942,N_13732,N_13778);
or U13943 (N_13943,N_13704,N_13731);
and U13944 (N_13944,N_13772,N_13795);
nand U13945 (N_13945,N_13785,N_13781);
xor U13946 (N_13946,N_13659,N_13711);
nor U13947 (N_13947,N_13711,N_13723);
nand U13948 (N_13948,N_13723,N_13780);
nor U13949 (N_13949,N_13616,N_13729);
xnor U13950 (N_13950,N_13649,N_13602);
and U13951 (N_13951,N_13731,N_13766);
xor U13952 (N_13952,N_13635,N_13716);
xor U13953 (N_13953,N_13651,N_13715);
nand U13954 (N_13954,N_13722,N_13768);
xor U13955 (N_13955,N_13784,N_13610);
xor U13956 (N_13956,N_13644,N_13615);
nor U13957 (N_13957,N_13668,N_13756);
and U13958 (N_13958,N_13740,N_13641);
nor U13959 (N_13959,N_13749,N_13621);
and U13960 (N_13960,N_13700,N_13652);
nand U13961 (N_13961,N_13646,N_13728);
and U13962 (N_13962,N_13720,N_13672);
and U13963 (N_13963,N_13703,N_13629);
xor U13964 (N_13964,N_13679,N_13743);
nor U13965 (N_13965,N_13614,N_13708);
nand U13966 (N_13966,N_13790,N_13620);
nand U13967 (N_13967,N_13756,N_13652);
xnor U13968 (N_13968,N_13726,N_13648);
nor U13969 (N_13969,N_13757,N_13794);
or U13970 (N_13970,N_13763,N_13641);
or U13971 (N_13971,N_13699,N_13689);
and U13972 (N_13972,N_13713,N_13614);
xnor U13973 (N_13973,N_13696,N_13672);
nor U13974 (N_13974,N_13628,N_13718);
nand U13975 (N_13975,N_13710,N_13781);
xnor U13976 (N_13976,N_13705,N_13794);
and U13977 (N_13977,N_13623,N_13667);
nand U13978 (N_13978,N_13713,N_13774);
nor U13979 (N_13979,N_13603,N_13788);
nor U13980 (N_13980,N_13634,N_13765);
nand U13981 (N_13981,N_13741,N_13740);
nand U13982 (N_13982,N_13679,N_13701);
nor U13983 (N_13983,N_13654,N_13712);
xor U13984 (N_13984,N_13755,N_13617);
xor U13985 (N_13985,N_13672,N_13709);
nor U13986 (N_13986,N_13601,N_13643);
nand U13987 (N_13987,N_13633,N_13754);
nor U13988 (N_13988,N_13607,N_13617);
or U13989 (N_13989,N_13687,N_13776);
nor U13990 (N_13990,N_13747,N_13660);
xnor U13991 (N_13991,N_13613,N_13689);
nand U13992 (N_13992,N_13761,N_13747);
xnor U13993 (N_13993,N_13673,N_13713);
nand U13994 (N_13994,N_13704,N_13705);
nand U13995 (N_13995,N_13718,N_13722);
xor U13996 (N_13996,N_13781,N_13601);
xnor U13997 (N_13997,N_13784,N_13686);
and U13998 (N_13998,N_13754,N_13679);
nand U13999 (N_13999,N_13621,N_13706);
xnor U14000 (N_14000,N_13998,N_13945);
nand U14001 (N_14001,N_13804,N_13852);
nor U14002 (N_14002,N_13824,N_13825);
or U14003 (N_14003,N_13978,N_13961);
nor U14004 (N_14004,N_13931,N_13964);
nor U14005 (N_14005,N_13848,N_13912);
and U14006 (N_14006,N_13937,N_13965);
nor U14007 (N_14007,N_13842,N_13935);
or U14008 (N_14008,N_13827,N_13882);
or U14009 (N_14009,N_13851,N_13969);
xnor U14010 (N_14010,N_13883,N_13806);
nand U14011 (N_14011,N_13843,N_13856);
xnor U14012 (N_14012,N_13909,N_13895);
nor U14013 (N_14013,N_13810,N_13854);
xor U14014 (N_14014,N_13832,N_13914);
nor U14015 (N_14015,N_13845,N_13836);
or U14016 (N_14016,N_13819,N_13923);
nor U14017 (N_14017,N_13812,N_13946);
nor U14018 (N_14018,N_13849,N_13947);
nand U14019 (N_14019,N_13943,N_13841);
xor U14020 (N_14020,N_13959,N_13877);
nor U14021 (N_14021,N_13902,N_13818);
nor U14022 (N_14022,N_13861,N_13980);
nand U14023 (N_14023,N_13846,N_13879);
nor U14024 (N_14024,N_13892,N_13899);
or U14025 (N_14025,N_13971,N_13829);
or U14026 (N_14026,N_13988,N_13904);
xnor U14027 (N_14027,N_13938,N_13976);
nor U14028 (N_14028,N_13839,N_13957);
nor U14029 (N_14029,N_13991,N_13894);
xor U14030 (N_14030,N_13887,N_13950);
nor U14031 (N_14031,N_13815,N_13928);
nand U14032 (N_14032,N_13990,N_13932);
nor U14033 (N_14033,N_13886,N_13996);
and U14034 (N_14034,N_13925,N_13910);
nor U14035 (N_14035,N_13906,N_13955);
nand U14036 (N_14036,N_13891,N_13911);
nor U14037 (N_14037,N_13995,N_13983);
nor U14038 (N_14038,N_13800,N_13908);
nand U14039 (N_14039,N_13954,N_13985);
and U14040 (N_14040,N_13967,N_13941);
xor U14041 (N_14041,N_13898,N_13801);
nand U14042 (N_14042,N_13913,N_13808);
nand U14043 (N_14043,N_13933,N_13835);
nor U14044 (N_14044,N_13916,N_13968);
or U14045 (N_14045,N_13974,N_13901);
nand U14046 (N_14046,N_13951,N_13949);
nor U14047 (N_14047,N_13830,N_13917);
nor U14048 (N_14048,N_13927,N_13807);
or U14049 (N_14049,N_13868,N_13867);
or U14050 (N_14050,N_13878,N_13837);
nor U14051 (N_14051,N_13940,N_13915);
xnor U14052 (N_14052,N_13885,N_13822);
and U14053 (N_14053,N_13855,N_13872);
and U14054 (N_14054,N_13926,N_13862);
xnor U14055 (N_14055,N_13817,N_13875);
and U14056 (N_14056,N_13920,N_13870);
or U14057 (N_14057,N_13874,N_13919);
and U14058 (N_14058,N_13942,N_13814);
or U14059 (N_14059,N_13864,N_13850);
xnor U14060 (N_14060,N_13813,N_13994);
and U14061 (N_14061,N_13805,N_13989);
or U14062 (N_14062,N_13860,N_13821);
nand U14063 (N_14063,N_13939,N_13953);
or U14064 (N_14064,N_13833,N_13809);
nor U14065 (N_14065,N_13958,N_13803);
nor U14066 (N_14066,N_13828,N_13962);
nor U14067 (N_14067,N_13963,N_13863);
nor U14068 (N_14068,N_13982,N_13858);
nor U14069 (N_14069,N_13979,N_13884);
and U14070 (N_14070,N_13922,N_13897);
nand U14071 (N_14071,N_13993,N_13973);
and U14072 (N_14072,N_13934,N_13929);
nand U14073 (N_14073,N_13888,N_13900);
nor U14074 (N_14074,N_13880,N_13890);
nor U14075 (N_14075,N_13987,N_13834);
and U14076 (N_14076,N_13966,N_13918);
and U14077 (N_14077,N_13986,N_13811);
nor U14078 (N_14078,N_13847,N_13992);
or U14079 (N_14079,N_13936,N_13840);
nor U14080 (N_14080,N_13873,N_13831);
nand U14081 (N_14081,N_13869,N_13997);
nor U14082 (N_14082,N_13970,N_13905);
nand U14083 (N_14083,N_13881,N_13820);
xnor U14084 (N_14084,N_13859,N_13865);
nor U14085 (N_14085,N_13921,N_13889);
nor U14086 (N_14086,N_13844,N_13981);
xnor U14087 (N_14087,N_13975,N_13952);
xor U14088 (N_14088,N_13896,N_13956);
or U14089 (N_14089,N_13903,N_13977);
nand U14090 (N_14090,N_13838,N_13972);
nor U14091 (N_14091,N_13816,N_13823);
or U14092 (N_14092,N_13802,N_13999);
or U14093 (N_14093,N_13930,N_13871);
and U14094 (N_14094,N_13893,N_13853);
or U14095 (N_14095,N_13984,N_13924);
and U14096 (N_14096,N_13960,N_13866);
nand U14097 (N_14097,N_13876,N_13948);
xnor U14098 (N_14098,N_13907,N_13826);
and U14099 (N_14099,N_13857,N_13944);
and U14100 (N_14100,N_13954,N_13850);
or U14101 (N_14101,N_13899,N_13997);
nor U14102 (N_14102,N_13804,N_13964);
nor U14103 (N_14103,N_13992,N_13801);
or U14104 (N_14104,N_13966,N_13871);
nand U14105 (N_14105,N_13886,N_13905);
or U14106 (N_14106,N_13938,N_13989);
nor U14107 (N_14107,N_13888,N_13953);
and U14108 (N_14108,N_13983,N_13879);
xnor U14109 (N_14109,N_13818,N_13952);
or U14110 (N_14110,N_13816,N_13900);
nor U14111 (N_14111,N_13872,N_13937);
and U14112 (N_14112,N_13845,N_13960);
xnor U14113 (N_14113,N_13929,N_13940);
xor U14114 (N_14114,N_13848,N_13802);
or U14115 (N_14115,N_13904,N_13867);
or U14116 (N_14116,N_13896,N_13930);
nand U14117 (N_14117,N_13916,N_13800);
xor U14118 (N_14118,N_13997,N_13951);
nand U14119 (N_14119,N_13857,N_13977);
xor U14120 (N_14120,N_13888,N_13854);
nor U14121 (N_14121,N_13998,N_13844);
nand U14122 (N_14122,N_13891,N_13871);
and U14123 (N_14123,N_13998,N_13889);
nor U14124 (N_14124,N_13936,N_13999);
and U14125 (N_14125,N_13831,N_13827);
nor U14126 (N_14126,N_13988,N_13946);
and U14127 (N_14127,N_13979,N_13829);
xor U14128 (N_14128,N_13952,N_13823);
or U14129 (N_14129,N_13891,N_13809);
or U14130 (N_14130,N_13949,N_13912);
or U14131 (N_14131,N_13982,N_13990);
xor U14132 (N_14132,N_13833,N_13835);
xor U14133 (N_14133,N_13956,N_13915);
nand U14134 (N_14134,N_13838,N_13883);
and U14135 (N_14135,N_13959,N_13847);
or U14136 (N_14136,N_13836,N_13879);
or U14137 (N_14137,N_13900,N_13889);
or U14138 (N_14138,N_13926,N_13825);
nand U14139 (N_14139,N_13997,N_13843);
nor U14140 (N_14140,N_13801,N_13857);
or U14141 (N_14141,N_13887,N_13834);
xnor U14142 (N_14142,N_13850,N_13874);
or U14143 (N_14143,N_13977,N_13976);
and U14144 (N_14144,N_13939,N_13863);
xor U14145 (N_14145,N_13946,N_13842);
nand U14146 (N_14146,N_13806,N_13981);
and U14147 (N_14147,N_13898,N_13888);
xor U14148 (N_14148,N_13832,N_13804);
xor U14149 (N_14149,N_13956,N_13916);
xnor U14150 (N_14150,N_13905,N_13975);
nor U14151 (N_14151,N_13865,N_13957);
nand U14152 (N_14152,N_13829,N_13955);
and U14153 (N_14153,N_13905,N_13994);
nand U14154 (N_14154,N_13928,N_13999);
nand U14155 (N_14155,N_13936,N_13881);
or U14156 (N_14156,N_13904,N_13991);
and U14157 (N_14157,N_13977,N_13922);
nor U14158 (N_14158,N_13865,N_13943);
xor U14159 (N_14159,N_13843,N_13887);
nor U14160 (N_14160,N_13834,N_13979);
and U14161 (N_14161,N_13872,N_13817);
nor U14162 (N_14162,N_13830,N_13927);
xor U14163 (N_14163,N_13942,N_13945);
and U14164 (N_14164,N_13877,N_13937);
and U14165 (N_14165,N_13819,N_13858);
xnor U14166 (N_14166,N_13883,N_13901);
and U14167 (N_14167,N_13969,N_13958);
nand U14168 (N_14168,N_13888,N_13837);
and U14169 (N_14169,N_13834,N_13866);
xnor U14170 (N_14170,N_13904,N_13816);
and U14171 (N_14171,N_13955,N_13919);
and U14172 (N_14172,N_13998,N_13851);
nand U14173 (N_14173,N_13958,N_13878);
nand U14174 (N_14174,N_13808,N_13892);
or U14175 (N_14175,N_13945,N_13889);
xor U14176 (N_14176,N_13819,N_13939);
xnor U14177 (N_14177,N_13983,N_13849);
and U14178 (N_14178,N_13862,N_13863);
nand U14179 (N_14179,N_13891,N_13956);
xnor U14180 (N_14180,N_13851,N_13861);
xnor U14181 (N_14181,N_13885,N_13898);
and U14182 (N_14182,N_13853,N_13943);
or U14183 (N_14183,N_13836,N_13875);
xor U14184 (N_14184,N_13952,N_13870);
xor U14185 (N_14185,N_13990,N_13824);
xnor U14186 (N_14186,N_13877,N_13972);
nor U14187 (N_14187,N_13827,N_13861);
nand U14188 (N_14188,N_13863,N_13895);
and U14189 (N_14189,N_13841,N_13935);
nand U14190 (N_14190,N_13961,N_13936);
nor U14191 (N_14191,N_13825,N_13802);
nor U14192 (N_14192,N_13813,N_13927);
nand U14193 (N_14193,N_13975,N_13928);
nand U14194 (N_14194,N_13974,N_13831);
and U14195 (N_14195,N_13926,N_13885);
nor U14196 (N_14196,N_13818,N_13978);
nor U14197 (N_14197,N_13924,N_13981);
nor U14198 (N_14198,N_13805,N_13824);
xnor U14199 (N_14199,N_13848,N_13990);
nand U14200 (N_14200,N_14062,N_14192);
and U14201 (N_14201,N_14015,N_14003);
and U14202 (N_14202,N_14004,N_14041);
nor U14203 (N_14203,N_14156,N_14180);
and U14204 (N_14204,N_14025,N_14154);
nand U14205 (N_14205,N_14103,N_14122);
nor U14206 (N_14206,N_14087,N_14105);
or U14207 (N_14207,N_14158,N_14165);
and U14208 (N_14208,N_14191,N_14001);
xnor U14209 (N_14209,N_14086,N_14173);
or U14210 (N_14210,N_14061,N_14104);
and U14211 (N_14211,N_14157,N_14076);
xor U14212 (N_14212,N_14161,N_14194);
and U14213 (N_14213,N_14054,N_14112);
nand U14214 (N_14214,N_14094,N_14106);
and U14215 (N_14215,N_14052,N_14159);
and U14216 (N_14216,N_14068,N_14029);
xnor U14217 (N_14217,N_14110,N_14189);
and U14218 (N_14218,N_14175,N_14117);
xor U14219 (N_14219,N_14126,N_14008);
xnor U14220 (N_14220,N_14199,N_14155);
and U14221 (N_14221,N_14160,N_14049);
nor U14222 (N_14222,N_14168,N_14066);
xor U14223 (N_14223,N_14114,N_14193);
xor U14224 (N_14224,N_14047,N_14034);
or U14225 (N_14225,N_14083,N_14053);
and U14226 (N_14226,N_14081,N_14151);
xnor U14227 (N_14227,N_14016,N_14065);
nor U14228 (N_14228,N_14116,N_14019);
and U14229 (N_14229,N_14095,N_14079);
or U14230 (N_14230,N_14013,N_14181);
or U14231 (N_14231,N_14098,N_14136);
and U14232 (N_14232,N_14051,N_14163);
and U14233 (N_14233,N_14190,N_14109);
and U14234 (N_14234,N_14072,N_14107);
nor U14235 (N_14235,N_14139,N_14028);
xnor U14236 (N_14236,N_14182,N_14042);
nor U14237 (N_14237,N_14164,N_14044);
and U14238 (N_14238,N_14125,N_14078);
and U14239 (N_14239,N_14134,N_14119);
xnor U14240 (N_14240,N_14070,N_14030);
or U14241 (N_14241,N_14091,N_14069);
nand U14242 (N_14242,N_14073,N_14185);
nor U14243 (N_14243,N_14142,N_14058);
or U14244 (N_14244,N_14057,N_14020);
and U14245 (N_14245,N_14133,N_14031);
xor U14246 (N_14246,N_14100,N_14021);
or U14247 (N_14247,N_14040,N_14184);
nand U14248 (N_14248,N_14082,N_14059);
and U14249 (N_14249,N_14179,N_14046);
xor U14250 (N_14250,N_14027,N_14012);
xnor U14251 (N_14251,N_14118,N_14166);
nand U14252 (N_14252,N_14140,N_14063);
nor U14253 (N_14253,N_14167,N_14036);
or U14254 (N_14254,N_14093,N_14129);
nand U14255 (N_14255,N_14141,N_14147);
or U14256 (N_14256,N_14014,N_14005);
nor U14257 (N_14257,N_14197,N_14026);
and U14258 (N_14258,N_14011,N_14131);
nor U14259 (N_14259,N_14032,N_14007);
or U14260 (N_14260,N_14077,N_14170);
and U14261 (N_14261,N_14002,N_14097);
nand U14262 (N_14262,N_14178,N_14085);
nor U14263 (N_14263,N_14138,N_14090);
nand U14264 (N_14264,N_14084,N_14121);
nor U14265 (N_14265,N_14045,N_14010);
and U14266 (N_14266,N_14128,N_14080);
or U14267 (N_14267,N_14006,N_14101);
nor U14268 (N_14268,N_14132,N_14102);
xor U14269 (N_14269,N_14064,N_14196);
xor U14270 (N_14270,N_14099,N_14187);
and U14271 (N_14271,N_14177,N_14171);
nor U14272 (N_14272,N_14035,N_14148);
nor U14273 (N_14273,N_14145,N_14198);
xnor U14274 (N_14274,N_14039,N_14037);
nand U14275 (N_14275,N_14000,N_14172);
nand U14276 (N_14276,N_14096,N_14043);
or U14277 (N_14277,N_14169,N_14195);
xnor U14278 (N_14278,N_14108,N_14137);
nand U14279 (N_14279,N_14018,N_14024);
or U14280 (N_14280,N_14023,N_14067);
or U14281 (N_14281,N_14115,N_14050);
nor U14282 (N_14282,N_14088,N_14038);
and U14283 (N_14283,N_14060,N_14146);
and U14284 (N_14284,N_14111,N_14113);
and U14285 (N_14285,N_14162,N_14149);
xor U14286 (N_14286,N_14188,N_14071);
or U14287 (N_14287,N_14153,N_14186);
xor U14288 (N_14288,N_14089,N_14176);
nor U14289 (N_14289,N_14120,N_14092);
nand U14290 (N_14290,N_14150,N_14055);
xnor U14291 (N_14291,N_14127,N_14056);
or U14292 (N_14292,N_14074,N_14009);
nor U14293 (N_14293,N_14152,N_14174);
nor U14294 (N_14294,N_14183,N_14124);
nand U14295 (N_14295,N_14144,N_14135);
nor U14296 (N_14296,N_14075,N_14022);
nor U14297 (N_14297,N_14017,N_14033);
or U14298 (N_14298,N_14130,N_14143);
nor U14299 (N_14299,N_14123,N_14048);
nor U14300 (N_14300,N_14142,N_14065);
xor U14301 (N_14301,N_14043,N_14100);
xor U14302 (N_14302,N_14002,N_14104);
nor U14303 (N_14303,N_14053,N_14019);
nor U14304 (N_14304,N_14157,N_14000);
nor U14305 (N_14305,N_14085,N_14167);
or U14306 (N_14306,N_14118,N_14175);
and U14307 (N_14307,N_14182,N_14097);
and U14308 (N_14308,N_14033,N_14035);
or U14309 (N_14309,N_14133,N_14100);
and U14310 (N_14310,N_14105,N_14096);
xnor U14311 (N_14311,N_14042,N_14121);
nor U14312 (N_14312,N_14050,N_14080);
xor U14313 (N_14313,N_14053,N_14090);
nand U14314 (N_14314,N_14044,N_14103);
or U14315 (N_14315,N_14025,N_14163);
or U14316 (N_14316,N_14132,N_14124);
nand U14317 (N_14317,N_14029,N_14120);
nand U14318 (N_14318,N_14073,N_14183);
nand U14319 (N_14319,N_14115,N_14049);
xor U14320 (N_14320,N_14088,N_14136);
nor U14321 (N_14321,N_14007,N_14033);
xor U14322 (N_14322,N_14050,N_14102);
and U14323 (N_14323,N_14003,N_14001);
and U14324 (N_14324,N_14042,N_14132);
nand U14325 (N_14325,N_14070,N_14171);
or U14326 (N_14326,N_14170,N_14063);
xor U14327 (N_14327,N_14034,N_14010);
or U14328 (N_14328,N_14079,N_14084);
or U14329 (N_14329,N_14057,N_14050);
or U14330 (N_14330,N_14068,N_14078);
nor U14331 (N_14331,N_14058,N_14079);
or U14332 (N_14332,N_14174,N_14025);
xor U14333 (N_14333,N_14071,N_14054);
nor U14334 (N_14334,N_14113,N_14086);
nor U14335 (N_14335,N_14191,N_14178);
or U14336 (N_14336,N_14055,N_14192);
nor U14337 (N_14337,N_14027,N_14118);
or U14338 (N_14338,N_14012,N_14114);
nand U14339 (N_14339,N_14150,N_14050);
nor U14340 (N_14340,N_14187,N_14014);
and U14341 (N_14341,N_14034,N_14042);
nand U14342 (N_14342,N_14146,N_14161);
and U14343 (N_14343,N_14023,N_14077);
nor U14344 (N_14344,N_14138,N_14159);
and U14345 (N_14345,N_14108,N_14156);
and U14346 (N_14346,N_14166,N_14020);
nor U14347 (N_14347,N_14007,N_14117);
nor U14348 (N_14348,N_14148,N_14107);
and U14349 (N_14349,N_14091,N_14158);
or U14350 (N_14350,N_14062,N_14052);
xnor U14351 (N_14351,N_14010,N_14016);
and U14352 (N_14352,N_14100,N_14140);
or U14353 (N_14353,N_14085,N_14109);
nand U14354 (N_14354,N_14055,N_14021);
xnor U14355 (N_14355,N_14119,N_14030);
or U14356 (N_14356,N_14197,N_14080);
or U14357 (N_14357,N_14034,N_14057);
and U14358 (N_14358,N_14162,N_14173);
xnor U14359 (N_14359,N_14069,N_14167);
nor U14360 (N_14360,N_14106,N_14184);
xor U14361 (N_14361,N_14126,N_14055);
nor U14362 (N_14362,N_14075,N_14174);
and U14363 (N_14363,N_14122,N_14014);
xnor U14364 (N_14364,N_14078,N_14177);
xnor U14365 (N_14365,N_14150,N_14093);
and U14366 (N_14366,N_14052,N_14046);
and U14367 (N_14367,N_14020,N_14181);
xor U14368 (N_14368,N_14172,N_14069);
or U14369 (N_14369,N_14155,N_14084);
xnor U14370 (N_14370,N_14183,N_14170);
nand U14371 (N_14371,N_14088,N_14059);
xnor U14372 (N_14372,N_14026,N_14024);
and U14373 (N_14373,N_14098,N_14104);
or U14374 (N_14374,N_14149,N_14116);
nor U14375 (N_14375,N_14111,N_14052);
nor U14376 (N_14376,N_14028,N_14196);
nand U14377 (N_14377,N_14133,N_14176);
nand U14378 (N_14378,N_14068,N_14062);
nand U14379 (N_14379,N_14179,N_14078);
and U14380 (N_14380,N_14054,N_14145);
nor U14381 (N_14381,N_14136,N_14148);
nor U14382 (N_14382,N_14155,N_14101);
nand U14383 (N_14383,N_14104,N_14166);
nor U14384 (N_14384,N_14066,N_14001);
xor U14385 (N_14385,N_14078,N_14123);
nand U14386 (N_14386,N_14141,N_14199);
xnor U14387 (N_14387,N_14027,N_14132);
and U14388 (N_14388,N_14166,N_14080);
nor U14389 (N_14389,N_14141,N_14129);
xnor U14390 (N_14390,N_14070,N_14129);
or U14391 (N_14391,N_14044,N_14072);
and U14392 (N_14392,N_14189,N_14158);
nor U14393 (N_14393,N_14069,N_14049);
and U14394 (N_14394,N_14051,N_14029);
xor U14395 (N_14395,N_14179,N_14016);
nor U14396 (N_14396,N_14075,N_14065);
xnor U14397 (N_14397,N_14053,N_14095);
nand U14398 (N_14398,N_14136,N_14172);
nor U14399 (N_14399,N_14086,N_14103);
or U14400 (N_14400,N_14336,N_14277);
xnor U14401 (N_14401,N_14241,N_14297);
and U14402 (N_14402,N_14389,N_14228);
nand U14403 (N_14403,N_14267,N_14239);
and U14404 (N_14404,N_14325,N_14318);
xor U14405 (N_14405,N_14375,N_14245);
xnor U14406 (N_14406,N_14327,N_14349);
nand U14407 (N_14407,N_14292,N_14324);
and U14408 (N_14408,N_14238,N_14398);
or U14409 (N_14409,N_14284,N_14202);
and U14410 (N_14410,N_14330,N_14334);
xnor U14411 (N_14411,N_14237,N_14272);
nand U14412 (N_14412,N_14328,N_14335);
xor U14413 (N_14413,N_14293,N_14259);
or U14414 (N_14414,N_14363,N_14366);
and U14415 (N_14415,N_14215,N_14354);
nand U14416 (N_14416,N_14299,N_14224);
or U14417 (N_14417,N_14344,N_14381);
xnor U14418 (N_14418,N_14214,N_14396);
and U14419 (N_14419,N_14343,N_14219);
nand U14420 (N_14420,N_14306,N_14337);
xor U14421 (N_14421,N_14294,N_14280);
nor U14422 (N_14422,N_14285,N_14218);
and U14423 (N_14423,N_14323,N_14394);
nor U14424 (N_14424,N_14244,N_14383);
and U14425 (N_14425,N_14281,N_14282);
xnor U14426 (N_14426,N_14377,N_14283);
and U14427 (N_14427,N_14257,N_14251);
nand U14428 (N_14428,N_14317,N_14248);
nor U14429 (N_14429,N_14311,N_14345);
and U14430 (N_14430,N_14268,N_14392);
or U14431 (N_14431,N_14258,N_14273);
nor U14432 (N_14432,N_14295,N_14221);
nor U14433 (N_14433,N_14376,N_14271);
xnor U14434 (N_14434,N_14379,N_14316);
or U14435 (N_14435,N_14359,N_14240);
or U14436 (N_14436,N_14395,N_14216);
nor U14437 (N_14437,N_14310,N_14233);
xnor U14438 (N_14438,N_14378,N_14230);
nand U14439 (N_14439,N_14367,N_14338);
nand U14440 (N_14440,N_14242,N_14321);
or U14441 (N_14441,N_14399,N_14225);
xnor U14442 (N_14442,N_14342,N_14264);
nand U14443 (N_14443,N_14305,N_14368);
nor U14444 (N_14444,N_14210,N_14390);
nand U14445 (N_14445,N_14351,N_14296);
nand U14446 (N_14446,N_14397,N_14226);
xnor U14447 (N_14447,N_14207,N_14331);
or U14448 (N_14448,N_14304,N_14200);
nor U14449 (N_14449,N_14320,N_14236);
or U14450 (N_14450,N_14278,N_14301);
and U14451 (N_14451,N_14246,N_14313);
and U14452 (N_14452,N_14300,N_14260);
and U14453 (N_14453,N_14235,N_14222);
nor U14454 (N_14454,N_14326,N_14266);
and U14455 (N_14455,N_14302,N_14208);
and U14456 (N_14456,N_14391,N_14234);
or U14457 (N_14457,N_14308,N_14333);
nand U14458 (N_14458,N_14357,N_14227);
nor U14459 (N_14459,N_14350,N_14322);
or U14460 (N_14460,N_14373,N_14384);
nor U14461 (N_14461,N_14358,N_14252);
or U14462 (N_14462,N_14370,N_14269);
nor U14463 (N_14463,N_14307,N_14303);
xnor U14464 (N_14464,N_14346,N_14347);
xnor U14465 (N_14465,N_14360,N_14348);
or U14466 (N_14466,N_14319,N_14388);
nand U14467 (N_14467,N_14231,N_14205);
nor U14468 (N_14468,N_14341,N_14380);
xor U14469 (N_14469,N_14209,N_14329);
nand U14470 (N_14470,N_14286,N_14365);
nand U14471 (N_14471,N_14362,N_14276);
and U14472 (N_14472,N_14374,N_14393);
and U14473 (N_14473,N_14289,N_14220);
nor U14474 (N_14474,N_14356,N_14232);
xor U14475 (N_14475,N_14386,N_14261);
xor U14476 (N_14476,N_14270,N_14217);
nor U14477 (N_14477,N_14265,N_14339);
or U14478 (N_14478,N_14352,N_14201);
nand U14479 (N_14479,N_14253,N_14262);
nor U14480 (N_14480,N_14291,N_14212);
xnor U14481 (N_14481,N_14371,N_14355);
and U14482 (N_14482,N_14247,N_14255);
nor U14483 (N_14483,N_14315,N_14361);
nor U14484 (N_14484,N_14287,N_14290);
nand U14485 (N_14485,N_14229,N_14314);
nand U14486 (N_14486,N_14206,N_14369);
nor U14487 (N_14487,N_14288,N_14256);
xnor U14488 (N_14488,N_14382,N_14372);
nand U14489 (N_14489,N_14223,N_14312);
and U14490 (N_14490,N_14387,N_14250);
or U14491 (N_14491,N_14243,N_14385);
xnor U14492 (N_14492,N_14279,N_14211);
or U14493 (N_14493,N_14274,N_14249);
nand U14494 (N_14494,N_14204,N_14213);
and U14495 (N_14495,N_14263,N_14254);
or U14496 (N_14496,N_14203,N_14353);
xor U14497 (N_14497,N_14364,N_14309);
or U14498 (N_14498,N_14340,N_14275);
nor U14499 (N_14499,N_14298,N_14332);
nor U14500 (N_14500,N_14230,N_14305);
or U14501 (N_14501,N_14250,N_14210);
and U14502 (N_14502,N_14337,N_14240);
or U14503 (N_14503,N_14315,N_14327);
xor U14504 (N_14504,N_14305,N_14306);
nor U14505 (N_14505,N_14217,N_14258);
nor U14506 (N_14506,N_14309,N_14259);
or U14507 (N_14507,N_14237,N_14326);
nand U14508 (N_14508,N_14392,N_14200);
or U14509 (N_14509,N_14339,N_14219);
xor U14510 (N_14510,N_14322,N_14223);
nand U14511 (N_14511,N_14299,N_14208);
xnor U14512 (N_14512,N_14255,N_14311);
xnor U14513 (N_14513,N_14310,N_14229);
nor U14514 (N_14514,N_14240,N_14276);
nor U14515 (N_14515,N_14395,N_14210);
nor U14516 (N_14516,N_14204,N_14252);
and U14517 (N_14517,N_14390,N_14297);
nor U14518 (N_14518,N_14210,N_14222);
and U14519 (N_14519,N_14221,N_14311);
nand U14520 (N_14520,N_14229,N_14353);
xnor U14521 (N_14521,N_14387,N_14346);
xnor U14522 (N_14522,N_14282,N_14241);
and U14523 (N_14523,N_14379,N_14381);
or U14524 (N_14524,N_14373,N_14306);
or U14525 (N_14525,N_14356,N_14282);
and U14526 (N_14526,N_14257,N_14263);
and U14527 (N_14527,N_14232,N_14373);
nor U14528 (N_14528,N_14260,N_14285);
or U14529 (N_14529,N_14365,N_14305);
or U14530 (N_14530,N_14253,N_14313);
nand U14531 (N_14531,N_14309,N_14396);
and U14532 (N_14532,N_14249,N_14352);
nand U14533 (N_14533,N_14270,N_14366);
nand U14534 (N_14534,N_14305,N_14242);
nor U14535 (N_14535,N_14375,N_14271);
or U14536 (N_14536,N_14273,N_14315);
nand U14537 (N_14537,N_14390,N_14393);
nand U14538 (N_14538,N_14234,N_14254);
nor U14539 (N_14539,N_14270,N_14285);
xnor U14540 (N_14540,N_14204,N_14229);
nor U14541 (N_14541,N_14266,N_14284);
or U14542 (N_14542,N_14279,N_14251);
nor U14543 (N_14543,N_14296,N_14200);
nor U14544 (N_14544,N_14275,N_14230);
and U14545 (N_14545,N_14362,N_14344);
and U14546 (N_14546,N_14213,N_14382);
and U14547 (N_14547,N_14274,N_14248);
xnor U14548 (N_14548,N_14317,N_14308);
or U14549 (N_14549,N_14201,N_14319);
and U14550 (N_14550,N_14236,N_14309);
nand U14551 (N_14551,N_14228,N_14303);
and U14552 (N_14552,N_14260,N_14339);
nand U14553 (N_14553,N_14266,N_14382);
xor U14554 (N_14554,N_14250,N_14347);
nand U14555 (N_14555,N_14364,N_14233);
nand U14556 (N_14556,N_14357,N_14336);
xnor U14557 (N_14557,N_14237,N_14228);
xnor U14558 (N_14558,N_14369,N_14397);
and U14559 (N_14559,N_14369,N_14260);
nand U14560 (N_14560,N_14314,N_14249);
nand U14561 (N_14561,N_14233,N_14223);
or U14562 (N_14562,N_14365,N_14310);
xor U14563 (N_14563,N_14316,N_14204);
xor U14564 (N_14564,N_14231,N_14221);
nor U14565 (N_14565,N_14369,N_14201);
nor U14566 (N_14566,N_14335,N_14298);
nand U14567 (N_14567,N_14364,N_14363);
nor U14568 (N_14568,N_14288,N_14304);
nor U14569 (N_14569,N_14266,N_14282);
nor U14570 (N_14570,N_14313,N_14372);
nand U14571 (N_14571,N_14385,N_14293);
or U14572 (N_14572,N_14323,N_14322);
xnor U14573 (N_14573,N_14308,N_14212);
nand U14574 (N_14574,N_14364,N_14291);
nor U14575 (N_14575,N_14277,N_14305);
nand U14576 (N_14576,N_14287,N_14383);
nor U14577 (N_14577,N_14386,N_14278);
or U14578 (N_14578,N_14237,N_14276);
nor U14579 (N_14579,N_14254,N_14259);
or U14580 (N_14580,N_14246,N_14264);
or U14581 (N_14581,N_14222,N_14386);
xnor U14582 (N_14582,N_14257,N_14304);
xnor U14583 (N_14583,N_14207,N_14283);
nand U14584 (N_14584,N_14234,N_14310);
and U14585 (N_14585,N_14336,N_14363);
or U14586 (N_14586,N_14320,N_14206);
nand U14587 (N_14587,N_14345,N_14331);
nor U14588 (N_14588,N_14274,N_14288);
nor U14589 (N_14589,N_14371,N_14314);
or U14590 (N_14590,N_14242,N_14261);
or U14591 (N_14591,N_14300,N_14297);
nand U14592 (N_14592,N_14291,N_14386);
xnor U14593 (N_14593,N_14253,N_14306);
and U14594 (N_14594,N_14236,N_14331);
and U14595 (N_14595,N_14308,N_14267);
nor U14596 (N_14596,N_14339,N_14350);
nor U14597 (N_14597,N_14354,N_14344);
or U14598 (N_14598,N_14287,N_14256);
nor U14599 (N_14599,N_14225,N_14267);
nand U14600 (N_14600,N_14420,N_14485);
or U14601 (N_14601,N_14502,N_14541);
or U14602 (N_14602,N_14446,N_14463);
xnor U14603 (N_14603,N_14483,N_14491);
or U14604 (N_14604,N_14560,N_14411);
xnor U14605 (N_14605,N_14469,N_14436);
or U14606 (N_14606,N_14460,N_14540);
nor U14607 (N_14607,N_14581,N_14416);
or U14608 (N_14608,N_14584,N_14578);
xnor U14609 (N_14609,N_14497,N_14415);
and U14610 (N_14610,N_14454,N_14537);
and U14611 (N_14611,N_14434,N_14533);
xnor U14612 (N_14612,N_14453,N_14574);
xnor U14613 (N_14613,N_14545,N_14448);
and U14614 (N_14614,N_14492,N_14473);
or U14615 (N_14615,N_14490,N_14400);
and U14616 (N_14616,N_14408,N_14464);
and U14617 (N_14617,N_14439,N_14573);
or U14618 (N_14618,N_14594,N_14542);
or U14619 (N_14619,N_14595,N_14539);
xor U14620 (N_14620,N_14481,N_14547);
xnor U14621 (N_14621,N_14557,N_14467);
or U14622 (N_14622,N_14493,N_14479);
and U14623 (N_14623,N_14474,N_14471);
or U14624 (N_14624,N_14546,N_14487);
and U14625 (N_14625,N_14429,N_14567);
and U14626 (N_14626,N_14597,N_14528);
xnor U14627 (N_14627,N_14449,N_14516);
xor U14628 (N_14628,N_14519,N_14402);
nor U14629 (N_14629,N_14520,N_14480);
and U14630 (N_14630,N_14455,N_14571);
and U14631 (N_14631,N_14518,N_14554);
xnor U14632 (N_14632,N_14532,N_14432);
nand U14633 (N_14633,N_14529,N_14424);
nor U14634 (N_14634,N_14462,N_14565);
nor U14635 (N_14635,N_14562,N_14538);
and U14636 (N_14636,N_14503,N_14419);
nand U14637 (N_14637,N_14468,N_14511);
nor U14638 (N_14638,N_14440,N_14409);
nor U14639 (N_14639,N_14501,N_14459);
nand U14640 (N_14640,N_14437,N_14450);
nand U14641 (N_14641,N_14580,N_14517);
xnor U14642 (N_14642,N_14593,N_14530);
and U14643 (N_14643,N_14552,N_14555);
nand U14644 (N_14644,N_14456,N_14401);
xnor U14645 (N_14645,N_14531,N_14451);
or U14646 (N_14646,N_14510,N_14404);
and U14647 (N_14647,N_14596,N_14412);
nor U14648 (N_14648,N_14452,N_14476);
or U14649 (N_14649,N_14553,N_14498);
nor U14650 (N_14650,N_14470,N_14442);
xor U14651 (N_14651,N_14522,N_14495);
xor U14652 (N_14652,N_14509,N_14421);
nand U14653 (N_14653,N_14582,N_14417);
nor U14654 (N_14654,N_14535,N_14556);
nand U14655 (N_14655,N_14489,N_14422);
xor U14656 (N_14656,N_14472,N_14423);
nand U14657 (N_14657,N_14587,N_14579);
xnor U14658 (N_14658,N_14465,N_14405);
nand U14659 (N_14659,N_14599,N_14443);
nand U14660 (N_14660,N_14575,N_14585);
nor U14661 (N_14661,N_14536,N_14568);
nand U14662 (N_14662,N_14403,N_14438);
nand U14663 (N_14663,N_14561,N_14457);
xor U14664 (N_14664,N_14407,N_14558);
or U14665 (N_14665,N_14410,N_14577);
and U14666 (N_14666,N_14505,N_14418);
nor U14667 (N_14667,N_14499,N_14583);
or U14668 (N_14668,N_14435,N_14447);
xor U14669 (N_14669,N_14482,N_14513);
nand U14670 (N_14670,N_14564,N_14592);
nor U14671 (N_14671,N_14486,N_14500);
nor U14672 (N_14672,N_14506,N_14461);
and U14673 (N_14673,N_14458,N_14572);
or U14674 (N_14674,N_14566,N_14444);
xnor U14675 (N_14675,N_14559,N_14433);
xor U14676 (N_14676,N_14523,N_14445);
and U14677 (N_14677,N_14441,N_14508);
and U14678 (N_14678,N_14524,N_14576);
xor U14679 (N_14679,N_14512,N_14543);
and U14680 (N_14680,N_14549,N_14430);
xnor U14681 (N_14681,N_14586,N_14428);
nand U14682 (N_14682,N_14504,N_14544);
and U14683 (N_14683,N_14591,N_14570);
nand U14684 (N_14684,N_14425,N_14526);
xor U14685 (N_14685,N_14477,N_14478);
nor U14686 (N_14686,N_14590,N_14488);
nand U14687 (N_14687,N_14551,N_14515);
nand U14688 (N_14688,N_14466,N_14534);
and U14689 (N_14689,N_14598,N_14494);
xnor U14690 (N_14690,N_14427,N_14475);
xnor U14691 (N_14691,N_14414,N_14525);
nand U14692 (N_14692,N_14413,N_14496);
xor U14693 (N_14693,N_14589,N_14514);
or U14694 (N_14694,N_14527,N_14521);
nor U14695 (N_14695,N_14406,N_14431);
and U14696 (N_14696,N_14507,N_14484);
nor U14697 (N_14697,N_14550,N_14563);
nor U14698 (N_14698,N_14569,N_14548);
xor U14699 (N_14699,N_14588,N_14426);
nand U14700 (N_14700,N_14410,N_14439);
nor U14701 (N_14701,N_14423,N_14547);
and U14702 (N_14702,N_14555,N_14508);
and U14703 (N_14703,N_14461,N_14469);
nor U14704 (N_14704,N_14576,N_14421);
or U14705 (N_14705,N_14466,N_14582);
or U14706 (N_14706,N_14576,N_14426);
or U14707 (N_14707,N_14534,N_14484);
xor U14708 (N_14708,N_14417,N_14510);
and U14709 (N_14709,N_14460,N_14403);
xnor U14710 (N_14710,N_14564,N_14555);
xnor U14711 (N_14711,N_14521,N_14454);
or U14712 (N_14712,N_14515,N_14469);
nor U14713 (N_14713,N_14584,N_14464);
or U14714 (N_14714,N_14562,N_14581);
xnor U14715 (N_14715,N_14475,N_14447);
or U14716 (N_14716,N_14531,N_14583);
nor U14717 (N_14717,N_14425,N_14592);
or U14718 (N_14718,N_14407,N_14501);
and U14719 (N_14719,N_14542,N_14545);
and U14720 (N_14720,N_14489,N_14437);
and U14721 (N_14721,N_14594,N_14565);
nand U14722 (N_14722,N_14546,N_14447);
and U14723 (N_14723,N_14588,N_14446);
or U14724 (N_14724,N_14445,N_14444);
and U14725 (N_14725,N_14586,N_14427);
nor U14726 (N_14726,N_14416,N_14568);
and U14727 (N_14727,N_14408,N_14451);
nand U14728 (N_14728,N_14431,N_14536);
or U14729 (N_14729,N_14570,N_14424);
nor U14730 (N_14730,N_14405,N_14434);
nor U14731 (N_14731,N_14596,N_14577);
xor U14732 (N_14732,N_14464,N_14451);
xor U14733 (N_14733,N_14447,N_14591);
nor U14734 (N_14734,N_14483,N_14593);
xnor U14735 (N_14735,N_14470,N_14587);
xnor U14736 (N_14736,N_14469,N_14416);
nor U14737 (N_14737,N_14438,N_14482);
xnor U14738 (N_14738,N_14574,N_14404);
and U14739 (N_14739,N_14476,N_14462);
nor U14740 (N_14740,N_14497,N_14417);
nor U14741 (N_14741,N_14505,N_14531);
nor U14742 (N_14742,N_14566,N_14520);
nand U14743 (N_14743,N_14497,N_14408);
nor U14744 (N_14744,N_14534,N_14554);
nand U14745 (N_14745,N_14572,N_14505);
nand U14746 (N_14746,N_14471,N_14548);
nor U14747 (N_14747,N_14513,N_14571);
or U14748 (N_14748,N_14417,N_14584);
nand U14749 (N_14749,N_14530,N_14513);
xnor U14750 (N_14750,N_14424,N_14574);
nor U14751 (N_14751,N_14486,N_14523);
nor U14752 (N_14752,N_14567,N_14457);
nor U14753 (N_14753,N_14494,N_14422);
xnor U14754 (N_14754,N_14488,N_14514);
xor U14755 (N_14755,N_14553,N_14514);
or U14756 (N_14756,N_14455,N_14407);
nor U14757 (N_14757,N_14412,N_14569);
and U14758 (N_14758,N_14532,N_14419);
nand U14759 (N_14759,N_14574,N_14400);
nor U14760 (N_14760,N_14415,N_14540);
nand U14761 (N_14761,N_14516,N_14455);
nor U14762 (N_14762,N_14508,N_14553);
nand U14763 (N_14763,N_14444,N_14542);
nor U14764 (N_14764,N_14527,N_14575);
nor U14765 (N_14765,N_14465,N_14534);
nand U14766 (N_14766,N_14435,N_14486);
nand U14767 (N_14767,N_14450,N_14500);
or U14768 (N_14768,N_14565,N_14596);
xnor U14769 (N_14769,N_14524,N_14457);
nor U14770 (N_14770,N_14483,N_14564);
nor U14771 (N_14771,N_14409,N_14517);
and U14772 (N_14772,N_14409,N_14486);
and U14773 (N_14773,N_14559,N_14427);
nor U14774 (N_14774,N_14449,N_14550);
and U14775 (N_14775,N_14515,N_14577);
xor U14776 (N_14776,N_14461,N_14507);
or U14777 (N_14777,N_14529,N_14589);
xor U14778 (N_14778,N_14450,N_14599);
nand U14779 (N_14779,N_14426,N_14418);
xor U14780 (N_14780,N_14427,N_14428);
nand U14781 (N_14781,N_14402,N_14496);
or U14782 (N_14782,N_14474,N_14599);
or U14783 (N_14783,N_14516,N_14404);
and U14784 (N_14784,N_14587,N_14441);
or U14785 (N_14785,N_14461,N_14439);
nor U14786 (N_14786,N_14401,N_14586);
xnor U14787 (N_14787,N_14402,N_14411);
and U14788 (N_14788,N_14559,N_14575);
or U14789 (N_14789,N_14431,N_14529);
xnor U14790 (N_14790,N_14477,N_14555);
or U14791 (N_14791,N_14540,N_14518);
or U14792 (N_14792,N_14474,N_14516);
and U14793 (N_14793,N_14571,N_14490);
and U14794 (N_14794,N_14445,N_14562);
or U14795 (N_14795,N_14519,N_14553);
or U14796 (N_14796,N_14458,N_14449);
nor U14797 (N_14797,N_14491,N_14553);
nor U14798 (N_14798,N_14434,N_14584);
nor U14799 (N_14799,N_14437,N_14513);
xor U14800 (N_14800,N_14743,N_14629);
or U14801 (N_14801,N_14645,N_14708);
and U14802 (N_14802,N_14658,N_14763);
nor U14803 (N_14803,N_14672,N_14607);
nand U14804 (N_14804,N_14682,N_14632);
nor U14805 (N_14805,N_14750,N_14783);
or U14806 (N_14806,N_14752,N_14730);
nand U14807 (N_14807,N_14664,N_14669);
xor U14808 (N_14808,N_14753,N_14720);
nand U14809 (N_14809,N_14751,N_14662);
xnor U14810 (N_14810,N_14697,N_14755);
or U14811 (N_14811,N_14670,N_14722);
nor U14812 (N_14812,N_14626,N_14636);
nand U14813 (N_14813,N_14721,N_14630);
nand U14814 (N_14814,N_14617,N_14698);
xnor U14815 (N_14815,N_14740,N_14719);
xnor U14816 (N_14816,N_14735,N_14631);
nand U14817 (N_14817,N_14627,N_14780);
nor U14818 (N_14818,N_14642,N_14649);
or U14819 (N_14819,N_14654,N_14709);
xnor U14820 (N_14820,N_14643,N_14726);
nor U14821 (N_14821,N_14683,N_14729);
nor U14822 (N_14822,N_14640,N_14603);
xnor U14823 (N_14823,N_14641,N_14711);
xnor U14824 (N_14824,N_14656,N_14684);
or U14825 (N_14825,N_14675,N_14718);
and U14826 (N_14826,N_14728,N_14702);
or U14827 (N_14827,N_14615,N_14772);
nor U14828 (N_14828,N_14717,N_14677);
xnor U14829 (N_14829,N_14621,N_14761);
or U14830 (N_14830,N_14614,N_14620);
or U14831 (N_14831,N_14745,N_14610);
nor U14832 (N_14832,N_14787,N_14765);
nand U14833 (N_14833,N_14706,N_14689);
and U14834 (N_14834,N_14657,N_14638);
xor U14835 (N_14835,N_14736,N_14668);
or U14836 (N_14836,N_14786,N_14696);
xnor U14837 (N_14837,N_14789,N_14609);
nand U14838 (N_14838,N_14754,N_14613);
xor U14839 (N_14839,N_14707,N_14798);
nand U14840 (N_14840,N_14681,N_14678);
or U14841 (N_14841,N_14602,N_14655);
xor U14842 (N_14842,N_14741,N_14616);
and U14843 (N_14843,N_14673,N_14608);
nor U14844 (N_14844,N_14701,N_14703);
nand U14845 (N_14845,N_14688,N_14785);
or U14846 (N_14846,N_14606,N_14674);
nor U14847 (N_14847,N_14666,N_14738);
nand U14848 (N_14848,N_14793,N_14650);
nor U14849 (N_14849,N_14625,N_14769);
nand U14850 (N_14850,N_14651,N_14747);
and U14851 (N_14851,N_14733,N_14790);
xor U14852 (N_14852,N_14797,N_14716);
nor U14853 (N_14853,N_14749,N_14796);
xor U14854 (N_14854,N_14756,N_14665);
or U14855 (N_14855,N_14639,N_14727);
nor U14856 (N_14856,N_14760,N_14795);
xnor U14857 (N_14857,N_14723,N_14634);
or U14858 (N_14858,N_14748,N_14676);
nand U14859 (N_14859,N_14660,N_14778);
or U14860 (N_14860,N_14794,N_14691);
or U14861 (N_14861,N_14724,N_14744);
and U14862 (N_14862,N_14799,N_14775);
and U14863 (N_14863,N_14746,N_14628);
nor U14864 (N_14864,N_14739,N_14771);
nand U14865 (N_14865,N_14604,N_14618);
nor U14866 (N_14866,N_14768,N_14646);
and U14867 (N_14867,N_14661,N_14762);
and U14868 (N_14868,N_14776,N_14653);
nand U14869 (N_14869,N_14791,N_14619);
nor U14870 (N_14870,N_14667,N_14659);
nand U14871 (N_14871,N_14671,N_14737);
nand U14872 (N_14872,N_14690,N_14757);
or U14873 (N_14873,N_14773,N_14770);
xor U14874 (N_14874,N_14679,N_14759);
or U14875 (N_14875,N_14622,N_14600);
and U14876 (N_14876,N_14652,N_14792);
and U14877 (N_14877,N_14637,N_14710);
and U14878 (N_14878,N_14734,N_14781);
nor U14879 (N_14879,N_14633,N_14725);
and U14880 (N_14880,N_14779,N_14695);
xor U14881 (N_14881,N_14700,N_14714);
and U14882 (N_14882,N_14731,N_14686);
or U14883 (N_14883,N_14732,N_14624);
xor U14884 (N_14884,N_14612,N_14764);
or U14885 (N_14885,N_14777,N_14713);
or U14886 (N_14886,N_14611,N_14693);
nand U14887 (N_14887,N_14774,N_14635);
nand U14888 (N_14888,N_14766,N_14647);
nand U14889 (N_14889,N_14715,N_14782);
nor U14890 (N_14890,N_14784,N_14758);
nand U14891 (N_14891,N_14742,N_14712);
nor U14892 (N_14892,N_14680,N_14663);
and U14893 (N_14893,N_14694,N_14705);
nor U14894 (N_14894,N_14601,N_14685);
nand U14895 (N_14895,N_14704,N_14692);
or U14896 (N_14896,N_14623,N_14788);
nand U14897 (N_14897,N_14644,N_14699);
xnor U14898 (N_14898,N_14767,N_14605);
and U14899 (N_14899,N_14648,N_14687);
and U14900 (N_14900,N_14706,N_14785);
and U14901 (N_14901,N_14626,N_14713);
and U14902 (N_14902,N_14789,N_14666);
nor U14903 (N_14903,N_14629,N_14762);
and U14904 (N_14904,N_14655,N_14786);
or U14905 (N_14905,N_14783,N_14678);
and U14906 (N_14906,N_14694,N_14601);
or U14907 (N_14907,N_14637,N_14685);
or U14908 (N_14908,N_14676,N_14756);
xnor U14909 (N_14909,N_14709,N_14729);
or U14910 (N_14910,N_14794,N_14653);
or U14911 (N_14911,N_14642,N_14672);
nor U14912 (N_14912,N_14712,N_14716);
and U14913 (N_14913,N_14698,N_14622);
nand U14914 (N_14914,N_14686,N_14726);
xnor U14915 (N_14915,N_14646,N_14679);
and U14916 (N_14916,N_14794,N_14722);
and U14917 (N_14917,N_14712,N_14646);
nor U14918 (N_14918,N_14717,N_14684);
or U14919 (N_14919,N_14733,N_14712);
nand U14920 (N_14920,N_14740,N_14761);
nand U14921 (N_14921,N_14680,N_14667);
nor U14922 (N_14922,N_14787,N_14694);
nand U14923 (N_14923,N_14738,N_14602);
and U14924 (N_14924,N_14695,N_14639);
xor U14925 (N_14925,N_14615,N_14726);
nand U14926 (N_14926,N_14614,N_14635);
xor U14927 (N_14927,N_14769,N_14621);
nor U14928 (N_14928,N_14717,N_14728);
nor U14929 (N_14929,N_14708,N_14669);
and U14930 (N_14930,N_14754,N_14603);
xnor U14931 (N_14931,N_14644,N_14757);
nor U14932 (N_14932,N_14627,N_14689);
and U14933 (N_14933,N_14694,N_14780);
and U14934 (N_14934,N_14717,N_14785);
and U14935 (N_14935,N_14604,N_14718);
nor U14936 (N_14936,N_14649,N_14765);
nand U14937 (N_14937,N_14731,N_14600);
xor U14938 (N_14938,N_14675,N_14769);
or U14939 (N_14939,N_14705,N_14680);
or U14940 (N_14940,N_14611,N_14761);
nor U14941 (N_14941,N_14703,N_14754);
xnor U14942 (N_14942,N_14707,N_14751);
or U14943 (N_14943,N_14760,N_14703);
nor U14944 (N_14944,N_14668,N_14672);
nand U14945 (N_14945,N_14732,N_14641);
nand U14946 (N_14946,N_14684,N_14640);
xnor U14947 (N_14947,N_14795,N_14692);
xor U14948 (N_14948,N_14712,N_14658);
nor U14949 (N_14949,N_14750,N_14729);
nor U14950 (N_14950,N_14605,N_14742);
nor U14951 (N_14951,N_14628,N_14735);
and U14952 (N_14952,N_14782,N_14795);
xor U14953 (N_14953,N_14654,N_14689);
nand U14954 (N_14954,N_14704,N_14650);
nand U14955 (N_14955,N_14785,N_14789);
xnor U14956 (N_14956,N_14746,N_14694);
or U14957 (N_14957,N_14724,N_14688);
nand U14958 (N_14958,N_14768,N_14610);
and U14959 (N_14959,N_14761,N_14626);
nor U14960 (N_14960,N_14757,N_14692);
nor U14961 (N_14961,N_14608,N_14630);
nor U14962 (N_14962,N_14655,N_14771);
and U14963 (N_14963,N_14647,N_14697);
xor U14964 (N_14964,N_14669,N_14705);
nand U14965 (N_14965,N_14720,N_14681);
and U14966 (N_14966,N_14662,N_14622);
nor U14967 (N_14967,N_14795,N_14749);
and U14968 (N_14968,N_14601,N_14754);
nor U14969 (N_14969,N_14775,N_14783);
and U14970 (N_14970,N_14655,N_14653);
nand U14971 (N_14971,N_14643,N_14758);
xnor U14972 (N_14972,N_14760,N_14793);
or U14973 (N_14973,N_14751,N_14609);
and U14974 (N_14974,N_14652,N_14675);
nor U14975 (N_14975,N_14607,N_14647);
or U14976 (N_14976,N_14627,N_14714);
or U14977 (N_14977,N_14707,N_14768);
or U14978 (N_14978,N_14647,N_14726);
xnor U14979 (N_14979,N_14778,N_14671);
nand U14980 (N_14980,N_14611,N_14755);
nand U14981 (N_14981,N_14675,N_14670);
nand U14982 (N_14982,N_14711,N_14694);
and U14983 (N_14983,N_14687,N_14606);
and U14984 (N_14984,N_14696,N_14690);
xnor U14985 (N_14985,N_14641,N_14785);
or U14986 (N_14986,N_14658,N_14605);
nand U14987 (N_14987,N_14722,N_14657);
nand U14988 (N_14988,N_14653,N_14698);
nor U14989 (N_14989,N_14784,N_14776);
nor U14990 (N_14990,N_14673,N_14791);
or U14991 (N_14991,N_14698,N_14747);
xnor U14992 (N_14992,N_14614,N_14725);
or U14993 (N_14993,N_14724,N_14715);
nand U14994 (N_14994,N_14668,N_14614);
and U14995 (N_14995,N_14633,N_14693);
xnor U14996 (N_14996,N_14674,N_14687);
xnor U14997 (N_14997,N_14746,N_14752);
nor U14998 (N_14998,N_14720,N_14601);
nand U14999 (N_14999,N_14762,N_14657);
and U15000 (N_15000,N_14982,N_14840);
or U15001 (N_15001,N_14912,N_14977);
nand U15002 (N_15002,N_14896,N_14957);
or U15003 (N_15003,N_14891,N_14954);
and U15004 (N_15004,N_14932,N_14828);
xnor U15005 (N_15005,N_14809,N_14919);
nor U15006 (N_15006,N_14878,N_14899);
nor U15007 (N_15007,N_14991,N_14830);
or U15008 (N_15008,N_14835,N_14881);
nor U15009 (N_15009,N_14858,N_14903);
nand U15010 (N_15010,N_14998,N_14975);
nor U15011 (N_15011,N_14940,N_14846);
nor U15012 (N_15012,N_14814,N_14851);
and U15013 (N_15013,N_14813,N_14883);
nand U15014 (N_15014,N_14887,N_14861);
nand U15015 (N_15015,N_14965,N_14870);
and U15016 (N_15016,N_14807,N_14923);
xor U15017 (N_15017,N_14911,N_14889);
nor U15018 (N_15018,N_14986,N_14852);
xnor U15019 (N_15019,N_14875,N_14926);
nor U15020 (N_15020,N_14948,N_14951);
xor U15021 (N_15021,N_14946,N_14880);
or U15022 (N_15022,N_14959,N_14906);
or U15023 (N_15023,N_14818,N_14990);
xor U15024 (N_15024,N_14824,N_14925);
or U15025 (N_15025,N_14964,N_14897);
nand U15026 (N_15026,N_14847,N_14869);
nand U15027 (N_15027,N_14812,N_14848);
nand U15028 (N_15028,N_14934,N_14928);
nand U15029 (N_15029,N_14850,N_14842);
nand U15030 (N_15030,N_14819,N_14958);
or U15031 (N_15031,N_14989,N_14803);
xor U15032 (N_15032,N_14826,N_14933);
or U15033 (N_15033,N_14987,N_14993);
or U15034 (N_15034,N_14973,N_14873);
or U15035 (N_15035,N_14862,N_14844);
nand U15036 (N_15036,N_14865,N_14909);
nand U15037 (N_15037,N_14985,N_14882);
and U15038 (N_15038,N_14963,N_14944);
xnor U15039 (N_15039,N_14931,N_14829);
nand U15040 (N_15040,N_14833,N_14856);
or U15041 (N_15041,N_14943,N_14902);
and U15042 (N_15042,N_14885,N_14930);
and U15043 (N_15043,N_14872,N_14811);
nand U15044 (N_15044,N_14997,N_14917);
xor U15045 (N_15045,N_14970,N_14994);
nand U15046 (N_15046,N_14960,N_14966);
nor U15047 (N_15047,N_14984,N_14901);
and U15048 (N_15048,N_14995,N_14927);
xnor U15049 (N_15049,N_14996,N_14821);
and U15050 (N_15050,N_14941,N_14810);
and U15051 (N_15051,N_14854,N_14894);
or U15052 (N_15052,N_14808,N_14999);
and U15053 (N_15053,N_14866,N_14949);
xor U15054 (N_15054,N_14815,N_14979);
or U15055 (N_15055,N_14859,N_14886);
or U15056 (N_15056,N_14841,N_14962);
or U15057 (N_15057,N_14893,N_14860);
nor U15058 (N_15058,N_14913,N_14825);
and U15059 (N_15059,N_14974,N_14904);
or U15060 (N_15060,N_14976,N_14969);
and U15061 (N_15061,N_14947,N_14898);
nand U15062 (N_15062,N_14950,N_14867);
or U15063 (N_15063,N_14879,N_14900);
and U15064 (N_15064,N_14980,N_14956);
xnor U15065 (N_15065,N_14817,N_14800);
and U15066 (N_15066,N_14955,N_14914);
nor U15067 (N_15067,N_14876,N_14924);
xnor U15068 (N_15068,N_14968,N_14961);
nand U15069 (N_15069,N_14849,N_14802);
xor U15070 (N_15070,N_14929,N_14857);
and U15071 (N_15071,N_14972,N_14945);
xnor U15072 (N_15072,N_14915,N_14806);
or U15073 (N_15073,N_14978,N_14804);
or U15074 (N_15074,N_14910,N_14922);
or U15075 (N_15075,N_14822,N_14936);
nor U15076 (N_15076,N_14992,N_14845);
or U15077 (N_15077,N_14871,N_14868);
nand U15078 (N_15078,N_14938,N_14983);
nand U15079 (N_15079,N_14839,N_14877);
and U15080 (N_15080,N_14939,N_14988);
and U15081 (N_15081,N_14953,N_14864);
and U15082 (N_15082,N_14853,N_14908);
nand U15083 (N_15083,N_14905,N_14920);
xnor U15084 (N_15084,N_14942,N_14937);
nand U15085 (N_15085,N_14836,N_14921);
nand U15086 (N_15086,N_14832,N_14907);
nor U15087 (N_15087,N_14918,N_14831);
nand U15088 (N_15088,N_14838,N_14837);
nand U15089 (N_15089,N_14874,N_14935);
nor U15090 (N_15090,N_14916,N_14827);
or U15091 (N_15091,N_14981,N_14863);
nand U15092 (N_15092,N_14823,N_14820);
and U15093 (N_15093,N_14967,N_14952);
xnor U15094 (N_15094,N_14884,N_14816);
nand U15095 (N_15095,N_14805,N_14843);
nand U15096 (N_15096,N_14890,N_14971);
and U15097 (N_15097,N_14834,N_14892);
nand U15098 (N_15098,N_14888,N_14895);
xnor U15099 (N_15099,N_14855,N_14801);
nor U15100 (N_15100,N_14802,N_14961);
or U15101 (N_15101,N_14874,N_14991);
xor U15102 (N_15102,N_14990,N_14807);
nand U15103 (N_15103,N_14821,N_14993);
or U15104 (N_15104,N_14941,N_14945);
and U15105 (N_15105,N_14985,N_14858);
xor U15106 (N_15106,N_14931,N_14827);
nor U15107 (N_15107,N_14925,N_14896);
xnor U15108 (N_15108,N_14979,N_14848);
and U15109 (N_15109,N_14830,N_14990);
or U15110 (N_15110,N_14873,N_14875);
or U15111 (N_15111,N_14998,N_14816);
xor U15112 (N_15112,N_14843,N_14895);
nand U15113 (N_15113,N_14916,N_14961);
and U15114 (N_15114,N_14896,N_14959);
nor U15115 (N_15115,N_14937,N_14944);
xor U15116 (N_15116,N_14905,N_14820);
xnor U15117 (N_15117,N_14930,N_14965);
or U15118 (N_15118,N_14834,N_14863);
or U15119 (N_15119,N_14811,N_14969);
nor U15120 (N_15120,N_14803,N_14908);
and U15121 (N_15121,N_14920,N_14856);
nand U15122 (N_15122,N_14924,N_14966);
nand U15123 (N_15123,N_14877,N_14972);
and U15124 (N_15124,N_14966,N_14979);
nor U15125 (N_15125,N_14849,N_14816);
and U15126 (N_15126,N_14993,N_14886);
xnor U15127 (N_15127,N_14866,N_14912);
nand U15128 (N_15128,N_14866,N_14880);
and U15129 (N_15129,N_14819,N_14919);
and U15130 (N_15130,N_14837,N_14859);
nand U15131 (N_15131,N_14974,N_14860);
nand U15132 (N_15132,N_14840,N_14870);
nor U15133 (N_15133,N_14912,N_14804);
xnor U15134 (N_15134,N_14806,N_14974);
or U15135 (N_15135,N_14825,N_14959);
nand U15136 (N_15136,N_14854,N_14939);
nand U15137 (N_15137,N_14985,N_14964);
nor U15138 (N_15138,N_14949,N_14876);
nor U15139 (N_15139,N_14890,N_14912);
nor U15140 (N_15140,N_14881,N_14811);
or U15141 (N_15141,N_14916,N_14877);
and U15142 (N_15142,N_14896,N_14863);
and U15143 (N_15143,N_14897,N_14909);
or U15144 (N_15144,N_14863,N_14883);
nand U15145 (N_15145,N_14848,N_14932);
nor U15146 (N_15146,N_14801,N_14979);
and U15147 (N_15147,N_14904,N_14895);
or U15148 (N_15148,N_14874,N_14865);
xnor U15149 (N_15149,N_14996,N_14999);
nor U15150 (N_15150,N_14827,N_14898);
nor U15151 (N_15151,N_14938,N_14927);
nand U15152 (N_15152,N_14995,N_14975);
or U15153 (N_15153,N_14910,N_14937);
or U15154 (N_15154,N_14826,N_14880);
nor U15155 (N_15155,N_14981,N_14979);
nor U15156 (N_15156,N_14814,N_14802);
nor U15157 (N_15157,N_14990,N_14984);
nor U15158 (N_15158,N_14826,N_14876);
xnor U15159 (N_15159,N_14851,N_14921);
nor U15160 (N_15160,N_14828,N_14929);
and U15161 (N_15161,N_14993,N_14819);
or U15162 (N_15162,N_14847,N_14972);
and U15163 (N_15163,N_14901,N_14849);
xor U15164 (N_15164,N_14900,N_14995);
nor U15165 (N_15165,N_14866,N_14913);
or U15166 (N_15166,N_14828,N_14853);
nor U15167 (N_15167,N_14987,N_14926);
nand U15168 (N_15168,N_14871,N_14886);
nand U15169 (N_15169,N_14938,N_14811);
nand U15170 (N_15170,N_14975,N_14941);
or U15171 (N_15171,N_14938,N_14974);
or U15172 (N_15172,N_14964,N_14915);
or U15173 (N_15173,N_14924,N_14807);
or U15174 (N_15174,N_14921,N_14969);
nand U15175 (N_15175,N_14956,N_14990);
xnor U15176 (N_15176,N_14986,N_14802);
or U15177 (N_15177,N_14906,N_14907);
and U15178 (N_15178,N_14979,N_14814);
nand U15179 (N_15179,N_14828,N_14999);
xnor U15180 (N_15180,N_14904,N_14896);
nor U15181 (N_15181,N_14890,N_14879);
and U15182 (N_15182,N_14920,N_14837);
or U15183 (N_15183,N_14824,N_14825);
xor U15184 (N_15184,N_14972,N_14906);
xnor U15185 (N_15185,N_14923,N_14934);
nor U15186 (N_15186,N_14843,N_14945);
xnor U15187 (N_15187,N_14837,N_14941);
or U15188 (N_15188,N_14991,N_14949);
xnor U15189 (N_15189,N_14918,N_14826);
or U15190 (N_15190,N_14992,N_14892);
xnor U15191 (N_15191,N_14990,N_14988);
and U15192 (N_15192,N_14906,N_14977);
xnor U15193 (N_15193,N_14936,N_14961);
nor U15194 (N_15194,N_14842,N_14920);
xor U15195 (N_15195,N_14987,N_14818);
or U15196 (N_15196,N_14885,N_14824);
xnor U15197 (N_15197,N_14832,N_14817);
nand U15198 (N_15198,N_14830,N_14850);
and U15199 (N_15199,N_14803,N_14874);
xor U15200 (N_15200,N_15173,N_15038);
or U15201 (N_15201,N_15082,N_15140);
nor U15202 (N_15202,N_15129,N_15064);
xnor U15203 (N_15203,N_15090,N_15161);
nor U15204 (N_15204,N_15124,N_15123);
xor U15205 (N_15205,N_15199,N_15126);
nor U15206 (N_15206,N_15174,N_15007);
nand U15207 (N_15207,N_15139,N_15097);
xnor U15208 (N_15208,N_15182,N_15115);
xnor U15209 (N_15209,N_15109,N_15025);
nor U15210 (N_15210,N_15148,N_15169);
or U15211 (N_15211,N_15177,N_15049);
and U15212 (N_15212,N_15046,N_15010);
and U15213 (N_15213,N_15145,N_15181);
xor U15214 (N_15214,N_15059,N_15119);
or U15215 (N_15215,N_15063,N_15144);
or U15216 (N_15216,N_15114,N_15078);
and U15217 (N_15217,N_15080,N_15015);
nor U15218 (N_15218,N_15089,N_15167);
xnor U15219 (N_15219,N_15093,N_15157);
xnor U15220 (N_15220,N_15088,N_15076);
xor U15221 (N_15221,N_15164,N_15155);
and U15222 (N_15222,N_15104,N_15185);
and U15223 (N_15223,N_15037,N_15122);
and U15224 (N_15224,N_15194,N_15081);
nand U15225 (N_15225,N_15047,N_15018);
or U15226 (N_15226,N_15055,N_15065);
xnor U15227 (N_15227,N_15006,N_15075);
nor U15228 (N_15228,N_15094,N_15153);
nor U15229 (N_15229,N_15100,N_15011);
and U15230 (N_15230,N_15019,N_15176);
xor U15231 (N_15231,N_15195,N_15067);
nand U15232 (N_15232,N_15004,N_15039);
and U15233 (N_15233,N_15077,N_15156);
nand U15234 (N_15234,N_15068,N_15092);
xnor U15235 (N_15235,N_15095,N_15186);
nand U15236 (N_15236,N_15151,N_15178);
or U15237 (N_15237,N_15134,N_15086);
xor U15238 (N_15238,N_15105,N_15052);
or U15239 (N_15239,N_15158,N_15184);
nor U15240 (N_15240,N_15131,N_15034);
xor U15241 (N_15241,N_15009,N_15137);
and U15242 (N_15242,N_15159,N_15027);
or U15243 (N_15243,N_15024,N_15172);
and U15244 (N_15244,N_15036,N_15111);
xor U15245 (N_15245,N_15026,N_15099);
nor U15246 (N_15246,N_15053,N_15168);
and U15247 (N_15247,N_15031,N_15060);
or U15248 (N_15248,N_15113,N_15147);
xor U15249 (N_15249,N_15187,N_15045);
or U15250 (N_15250,N_15069,N_15012);
nand U15251 (N_15251,N_15020,N_15141);
nor U15252 (N_15252,N_15127,N_15021);
nand U15253 (N_15253,N_15190,N_15016);
or U15254 (N_15254,N_15183,N_15170);
xnor U15255 (N_15255,N_15035,N_15149);
or U15256 (N_15256,N_15091,N_15056);
nand U15257 (N_15257,N_15108,N_15061);
nor U15258 (N_15258,N_15058,N_15180);
nor U15259 (N_15259,N_15192,N_15085);
xnor U15260 (N_15260,N_15198,N_15118);
and U15261 (N_15261,N_15022,N_15073);
nor U15262 (N_15262,N_15101,N_15003);
xor U15263 (N_15263,N_15128,N_15146);
or U15264 (N_15264,N_15107,N_15001);
nor U15265 (N_15265,N_15032,N_15071);
xnor U15266 (N_15266,N_15166,N_15130);
xor U15267 (N_15267,N_15057,N_15066);
xnor U15268 (N_15268,N_15084,N_15112);
nor U15269 (N_15269,N_15098,N_15013);
or U15270 (N_15270,N_15005,N_15029);
nand U15271 (N_15271,N_15048,N_15162);
xor U15272 (N_15272,N_15040,N_15044);
and U15273 (N_15273,N_15138,N_15103);
and U15274 (N_15274,N_15041,N_15179);
nand U15275 (N_15275,N_15121,N_15165);
nand U15276 (N_15276,N_15117,N_15062);
and U15277 (N_15277,N_15175,N_15125);
or U15278 (N_15278,N_15028,N_15196);
xor U15279 (N_15279,N_15023,N_15030);
and U15280 (N_15280,N_15171,N_15154);
xnor U15281 (N_15281,N_15106,N_15096);
or U15282 (N_15282,N_15132,N_15017);
nor U15283 (N_15283,N_15083,N_15143);
nand U15284 (N_15284,N_15120,N_15191);
and U15285 (N_15285,N_15150,N_15163);
nor U15286 (N_15286,N_15000,N_15142);
nand U15287 (N_15287,N_15002,N_15043);
nand U15288 (N_15288,N_15133,N_15110);
or U15289 (N_15289,N_15050,N_15054);
or U15290 (N_15290,N_15136,N_15193);
nor U15291 (N_15291,N_15072,N_15160);
and U15292 (N_15292,N_15189,N_15102);
and U15293 (N_15293,N_15079,N_15188);
xnor U15294 (N_15294,N_15033,N_15135);
and U15295 (N_15295,N_15197,N_15014);
or U15296 (N_15296,N_15074,N_15070);
xor U15297 (N_15297,N_15152,N_15116);
and U15298 (N_15298,N_15042,N_15087);
nand U15299 (N_15299,N_15051,N_15008);
or U15300 (N_15300,N_15182,N_15102);
nor U15301 (N_15301,N_15153,N_15136);
nor U15302 (N_15302,N_15006,N_15077);
xnor U15303 (N_15303,N_15150,N_15025);
xnor U15304 (N_15304,N_15020,N_15118);
nor U15305 (N_15305,N_15032,N_15000);
nor U15306 (N_15306,N_15013,N_15047);
nand U15307 (N_15307,N_15140,N_15108);
nor U15308 (N_15308,N_15071,N_15159);
xnor U15309 (N_15309,N_15198,N_15089);
xnor U15310 (N_15310,N_15187,N_15190);
nand U15311 (N_15311,N_15039,N_15128);
nor U15312 (N_15312,N_15181,N_15162);
nand U15313 (N_15313,N_15176,N_15051);
nor U15314 (N_15314,N_15029,N_15049);
or U15315 (N_15315,N_15015,N_15049);
nand U15316 (N_15316,N_15091,N_15024);
nand U15317 (N_15317,N_15194,N_15050);
or U15318 (N_15318,N_15030,N_15067);
nand U15319 (N_15319,N_15182,N_15192);
nor U15320 (N_15320,N_15108,N_15016);
or U15321 (N_15321,N_15115,N_15199);
or U15322 (N_15322,N_15079,N_15099);
or U15323 (N_15323,N_15041,N_15089);
or U15324 (N_15324,N_15061,N_15071);
and U15325 (N_15325,N_15141,N_15112);
nand U15326 (N_15326,N_15127,N_15029);
nor U15327 (N_15327,N_15178,N_15078);
or U15328 (N_15328,N_15125,N_15027);
nand U15329 (N_15329,N_15069,N_15134);
nand U15330 (N_15330,N_15082,N_15192);
xnor U15331 (N_15331,N_15178,N_15003);
and U15332 (N_15332,N_15014,N_15189);
xor U15333 (N_15333,N_15168,N_15162);
and U15334 (N_15334,N_15160,N_15019);
nand U15335 (N_15335,N_15002,N_15165);
xor U15336 (N_15336,N_15072,N_15081);
or U15337 (N_15337,N_15104,N_15095);
nand U15338 (N_15338,N_15010,N_15173);
and U15339 (N_15339,N_15085,N_15073);
and U15340 (N_15340,N_15105,N_15185);
xnor U15341 (N_15341,N_15083,N_15069);
and U15342 (N_15342,N_15073,N_15113);
xor U15343 (N_15343,N_15001,N_15126);
and U15344 (N_15344,N_15180,N_15145);
or U15345 (N_15345,N_15107,N_15119);
nand U15346 (N_15346,N_15158,N_15014);
nand U15347 (N_15347,N_15117,N_15147);
and U15348 (N_15348,N_15141,N_15176);
nand U15349 (N_15349,N_15086,N_15188);
or U15350 (N_15350,N_15123,N_15142);
xnor U15351 (N_15351,N_15127,N_15080);
xor U15352 (N_15352,N_15185,N_15080);
nor U15353 (N_15353,N_15159,N_15092);
and U15354 (N_15354,N_15096,N_15101);
nand U15355 (N_15355,N_15097,N_15140);
or U15356 (N_15356,N_15018,N_15095);
or U15357 (N_15357,N_15165,N_15148);
nand U15358 (N_15358,N_15069,N_15011);
or U15359 (N_15359,N_15142,N_15169);
xnor U15360 (N_15360,N_15067,N_15092);
xnor U15361 (N_15361,N_15060,N_15015);
nor U15362 (N_15362,N_15151,N_15023);
and U15363 (N_15363,N_15087,N_15182);
nor U15364 (N_15364,N_15010,N_15054);
or U15365 (N_15365,N_15037,N_15117);
or U15366 (N_15366,N_15165,N_15038);
and U15367 (N_15367,N_15181,N_15152);
and U15368 (N_15368,N_15170,N_15028);
or U15369 (N_15369,N_15104,N_15088);
nor U15370 (N_15370,N_15087,N_15121);
or U15371 (N_15371,N_15024,N_15049);
xnor U15372 (N_15372,N_15091,N_15182);
nor U15373 (N_15373,N_15183,N_15074);
nand U15374 (N_15374,N_15075,N_15048);
or U15375 (N_15375,N_15059,N_15072);
nand U15376 (N_15376,N_15196,N_15109);
or U15377 (N_15377,N_15144,N_15108);
or U15378 (N_15378,N_15193,N_15029);
nand U15379 (N_15379,N_15141,N_15052);
nor U15380 (N_15380,N_15001,N_15078);
or U15381 (N_15381,N_15084,N_15072);
and U15382 (N_15382,N_15019,N_15148);
xnor U15383 (N_15383,N_15160,N_15045);
xor U15384 (N_15384,N_15124,N_15051);
xor U15385 (N_15385,N_15115,N_15015);
xor U15386 (N_15386,N_15198,N_15131);
nor U15387 (N_15387,N_15044,N_15019);
xor U15388 (N_15388,N_15023,N_15090);
and U15389 (N_15389,N_15089,N_15134);
or U15390 (N_15390,N_15094,N_15115);
and U15391 (N_15391,N_15175,N_15152);
xnor U15392 (N_15392,N_15051,N_15030);
and U15393 (N_15393,N_15087,N_15011);
and U15394 (N_15394,N_15144,N_15001);
nand U15395 (N_15395,N_15015,N_15174);
nor U15396 (N_15396,N_15152,N_15080);
and U15397 (N_15397,N_15036,N_15123);
and U15398 (N_15398,N_15110,N_15103);
nand U15399 (N_15399,N_15114,N_15035);
xnor U15400 (N_15400,N_15268,N_15265);
nor U15401 (N_15401,N_15382,N_15273);
or U15402 (N_15402,N_15290,N_15235);
nand U15403 (N_15403,N_15215,N_15259);
xnor U15404 (N_15404,N_15335,N_15375);
and U15405 (N_15405,N_15327,N_15230);
xnor U15406 (N_15406,N_15251,N_15261);
nor U15407 (N_15407,N_15318,N_15253);
or U15408 (N_15408,N_15336,N_15312);
or U15409 (N_15409,N_15281,N_15274);
nand U15410 (N_15410,N_15302,N_15288);
nor U15411 (N_15411,N_15324,N_15287);
or U15412 (N_15412,N_15246,N_15376);
and U15413 (N_15413,N_15262,N_15227);
nand U15414 (N_15414,N_15284,N_15283);
and U15415 (N_15415,N_15393,N_15206);
or U15416 (N_15416,N_15322,N_15285);
or U15417 (N_15417,N_15263,N_15264);
xnor U15418 (N_15418,N_15347,N_15388);
and U15419 (N_15419,N_15398,N_15236);
nand U15420 (N_15420,N_15221,N_15249);
or U15421 (N_15421,N_15257,N_15344);
and U15422 (N_15422,N_15389,N_15357);
nor U15423 (N_15423,N_15291,N_15316);
xnor U15424 (N_15424,N_15373,N_15297);
nand U15425 (N_15425,N_15223,N_15208);
xor U15426 (N_15426,N_15224,N_15229);
and U15427 (N_15427,N_15279,N_15201);
and U15428 (N_15428,N_15352,N_15305);
xnor U15429 (N_15429,N_15346,N_15295);
xor U15430 (N_15430,N_15314,N_15379);
xor U15431 (N_15431,N_15372,N_15212);
xor U15432 (N_15432,N_15228,N_15300);
nor U15433 (N_15433,N_15315,N_15359);
or U15434 (N_15434,N_15204,N_15304);
nand U15435 (N_15435,N_15396,N_15330);
nor U15436 (N_15436,N_15354,N_15231);
or U15437 (N_15437,N_15267,N_15394);
or U15438 (N_15438,N_15320,N_15337);
and U15439 (N_15439,N_15205,N_15341);
or U15440 (N_15440,N_15366,N_15244);
and U15441 (N_15441,N_15241,N_15343);
or U15442 (N_15442,N_15210,N_15216);
nand U15443 (N_15443,N_15385,N_15226);
nor U15444 (N_15444,N_15321,N_15238);
xor U15445 (N_15445,N_15313,N_15217);
nor U15446 (N_15446,N_15219,N_15319);
or U15447 (N_15447,N_15270,N_15367);
nor U15448 (N_15448,N_15349,N_15202);
nand U15449 (N_15449,N_15271,N_15239);
xnor U15450 (N_15450,N_15399,N_15334);
nand U15451 (N_15451,N_15277,N_15339);
nand U15452 (N_15452,N_15350,N_15325);
nor U15453 (N_15453,N_15387,N_15390);
and U15454 (N_15454,N_15381,N_15361);
and U15455 (N_15455,N_15275,N_15363);
nor U15456 (N_15456,N_15333,N_15384);
or U15457 (N_15457,N_15243,N_15329);
xnor U15458 (N_15458,N_15345,N_15266);
nand U15459 (N_15459,N_15232,N_15293);
or U15460 (N_15460,N_15342,N_15269);
and U15461 (N_15461,N_15328,N_15323);
and U15462 (N_15462,N_15258,N_15252);
xor U15463 (N_15463,N_15303,N_15391);
or U15464 (N_15464,N_15256,N_15247);
xor U15465 (N_15465,N_15272,N_15218);
and U15466 (N_15466,N_15207,N_15368);
nor U15467 (N_15467,N_15395,N_15209);
and U15468 (N_15468,N_15296,N_15356);
nor U15469 (N_15469,N_15237,N_15242);
xor U15470 (N_15470,N_15308,N_15317);
and U15471 (N_15471,N_15254,N_15289);
and U15472 (N_15472,N_15378,N_15220);
nor U15473 (N_15473,N_15260,N_15294);
xor U15474 (N_15474,N_15355,N_15338);
nand U15475 (N_15475,N_15280,N_15306);
or U15476 (N_15476,N_15301,N_15309);
nand U15477 (N_15477,N_15370,N_15200);
nor U15478 (N_15478,N_15362,N_15234);
nand U15479 (N_15479,N_15358,N_15351);
xor U15480 (N_15480,N_15326,N_15282);
xor U15481 (N_15481,N_15392,N_15240);
nand U15482 (N_15482,N_15276,N_15203);
xnor U15483 (N_15483,N_15371,N_15307);
or U15484 (N_15484,N_15311,N_15245);
nor U15485 (N_15485,N_15369,N_15250);
nor U15486 (N_15486,N_15248,N_15386);
nand U15487 (N_15487,N_15225,N_15380);
and U15488 (N_15488,N_15340,N_15299);
and U15489 (N_15489,N_15348,N_15364);
nand U15490 (N_15490,N_15397,N_15233);
and U15491 (N_15491,N_15292,N_15332);
xnor U15492 (N_15492,N_15298,N_15374);
nand U15493 (N_15493,N_15353,N_15278);
and U15494 (N_15494,N_15360,N_15331);
and U15495 (N_15495,N_15255,N_15213);
or U15496 (N_15496,N_15383,N_15377);
or U15497 (N_15497,N_15222,N_15365);
nand U15498 (N_15498,N_15310,N_15286);
and U15499 (N_15499,N_15211,N_15214);
xnor U15500 (N_15500,N_15349,N_15317);
nand U15501 (N_15501,N_15258,N_15321);
and U15502 (N_15502,N_15388,N_15297);
and U15503 (N_15503,N_15287,N_15205);
or U15504 (N_15504,N_15296,N_15226);
or U15505 (N_15505,N_15287,N_15348);
nand U15506 (N_15506,N_15301,N_15311);
and U15507 (N_15507,N_15372,N_15315);
xnor U15508 (N_15508,N_15361,N_15396);
nand U15509 (N_15509,N_15316,N_15397);
and U15510 (N_15510,N_15217,N_15322);
nor U15511 (N_15511,N_15255,N_15378);
and U15512 (N_15512,N_15233,N_15330);
nand U15513 (N_15513,N_15329,N_15267);
nand U15514 (N_15514,N_15322,N_15206);
xnor U15515 (N_15515,N_15363,N_15217);
or U15516 (N_15516,N_15278,N_15305);
and U15517 (N_15517,N_15304,N_15365);
or U15518 (N_15518,N_15357,N_15201);
and U15519 (N_15519,N_15262,N_15276);
xnor U15520 (N_15520,N_15331,N_15267);
or U15521 (N_15521,N_15227,N_15304);
xnor U15522 (N_15522,N_15387,N_15332);
or U15523 (N_15523,N_15259,N_15278);
nor U15524 (N_15524,N_15318,N_15269);
and U15525 (N_15525,N_15320,N_15392);
xnor U15526 (N_15526,N_15237,N_15327);
nor U15527 (N_15527,N_15384,N_15219);
nor U15528 (N_15528,N_15228,N_15376);
nand U15529 (N_15529,N_15256,N_15333);
nand U15530 (N_15530,N_15349,N_15354);
or U15531 (N_15531,N_15240,N_15216);
nor U15532 (N_15532,N_15298,N_15334);
nand U15533 (N_15533,N_15371,N_15321);
nor U15534 (N_15534,N_15329,N_15278);
nor U15535 (N_15535,N_15319,N_15273);
nand U15536 (N_15536,N_15399,N_15249);
nand U15537 (N_15537,N_15327,N_15221);
or U15538 (N_15538,N_15286,N_15222);
xor U15539 (N_15539,N_15304,N_15359);
and U15540 (N_15540,N_15222,N_15303);
nand U15541 (N_15541,N_15248,N_15317);
xnor U15542 (N_15542,N_15395,N_15380);
and U15543 (N_15543,N_15251,N_15244);
and U15544 (N_15544,N_15289,N_15258);
or U15545 (N_15545,N_15262,N_15351);
or U15546 (N_15546,N_15308,N_15328);
or U15547 (N_15547,N_15246,N_15249);
nor U15548 (N_15548,N_15226,N_15307);
nor U15549 (N_15549,N_15293,N_15279);
xor U15550 (N_15550,N_15236,N_15241);
nor U15551 (N_15551,N_15276,N_15258);
and U15552 (N_15552,N_15360,N_15335);
nor U15553 (N_15553,N_15277,N_15239);
nor U15554 (N_15554,N_15267,N_15366);
nor U15555 (N_15555,N_15335,N_15256);
nor U15556 (N_15556,N_15336,N_15268);
xnor U15557 (N_15557,N_15398,N_15291);
and U15558 (N_15558,N_15327,N_15296);
nand U15559 (N_15559,N_15378,N_15235);
xor U15560 (N_15560,N_15249,N_15245);
and U15561 (N_15561,N_15398,N_15333);
nand U15562 (N_15562,N_15357,N_15364);
and U15563 (N_15563,N_15245,N_15239);
nor U15564 (N_15564,N_15254,N_15394);
and U15565 (N_15565,N_15293,N_15312);
xor U15566 (N_15566,N_15376,N_15308);
xnor U15567 (N_15567,N_15219,N_15397);
and U15568 (N_15568,N_15325,N_15305);
xnor U15569 (N_15569,N_15315,N_15348);
nand U15570 (N_15570,N_15340,N_15390);
and U15571 (N_15571,N_15220,N_15219);
nor U15572 (N_15572,N_15245,N_15204);
xor U15573 (N_15573,N_15348,N_15220);
or U15574 (N_15574,N_15284,N_15353);
nor U15575 (N_15575,N_15280,N_15248);
or U15576 (N_15576,N_15279,N_15270);
or U15577 (N_15577,N_15388,N_15308);
nor U15578 (N_15578,N_15205,N_15272);
nor U15579 (N_15579,N_15276,N_15252);
nand U15580 (N_15580,N_15253,N_15384);
and U15581 (N_15581,N_15357,N_15286);
nand U15582 (N_15582,N_15396,N_15344);
xnor U15583 (N_15583,N_15272,N_15270);
xor U15584 (N_15584,N_15252,N_15230);
xnor U15585 (N_15585,N_15393,N_15311);
nand U15586 (N_15586,N_15358,N_15390);
nor U15587 (N_15587,N_15314,N_15397);
and U15588 (N_15588,N_15303,N_15272);
or U15589 (N_15589,N_15204,N_15297);
xnor U15590 (N_15590,N_15345,N_15222);
nand U15591 (N_15591,N_15391,N_15383);
or U15592 (N_15592,N_15335,N_15338);
or U15593 (N_15593,N_15329,N_15358);
nand U15594 (N_15594,N_15354,N_15303);
nand U15595 (N_15595,N_15364,N_15216);
nor U15596 (N_15596,N_15361,N_15384);
and U15597 (N_15597,N_15298,N_15265);
and U15598 (N_15598,N_15262,N_15286);
nand U15599 (N_15599,N_15213,N_15368);
or U15600 (N_15600,N_15538,N_15490);
or U15601 (N_15601,N_15426,N_15500);
or U15602 (N_15602,N_15529,N_15461);
nand U15603 (N_15603,N_15484,N_15497);
xnor U15604 (N_15604,N_15504,N_15452);
nor U15605 (N_15605,N_15425,N_15496);
nand U15606 (N_15606,N_15480,N_15405);
nor U15607 (N_15607,N_15511,N_15568);
nor U15608 (N_15608,N_15553,N_15444);
nand U15609 (N_15609,N_15411,N_15508);
and U15610 (N_15610,N_15423,N_15558);
or U15611 (N_15611,N_15531,N_15533);
and U15612 (N_15612,N_15437,N_15416);
nand U15613 (N_15613,N_15474,N_15576);
nor U15614 (N_15614,N_15495,N_15563);
and U15615 (N_15615,N_15445,N_15441);
and U15616 (N_15616,N_15435,N_15582);
xnor U15617 (N_15617,N_15488,N_15560);
or U15618 (N_15618,N_15578,N_15525);
and U15619 (N_15619,N_15583,N_15595);
or U15620 (N_15620,N_15551,N_15400);
nor U15621 (N_15621,N_15467,N_15570);
nand U15622 (N_15622,N_15465,N_15516);
nand U15623 (N_15623,N_15564,N_15569);
nand U15624 (N_15624,N_15572,N_15459);
and U15625 (N_15625,N_15527,N_15584);
xor U15626 (N_15626,N_15442,N_15440);
nor U15627 (N_15627,N_15518,N_15540);
nand U15628 (N_15628,N_15438,N_15580);
or U15629 (N_15629,N_15422,N_15526);
xnor U15630 (N_15630,N_15589,N_15514);
nand U15631 (N_15631,N_15544,N_15520);
xnor U15632 (N_15632,N_15434,N_15433);
and U15633 (N_15633,N_15519,N_15450);
nor U15634 (N_15634,N_15460,N_15468);
nand U15635 (N_15635,N_15457,N_15528);
nor U15636 (N_15636,N_15436,N_15509);
nor U15637 (N_15637,N_15403,N_15477);
and U15638 (N_15638,N_15594,N_15464);
nand U15639 (N_15639,N_15499,N_15547);
and U15640 (N_15640,N_15566,N_15507);
nor U15641 (N_15641,N_15409,N_15552);
xnor U15642 (N_15642,N_15453,N_15493);
and U15643 (N_15643,N_15410,N_15565);
xnor U15644 (N_15644,N_15574,N_15414);
nand U15645 (N_15645,N_15503,N_15542);
or U15646 (N_15646,N_15485,N_15458);
nor U15647 (N_15647,N_15590,N_15408);
and U15648 (N_15648,N_15418,N_15536);
nand U15649 (N_15649,N_15449,N_15556);
or U15650 (N_15650,N_15479,N_15428);
nand U15651 (N_15651,N_15567,N_15539);
nor U15652 (N_15652,N_15413,N_15489);
nand U15653 (N_15653,N_15475,N_15546);
nand U15654 (N_15654,N_15482,N_15406);
nand U15655 (N_15655,N_15419,N_15439);
and U15656 (N_15656,N_15454,N_15585);
nand U15657 (N_15657,N_15501,N_15549);
or U15658 (N_15658,N_15506,N_15517);
xnor U15659 (N_15659,N_15535,N_15471);
xor U15660 (N_15660,N_15463,N_15559);
and U15661 (N_15661,N_15447,N_15543);
nand U15662 (N_15662,N_15402,N_15532);
nand U15663 (N_15663,N_15462,N_15581);
or U15664 (N_15664,N_15513,N_15550);
or U15665 (N_15665,N_15466,N_15591);
nand U15666 (N_15666,N_15427,N_15541);
nor U15667 (N_15667,N_15555,N_15573);
and U15668 (N_15668,N_15492,N_15598);
xor U15669 (N_15669,N_15545,N_15421);
nor U15670 (N_15670,N_15486,N_15469);
xor U15671 (N_15671,N_15478,N_15483);
or U15672 (N_15672,N_15456,N_15523);
or U15673 (N_15673,N_15491,N_15472);
and U15674 (N_15674,N_15571,N_15432);
nand U15675 (N_15675,N_15424,N_15522);
or U15676 (N_15676,N_15502,N_15505);
xor U15677 (N_15677,N_15455,N_15407);
nand U15678 (N_15678,N_15596,N_15448);
nor U15679 (N_15679,N_15412,N_15430);
nor U15680 (N_15680,N_15443,N_15446);
or U15681 (N_15681,N_15548,N_15473);
or U15682 (N_15682,N_15404,N_15415);
and U15683 (N_15683,N_15431,N_15579);
or U15684 (N_15684,N_15524,N_15537);
xor U15685 (N_15685,N_15451,N_15593);
or U15686 (N_15686,N_15586,N_15599);
or U15687 (N_15687,N_15476,N_15494);
and U15688 (N_15688,N_15588,N_15417);
nor U15689 (N_15689,N_15562,N_15512);
or U15690 (N_15690,N_15561,N_15470);
nor U15691 (N_15691,N_15530,N_15554);
nor U15692 (N_15692,N_15515,N_15575);
xnor U15693 (N_15693,N_15481,N_15521);
and U15694 (N_15694,N_15487,N_15577);
nand U15695 (N_15695,N_15420,N_15592);
nand U15696 (N_15696,N_15597,N_15587);
nor U15697 (N_15697,N_15498,N_15510);
or U15698 (N_15698,N_15534,N_15401);
xnor U15699 (N_15699,N_15429,N_15557);
and U15700 (N_15700,N_15497,N_15409);
or U15701 (N_15701,N_15478,N_15516);
xor U15702 (N_15702,N_15477,N_15418);
nor U15703 (N_15703,N_15577,N_15451);
xnor U15704 (N_15704,N_15515,N_15535);
xor U15705 (N_15705,N_15557,N_15520);
or U15706 (N_15706,N_15471,N_15565);
nand U15707 (N_15707,N_15550,N_15414);
nand U15708 (N_15708,N_15481,N_15598);
nor U15709 (N_15709,N_15518,N_15534);
or U15710 (N_15710,N_15457,N_15594);
or U15711 (N_15711,N_15581,N_15580);
nand U15712 (N_15712,N_15502,N_15489);
xnor U15713 (N_15713,N_15431,N_15549);
and U15714 (N_15714,N_15585,N_15521);
or U15715 (N_15715,N_15569,N_15465);
nor U15716 (N_15716,N_15471,N_15537);
nor U15717 (N_15717,N_15581,N_15415);
or U15718 (N_15718,N_15522,N_15409);
xor U15719 (N_15719,N_15414,N_15427);
nand U15720 (N_15720,N_15428,N_15539);
nand U15721 (N_15721,N_15401,N_15438);
nand U15722 (N_15722,N_15591,N_15421);
and U15723 (N_15723,N_15515,N_15470);
or U15724 (N_15724,N_15524,N_15595);
nor U15725 (N_15725,N_15532,N_15460);
or U15726 (N_15726,N_15590,N_15556);
nand U15727 (N_15727,N_15462,N_15550);
nand U15728 (N_15728,N_15580,N_15562);
xnor U15729 (N_15729,N_15480,N_15526);
nor U15730 (N_15730,N_15509,N_15470);
and U15731 (N_15731,N_15599,N_15445);
nor U15732 (N_15732,N_15580,N_15515);
nand U15733 (N_15733,N_15471,N_15440);
nand U15734 (N_15734,N_15586,N_15400);
nor U15735 (N_15735,N_15573,N_15425);
xor U15736 (N_15736,N_15508,N_15538);
nor U15737 (N_15737,N_15405,N_15543);
nor U15738 (N_15738,N_15578,N_15481);
xnor U15739 (N_15739,N_15563,N_15447);
xnor U15740 (N_15740,N_15569,N_15407);
nand U15741 (N_15741,N_15534,N_15565);
or U15742 (N_15742,N_15548,N_15438);
xor U15743 (N_15743,N_15561,N_15430);
or U15744 (N_15744,N_15596,N_15547);
or U15745 (N_15745,N_15414,N_15460);
nand U15746 (N_15746,N_15560,N_15433);
xnor U15747 (N_15747,N_15511,N_15453);
nand U15748 (N_15748,N_15419,N_15595);
or U15749 (N_15749,N_15414,N_15523);
or U15750 (N_15750,N_15440,N_15447);
and U15751 (N_15751,N_15504,N_15473);
nand U15752 (N_15752,N_15552,N_15443);
or U15753 (N_15753,N_15519,N_15548);
nor U15754 (N_15754,N_15487,N_15436);
or U15755 (N_15755,N_15566,N_15533);
nor U15756 (N_15756,N_15499,N_15579);
or U15757 (N_15757,N_15576,N_15508);
or U15758 (N_15758,N_15491,N_15541);
or U15759 (N_15759,N_15566,N_15412);
nand U15760 (N_15760,N_15444,N_15492);
nor U15761 (N_15761,N_15579,N_15509);
nand U15762 (N_15762,N_15568,N_15464);
nand U15763 (N_15763,N_15484,N_15596);
and U15764 (N_15764,N_15567,N_15443);
nand U15765 (N_15765,N_15427,N_15488);
xor U15766 (N_15766,N_15424,N_15407);
and U15767 (N_15767,N_15528,N_15443);
nand U15768 (N_15768,N_15432,N_15541);
nor U15769 (N_15769,N_15481,N_15586);
nand U15770 (N_15770,N_15599,N_15526);
nand U15771 (N_15771,N_15423,N_15402);
xor U15772 (N_15772,N_15425,N_15514);
nand U15773 (N_15773,N_15499,N_15563);
nor U15774 (N_15774,N_15472,N_15559);
or U15775 (N_15775,N_15448,N_15572);
nor U15776 (N_15776,N_15550,N_15589);
xor U15777 (N_15777,N_15424,N_15528);
nor U15778 (N_15778,N_15498,N_15473);
and U15779 (N_15779,N_15565,N_15505);
xnor U15780 (N_15780,N_15445,N_15581);
and U15781 (N_15781,N_15518,N_15501);
nand U15782 (N_15782,N_15590,N_15432);
nand U15783 (N_15783,N_15537,N_15585);
and U15784 (N_15784,N_15562,N_15400);
or U15785 (N_15785,N_15418,N_15414);
nor U15786 (N_15786,N_15553,N_15464);
or U15787 (N_15787,N_15593,N_15467);
and U15788 (N_15788,N_15522,N_15597);
nand U15789 (N_15789,N_15515,N_15412);
nor U15790 (N_15790,N_15560,N_15473);
or U15791 (N_15791,N_15466,N_15563);
or U15792 (N_15792,N_15498,N_15553);
or U15793 (N_15793,N_15533,N_15485);
nand U15794 (N_15794,N_15504,N_15435);
nand U15795 (N_15795,N_15474,N_15545);
nor U15796 (N_15796,N_15441,N_15474);
nand U15797 (N_15797,N_15574,N_15483);
and U15798 (N_15798,N_15568,N_15423);
nor U15799 (N_15799,N_15549,N_15565);
nor U15800 (N_15800,N_15663,N_15768);
nand U15801 (N_15801,N_15681,N_15746);
and U15802 (N_15802,N_15719,N_15658);
nor U15803 (N_15803,N_15718,N_15694);
or U15804 (N_15804,N_15741,N_15730);
xnor U15805 (N_15805,N_15779,N_15795);
and U15806 (N_15806,N_15636,N_15641);
nand U15807 (N_15807,N_15733,N_15600);
nand U15808 (N_15808,N_15610,N_15618);
nand U15809 (N_15809,N_15764,N_15790);
or U15810 (N_15810,N_15762,N_15706);
nand U15811 (N_15811,N_15672,N_15725);
and U15812 (N_15812,N_15674,N_15700);
or U15813 (N_15813,N_15697,N_15684);
or U15814 (N_15814,N_15666,N_15716);
and U15815 (N_15815,N_15703,N_15747);
nor U15816 (N_15816,N_15606,N_15792);
and U15817 (N_15817,N_15794,N_15758);
nand U15818 (N_15818,N_15757,N_15776);
and U15819 (N_15819,N_15671,N_15749);
and U15820 (N_15820,N_15710,N_15637);
xnor U15821 (N_15821,N_15685,N_15767);
nand U15822 (N_15822,N_15754,N_15686);
nor U15823 (N_15823,N_15717,N_15755);
xor U15824 (N_15824,N_15711,N_15714);
nand U15825 (N_15825,N_15727,N_15739);
nand U15826 (N_15826,N_15683,N_15699);
nor U15827 (N_15827,N_15766,N_15744);
xnor U15828 (N_15828,N_15645,N_15750);
nor U15829 (N_15829,N_15653,N_15784);
and U15830 (N_15830,N_15709,N_15652);
nor U15831 (N_15831,N_15630,N_15634);
and U15832 (N_15832,N_15665,N_15635);
nand U15833 (N_15833,N_15676,N_15662);
and U15834 (N_15834,N_15705,N_15695);
or U15835 (N_15835,N_15715,N_15756);
xor U15836 (N_15836,N_15673,N_15793);
nor U15837 (N_15837,N_15609,N_15669);
or U15838 (N_15838,N_15798,N_15614);
xor U15839 (N_15839,N_15737,N_15632);
and U15840 (N_15840,N_15707,N_15661);
nor U15841 (N_15841,N_15704,N_15769);
or U15842 (N_15842,N_15690,N_15628);
nand U15843 (N_15843,N_15616,N_15724);
or U15844 (N_15844,N_15603,N_15778);
and U15845 (N_15845,N_15657,N_15722);
nor U15846 (N_15846,N_15738,N_15740);
xnor U15847 (N_15847,N_15745,N_15799);
nand U15848 (N_15848,N_15786,N_15698);
xor U15849 (N_15849,N_15633,N_15639);
or U15850 (N_15850,N_15638,N_15659);
nand U15851 (N_15851,N_15611,N_15734);
xor U15852 (N_15852,N_15787,N_15613);
nand U15853 (N_15853,N_15789,N_15687);
nor U15854 (N_15854,N_15677,N_15728);
and U15855 (N_15855,N_15732,N_15751);
or U15856 (N_15856,N_15693,N_15627);
or U15857 (N_15857,N_15660,N_15688);
nand U15858 (N_15858,N_15775,N_15650);
or U15859 (N_15859,N_15770,N_15691);
xnor U15860 (N_15860,N_15656,N_15651);
and U15861 (N_15861,N_15712,N_15612);
nand U15862 (N_15862,N_15605,N_15623);
xnor U15863 (N_15863,N_15743,N_15644);
and U15864 (N_15864,N_15620,N_15781);
xnor U15865 (N_15865,N_15782,N_15689);
and U15866 (N_15866,N_15742,N_15604);
or U15867 (N_15867,N_15675,N_15615);
xnor U15868 (N_15868,N_15680,N_15648);
xnor U15869 (N_15869,N_15621,N_15602);
xor U15870 (N_15870,N_15708,N_15731);
nor U15871 (N_15871,N_15780,N_15622);
nand U15872 (N_15872,N_15617,N_15679);
or U15873 (N_15873,N_15692,N_15774);
nor U15874 (N_15874,N_15682,N_15735);
or U15875 (N_15875,N_15696,N_15643);
xor U15876 (N_15876,N_15720,N_15753);
or U15877 (N_15877,N_15752,N_15601);
or U15878 (N_15878,N_15625,N_15721);
and U15879 (N_15879,N_15759,N_15629);
xor U15880 (N_15880,N_15649,N_15797);
nand U15881 (N_15881,N_15702,N_15788);
and U15882 (N_15882,N_15726,N_15667);
nand U15883 (N_15883,N_15748,N_15761);
or U15884 (N_15884,N_15646,N_15771);
nor U15885 (N_15885,N_15701,N_15642);
nor U15886 (N_15886,N_15668,N_15777);
or U15887 (N_15887,N_15713,N_15640);
and U15888 (N_15888,N_15619,N_15729);
xnor U15889 (N_15889,N_15723,N_15626);
or U15890 (N_15890,N_15760,N_15736);
xor U15891 (N_15891,N_15763,N_15783);
xnor U15892 (N_15892,N_15785,N_15647);
or U15893 (N_15893,N_15655,N_15624);
or U15894 (N_15894,N_15654,N_15772);
nand U15895 (N_15895,N_15607,N_15631);
and U15896 (N_15896,N_15773,N_15796);
xnor U15897 (N_15897,N_15791,N_15765);
and U15898 (N_15898,N_15678,N_15670);
xor U15899 (N_15899,N_15608,N_15664);
xor U15900 (N_15900,N_15614,N_15678);
xnor U15901 (N_15901,N_15665,N_15694);
nor U15902 (N_15902,N_15678,N_15694);
nor U15903 (N_15903,N_15646,N_15715);
and U15904 (N_15904,N_15785,N_15679);
nand U15905 (N_15905,N_15777,N_15702);
or U15906 (N_15906,N_15665,N_15699);
xor U15907 (N_15907,N_15791,N_15783);
xnor U15908 (N_15908,N_15712,N_15756);
xor U15909 (N_15909,N_15622,N_15703);
and U15910 (N_15910,N_15706,N_15774);
nor U15911 (N_15911,N_15727,N_15671);
nor U15912 (N_15912,N_15606,N_15765);
nor U15913 (N_15913,N_15607,N_15753);
xnor U15914 (N_15914,N_15751,N_15783);
xnor U15915 (N_15915,N_15651,N_15728);
xnor U15916 (N_15916,N_15699,N_15693);
xnor U15917 (N_15917,N_15647,N_15651);
xor U15918 (N_15918,N_15776,N_15700);
nor U15919 (N_15919,N_15685,N_15664);
or U15920 (N_15920,N_15612,N_15774);
nand U15921 (N_15921,N_15612,N_15667);
and U15922 (N_15922,N_15691,N_15750);
or U15923 (N_15923,N_15684,N_15768);
and U15924 (N_15924,N_15718,N_15684);
and U15925 (N_15925,N_15700,N_15729);
nand U15926 (N_15926,N_15747,N_15671);
xnor U15927 (N_15927,N_15768,N_15631);
or U15928 (N_15928,N_15605,N_15625);
or U15929 (N_15929,N_15656,N_15685);
and U15930 (N_15930,N_15653,N_15712);
nand U15931 (N_15931,N_15746,N_15766);
or U15932 (N_15932,N_15635,N_15769);
nor U15933 (N_15933,N_15789,N_15738);
or U15934 (N_15934,N_15609,N_15668);
nand U15935 (N_15935,N_15739,N_15632);
or U15936 (N_15936,N_15608,N_15708);
nor U15937 (N_15937,N_15766,N_15683);
and U15938 (N_15938,N_15762,N_15643);
and U15939 (N_15939,N_15626,N_15726);
nor U15940 (N_15940,N_15676,N_15611);
xor U15941 (N_15941,N_15753,N_15614);
and U15942 (N_15942,N_15762,N_15780);
nor U15943 (N_15943,N_15684,N_15714);
or U15944 (N_15944,N_15714,N_15687);
or U15945 (N_15945,N_15620,N_15704);
nor U15946 (N_15946,N_15686,N_15731);
nand U15947 (N_15947,N_15762,N_15642);
and U15948 (N_15948,N_15726,N_15659);
and U15949 (N_15949,N_15644,N_15709);
and U15950 (N_15950,N_15701,N_15706);
or U15951 (N_15951,N_15615,N_15764);
xor U15952 (N_15952,N_15691,N_15607);
nor U15953 (N_15953,N_15609,N_15652);
xnor U15954 (N_15954,N_15687,N_15796);
nor U15955 (N_15955,N_15683,N_15739);
nand U15956 (N_15956,N_15796,N_15788);
nor U15957 (N_15957,N_15696,N_15652);
nor U15958 (N_15958,N_15725,N_15681);
or U15959 (N_15959,N_15616,N_15645);
and U15960 (N_15960,N_15701,N_15724);
nor U15961 (N_15961,N_15602,N_15642);
nor U15962 (N_15962,N_15744,N_15694);
and U15963 (N_15963,N_15774,N_15733);
or U15964 (N_15964,N_15628,N_15629);
and U15965 (N_15965,N_15746,N_15754);
and U15966 (N_15966,N_15641,N_15766);
xor U15967 (N_15967,N_15641,N_15773);
or U15968 (N_15968,N_15697,N_15736);
xnor U15969 (N_15969,N_15668,N_15673);
nand U15970 (N_15970,N_15637,N_15682);
or U15971 (N_15971,N_15755,N_15685);
or U15972 (N_15972,N_15616,N_15658);
or U15973 (N_15973,N_15704,N_15787);
or U15974 (N_15974,N_15726,N_15665);
nand U15975 (N_15975,N_15620,N_15648);
and U15976 (N_15976,N_15773,N_15749);
nor U15977 (N_15977,N_15611,N_15617);
nand U15978 (N_15978,N_15608,N_15755);
xor U15979 (N_15979,N_15616,N_15687);
nand U15980 (N_15980,N_15763,N_15689);
nand U15981 (N_15981,N_15750,N_15672);
xor U15982 (N_15982,N_15738,N_15696);
or U15983 (N_15983,N_15764,N_15756);
or U15984 (N_15984,N_15742,N_15797);
xor U15985 (N_15985,N_15752,N_15724);
nor U15986 (N_15986,N_15718,N_15687);
or U15987 (N_15987,N_15618,N_15764);
or U15988 (N_15988,N_15713,N_15652);
or U15989 (N_15989,N_15772,N_15683);
or U15990 (N_15990,N_15704,N_15746);
or U15991 (N_15991,N_15601,N_15617);
and U15992 (N_15992,N_15737,N_15643);
nand U15993 (N_15993,N_15695,N_15617);
nand U15994 (N_15994,N_15753,N_15708);
or U15995 (N_15995,N_15737,N_15639);
or U15996 (N_15996,N_15625,N_15743);
xnor U15997 (N_15997,N_15698,N_15619);
and U15998 (N_15998,N_15644,N_15786);
or U15999 (N_15999,N_15676,N_15691);
or U16000 (N_16000,N_15877,N_15892);
nor U16001 (N_16001,N_15869,N_15928);
nand U16002 (N_16002,N_15978,N_15826);
and U16003 (N_16003,N_15974,N_15980);
and U16004 (N_16004,N_15906,N_15889);
nand U16005 (N_16005,N_15881,N_15846);
xor U16006 (N_16006,N_15950,N_15902);
xor U16007 (N_16007,N_15861,N_15835);
nand U16008 (N_16008,N_15952,N_15927);
nor U16009 (N_16009,N_15864,N_15991);
and U16010 (N_16010,N_15862,N_15893);
nor U16011 (N_16011,N_15988,N_15924);
or U16012 (N_16012,N_15853,N_15936);
nand U16013 (N_16013,N_15838,N_15815);
nor U16014 (N_16014,N_15866,N_15807);
or U16015 (N_16015,N_15970,N_15941);
or U16016 (N_16016,N_15883,N_15964);
and U16017 (N_16017,N_15983,N_15863);
nand U16018 (N_16018,N_15871,N_15872);
nor U16019 (N_16019,N_15804,N_15868);
or U16020 (N_16020,N_15934,N_15831);
and U16021 (N_16021,N_15987,N_15840);
or U16022 (N_16022,N_15856,N_15873);
xor U16023 (N_16023,N_15982,N_15947);
and U16024 (N_16024,N_15806,N_15848);
nand U16025 (N_16025,N_15801,N_15904);
xor U16026 (N_16026,N_15810,N_15986);
xor U16027 (N_16027,N_15901,N_15922);
nor U16028 (N_16028,N_15851,N_15805);
or U16029 (N_16029,N_15921,N_15944);
and U16030 (N_16030,N_15968,N_15899);
nand U16031 (N_16031,N_15992,N_15809);
xor U16032 (N_16032,N_15819,N_15857);
nand U16033 (N_16033,N_15898,N_15914);
nor U16034 (N_16034,N_15832,N_15984);
xor U16035 (N_16035,N_15940,N_15976);
nor U16036 (N_16036,N_15884,N_15960);
or U16037 (N_16037,N_15963,N_15993);
nor U16038 (N_16038,N_15937,N_15829);
and U16039 (N_16039,N_15814,N_15843);
or U16040 (N_16040,N_15979,N_15996);
nor U16041 (N_16041,N_15839,N_15823);
or U16042 (N_16042,N_15966,N_15985);
nor U16043 (N_16043,N_15948,N_15828);
nor U16044 (N_16044,N_15894,N_15890);
nor U16045 (N_16045,N_15958,N_15972);
nand U16046 (N_16046,N_15916,N_15926);
or U16047 (N_16047,N_15989,N_15885);
xnor U16048 (N_16048,N_15929,N_15808);
xor U16049 (N_16049,N_15850,N_15855);
and U16050 (N_16050,N_15879,N_15908);
and U16051 (N_16051,N_15931,N_15887);
and U16052 (N_16052,N_15859,N_15802);
nand U16053 (N_16053,N_15847,N_15897);
and U16054 (N_16054,N_15946,N_15896);
or U16055 (N_16055,N_15917,N_15943);
nor U16056 (N_16056,N_15822,N_15827);
xor U16057 (N_16057,N_15803,N_15800);
or U16058 (N_16058,N_15874,N_15930);
nor U16059 (N_16059,N_15938,N_15878);
nand U16060 (N_16060,N_15997,N_15969);
or U16061 (N_16061,N_15965,N_15844);
xnor U16062 (N_16062,N_15836,N_15867);
xor U16063 (N_16063,N_15860,N_15951);
nand U16064 (N_16064,N_15918,N_15820);
xor U16065 (N_16065,N_15812,N_15957);
nand U16066 (N_16066,N_15971,N_15995);
nor U16067 (N_16067,N_15923,N_15911);
and U16068 (N_16068,N_15811,N_15813);
and U16069 (N_16069,N_15870,N_15824);
nor U16070 (N_16070,N_15932,N_15949);
nand U16071 (N_16071,N_15903,N_15888);
nor U16072 (N_16072,N_15919,N_15962);
nor U16073 (N_16073,N_15880,N_15909);
xnor U16074 (N_16074,N_15912,N_15865);
and U16075 (N_16075,N_15852,N_15998);
xnor U16076 (N_16076,N_15900,N_15834);
or U16077 (N_16077,N_15913,N_15994);
and U16078 (N_16078,N_15954,N_15977);
nand U16079 (N_16079,N_15961,N_15830);
or U16080 (N_16080,N_15945,N_15915);
nor U16081 (N_16081,N_15895,N_15876);
xor U16082 (N_16082,N_15833,N_15999);
nand U16083 (N_16083,N_15925,N_15849);
or U16084 (N_16084,N_15953,N_15841);
and U16085 (N_16085,N_15967,N_15935);
or U16086 (N_16086,N_15858,N_15959);
nor U16087 (N_16087,N_15875,N_15981);
or U16088 (N_16088,N_15920,N_15933);
nand U16089 (N_16089,N_15990,N_15973);
or U16090 (N_16090,N_15956,N_15942);
nand U16091 (N_16091,N_15907,N_15845);
nor U16092 (N_16092,N_15905,N_15825);
nor U16093 (N_16093,N_15816,N_15837);
or U16094 (N_16094,N_15886,N_15882);
nand U16095 (N_16095,N_15842,N_15891);
nand U16096 (N_16096,N_15910,N_15854);
or U16097 (N_16097,N_15975,N_15939);
nor U16098 (N_16098,N_15955,N_15817);
and U16099 (N_16099,N_15818,N_15821);
and U16100 (N_16100,N_15855,N_15963);
nor U16101 (N_16101,N_15956,N_15978);
xnor U16102 (N_16102,N_15990,N_15859);
or U16103 (N_16103,N_15913,N_15990);
xor U16104 (N_16104,N_15953,N_15804);
nand U16105 (N_16105,N_15907,N_15818);
xor U16106 (N_16106,N_15925,N_15913);
nand U16107 (N_16107,N_15800,N_15992);
nand U16108 (N_16108,N_15942,N_15958);
nor U16109 (N_16109,N_15977,N_15933);
xnor U16110 (N_16110,N_15895,N_15822);
or U16111 (N_16111,N_15842,N_15846);
nand U16112 (N_16112,N_15890,N_15816);
nor U16113 (N_16113,N_15831,N_15989);
nand U16114 (N_16114,N_15953,N_15873);
and U16115 (N_16115,N_15918,N_15911);
nor U16116 (N_16116,N_15800,N_15887);
xor U16117 (N_16117,N_15840,N_15899);
xor U16118 (N_16118,N_15965,N_15932);
and U16119 (N_16119,N_15961,N_15901);
nand U16120 (N_16120,N_15894,N_15959);
nor U16121 (N_16121,N_15987,N_15982);
and U16122 (N_16122,N_15967,N_15831);
nor U16123 (N_16123,N_15930,N_15839);
and U16124 (N_16124,N_15825,N_15820);
xnor U16125 (N_16125,N_15849,N_15953);
xnor U16126 (N_16126,N_15881,N_15997);
nor U16127 (N_16127,N_15894,N_15952);
nand U16128 (N_16128,N_15881,N_15834);
xor U16129 (N_16129,N_15943,N_15807);
nand U16130 (N_16130,N_15911,N_15848);
and U16131 (N_16131,N_15810,N_15998);
xor U16132 (N_16132,N_15889,N_15908);
and U16133 (N_16133,N_15952,N_15881);
nor U16134 (N_16134,N_15975,N_15956);
and U16135 (N_16135,N_15881,N_15988);
nand U16136 (N_16136,N_15830,N_15917);
or U16137 (N_16137,N_15833,N_15899);
xnor U16138 (N_16138,N_15869,N_15891);
xnor U16139 (N_16139,N_15849,N_15996);
nand U16140 (N_16140,N_15819,N_15910);
nor U16141 (N_16141,N_15898,N_15961);
and U16142 (N_16142,N_15884,N_15996);
nand U16143 (N_16143,N_15804,N_15876);
and U16144 (N_16144,N_15979,N_15940);
xnor U16145 (N_16145,N_15865,N_15856);
and U16146 (N_16146,N_15953,N_15900);
xnor U16147 (N_16147,N_15935,N_15806);
xnor U16148 (N_16148,N_15994,N_15866);
nor U16149 (N_16149,N_15997,N_15838);
nand U16150 (N_16150,N_15941,N_15884);
or U16151 (N_16151,N_15865,N_15868);
xnor U16152 (N_16152,N_15888,N_15841);
xnor U16153 (N_16153,N_15987,N_15992);
nor U16154 (N_16154,N_15978,N_15992);
and U16155 (N_16155,N_15888,N_15943);
nor U16156 (N_16156,N_15973,N_15886);
and U16157 (N_16157,N_15935,N_15837);
or U16158 (N_16158,N_15998,N_15863);
or U16159 (N_16159,N_15906,N_15898);
nor U16160 (N_16160,N_15879,N_15860);
nand U16161 (N_16161,N_15960,N_15919);
or U16162 (N_16162,N_15856,N_15806);
nor U16163 (N_16163,N_15942,N_15891);
xnor U16164 (N_16164,N_15931,N_15922);
nor U16165 (N_16165,N_15981,N_15910);
nand U16166 (N_16166,N_15905,N_15857);
xor U16167 (N_16167,N_15917,N_15827);
xnor U16168 (N_16168,N_15969,N_15804);
nor U16169 (N_16169,N_15928,N_15953);
nor U16170 (N_16170,N_15879,N_15949);
or U16171 (N_16171,N_15824,N_15844);
xnor U16172 (N_16172,N_15916,N_15851);
nand U16173 (N_16173,N_15915,N_15989);
and U16174 (N_16174,N_15984,N_15888);
and U16175 (N_16175,N_15954,N_15922);
xor U16176 (N_16176,N_15804,N_15806);
nand U16177 (N_16177,N_15869,N_15988);
and U16178 (N_16178,N_15865,N_15811);
xor U16179 (N_16179,N_15922,N_15972);
and U16180 (N_16180,N_15899,N_15888);
nor U16181 (N_16181,N_15904,N_15824);
xor U16182 (N_16182,N_15946,N_15884);
or U16183 (N_16183,N_15883,N_15864);
nor U16184 (N_16184,N_15876,N_15913);
or U16185 (N_16185,N_15981,N_15959);
nand U16186 (N_16186,N_15917,N_15983);
or U16187 (N_16187,N_15959,N_15860);
xor U16188 (N_16188,N_15848,N_15886);
nand U16189 (N_16189,N_15855,N_15991);
and U16190 (N_16190,N_15866,N_15812);
nor U16191 (N_16191,N_15909,N_15806);
and U16192 (N_16192,N_15942,N_15824);
nand U16193 (N_16193,N_15909,N_15889);
nor U16194 (N_16194,N_15850,N_15965);
or U16195 (N_16195,N_15862,N_15963);
nand U16196 (N_16196,N_15831,N_15907);
or U16197 (N_16197,N_15896,N_15803);
xnor U16198 (N_16198,N_15830,N_15862);
nand U16199 (N_16199,N_15802,N_15965);
or U16200 (N_16200,N_16016,N_16035);
xor U16201 (N_16201,N_16188,N_16191);
xor U16202 (N_16202,N_16066,N_16128);
xor U16203 (N_16203,N_16182,N_16070);
xnor U16204 (N_16204,N_16040,N_16112);
or U16205 (N_16205,N_16093,N_16084);
xor U16206 (N_16206,N_16168,N_16021);
nand U16207 (N_16207,N_16079,N_16046);
xnor U16208 (N_16208,N_16174,N_16115);
xnor U16209 (N_16209,N_16090,N_16001);
and U16210 (N_16210,N_16183,N_16005);
or U16211 (N_16211,N_16071,N_16013);
xnor U16212 (N_16212,N_16012,N_16122);
xor U16213 (N_16213,N_16080,N_16136);
nand U16214 (N_16214,N_16078,N_16042);
xor U16215 (N_16215,N_16027,N_16109);
and U16216 (N_16216,N_16176,N_16131);
and U16217 (N_16217,N_16096,N_16055);
nor U16218 (N_16218,N_16197,N_16147);
xnor U16219 (N_16219,N_16065,N_16107);
xor U16220 (N_16220,N_16097,N_16024);
or U16221 (N_16221,N_16152,N_16148);
nand U16222 (N_16222,N_16150,N_16099);
and U16223 (N_16223,N_16199,N_16022);
xnor U16224 (N_16224,N_16015,N_16083);
xnor U16225 (N_16225,N_16155,N_16076);
or U16226 (N_16226,N_16139,N_16129);
xor U16227 (N_16227,N_16077,N_16019);
xnor U16228 (N_16228,N_16198,N_16048);
and U16229 (N_16229,N_16008,N_16039);
and U16230 (N_16230,N_16142,N_16043);
xor U16231 (N_16231,N_16069,N_16081);
xnor U16232 (N_16232,N_16140,N_16087);
and U16233 (N_16233,N_16153,N_16061);
or U16234 (N_16234,N_16116,N_16181);
and U16235 (N_16235,N_16169,N_16104);
nand U16236 (N_16236,N_16151,N_16092);
or U16237 (N_16237,N_16003,N_16089);
nor U16238 (N_16238,N_16082,N_16075);
and U16239 (N_16239,N_16117,N_16054);
xnor U16240 (N_16240,N_16184,N_16178);
xnor U16241 (N_16241,N_16127,N_16007);
nand U16242 (N_16242,N_16049,N_16185);
nor U16243 (N_16243,N_16121,N_16187);
xnor U16244 (N_16244,N_16144,N_16111);
nand U16245 (N_16245,N_16051,N_16026);
nor U16246 (N_16246,N_16073,N_16118);
and U16247 (N_16247,N_16165,N_16108);
or U16248 (N_16248,N_16011,N_16137);
and U16249 (N_16249,N_16159,N_16124);
xor U16250 (N_16250,N_16172,N_16130);
and U16251 (N_16251,N_16031,N_16037);
xnor U16252 (N_16252,N_16018,N_16004);
nand U16253 (N_16253,N_16041,N_16047);
xor U16254 (N_16254,N_16056,N_16038);
nor U16255 (N_16255,N_16158,N_16120);
nor U16256 (N_16256,N_16006,N_16103);
nor U16257 (N_16257,N_16044,N_16045);
nor U16258 (N_16258,N_16098,N_16002);
or U16259 (N_16259,N_16063,N_16141);
or U16260 (N_16260,N_16062,N_16101);
or U16261 (N_16261,N_16017,N_16189);
and U16262 (N_16262,N_16032,N_16057);
nor U16263 (N_16263,N_16023,N_16170);
or U16264 (N_16264,N_16146,N_16171);
or U16265 (N_16265,N_16190,N_16053);
and U16266 (N_16266,N_16033,N_16113);
nand U16267 (N_16267,N_16157,N_16068);
and U16268 (N_16268,N_16064,N_16134);
xor U16269 (N_16269,N_16058,N_16143);
or U16270 (N_16270,N_16163,N_16192);
xor U16271 (N_16271,N_16138,N_16166);
or U16272 (N_16272,N_16132,N_16059);
nand U16273 (N_16273,N_16102,N_16194);
and U16274 (N_16274,N_16028,N_16162);
or U16275 (N_16275,N_16010,N_16156);
or U16276 (N_16276,N_16014,N_16180);
xor U16277 (N_16277,N_16074,N_16105);
nand U16278 (N_16278,N_16034,N_16052);
or U16279 (N_16279,N_16025,N_16095);
xnor U16280 (N_16280,N_16029,N_16186);
or U16281 (N_16281,N_16125,N_16196);
xor U16282 (N_16282,N_16020,N_16114);
or U16283 (N_16283,N_16036,N_16193);
xnor U16284 (N_16284,N_16060,N_16145);
xnor U16285 (N_16285,N_16167,N_16091);
and U16286 (N_16286,N_16173,N_16135);
or U16287 (N_16287,N_16094,N_16009);
nand U16288 (N_16288,N_16000,N_16100);
or U16289 (N_16289,N_16164,N_16119);
xor U16290 (N_16290,N_16123,N_16149);
and U16291 (N_16291,N_16088,N_16067);
and U16292 (N_16292,N_16106,N_16086);
and U16293 (N_16293,N_16195,N_16177);
nor U16294 (N_16294,N_16160,N_16126);
or U16295 (N_16295,N_16072,N_16110);
xor U16296 (N_16296,N_16085,N_16179);
xor U16297 (N_16297,N_16133,N_16050);
nand U16298 (N_16298,N_16154,N_16161);
nand U16299 (N_16299,N_16030,N_16175);
xor U16300 (N_16300,N_16088,N_16092);
nand U16301 (N_16301,N_16000,N_16048);
xnor U16302 (N_16302,N_16076,N_16011);
xnor U16303 (N_16303,N_16047,N_16071);
xor U16304 (N_16304,N_16022,N_16128);
xnor U16305 (N_16305,N_16171,N_16113);
and U16306 (N_16306,N_16051,N_16136);
nand U16307 (N_16307,N_16170,N_16110);
nor U16308 (N_16308,N_16109,N_16107);
nor U16309 (N_16309,N_16129,N_16173);
and U16310 (N_16310,N_16051,N_16133);
nor U16311 (N_16311,N_16163,N_16148);
nand U16312 (N_16312,N_16174,N_16015);
xor U16313 (N_16313,N_16049,N_16072);
nor U16314 (N_16314,N_16076,N_16017);
or U16315 (N_16315,N_16107,N_16139);
nor U16316 (N_16316,N_16129,N_16149);
nor U16317 (N_16317,N_16140,N_16062);
nand U16318 (N_16318,N_16159,N_16033);
nand U16319 (N_16319,N_16037,N_16075);
or U16320 (N_16320,N_16096,N_16051);
xor U16321 (N_16321,N_16116,N_16033);
or U16322 (N_16322,N_16094,N_16077);
nor U16323 (N_16323,N_16093,N_16128);
xor U16324 (N_16324,N_16048,N_16017);
or U16325 (N_16325,N_16156,N_16105);
xnor U16326 (N_16326,N_16183,N_16154);
nand U16327 (N_16327,N_16110,N_16119);
and U16328 (N_16328,N_16050,N_16137);
and U16329 (N_16329,N_16121,N_16174);
nand U16330 (N_16330,N_16034,N_16057);
or U16331 (N_16331,N_16114,N_16177);
xor U16332 (N_16332,N_16057,N_16072);
xor U16333 (N_16333,N_16192,N_16135);
and U16334 (N_16334,N_16117,N_16176);
nand U16335 (N_16335,N_16125,N_16111);
nand U16336 (N_16336,N_16031,N_16092);
xnor U16337 (N_16337,N_16059,N_16131);
or U16338 (N_16338,N_16010,N_16092);
nand U16339 (N_16339,N_16118,N_16197);
nand U16340 (N_16340,N_16086,N_16051);
xor U16341 (N_16341,N_16132,N_16015);
nor U16342 (N_16342,N_16099,N_16163);
or U16343 (N_16343,N_16135,N_16026);
or U16344 (N_16344,N_16086,N_16058);
or U16345 (N_16345,N_16141,N_16008);
nand U16346 (N_16346,N_16186,N_16136);
and U16347 (N_16347,N_16063,N_16136);
and U16348 (N_16348,N_16051,N_16163);
or U16349 (N_16349,N_16170,N_16153);
nand U16350 (N_16350,N_16066,N_16136);
nor U16351 (N_16351,N_16011,N_16179);
nand U16352 (N_16352,N_16163,N_16012);
xor U16353 (N_16353,N_16011,N_16095);
nand U16354 (N_16354,N_16037,N_16120);
nand U16355 (N_16355,N_16149,N_16179);
or U16356 (N_16356,N_16038,N_16165);
and U16357 (N_16357,N_16022,N_16056);
nor U16358 (N_16358,N_16026,N_16090);
nor U16359 (N_16359,N_16071,N_16028);
or U16360 (N_16360,N_16131,N_16182);
and U16361 (N_16361,N_16113,N_16096);
nor U16362 (N_16362,N_16196,N_16075);
or U16363 (N_16363,N_16024,N_16125);
xor U16364 (N_16364,N_16082,N_16018);
and U16365 (N_16365,N_16139,N_16096);
or U16366 (N_16366,N_16154,N_16104);
nand U16367 (N_16367,N_16156,N_16124);
or U16368 (N_16368,N_16049,N_16066);
xor U16369 (N_16369,N_16082,N_16004);
nor U16370 (N_16370,N_16180,N_16123);
nand U16371 (N_16371,N_16194,N_16021);
nor U16372 (N_16372,N_16178,N_16082);
nor U16373 (N_16373,N_16161,N_16187);
nor U16374 (N_16374,N_16069,N_16000);
xor U16375 (N_16375,N_16057,N_16187);
and U16376 (N_16376,N_16175,N_16195);
nor U16377 (N_16377,N_16056,N_16010);
and U16378 (N_16378,N_16012,N_16099);
nand U16379 (N_16379,N_16007,N_16110);
nor U16380 (N_16380,N_16029,N_16160);
nor U16381 (N_16381,N_16162,N_16055);
and U16382 (N_16382,N_16074,N_16164);
or U16383 (N_16383,N_16018,N_16031);
nand U16384 (N_16384,N_16049,N_16002);
and U16385 (N_16385,N_16130,N_16036);
nor U16386 (N_16386,N_16188,N_16066);
nor U16387 (N_16387,N_16060,N_16067);
nor U16388 (N_16388,N_16032,N_16060);
and U16389 (N_16389,N_16039,N_16178);
nand U16390 (N_16390,N_16134,N_16194);
xor U16391 (N_16391,N_16136,N_16075);
nor U16392 (N_16392,N_16014,N_16053);
or U16393 (N_16393,N_16060,N_16134);
xnor U16394 (N_16394,N_16107,N_16160);
and U16395 (N_16395,N_16143,N_16059);
nor U16396 (N_16396,N_16101,N_16076);
nor U16397 (N_16397,N_16160,N_16188);
nor U16398 (N_16398,N_16089,N_16061);
or U16399 (N_16399,N_16166,N_16173);
nor U16400 (N_16400,N_16253,N_16205);
or U16401 (N_16401,N_16355,N_16319);
or U16402 (N_16402,N_16219,N_16228);
nand U16403 (N_16403,N_16252,N_16328);
nand U16404 (N_16404,N_16398,N_16327);
or U16405 (N_16405,N_16290,N_16275);
xnor U16406 (N_16406,N_16399,N_16394);
xor U16407 (N_16407,N_16236,N_16210);
or U16408 (N_16408,N_16229,N_16391);
and U16409 (N_16409,N_16304,N_16294);
nor U16410 (N_16410,N_16324,N_16350);
nor U16411 (N_16411,N_16222,N_16249);
or U16412 (N_16412,N_16237,N_16216);
nor U16413 (N_16413,N_16346,N_16357);
nor U16414 (N_16414,N_16367,N_16339);
nor U16415 (N_16415,N_16248,N_16352);
nor U16416 (N_16416,N_16246,N_16333);
and U16417 (N_16417,N_16227,N_16341);
nand U16418 (N_16418,N_16315,N_16306);
and U16419 (N_16419,N_16348,N_16250);
and U16420 (N_16420,N_16258,N_16272);
or U16421 (N_16421,N_16347,N_16207);
xor U16422 (N_16422,N_16279,N_16329);
or U16423 (N_16423,N_16376,N_16266);
and U16424 (N_16424,N_16254,N_16390);
nor U16425 (N_16425,N_16349,N_16225);
and U16426 (N_16426,N_16280,N_16221);
or U16427 (N_16427,N_16395,N_16365);
or U16428 (N_16428,N_16300,N_16383);
nor U16429 (N_16429,N_16309,N_16342);
nor U16430 (N_16430,N_16372,N_16358);
nand U16431 (N_16431,N_16220,N_16388);
or U16432 (N_16432,N_16316,N_16270);
nor U16433 (N_16433,N_16244,N_16359);
nand U16434 (N_16434,N_16223,N_16289);
xnor U16435 (N_16435,N_16240,N_16230);
or U16436 (N_16436,N_16344,N_16337);
nor U16437 (N_16437,N_16392,N_16307);
nand U16438 (N_16438,N_16296,N_16260);
and U16439 (N_16439,N_16369,N_16318);
and U16440 (N_16440,N_16354,N_16206);
nand U16441 (N_16441,N_16202,N_16314);
nand U16442 (N_16442,N_16233,N_16310);
nand U16443 (N_16443,N_16321,N_16269);
xnor U16444 (N_16444,N_16259,N_16345);
nand U16445 (N_16445,N_16375,N_16385);
nand U16446 (N_16446,N_16380,N_16256);
or U16447 (N_16447,N_16283,N_16261);
or U16448 (N_16448,N_16238,N_16325);
xor U16449 (N_16449,N_16317,N_16288);
nand U16450 (N_16450,N_16282,N_16331);
and U16451 (N_16451,N_16200,N_16277);
nand U16452 (N_16452,N_16281,N_16332);
nand U16453 (N_16453,N_16245,N_16215);
or U16454 (N_16454,N_16305,N_16268);
or U16455 (N_16455,N_16379,N_16242);
xor U16456 (N_16456,N_16322,N_16389);
nand U16457 (N_16457,N_16298,N_16276);
and U16458 (N_16458,N_16330,N_16263);
nor U16459 (N_16459,N_16364,N_16387);
nor U16460 (N_16460,N_16235,N_16217);
and U16461 (N_16461,N_16368,N_16373);
nor U16462 (N_16462,N_16293,N_16326);
nor U16463 (N_16463,N_16381,N_16287);
and U16464 (N_16464,N_16214,N_16213);
xnor U16465 (N_16465,N_16301,N_16299);
and U16466 (N_16466,N_16336,N_16371);
and U16467 (N_16467,N_16302,N_16320);
or U16468 (N_16468,N_16335,N_16377);
and U16469 (N_16469,N_16363,N_16267);
and U16470 (N_16470,N_16334,N_16312);
and U16471 (N_16471,N_16311,N_16286);
or U16472 (N_16472,N_16343,N_16247);
nand U16473 (N_16473,N_16351,N_16255);
nor U16474 (N_16474,N_16384,N_16204);
xnor U16475 (N_16475,N_16356,N_16386);
xnor U16476 (N_16476,N_16209,N_16360);
and U16477 (N_16477,N_16284,N_16212);
or U16478 (N_16478,N_16303,N_16285);
xnor U16479 (N_16479,N_16338,N_16361);
or U16480 (N_16480,N_16232,N_16340);
or U16481 (N_16481,N_16234,N_16274);
xnor U16482 (N_16482,N_16378,N_16224);
xor U16483 (N_16483,N_16264,N_16366);
nand U16484 (N_16484,N_16295,N_16292);
or U16485 (N_16485,N_16201,N_16226);
nor U16486 (N_16486,N_16374,N_16291);
nand U16487 (N_16487,N_16396,N_16271);
nor U16488 (N_16488,N_16218,N_16313);
and U16489 (N_16489,N_16308,N_16211);
or U16490 (N_16490,N_16239,N_16231);
nand U16491 (N_16491,N_16251,N_16278);
nand U16492 (N_16492,N_16362,N_16370);
xnor U16493 (N_16493,N_16265,N_16297);
nor U16494 (N_16494,N_16203,N_16397);
nor U16495 (N_16495,N_16257,N_16243);
nor U16496 (N_16496,N_16241,N_16393);
xor U16497 (N_16497,N_16208,N_16273);
nand U16498 (N_16498,N_16323,N_16262);
and U16499 (N_16499,N_16353,N_16382);
or U16500 (N_16500,N_16395,N_16252);
and U16501 (N_16501,N_16274,N_16310);
and U16502 (N_16502,N_16238,N_16350);
or U16503 (N_16503,N_16208,N_16366);
xor U16504 (N_16504,N_16316,N_16268);
nor U16505 (N_16505,N_16328,N_16216);
nor U16506 (N_16506,N_16218,N_16201);
and U16507 (N_16507,N_16312,N_16380);
or U16508 (N_16508,N_16399,N_16376);
nor U16509 (N_16509,N_16282,N_16225);
xnor U16510 (N_16510,N_16306,N_16211);
nand U16511 (N_16511,N_16396,N_16287);
and U16512 (N_16512,N_16229,N_16308);
nand U16513 (N_16513,N_16249,N_16311);
or U16514 (N_16514,N_16382,N_16389);
or U16515 (N_16515,N_16286,N_16248);
nand U16516 (N_16516,N_16332,N_16226);
nor U16517 (N_16517,N_16281,N_16231);
xnor U16518 (N_16518,N_16306,N_16319);
nand U16519 (N_16519,N_16280,N_16340);
and U16520 (N_16520,N_16252,N_16380);
nor U16521 (N_16521,N_16344,N_16306);
nand U16522 (N_16522,N_16215,N_16200);
and U16523 (N_16523,N_16212,N_16229);
xnor U16524 (N_16524,N_16387,N_16373);
or U16525 (N_16525,N_16288,N_16302);
xnor U16526 (N_16526,N_16346,N_16394);
or U16527 (N_16527,N_16205,N_16365);
and U16528 (N_16528,N_16316,N_16343);
and U16529 (N_16529,N_16359,N_16270);
nor U16530 (N_16530,N_16357,N_16335);
xnor U16531 (N_16531,N_16288,N_16224);
xor U16532 (N_16532,N_16352,N_16341);
xnor U16533 (N_16533,N_16350,N_16281);
nand U16534 (N_16534,N_16272,N_16283);
and U16535 (N_16535,N_16359,N_16280);
nor U16536 (N_16536,N_16325,N_16270);
nand U16537 (N_16537,N_16331,N_16353);
nand U16538 (N_16538,N_16217,N_16280);
xnor U16539 (N_16539,N_16239,N_16326);
and U16540 (N_16540,N_16209,N_16362);
nor U16541 (N_16541,N_16225,N_16394);
nor U16542 (N_16542,N_16270,N_16252);
and U16543 (N_16543,N_16354,N_16314);
xnor U16544 (N_16544,N_16209,N_16314);
nor U16545 (N_16545,N_16215,N_16213);
or U16546 (N_16546,N_16338,N_16355);
nand U16547 (N_16547,N_16331,N_16351);
nand U16548 (N_16548,N_16204,N_16334);
nand U16549 (N_16549,N_16382,N_16392);
nor U16550 (N_16550,N_16284,N_16369);
nand U16551 (N_16551,N_16345,N_16358);
and U16552 (N_16552,N_16363,N_16389);
nand U16553 (N_16553,N_16259,N_16275);
or U16554 (N_16554,N_16307,N_16342);
xor U16555 (N_16555,N_16332,N_16254);
xor U16556 (N_16556,N_16210,N_16288);
nand U16557 (N_16557,N_16217,N_16207);
nor U16558 (N_16558,N_16311,N_16389);
nand U16559 (N_16559,N_16222,N_16251);
xor U16560 (N_16560,N_16335,N_16231);
xnor U16561 (N_16561,N_16367,N_16265);
and U16562 (N_16562,N_16239,N_16307);
and U16563 (N_16563,N_16326,N_16211);
or U16564 (N_16564,N_16223,N_16207);
nand U16565 (N_16565,N_16274,N_16390);
xor U16566 (N_16566,N_16202,N_16236);
nand U16567 (N_16567,N_16236,N_16353);
xnor U16568 (N_16568,N_16356,N_16214);
nor U16569 (N_16569,N_16243,N_16385);
nor U16570 (N_16570,N_16215,N_16371);
xor U16571 (N_16571,N_16207,N_16284);
nor U16572 (N_16572,N_16288,N_16366);
and U16573 (N_16573,N_16395,N_16205);
and U16574 (N_16574,N_16281,N_16207);
or U16575 (N_16575,N_16226,N_16346);
or U16576 (N_16576,N_16223,N_16385);
xor U16577 (N_16577,N_16396,N_16377);
nor U16578 (N_16578,N_16351,N_16328);
nor U16579 (N_16579,N_16257,N_16308);
or U16580 (N_16580,N_16366,N_16222);
and U16581 (N_16581,N_16217,N_16252);
nand U16582 (N_16582,N_16331,N_16325);
nor U16583 (N_16583,N_16327,N_16235);
nor U16584 (N_16584,N_16351,N_16226);
nand U16585 (N_16585,N_16302,N_16286);
xor U16586 (N_16586,N_16343,N_16275);
nand U16587 (N_16587,N_16369,N_16289);
or U16588 (N_16588,N_16262,N_16383);
nand U16589 (N_16589,N_16379,N_16332);
nor U16590 (N_16590,N_16326,N_16209);
nand U16591 (N_16591,N_16363,N_16315);
nand U16592 (N_16592,N_16251,N_16297);
or U16593 (N_16593,N_16338,N_16339);
or U16594 (N_16594,N_16318,N_16281);
xnor U16595 (N_16595,N_16240,N_16316);
xnor U16596 (N_16596,N_16247,N_16279);
nand U16597 (N_16597,N_16335,N_16340);
nor U16598 (N_16598,N_16328,N_16204);
and U16599 (N_16599,N_16259,N_16279);
and U16600 (N_16600,N_16562,N_16422);
and U16601 (N_16601,N_16490,N_16484);
nor U16602 (N_16602,N_16525,N_16450);
nand U16603 (N_16603,N_16441,N_16594);
nand U16604 (N_16604,N_16488,N_16469);
or U16605 (N_16605,N_16546,N_16555);
or U16606 (N_16606,N_16438,N_16414);
and U16607 (N_16607,N_16457,N_16462);
xnor U16608 (N_16608,N_16405,N_16565);
nand U16609 (N_16609,N_16553,N_16548);
and U16610 (N_16610,N_16410,N_16489);
and U16611 (N_16611,N_16505,N_16478);
nor U16612 (N_16612,N_16411,N_16467);
or U16613 (N_16613,N_16509,N_16573);
or U16614 (N_16614,N_16471,N_16402);
and U16615 (N_16615,N_16420,N_16449);
xnor U16616 (N_16616,N_16453,N_16595);
nor U16617 (N_16617,N_16585,N_16495);
nand U16618 (N_16618,N_16445,N_16591);
nor U16619 (N_16619,N_16506,N_16432);
nand U16620 (N_16620,N_16530,N_16434);
xor U16621 (N_16621,N_16512,N_16482);
nor U16622 (N_16622,N_16480,N_16468);
nor U16623 (N_16623,N_16412,N_16475);
and U16624 (N_16624,N_16584,N_16401);
nand U16625 (N_16625,N_16447,N_16544);
or U16626 (N_16626,N_16421,N_16566);
xor U16627 (N_16627,N_16427,N_16425);
nor U16628 (N_16628,N_16452,N_16472);
and U16629 (N_16629,N_16523,N_16575);
or U16630 (N_16630,N_16520,N_16581);
or U16631 (N_16631,N_16424,N_16550);
nand U16632 (N_16632,N_16460,N_16400);
or U16633 (N_16633,N_16458,N_16564);
or U16634 (N_16634,N_16500,N_16580);
nor U16635 (N_16635,N_16470,N_16514);
or U16636 (N_16636,N_16487,N_16536);
or U16637 (N_16637,N_16503,N_16563);
and U16638 (N_16638,N_16527,N_16597);
xnor U16639 (N_16639,N_16493,N_16552);
nand U16640 (N_16640,N_16476,N_16504);
xor U16641 (N_16641,N_16596,N_16443);
or U16642 (N_16642,N_16403,N_16539);
and U16643 (N_16643,N_16494,N_16404);
or U16644 (N_16644,N_16570,N_16446);
and U16645 (N_16645,N_16513,N_16474);
nor U16646 (N_16646,N_16592,N_16454);
xnor U16647 (N_16647,N_16588,N_16524);
nor U16648 (N_16648,N_16444,N_16463);
nand U16649 (N_16649,N_16541,N_16549);
nor U16650 (N_16650,N_16423,N_16417);
nand U16651 (N_16651,N_16587,N_16416);
or U16652 (N_16652,N_16517,N_16574);
nor U16653 (N_16653,N_16464,N_16593);
and U16654 (N_16654,N_16531,N_16406);
nor U16655 (N_16655,N_16477,N_16521);
and U16656 (N_16656,N_16571,N_16538);
or U16657 (N_16657,N_16485,N_16577);
or U16658 (N_16658,N_16507,N_16455);
nor U16659 (N_16659,N_16543,N_16598);
nand U16660 (N_16660,N_16583,N_16437);
and U16661 (N_16661,N_16408,N_16481);
nand U16662 (N_16662,N_16599,N_16576);
xor U16663 (N_16663,N_16409,N_16483);
nand U16664 (N_16664,N_16542,N_16511);
or U16665 (N_16665,N_16526,N_16442);
nor U16666 (N_16666,N_16499,N_16569);
xor U16667 (N_16667,N_16433,N_16491);
or U16668 (N_16668,N_16529,N_16486);
nand U16669 (N_16669,N_16501,N_16498);
or U16670 (N_16670,N_16429,N_16451);
nand U16671 (N_16671,N_16461,N_16540);
or U16672 (N_16672,N_16473,N_16435);
xor U16673 (N_16673,N_16413,N_16436);
and U16674 (N_16674,N_16439,N_16519);
xnor U16675 (N_16675,N_16567,N_16558);
xnor U16676 (N_16676,N_16545,N_16533);
nor U16677 (N_16677,N_16448,N_16516);
and U16678 (N_16678,N_16518,N_16492);
nand U16679 (N_16679,N_16534,N_16415);
and U16680 (N_16680,N_16465,N_16586);
nand U16681 (N_16681,N_16561,N_16407);
xnor U16682 (N_16682,N_16496,N_16551);
and U16683 (N_16683,N_16532,N_16572);
or U16684 (N_16684,N_16426,N_16508);
xnor U16685 (N_16685,N_16537,N_16559);
or U16686 (N_16686,N_16554,N_16419);
xor U16687 (N_16687,N_16431,N_16560);
nor U16688 (N_16688,N_16547,N_16515);
xor U16689 (N_16689,N_16578,N_16428);
or U16690 (N_16690,N_16466,N_16497);
and U16691 (N_16691,N_16557,N_16459);
xor U16692 (N_16692,N_16418,N_16556);
nand U16693 (N_16693,N_16528,N_16589);
or U16694 (N_16694,N_16579,N_16582);
nor U16695 (N_16695,N_16479,N_16568);
xnor U16696 (N_16696,N_16535,N_16510);
xor U16697 (N_16697,N_16590,N_16502);
xnor U16698 (N_16698,N_16456,N_16430);
or U16699 (N_16699,N_16522,N_16440);
nor U16700 (N_16700,N_16449,N_16490);
nor U16701 (N_16701,N_16402,N_16558);
or U16702 (N_16702,N_16542,N_16597);
or U16703 (N_16703,N_16495,N_16510);
xnor U16704 (N_16704,N_16493,N_16502);
nor U16705 (N_16705,N_16573,N_16533);
nand U16706 (N_16706,N_16425,N_16497);
xnor U16707 (N_16707,N_16558,N_16570);
xnor U16708 (N_16708,N_16590,N_16554);
nand U16709 (N_16709,N_16489,N_16588);
nand U16710 (N_16710,N_16446,N_16457);
nand U16711 (N_16711,N_16422,N_16516);
nor U16712 (N_16712,N_16444,N_16509);
xor U16713 (N_16713,N_16547,N_16469);
or U16714 (N_16714,N_16413,N_16586);
xor U16715 (N_16715,N_16406,N_16566);
or U16716 (N_16716,N_16560,N_16598);
nor U16717 (N_16717,N_16561,N_16535);
and U16718 (N_16718,N_16452,N_16572);
xor U16719 (N_16719,N_16501,N_16441);
nand U16720 (N_16720,N_16548,N_16510);
nor U16721 (N_16721,N_16551,N_16413);
xnor U16722 (N_16722,N_16509,N_16524);
or U16723 (N_16723,N_16560,N_16414);
nand U16724 (N_16724,N_16551,N_16429);
and U16725 (N_16725,N_16569,N_16564);
nand U16726 (N_16726,N_16469,N_16436);
or U16727 (N_16727,N_16508,N_16475);
or U16728 (N_16728,N_16588,N_16513);
nor U16729 (N_16729,N_16417,N_16586);
xor U16730 (N_16730,N_16526,N_16543);
xnor U16731 (N_16731,N_16582,N_16540);
nor U16732 (N_16732,N_16598,N_16444);
nand U16733 (N_16733,N_16568,N_16572);
nor U16734 (N_16734,N_16551,N_16411);
xor U16735 (N_16735,N_16427,N_16441);
xnor U16736 (N_16736,N_16498,N_16580);
nand U16737 (N_16737,N_16427,N_16500);
xor U16738 (N_16738,N_16430,N_16536);
nor U16739 (N_16739,N_16502,N_16589);
and U16740 (N_16740,N_16417,N_16415);
or U16741 (N_16741,N_16533,N_16477);
nor U16742 (N_16742,N_16504,N_16561);
and U16743 (N_16743,N_16587,N_16409);
and U16744 (N_16744,N_16524,N_16447);
and U16745 (N_16745,N_16497,N_16597);
and U16746 (N_16746,N_16468,N_16441);
or U16747 (N_16747,N_16452,N_16545);
and U16748 (N_16748,N_16416,N_16564);
and U16749 (N_16749,N_16483,N_16592);
or U16750 (N_16750,N_16400,N_16582);
xnor U16751 (N_16751,N_16414,N_16597);
and U16752 (N_16752,N_16504,N_16540);
or U16753 (N_16753,N_16570,N_16571);
or U16754 (N_16754,N_16478,N_16501);
and U16755 (N_16755,N_16519,N_16569);
and U16756 (N_16756,N_16597,N_16579);
or U16757 (N_16757,N_16420,N_16592);
or U16758 (N_16758,N_16553,N_16468);
nor U16759 (N_16759,N_16575,N_16553);
nand U16760 (N_16760,N_16475,N_16515);
nand U16761 (N_16761,N_16502,N_16481);
or U16762 (N_16762,N_16541,N_16565);
or U16763 (N_16763,N_16549,N_16451);
nor U16764 (N_16764,N_16409,N_16462);
or U16765 (N_16765,N_16485,N_16509);
nor U16766 (N_16766,N_16461,N_16597);
xnor U16767 (N_16767,N_16427,N_16596);
nand U16768 (N_16768,N_16420,N_16474);
nor U16769 (N_16769,N_16524,N_16551);
nor U16770 (N_16770,N_16422,N_16508);
or U16771 (N_16771,N_16587,N_16533);
and U16772 (N_16772,N_16589,N_16407);
and U16773 (N_16773,N_16523,N_16497);
xnor U16774 (N_16774,N_16491,N_16414);
or U16775 (N_16775,N_16570,N_16479);
nor U16776 (N_16776,N_16535,N_16576);
and U16777 (N_16777,N_16472,N_16443);
xor U16778 (N_16778,N_16557,N_16408);
nand U16779 (N_16779,N_16502,N_16435);
nor U16780 (N_16780,N_16489,N_16587);
and U16781 (N_16781,N_16423,N_16559);
or U16782 (N_16782,N_16583,N_16567);
nor U16783 (N_16783,N_16567,N_16560);
and U16784 (N_16784,N_16503,N_16479);
nand U16785 (N_16785,N_16566,N_16594);
xnor U16786 (N_16786,N_16451,N_16490);
and U16787 (N_16787,N_16526,N_16469);
nand U16788 (N_16788,N_16552,N_16439);
or U16789 (N_16789,N_16443,N_16575);
or U16790 (N_16790,N_16521,N_16424);
or U16791 (N_16791,N_16508,N_16527);
or U16792 (N_16792,N_16568,N_16513);
xor U16793 (N_16793,N_16495,N_16451);
nor U16794 (N_16794,N_16574,N_16514);
nor U16795 (N_16795,N_16483,N_16449);
and U16796 (N_16796,N_16524,N_16565);
nor U16797 (N_16797,N_16428,N_16519);
and U16798 (N_16798,N_16446,N_16581);
nor U16799 (N_16799,N_16441,N_16475);
nor U16800 (N_16800,N_16621,N_16638);
xor U16801 (N_16801,N_16766,N_16759);
and U16802 (N_16802,N_16649,N_16721);
nand U16803 (N_16803,N_16637,N_16755);
nand U16804 (N_16804,N_16767,N_16798);
nand U16805 (N_16805,N_16738,N_16666);
or U16806 (N_16806,N_16752,N_16672);
xor U16807 (N_16807,N_16778,N_16760);
and U16808 (N_16808,N_16648,N_16670);
xor U16809 (N_16809,N_16761,N_16770);
or U16810 (N_16810,N_16754,N_16697);
xnor U16811 (N_16811,N_16714,N_16731);
nand U16812 (N_16812,N_16723,N_16622);
and U16813 (N_16813,N_16630,N_16611);
xor U16814 (N_16814,N_16785,N_16600);
and U16815 (N_16815,N_16702,N_16654);
or U16816 (N_16816,N_16665,N_16628);
nand U16817 (N_16817,N_16707,N_16765);
nand U16818 (N_16818,N_16633,N_16711);
nand U16819 (N_16819,N_16722,N_16613);
or U16820 (N_16820,N_16797,N_16753);
or U16821 (N_16821,N_16701,N_16604);
nand U16822 (N_16822,N_16744,N_16684);
or U16823 (N_16823,N_16642,N_16641);
xnor U16824 (N_16824,N_16605,N_16706);
nor U16825 (N_16825,N_16616,N_16615);
and U16826 (N_16826,N_16758,N_16653);
or U16827 (N_16827,N_16676,N_16788);
xnor U16828 (N_16828,N_16655,N_16712);
nor U16829 (N_16829,N_16631,N_16678);
nor U16830 (N_16830,N_16779,N_16728);
and U16831 (N_16831,N_16787,N_16750);
xnor U16832 (N_16832,N_16720,N_16727);
nand U16833 (N_16833,N_16632,N_16689);
xnor U16834 (N_16834,N_16775,N_16749);
and U16835 (N_16835,N_16606,N_16704);
nand U16836 (N_16836,N_16736,N_16743);
xnor U16837 (N_16837,N_16624,N_16674);
xnor U16838 (N_16838,N_16773,N_16667);
and U16839 (N_16839,N_16786,N_16636);
nand U16840 (N_16840,N_16740,N_16601);
and U16841 (N_16841,N_16780,N_16612);
nor U16842 (N_16842,N_16725,N_16635);
or U16843 (N_16843,N_16726,N_16662);
and U16844 (N_16844,N_16677,N_16686);
or U16845 (N_16845,N_16643,N_16629);
nor U16846 (N_16846,N_16647,N_16791);
or U16847 (N_16847,N_16732,N_16781);
nand U16848 (N_16848,N_16739,N_16793);
and U16849 (N_16849,N_16699,N_16695);
or U16850 (N_16850,N_16717,N_16730);
and U16851 (N_16851,N_16713,N_16658);
nand U16852 (N_16852,N_16768,N_16627);
and U16853 (N_16853,N_16683,N_16757);
nand U16854 (N_16854,N_16789,N_16692);
and U16855 (N_16855,N_16792,N_16774);
and U16856 (N_16856,N_16682,N_16603);
xnor U16857 (N_16857,N_16777,N_16652);
or U16858 (N_16858,N_16639,N_16708);
and U16859 (N_16859,N_16783,N_16742);
nor U16860 (N_16860,N_16657,N_16688);
and U16861 (N_16861,N_16718,N_16607);
nor U16862 (N_16862,N_16705,N_16659);
and U16863 (N_16863,N_16681,N_16764);
nand U16864 (N_16864,N_16782,N_16769);
nand U16865 (N_16865,N_16763,N_16790);
xnor U16866 (N_16866,N_16645,N_16733);
nand U16867 (N_16867,N_16719,N_16656);
or U16868 (N_16868,N_16673,N_16693);
nor U16869 (N_16869,N_16623,N_16784);
nor U16870 (N_16870,N_16651,N_16646);
nor U16871 (N_16871,N_16698,N_16703);
nor U16872 (N_16872,N_16650,N_16614);
or U16873 (N_16873,N_16669,N_16617);
and U16874 (N_16874,N_16735,N_16634);
or U16875 (N_16875,N_16729,N_16710);
nor U16876 (N_16876,N_16675,N_16687);
nor U16877 (N_16877,N_16746,N_16619);
and U16878 (N_16878,N_16794,N_16771);
and U16879 (N_16879,N_16608,N_16679);
and U16880 (N_16880,N_16747,N_16795);
or U16881 (N_16881,N_16762,N_16625);
nand U16882 (N_16882,N_16796,N_16626);
nand U16883 (N_16883,N_16724,N_16694);
nand U16884 (N_16884,N_16734,N_16716);
xnor U16885 (N_16885,N_16660,N_16644);
nand U16886 (N_16886,N_16685,N_16756);
and U16887 (N_16887,N_16663,N_16741);
nor U16888 (N_16888,N_16696,N_16709);
nor U16889 (N_16889,N_16664,N_16751);
or U16890 (N_16890,N_16748,N_16690);
nor U16891 (N_16891,N_16700,N_16715);
or U16892 (N_16892,N_16691,N_16640);
nand U16893 (N_16893,N_16737,N_16799);
nor U16894 (N_16894,N_16618,N_16609);
nor U16895 (N_16895,N_16776,N_16671);
or U16896 (N_16896,N_16610,N_16772);
xnor U16897 (N_16897,N_16620,N_16668);
or U16898 (N_16898,N_16602,N_16661);
nor U16899 (N_16899,N_16745,N_16680);
nor U16900 (N_16900,N_16637,N_16739);
xor U16901 (N_16901,N_16791,N_16626);
and U16902 (N_16902,N_16699,N_16779);
nor U16903 (N_16903,N_16647,N_16671);
xor U16904 (N_16904,N_16790,N_16723);
nand U16905 (N_16905,N_16652,N_16617);
nand U16906 (N_16906,N_16608,N_16658);
and U16907 (N_16907,N_16740,N_16788);
xnor U16908 (N_16908,N_16719,N_16612);
nor U16909 (N_16909,N_16721,N_16618);
nor U16910 (N_16910,N_16793,N_16663);
or U16911 (N_16911,N_16669,N_16786);
or U16912 (N_16912,N_16651,N_16685);
and U16913 (N_16913,N_16635,N_16744);
xnor U16914 (N_16914,N_16643,N_16746);
nor U16915 (N_16915,N_16790,N_16743);
nor U16916 (N_16916,N_16717,N_16637);
and U16917 (N_16917,N_16636,N_16614);
and U16918 (N_16918,N_16779,N_16619);
or U16919 (N_16919,N_16706,N_16689);
or U16920 (N_16920,N_16654,N_16774);
nand U16921 (N_16921,N_16751,N_16690);
nand U16922 (N_16922,N_16688,N_16721);
or U16923 (N_16923,N_16665,N_16752);
nand U16924 (N_16924,N_16621,N_16774);
nand U16925 (N_16925,N_16739,N_16745);
nand U16926 (N_16926,N_16693,N_16652);
xnor U16927 (N_16927,N_16769,N_16735);
xnor U16928 (N_16928,N_16626,N_16619);
and U16929 (N_16929,N_16755,N_16673);
or U16930 (N_16930,N_16711,N_16768);
and U16931 (N_16931,N_16681,N_16709);
nand U16932 (N_16932,N_16747,N_16708);
nor U16933 (N_16933,N_16713,N_16764);
xnor U16934 (N_16934,N_16771,N_16680);
nand U16935 (N_16935,N_16695,N_16790);
or U16936 (N_16936,N_16778,N_16697);
nor U16937 (N_16937,N_16694,N_16717);
xor U16938 (N_16938,N_16668,N_16782);
and U16939 (N_16939,N_16616,N_16649);
nor U16940 (N_16940,N_16619,N_16664);
nand U16941 (N_16941,N_16728,N_16609);
xor U16942 (N_16942,N_16737,N_16630);
nand U16943 (N_16943,N_16734,N_16681);
and U16944 (N_16944,N_16654,N_16655);
and U16945 (N_16945,N_16652,N_16779);
nor U16946 (N_16946,N_16687,N_16782);
and U16947 (N_16947,N_16794,N_16701);
nand U16948 (N_16948,N_16767,N_16632);
nor U16949 (N_16949,N_16723,N_16780);
and U16950 (N_16950,N_16664,N_16749);
and U16951 (N_16951,N_16692,N_16612);
nor U16952 (N_16952,N_16623,N_16619);
and U16953 (N_16953,N_16657,N_16749);
and U16954 (N_16954,N_16688,N_16690);
nand U16955 (N_16955,N_16691,N_16656);
and U16956 (N_16956,N_16746,N_16679);
and U16957 (N_16957,N_16794,N_16639);
nand U16958 (N_16958,N_16775,N_16606);
nor U16959 (N_16959,N_16794,N_16797);
nand U16960 (N_16960,N_16735,N_16626);
xor U16961 (N_16961,N_16668,N_16670);
xnor U16962 (N_16962,N_16703,N_16677);
nor U16963 (N_16963,N_16606,N_16767);
or U16964 (N_16964,N_16675,N_16790);
xor U16965 (N_16965,N_16647,N_16633);
or U16966 (N_16966,N_16700,N_16613);
nand U16967 (N_16967,N_16626,N_16702);
or U16968 (N_16968,N_16615,N_16651);
and U16969 (N_16969,N_16680,N_16741);
nand U16970 (N_16970,N_16630,N_16729);
or U16971 (N_16971,N_16767,N_16666);
and U16972 (N_16972,N_16736,N_16652);
or U16973 (N_16973,N_16726,N_16711);
xor U16974 (N_16974,N_16733,N_16737);
xnor U16975 (N_16975,N_16605,N_16649);
nand U16976 (N_16976,N_16727,N_16675);
xor U16977 (N_16977,N_16617,N_16719);
or U16978 (N_16978,N_16797,N_16754);
nor U16979 (N_16979,N_16665,N_16794);
nor U16980 (N_16980,N_16668,N_16719);
and U16981 (N_16981,N_16720,N_16705);
or U16982 (N_16982,N_16744,N_16633);
nor U16983 (N_16983,N_16688,N_16741);
xor U16984 (N_16984,N_16673,N_16664);
nand U16985 (N_16985,N_16709,N_16608);
or U16986 (N_16986,N_16611,N_16786);
nor U16987 (N_16987,N_16662,N_16748);
and U16988 (N_16988,N_16676,N_16637);
or U16989 (N_16989,N_16772,N_16602);
and U16990 (N_16990,N_16776,N_16719);
nor U16991 (N_16991,N_16729,N_16673);
nor U16992 (N_16992,N_16686,N_16710);
or U16993 (N_16993,N_16636,N_16731);
or U16994 (N_16994,N_16772,N_16754);
and U16995 (N_16995,N_16751,N_16676);
nor U16996 (N_16996,N_16602,N_16625);
or U16997 (N_16997,N_16784,N_16700);
nor U16998 (N_16998,N_16703,N_16622);
nand U16999 (N_16999,N_16718,N_16730);
nor U17000 (N_17000,N_16970,N_16875);
nor U17001 (N_17001,N_16831,N_16833);
and U17002 (N_17002,N_16899,N_16843);
nand U17003 (N_17003,N_16826,N_16835);
nand U17004 (N_17004,N_16964,N_16952);
nand U17005 (N_17005,N_16902,N_16834);
nor U17006 (N_17006,N_16914,N_16983);
nand U17007 (N_17007,N_16838,N_16823);
xnor U17008 (N_17008,N_16987,N_16904);
and U17009 (N_17009,N_16820,N_16865);
xnor U17010 (N_17010,N_16830,N_16901);
nand U17011 (N_17011,N_16848,N_16859);
nor U17012 (N_17012,N_16888,N_16981);
or U17013 (N_17013,N_16857,N_16920);
nor U17014 (N_17014,N_16965,N_16984);
nand U17015 (N_17015,N_16938,N_16819);
nand U17016 (N_17016,N_16947,N_16809);
and U17017 (N_17017,N_16844,N_16876);
or U17018 (N_17018,N_16894,N_16956);
or U17019 (N_17019,N_16852,N_16821);
nand U17020 (N_17020,N_16842,N_16851);
and U17021 (N_17021,N_16884,N_16994);
or U17022 (N_17022,N_16971,N_16801);
xnor U17023 (N_17023,N_16871,N_16988);
or U17024 (N_17024,N_16997,N_16817);
or U17025 (N_17025,N_16944,N_16934);
xor U17026 (N_17026,N_16870,N_16898);
and U17027 (N_17027,N_16960,N_16961);
and U17028 (N_17028,N_16913,N_16966);
nor U17029 (N_17029,N_16845,N_16918);
xor U17030 (N_17030,N_16977,N_16837);
xnor U17031 (N_17031,N_16919,N_16878);
nor U17032 (N_17032,N_16939,N_16963);
nor U17033 (N_17033,N_16962,N_16974);
nand U17034 (N_17034,N_16999,N_16883);
or U17035 (N_17035,N_16957,N_16800);
nand U17036 (N_17036,N_16840,N_16812);
nor U17037 (N_17037,N_16975,N_16815);
xnor U17038 (N_17038,N_16985,N_16923);
nand U17039 (N_17039,N_16846,N_16850);
and U17040 (N_17040,N_16839,N_16805);
nand U17041 (N_17041,N_16824,N_16935);
or U17042 (N_17042,N_16916,N_16982);
xor U17043 (N_17043,N_16877,N_16802);
xnor U17044 (N_17044,N_16853,N_16980);
or U17045 (N_17045,N_16861,N_16867);
nor U17046 (N_17046,N_16841,N_16893);
xor U17047 (N_17047,N_16995,N_16807);
or U17048 (N_17048,N_16932,N_16973);
nor U17049 (N_17049,N_16906,N_16949);
xnor U17050 (N_17050,N_16872,N_16889);
nand U17051 (N_17051,N_16813,N_16921);
xnor U17052 (N_17052,N_16863,N_16940);
nand U17053 (N_17053,N_16900,N_16911);
or U17054 (N_17054,N_16903,N_16879);
and U17055 (N_17055,N_16836,N_16972);
nand U17056 (N_17056,N_16990,N_16860);
nand U17057 (N_17057,N_16953,N_16895);
nor U17058 (N_17058,N_16862,N_16897);
and U17059 (N_17059,N_16978,N_16856);
xnor U17060 (N_17060,N_16885,N_16882);
and U17061 (N_17061,N_16874,N_16854);
nand U17062 (N_17062,N_16814,N_16991);
and U17063 (N_17063,N_16890,N_16955);
or U17064 (N_17064,N_16909,N_16958);
xnor U17065 (N_17065,N_16891,N_16954);
nand U17066 (N_17066,N_16989,N_16931);
or U17067 (N_17067,N_16950,N_16942);
xnor U17068 (N_17068,N_16868,N_16855);
and U17069 (N_17069,N_16908,N_16986);
nand U17070 (N_17070,N_16976,N_16930);
nor U17071 (N_17071,N_16943,N_16925);
and U17072 (N_17072,N_16892,N_16946);
nand U17073 (N_17073,N_16948,N_16886);
or U17074 (N_17074,N_16912,N_16945);
xnor U17075 (N_17075,N_16880,N_16896);
nor U17076 (N_17076,N_16869,N_16905);
or U17077 (N_17077,N_16832,N_16887);
and U17078 (N_17078,N_16910,N_16858);
nor U17079 (N_17079,N_16998,N_16825);
or U17080 (N_17080,N_16967,N_16849);
nand U17081 (N_17081,N_16808,N_16827);
xnor U17082 (N_17082,N_16941,N_16866);
nand U17083 (N_17083,N_16873,N_16822);
or U17084 (N_17084,N_16933,N_16951);
nand U17085 (N_17085,N_16993,N_16936);
or U17086 (N_17086,N_16806,N_16927);
and U17087 (N_17087,N_16937,N_16959);
nor U17088 (N_17088,N_16864,N_16992);
xor U17089 (N_17089,N_16969,N_16818);
and U17090 (N_17090,N_16829,N_16924);
or U17091 (N_17091,N_16922,N_16804);
nor U17092 (N_17092,N_16926,N_16928);
or U17093 (N_17093,N_16810,N_16996);
or U17094 (N_17094,N_16881,N_16917);
or U17095 (N_17095,N_16847,N_16907);
nor U17096 (N_17096,N_16915,N_16828);
nor U17097 (N_17097,N_16816,N_16803);
nor U17098 (N_17098,N_16979,N_16968);
or U17099 (N_17099,N_16811,N_16929);
nor U17100 (N_17100,N_16953,N_16833);
nand U17101 (N_17101,N_16909,N_16841);
nor U17102 (N_17102,N_16816,N_16818);
xnor U17103 (N_17103,N_16814,N_16938);
nor U17104 (N_17104,N_16962,N_16938);
and U17105 (N_17105,N_16900,N_16950);
xnor U17106 (N_17106,N_16872,N_16958);
and U17107 (N_17107,N_16984,N_16944);
xor U17108 (N_17108,N_16888,N_16997);
nor U17109 (N_17109,N_16863,N_16861);
and U17110 (N_17110,N_16848,N_16864);
or U17111 (N_17111,N_16923,N_16832);
nand U17112 (N_17112,N_16960,N_16840);
xnor U17113 (N_17113,N_16931,N_16832);
and U17114 (N_17114,N_16818,N_16900);
and U17115 (N_17115,N_16973,N_16850);
xnor U17116 (N_17116,N_16881,N_16820);
nor U17117 (N_17117,N_16805,N_16853);
and U17118 (N_17118,N_16939,N_16834);
xnor U17119 (N_17119,N_16920,N_16975);
or U17120 (N_17120,N_16996,N_16871);
nor U17121 (N_17121,N_16808,N_16851);
nor U17122 (N_17122,N_16859,N_16875);
or U17123 (N_17123,N_16899,N_16903);
nand U17124 (N_17124,N_16816,N_16842);
nor U17125 (N_17125,N_16935,N_16918);
xor U17126 (N_17126,N_16805,N_16852);
and U17127 (N_17127,N_16936,N_16825);
nand U17128 (N_17128,N_16887,N_16868);
nand U17129 (N_17129,N_16835,N_16906);
or U17130 (N_17130,N_16944,N_16901);
nand U17131 (N_17131,N_16839,N_16981);
and U17132 (N_17132,N_16813,N_16935);
nor U17133 (N_17133,N_16948,N_16850);
or U17134 (N_17134,N_16978,N_16886);
xor U17135 (N_17135,N_16844,N_16826);
and U17136 (N_17136,N_16981,N_16935);
and U17137 (N_17137,N_16986,N_16845);
xnor U17138 (N_17138,N_16962,N_16822);
nand U17139 (N_17139,N_16835,N_16932);
or U17140 (N_17140,N_16928,N_16848);
nand U17141 (N_17141,N_16926,N_16853);
or U17142 (N_17142,N_16803,N_16927);
nor U17143 (N_17143,N_16919,N_16974);
and U17144 (N_17144,N_16952,N_16993);
xor U17145 (N_17145,N_16980,N_16983);
nand U17146 (N_17146,N_16924,N_16995);
nor U17147 (N_17147,N_16815,N_16881);
xnor U17148 (N_17148,N_16843,N_16981);
xnor U17149 (N_17149,N_16951,N_16983);
nor U17150 (N_17150,N_16918,N_16943);
or U17151 (N_17151,N_16837,N_16827);
or U17152 (N_17152,N_16906,N_16927);
and U17153 (N_17153,N_16926,N_16962);
or U17154 (N_17154,N_16897,N_16969);
nor U17155 (N_17155,N_16961,N_16903);
nand U17156 (N_17156,N_16837,N_16872);
nor U17157 (N_17157,N_16926,N_16831);
and U17158 (N_17158,N_16929,N_16965);
xor U17159 (N_17159,N_16883,N_16871);
nand U17160 (N_17160,N_16920,N_16846);
xnor U17161 (N_17161,N_16971,N_16827);
nand U17162 (N_17162,N_16999,N_16870);
nand U17163 (N_17163,N_16837,N_16904);
nand U17164 (N_17164,N_16874,N_16809);
or U17165 (N_17165,N_16942,N_16889);
nor U17166 (N_17166,N_16964,N_16826);
nor U17167 (N_17167,N_16892,N_16872);
or U17168 (N_17168,N_16904,N_16917);
nor U17169 (N_17169,N_16979,N_16962);
nor U17170 (N_17170,N_16904,N_16951);
nand U17171 (N_17171,N_16893,N_16852);
nand U17172 (N_17172,N_16958,N_16876);
nor U17173 (N_17173,N_16865,N_16926);
xor U17174 (N_17174,N_16949,N_16899);
and U17175 (N_17175,N_16915,N_16988);
nor U17176 (N_17176,N_16990,N_16867);
and U17177 (N_17177,N_16827,N_16864);
or U17178 (N_17178,N_16898,N_16834);
nand U17179 (N_17179,N_16972,N_16868);
nand U17180 (N_17180,N_16849,N_16900);
nor U17181 (N_17181,N_16948,N_16963);
and U17182 (N_17182,N_16851,N_16829);
nor U17183 (N_17183,N_16989,N_16990);
and U17184 (N_17184,N_16921,N_16981);
or U17185 (N_17185,N_16838,N_16834);
nor U17186 (N_17186,N_16856,N_16857);
and U17187 (N_17187,N_16987,N_16853);
and U17188 (N_17188,N_16866,N_16959);
nand U17189 (N_17189,N_16986,N_16993);
or U17190 (N_17190,N_16887,N_16930);
or U17191 (N_17191,N_16858,N_16870);
or U17192 (N_17192,N_16943,N_16965);
or U17193 (N_17193,N_16857,N_16837);
or U17194 (N_17194,N_16861,N_16999);
nor U17195 (N_17195,N_16963,N_16982);
and U17196 (N_17196,N_16843,N_16907);
or U17197 (N_17197,N_16977,N_16920);
and U17198 (N_17198,N_16821,N_16908);
xnor U17199 (N_17199,N_16974,N_16816);
or U17200 (N_17200,N_17043,N_17113);
nand U17201 (N_17201,N_17088,N_17186);
or U17202 (N_17202,N_17000,N_17152);
xor U17203 (N_17203,N_17101,N_17036);
and U17204 (N_17204,N_17137,N_17158);
xor U17205 (N_17205,N_17071,N_17098);
and U17206 (N_17206,N_17061,N_17155);
or U17207 (N_17207,N_17078,N_17162);
xnor U17208 (N_17208,N_17080,N_17034);
xnor U17209 (N_17209,N_17131,N_17119);
nor U17210 (N_17210,N_17191,N_17044);
nor U17211 (N_17211,N_17074,N_17125);
nor U17212 (N_17212,N_17116,N_17025);
nor U17213 (N_17213,N_17070,N_17083);
or U17214 (N_17214,N_17195,N_17163);
and U17215 (N_17215,N_17005,N_17149);
xnor U17216 (N_17216,N_17094,N_17003);
nor U17217 (N_17217,N_17157,N_17147);
nand U17218 (N_17218,N_17124,N_17004);
and U17219 (N_17219,N_17050,N_17148);
and U17220 (N_17220,N_17140,N_17171);
nand U17221 (N_17221,N_17129,N_17198);
and U17222 (N_17222,N_17045,N_17072);
nor U17223 (N_17223,N_17188,N_17082);
nand U17224 (N_17224,N_17159,N_17011);
or U17225 (N_17225,N_17096,N_17118);
and U17226 (N_17226,N_17182,N_17102);
or U17227 (N_17227,N_17023,N_17064);
xnor U17228 (N_17228,N_17151,N_17130);
nand U17229 (N_17229,N_17189,N_17062);
or U17230 (N_17230,N_17041,N_17087);
nand U17231 (N_17231,N_17017,N_17046);
xor U17232 (N_17232,N_17079,N_17166);
nand U17233 (N_17233,N_17056,N_17136);
xor U17234 (N_17234,N_17144,N_17154);
and U17235 (N_17235,N_17066,N_17052);
or U17236 (N_17236,N_17057,N_17018);
nand U17237 (N_17237,N_17197,N_17109);
nor U17238 (N_17238,N_17123,N_17134);
and U17239 (N_17239,N_17037,N_17160);
nor U17240 (N_17240,N_17103,N_17180);
or U17241 (N_17241,N_17038,N_17165);
or U17242 (N_17242,N_17002,N_17183);
nor U17243 (N_17243,N_17133,N_17107);
and U17244 (N_17244,N_17019,N_17048);
and U17245 (N_17245,N_17010,N_17001);
nand U17246 (N_17246,N_17039,N_17091);
and U17247 (N_17247,N_17168,N_17111);
and U17248 (N_17248,N_17065,N_17053);
xnor U17249 (N_17249,N_17084,N_17106);
and U17250 (N_17250,N_17179,N_17100);
or U17251 (N_17251,N_17187,N_17150);
xor U17252 (N_17252,N_17112,N_17090);
or U17253 (N_17253,N_17051,N_17086);
and U17254 (N_17254,N_17095,N_17135);
xor U17255 (N_17255,N_17073,N_17059);
xor U17256 (N_17256,N_17169,N_17022);
and U17257 (N_17257,N_17027,N_17193);
nor U17258 (N_17258,N_17175,N_17035);
or U17259 (N_17259,N_17015,N_17199);
nand U17260 (N_17260,N_17049,N_17146);
xor U17261 (N_17261,N_17194,N_17190);
xnor U17262 (N_17262,N_17054,N_17172);
and U17263 (N_17263,N_17026,N_17012);
nand U17264 (N_17264,N_17164,N_17170);
and U17265 (N_17265,N_17081,N_17121);
xor U17266 (N_17266,N_17063,N_17060);
and U17267 (N_17267,N_17132,N_17007);
nor U17268 (N_17268,N_17127,N_17181);
and U17269 (N_17269,N_17141,N_17128);
nand U17270 (N_17270,N_17058,N_17099);
or U17271 (N_17271,N_17120,N_17177);
or U17272 (N_17272,N_17196,N_17126);
xnor U17273 (N_17273,N_17085,N_17092);
nor U17274 (N_17274,N_17031,N_17047);
xnor U17275 (N_17275,N_17068,N_17076);
nand U17276 (N_17276,N_17016,N_17069);
nor U17277 (N_17277,N_17161,N_17077);
nor U17278 (N_17278,N_17021,N_17032);
nand U17279 (N_17279,N_17153,N_17139);
xor U17280 (N_17280,N_17145,N_17156);
or U17281 (N_17281,N_17040,N_17115);
xor U17282 (N_17282,N_17093,N_17110);
nand U17283 (N_17283,N_17097,N_17067);
or U17284 (N_17284,N_17089,N_17138);
nand U17285 (N_17285,N_17075,N_17013);
nand U17286 (N_17286,N_17185,N_17114);
nor U17287 (N_17287,N_17009,N_17108);
nor U17288 (N_17288,N_17105,N_17143);
nor U17289 (N_17289,N_17028,N_17042);
xor U17290 (N_17290,N_17030,N_17006);
xnor U17291 (N_17291,N_17033,N_17008);
nor U17292 (N_17292,N_17020,N_17173);
or U17293 (N_17293,N_17104,N_17142);
xnor U17294 (N_17294,N_17055,N_17117);
or U17295 (N_17295,N_17029,N_17178);
or U17296 (N_17296,N_17184,N_17024);
or U17297 (N_17297,N_17192,N_17014);
nand U17298 (N_17298,N_17167,N_17174);
or U17299 (N_17299,N_17122,N_17176);
and U17300 (N_17300,N_17136,N_17118);
or U17301 (N_17301,N_17029,N_17193);
nor U17302 (N_17302,N_17054,N_17104);
and U17303 (N_17303,N_17117,N_17142);
nor U17304 (N_17304,N_17043,N_17008);
xor U17305 (N_17305,N_17075,N_17156);
or U17306 (N_17306,N_17016,N_17122);
or U17307 (N_17307,N_17160,N_17178);
or U17308 (N_17308,N_17003,N_17095);
nor U17309 (N_17309,N_17100,N_17182);
nor U17310 (N_17310,N_17021,N_17030);
nor U17311 (N_17311,N_17184,N_17032);
nor U17312 (N_17312,N_17047,N_17072);
nand U17313 (N_17313,N_17196,N_17173);
nor U17314 (N_17314,N_17095,N_17142);
nand U17315 (N_17315,N_17082,N_17155);
nor U17316 (N_17316,N_17096,N_17123);
and U17317 (N_17317,N_17185,N_17118);
nor U17318 (N_17318,N_17051,N_17113);
and U17319 (N_17319,N_17118,N_17179);
nor U17320 (N_17320,N_17104,N_17199);
and U17321 (N_17321,N_17157,N_17143);
nor U17322 (N_17322,N_17156,N_17183);
nand U17323 (N_17323,N_17096,N_17053);
nor U17324 (N_17324,N_17024,N_17050);
nor U17325 (N_17325,N_17004,N_17088);
and U17326 (N_17326,N_17130,N_17038);
or U17327 (N_17327,N_17117,N_17060);
or U17328 (N_17328,N_17021,N_17133);
and U17329 (N_17329,N_17173,N_17084);
nand U17330 (N_17330,N_17136,N_17109);
nand U17331 (N_17331,N_17075,N_17143);
or U17332 (N_17332,N_17138,N_17182);
or U17333 (N_17333,N_17001,N_17021);
or U17334 (N_17334,N_17095,N_17046);
xnor U17335 (N_17335,N_17078,N_17199);
nor U17336 (N_17336,N_17150,N_17065);
or U17337 (N_17337,N_17186,N_17061);
xor U17338 (N_17338,N_17159,N_17071);
nand U17339 (N_17339,N_17169,N_17093);
xnor U17340 (N_17340,N_17135,N_17130);
nand U17341 (N_17341,N_17089,N_17035);
nor U17342 (N_17342,N_17098,N_17182);
nand U17343 (N_17343,N_17105,N_17179);
or U17344 (N_17344,N_17194,N_17114);
nand U17345 (N_17345,N_17123,N_17111);
nor U17346 (N_17346,N_17186,N_17022);
xnor U17347 (N_17347,N_17170,N_17163);
and U17348 (N_17348,N_17073,N_17089);
and U17349 (N_17349,N_17048,N_17107);
nor U17350 (N_17350,N_17056,N_17169);
or U17351 (N_17351,N_17199,N_17032);
nand U17352 (N_17352,N_17185,N_17188);
xor U17353 (N_17353,N_17072,N_17151);
xor U17354 (N_17354,N_17173,N_17170);
or U17355 (N_17355,N_17056,N_17110);
nor U17356 (N_17356,N_17175,N_17099);
or U17357 (N_17357,N_17177,N_17143);
nor U17358 (N_17358,N_17115,N_17100);
or U17359 (N_17359,N_17016,N_17084);
nand U17360 (N_17360,N_17064,N_17159);
or U17361 (N_17361,N_17087,N_17039);
nand U17362 (N_17362,N_17135,N_17101);
nor U17363 (N_17363,N_17042,N_17089);
nor U17364 (N_17364,N_17106,N_17139);
xor U17365 (N_17365,N_17185,N_17067);
nand U17366 (N_17366,N_17073,N_17054);
nor U17367 (N_17367,N_17039,N_17097);
nor U17368 (N_17368,N_17082,N_17169);
or U17369 (N_17369,N_17074,N_17031);
nor U17370 (N_17370,N_17145,N_17042);
nor U17371 (N_17371,N_17001,N_17006);
xor U17372 (N_17372,N_17071,N_17117);
or U17373 (N_17373,N_17094,N_17112);
nor U17374 (N_17374,N_17048,N_17051);
xnor U17375 (N_17375,N_17055,N_17050);
nand U17376 (N_17376,N_17062,N_17049);
nor U17377 (N_17377,N_17019,N_17044);
xor U17378 (N_17378,N_17022,N_17007);
xor U17379 (N_17379,N_17027,N_17146);
or U17380 (N_17380,N_17002,N_17095);
or U17381 (N_17381,N_17198,N_17181);
or U17382 (N_17382,N_17018,N_17056);
nor U17383 (N_17383,N_17049,N_17149);
and U17384 (N_17384,N_17028,N_17129);
or U17385 (N_17385,N_17140,N_17161);
and U17386 (N_17386,N_17156,N_17070);
and U17387 (N_17387,N_17005,N_17063);
and U17388 (N_17388,N_17092,N_17104);
nor U17389 (N_17389,N_17191,N_17092);
or U17390 (N_17390,N_17060,N_17064);
nor U17391 (N_17391,N_17143,N_17059);
or U17392 (N_17392,N_17095,N_17035);
nand U17393 (N_17393,N_17130,N_17129);
xnor U17394 (N_17394,N_17001,N_17051);
xnor U17395 (N_17395,N_17043,N_17100);
xnor U17396 (N_17396,N_17091,N_17045);
nor U17397 (N_17397,N_17075,N_17054);
or U17398 (N_17398,N_17114,N_17181);
and U17399 (N_17399,N_17130,N_17118);
and U17400 (N_17400,N_17385,N_17371);
nor U17401 (N_17401,N_17213,N_17286);
and U17402 (N_17402,N_17285,N_17264);
or U17403 (N_17403,N_17250,N_17211);
nor U17404 (N_17404,N_17360,N_17335);
nor U17405 (N_17405,N_17353,N_17221);
and U17406 (N_17406,N_17332,N_17295);
nand U17407 (N_17407,N_17322,N_17337);
nor U17408 (N_17408,N_17325,N_17282);
nor U17409 (N_17409,N_17293,N_17363);
nand U17410 (N_17410,N_17336,N_17222);
or U17411 (N_17411,N_17330,N_17212);
nor U17412 (N_17412,N_17254,N_17237);
nand U17413 (N_17413,N_17260,N_17326);
nand U17414 (N_17414,N_17201,N_17305);
nor U17415 (N_17415,N_17344,N_17262);
xor U17416 (N_17416,N_17359,N_17376);
nand U17417 (N_17417,N_17239,N_17299);
nand U17418 (N_17418,N_17381,N_17346);
or U17419 (N_17419,N_17288,N_17358);
nor U17420 (N_17420,N_17297,N_17296);
xnor U17421 (N_17421,N_17320,N_17272);
and U17422 (N_17422,N_17374,N_17321);
nand U17423 (N_17423,N_17343,N_17224);
xnor U17424 (N_17424,N_17246,N_17352);
or U17425 (N_17425,N_17279,N_17303);
nor U17426 (N_17426,N_17277,N_17365);
nor U17427 (N_17427,N_17313,N_17227);
nor U17428 (N_17428,N_17284,N_17348);
nor U17429 (N_17429,N_17240,N_17347);
xnor U17430 (N_17430,N_17364,N_17256);
nor U17431 (N_17431,N_17281,N_17234);
or U17432 (N_17432,N_17208,N_17215);
nor U17433 (N_17433,N_17290,N_17306);
xor U17434 (N_17434,N_17219,N_17382);
xor U17435 (N_17435,N_17311,N_17386);
and U17436 (N_17436,N_17251,N_17380);
and U17437 (N_17437,N_17309,N_17276);
nand U17438 (N_17438,N_17389,N_17245);
nor U17439 (N_17439,N_17228,N_17257);
xor U17440 (N_17440,N_17274,N_17216);
nor U17441 (N_17441,N_17368,N_17298);
nand U17442 (N_17442,N_17247,N_17369);
nor U17443 (N_17443,N_17283,N_17340);
nor U17444 (N_17444,N_17204,N_17307);
or U17445 (N_17445,N_17200,N_17384);
nand U17446 (N_17446,N_17339,N_17361);
or U17447 (N_17447,N_17235,N_17367);
or U17448 (N_17448,N_17202,N_17327);
or U17449 (N_17449,N_17362,N_17357);
or U17450 (N_17450,N_17230,N_17248);
and U17451 (N_17451,N_17207,N_17271);
and U17452 (N_17452,N_17214,N_17300);
nor U17453 (N_17453,N_17310,N_17378);
or U17454 (N_17454,N_17255,N_17258);
nand U17455 (N_17455,N_17315,N_17377);
or U17456 (N_17456,N_17291,N_17263);
nand U17457 (N_17457,N_17398,N_17223);
nor U17458 (N_17458,N_17232,N_17231);
xnor U17459 (N_17459,N_17354,N_17203);
xnor U17460 (N_17460,N_17217,N_17289);
nor U17461 (N_17461,N_17233,N_17273);
and U17462 (N_17462,N_17243,N_17292);
nor U17463 (N_17463,N_17308,N_17395);
xor U17464 (N_17464,N_17314,N_17205);
xnor U17465 (N_17465,N_17275,N_17316);
nor U17466 (N_17466,N_17345,N_17270);
nand U17467 (N_17467,N_17370,N_17261);
xor U17468 (N_17468,N_17375,N_17323);
xnor U17469 (N_17469,N_17333,N_17393);
xnor U17470 (N_17470,N_17220,N_17253);
nor U17471 (N_17471,N_17366,N_17387);
and U17472 (N_17472,N_17209,N_17287);
nand U17473 (N_17473,N_17338,N_17210);
nand U17474 (N_17474,N_17280,N_17350);
and U17475 (N_17475,N_17331,N_17356);
and U17476 (N_17476,N_17278,N_17266);
nor U17477 (N_17477,N_17392,N_17324);
nand U17478 (N_17478,N_17206,N_17229);
nand U17479 (N_17479,N_17341,N_17294);
or U17480 (N_17480,N_17267,N_17312);
xor U17481 (N_17481,N_17319,N_17342);
nor U17482 (N_17482,N_17351,N_17249);
xor U17483 (N_17483,N_17259,N_17349);
nor U17484 (N_17484,N_17372,N_17328);
or U17485 (N_17485,N_17268,N_17383);
nor U17486 (N_17486,N_17396,N_17218);
and U17487 (N_17487,N_17317,N_17242);
or U17488 (N_17488,N_17391,N_17236);
nand U17489 (N_17489,N_17373,N_17399);
xnor U17490 (N_17490,N_17265,N_17379);
or U17491 (N_17491,N_17241,N_17394);
or U17492 (N_17492,N_17318,N_17355);
nor U17493 (N_17493,N_17301,N_17226);
xor U17494 (N_17494,N_17244,N_17252);
nand U17495 (N_17495,N_17269,N_17388);
and U17496 (N_17496,N_17334,N_17390);
xor U17497 (N_17497,N_17304,N_17225);
xor U17498 (N_17498,N_17238,N_17302);
nor U17499 (N_17499,N_17329,N_17397);
and U17500 (N_17500,N_17202,N_17282);
nor U17501 (N_17501,N_17300,N_17256);
xnor U17502 (N_17502,N_17254,N_17284);
or U17503 (N_17503,N_17216,N_17397);
nor U17504 (N_17504,N_17284,N_17278);
nand U17505 (N_17505,N_17386,N_17394);
nor U17506 (N_17506,N_17360,N_17292);
xor U17507 (N_17507,N_17318,N_17278);
nand U17508 (N_17508,N_17299,N_17358);
and U17509 (N_17509,N_17296,N_17234);
or U17510 (N_17510,N_17259,N_17373);
or U17511 (N_17511,N_17203,N_17313);
nand U17512 (N_17512,N_17326,N_17338);
xnor U17513 (N_17513,N_17250,N_17319);
xor U17514 (N_17514,N_17335,N_17229);
xnor U17515 (N_17515,N_17383,N_17223);
xor U17516 (N_17516,N_17296,N_17336);
nand U17517 (N_17517,N_17295,N_17330);
or U17518 (N_17518,N_17317,N_17324);
nand U17519 (N_17519,N_17326,N_17270);
xor U17520 (N_17520,N_17360,N_17240);
nand U17521 (N_17521,N_17369,N_17306);
nand U17522 (N_17522,N_17266,N_17300);
nor U17523 (N_17523,N_17247,N_17353);
and U17524 (N_17524,N_17359,N_17354);
or U17525 (N_17525,N_17358,N_17337);
nand U17526 (N_17526,N_17362,N_17324);
or U17527 (N_17527,N_17375,N_17339);
or U17528 (N_17528,N_17236,N_17307);
nor U17529 (N_17529,N_17328,N_17256);
nor U17530 (N_17530,N_17283,N_17307);
nor U17531 (N_17531,N_17338,N_17308);
nor U17532 (N_17532,N_17242,N_17209);
nor U17533 (N_17533,N_17380,N_17295);
nor U17534 (N_17534,N_17346,N_17297);
nor U17535 (N_17535,N_17317,N_17375);
xnor U17536 (N_17536,N_17234,N_17384);
xor U17537 (N_17537,N_17212,N_17340);
xnor U17538 (N_17538,N_17372,N_17316);
nor U17539 (N_17539,N_17273,N_17297);
and U17540 (N_17540,N_17210,N_17396);
nand U17541 (N_17541,N_17377,N_17273);
and U17542 (N_17542,N_17200,N_17386);
nand U17543 (N_17543,N_17228,N_17331);
and U17544 (N_17544,N_17203,N_17340);
nor U17545 (N_17545,N_17201,N_17351);
and U17546 (N_17546,N_17359,N_17300);
or U17547 (N_17547,N_17320,N_17225);
nor U17548 (N_17548,N_17220,N_17379);
or U17549 (N_17549,N_17287,N_17230);
nor U17550 (N_17550,N_17257,N_17309);
or U17551 (N_17551,N_17251,N_17375);
xnor U17552 (N_17552,N_17275,N_17359);
and U17553 (N_17553,N_17254,N_17326);
nor U17554 (N_17554,N_17335,N_17302);
xor U17555 (N_17555,N_17200,N_17212);
or U17556 (N_17556,N_17314,N_17250);
or U17557 (N_17557,N_17286,N_17316);
nand U17558 (N_17558,N_17381,N_17214);
or U17559 (N_17559,N_17371,N_17246);
xnor U17560 (N_17560,N_17216,N_17321);
xor U17561 (N_17561,N_17359,N_17331);
and U17562 (N_17562,N_17235,N_17290);
and U17563 (N_17563,N_17255,N_17219);
or U17564 (N_17564,N_17322,N_17315);
xor U17565 (N_17565,N_17215,N_17298);
nand U17566 (N_17566,N_17248,N_17352);
and U17567 (N_17567,N_17238,N_17213);
nor U17568 (N_17568,N_17249,N_17377);
and U17569 (N_17569,N_17255,N_17322);
or U17570 (N_17570,N_17335,N_17213);
xor U17571 (N_17571,N_17320,N_17299);
nor U17572 (N_17572,N_17211,N_17263);
xnor U17573 (N_17573,N_17221,N_17345);
xor U17574 (N_17574,N_17292,N_17247);
xor U17575 (N_17575,N_17253,N_17227);
and U17576 (N_17576,N_17337,N_17295);
xor U17577 (N_17577,N_17304,N_17296);
nand U17578 (N_17578,N_17370,N_17251);
or U17579 (N_17579,N_17325,N_17226);
or U17580 (N_17580,N_17249,N_17352);
xnor U17581 (N_17581,N_17393,N_17319);
and U17582 (N_17582,N_17392,N_17343);
xnor U17583 (N_17583,N_17358,N_17295);
nand U17584 (N_17584,N_17364,N_17260);
nor U17585 (N_17585,N_17384,N_17319);
and U17586 (N_17586,N_17260,N_17250);
or U17587 (N_17587,N_17381,N_17212);
nor U17588 (N_17588,N_17334,N_17200);
nor U17589 (N_17589,N_17268,N_17314);
xnor U17590 (N_17590,N_17202,N_17284);
and U17591 (N_17591,N_17332,N_17230);
and U17592 (N_17592,N_17315,N_17229);
and U17593 (N_17593,N_17310,N_17398);
or U17594 (N_17594,N_17379,N_17307);
or U17595 (N_17595,N_17286,N_17276);
nor U17596 (N_17596,N_17365,N_17370);
nand U17597 (N_17597,N_17234,N_17290);
xor U17598 (N_17598,N_17348,N_17249);
xor U17599 (N_17599,N_17220,N_17308);
and U17600 (N_17600,N_17415,N_17411);
or U17601 (N_17601,N_17571,N_17522);
xnor U17602 (N_17602,N_17479,N_17421);
xnor U17603 (N_17603,N_17436,N_17561);
xnor U17604 (N_17604,N_17449,N_17408);
and U17605 (N_17605,N_17562,N_17472);
xor U17606 (N_17606,N_17448,N_17577);
and U17607 (N_17607,N_17566,N_17503);
or U17608 (N_17608,N_17550,N_17535);
nand U17609 (N_17609,N_17445,N_17513);
or U17610 (N_17610,N_17546,N_17490);
nor U17611 (N_17611,N_17426,N_17560);
or U17612 (N_17612,N_17502,N_17567);
and U17613 (N_17613,N_17570,N_17494);
xor U17614 (N_17614,N_17478,N_17425);
nor U17615 (N_17615,N_17439,N_17515);
xnor U17616 (N_17616,N_17552,N_17540);
xor U17617 (N_17617,N_17446,N_17589);
or U17618 (N_17618,N_17419,N_17451);
xnor U17619 (N_17619,N_17491,N_17469);
xor U17620 (N_17620,N_17576,N_17558);
nand U17621 (N_17621,N_17548,N_17453);
xnor U17622 (N_17622,N_17466,N_17519);
nand U17623 (N_17623,N_17420,N_17534);
and U17624 (N_17624,N_17578,N_17594);
and U17625 (N_17625,N_17433,N_17518);
or U17626 (N_17626,N_17512,N_17542);
nand U17627 (N_17627,N_17477,N_17444);
and U17628 (N_17628,N_17409,N_17596);
and U17629 (N_17629,N_17559,N_17508);
nand U17630 (N_17630,N_17405,N_17592);
or U17631 (N_17631,N_17460,N_17468);
and U17632 (N_17632,N_17401,N_17556);
or U17633 (N_17633,N_17450,N_17431);
and U17634 (N_17634,N_17483,N_17489);
and U17635 (N_17635,N_17467,N_17569);
and U17636 (N_17636,N_17572,N_17418);
nor U17637 (N_17637,N_17551,N_17510);
or U17638 (N_17638,N_17543,N_17525);
or U17639 (N_17639,N_17523,N_17485);
and U17640 (N_17640,N_17574,N_17435);
or U17641 (N_17641,N_17443,N_17511);
xnor U17642 (N_17642,N_17538,N_17595);
and U17643 (N_17643,N_17529,N_17524);
or U17644 (N_17644,N_17553,N_17459);
and U17645 (N_17645,N_17456,N_17410);
nor U17646 (N_17646,N_17586,N_17424);
nor U17647 (N_17647,N_17416,N_17434);
nand U17648 (N_17648,N_17520,N_17585);
nor U17649 (N_17649,N_17563,N_17430);
xor U17650 (N_17650,N_17590,N_17579);
xnor U17651 (N_17651,N_17598,N_17476);
or U17652 (N_17652,N_17500,N_17593);
nor U17653 (N_17653,N_17537,N_17464);
nor U17654 (N_17654,N_17432,N_17454);
and U17655 (N_17655,N_17487,N_17549);
xor U17656 (N_17656,N_17514,N_17533);
nand U17657 (N_17657,N_17547,N_17565);
and U17658 (N_17658,N_17564,N_17582);
xor U17659 (N_17659,N_17455,N_17597);
nor U17660 (N_17660,N_17499,N_17437);
xor U17661 (N_17661,N_17539,N_17497);
and U17662 (N_17662,N_17527,N_17555);
nand U17663 (N_17663,N_17473,N_17428);
and U17664 (N_17664,N_17544,N_17587);
nand U17665 (N_17665,N_17442,N_17471);
and U17666 (N_17666,N_17495,N_17554);
or U17667 (N_17667,N_17498,N_17532);
or U17668 (N_17668,N_17493,N_17438);
or U17669 (N_17669,N_17412,N_17517);
or U17670 (N_17670,N_17584,N_17458);
xor U17671 (N_17671,N_17530,N_17557);
nor U17672 (N_17672,N_17407,N_17504);
xor U17673 (N_17673,N_17440,N_17526);
nor U17674 (N_17674,N_17447,N_17536);
xor U17675 (N_17675,N_17481,N_17452);
nand U17676 (N_17676,N_17531,N_17583);
or U17677 (N_17677,N_17492,N_17465);
nand U17678 (N_17678,N_17591,N_17400);
nand U17679 (N_17679,N_17528,N_17462);
or U17680 (N_17680,N_17470,N_17506);
and U17681 (N_17681,N_17402,N_17541);
and U17682 (N_17682,N_17423,N_17457);
or U17683 (N_17683,N_17588,N_17568);
and U17684 (N_17684,N_17509,N_17427);
and U17685 (N_17685,N_17496,N_17545);
nor U17686 (N_17686,N_17575,N_17429);
xor U17687 (N_17687,N_17488,N_17573);
and U17688 (N_17688,N_17413,N_17581);
or U17689 (N_17689,N_17475,N_17484);
xnor U17690 (N_17690,N_17599,N_17404);
nor U17691 (N_17691,N_17414,N_17417);
nor U17692 (N_17692,N_17474,N_17486);
and U17693 (N_17693,N_17403,N_17461);
or U17694 (N_17694,N_17521,N_17422);
nor U17695 (N_17695,N_17507,N_17501);
and U17696 (N_17696,N_17406,N_17516);
xnor U17697 (N_17697,N_17441,N_17480);
nor U17698 (N_17698,N_17580,N_17463);
or U17699 (N_17699,N_17505,N_17482);
or U17700 (N_17700,N_17480,N_17434);
or U17701 (N_17701,N_17445,N_17544);
and U17702 (N_17702,N_17413,N_17473);
or U17703 (N_17703,N_17411,N_17544);
nand U17704 (N_17704,N_17557,N_17549);
or U17705 (N_17705,N_17507,N_17497);
or U17706 (N_17706,N_17525,N_17545);
nor U17707 (N_17707,N_17422,N_17523);
and U17708 (N_17708,N_17517,N_17409);
nand U17709 (N_17709,N_17488,N_17457);
nor U17710 (N_17710,N_17555,N_17584);
or U17711 (N_17711,N_17587,N_17427);
and U17712 (N_17712,N_17574,N_17508);
xor U17713 (N_17713,N_17597,N_17430);
and U17714 (N_17714,N_17427,N_17554);
and U17715 (N_17715,N_17518,N_17429);
and U17716 (N_17716,N_17526,N_17523);
or U17717 (N_17717,N_17548,N_17566);
or U17718 (N_17718,N_17470,N_17521);
or U17719 (N_17719,N_17495,N_17500);
and U17720 (N_17720,N_17414,N_17507);
or U17721 (N_17721,N_17433,N_17456);
nand U17722 (N_17722,N_17571,N_17589);
or U17723 (N_17723,N_17476,N_17409);
xnor U17724 (N_17724,N_17455,N_17539);
and U17725 (N_17725,N_17515,N_17403);
nor U17726 (N_17726,N_17592,N_17424);
nor U17727 (N_17727,N_17505,N_17592);
xnor U17728 (N_17728,N_17577,N_17507);
nand U17729 (N_17729,N_17518,N_17503);
nor U17730 (N_17730,N_17550,N_17544);
and U17731 (N_17731,N_17422,N_17441);
or U17732 (N_17732,N_17568,N_17401);
and U17733 (N_17733,N_17417,N_17509);
and U17734 (N_17734,N_17558,N_17565);
nand U17735 (N_17735,N_17585,N_17566);
or U17736 (N_17736,N_17561,N_17463);
nor U17737 (N_17737,N_17585,N_17572);
or U17738 (N_17738,N_17541,N_17424);
xor U17739 (N_17739,N_17530,N_17559);
nand U17740 (N_17740,N_17493,N_17437);
nand U17741 (N_17741,N_17478,N_17428);
xor U17742 (N_17742,N_17408,N_17573);
xnor U17743 (N_17743,N_17404,N_17562);
or U17744 (N_17744,N_17571,N_17501);
nand U17745 (N_17745,N_17523,N_17443);
nand U17746 (N_17746,N_17407,N_17408);
xor U17747 (N_17747,N_17422,N_17453);
nor U17748 (N_17748,N_17506,N_17416);
and U17749 (N_17749,N_17443,N_17538);
xor U17750 (N_17750,N_17542,N_17555);
nand U17751 (N_17751,N_17533,N_17499);
nand U17752 (N_17752,N_17570,N_17437);
xor U17753 (N_17753,N_17443,N_17501);
nor U17754 (N_17754,N_17556,N_17578);
xor U17755 (N_17755,N_17495,N_17570);
or U17756 (N_17756,N_17540,N_17500);
xor U17757 (N_17757,N_17457,N_17427);
nor U17758 (N_17758,N_17573,N_17475);
xnor U17759 (N_17759,N_17468,N_17471);
nand U17760 (N_17760,N_17546,N_17565);
and U17761 (N_17761,N_17442,N_17523);
and U17762 (N_17762,N_17486,N_17569);
nor U17763 (N_17763,N_17534,N_17481);
or U17764 (N_17764,N_17563,N_17496);
or U17765 (N_17765,N_17408,N_17474);
or U17766 (N_17766,N_17424,N_17419);
xnor U17767 (N_17767,N_17540,N_17454);
nand U17768 (N_17768,N_17578,N_17480);
or U17769 (N_17769,N_17589,N_17481);
xor U17770 (N_17770,N_17408,N_17443);
and U17771 (N_17771,N_17550,N_17449);
xor U17772 (N_17772,N_17412,N_17580);
nor U17773 (N_17773,N_17565,N_17400);
xnor U17774 (N_17774,N_17464,N_17414);
or U17775 (N_17775,N_17490,N_17515);
and U17776 (N_17776,N_17402,N_17469);
nand U17777 (N_17777,N_17584,N_17401);
nand U17778 (N_17778,N_17579,N_17425);
xor U17779 (N_17779,N_17406,N_17571);
nor U17780 (N_17780,N_17483,N_17545);
and U17781 (N_17781,N_17485,N_17579);
nor U17782 (N_17782,N_17544,N_17554);
and U17783 (N_17783,N_17460,N_17457);
nand U17784 (N_17784,N_17461,N_17512);
and U17785 (N_17785,N_17496,N_17477);
and U17786 (N_17786,N_17414,N_17420);
nand U17787 (N_17787,N_17506,N_17497);
nor U17788 (N_17788,N_17417,N_17449);
xnor U17789 (N_17789,N_17494,N_17428);
nor U17790 (N_17790,N_17429,N_17524);
nand U17791 (N_17791,N_17431,N_17453);
nand U17792 (N_17792,N_17549,N_17449);
xor U17793 (N_17793,N_17590,N_17526);
or U17794 (N_17794,N_17496,N_17485);
nand U17795 (N_17795,N_17510,N_17403);
and U17796 (N_17796,N_17516,N_17506);
or U17797 (N_17797,N_17425,N_17555);
and U17798 (N_17798,N_17490,N_17554);
or U17799 (N_17799,N_17494,N_17584);
xor U17800 (N_17800,N_17706,N_17761);
xor U17801 (N_17801,N_17793,N_17626);
and U17802 (N_17802,N_17772,N_17658);
and U17803 (N_17803,N_17775,N_17600);
nand U17804 (N_17804,N_17750,N_17625);
nor U17805 (N_17805,N_17640,N_17756);
xor U17806 (N_17806,N_17684,N_17673);
xor U17807 (N_17807,N_17783,N_17691);
nor U17808 (N_17808,N_17650,N_17721);
nand U17809 (N_17809,N_17611,N_17733);
and U17810 (N_17810,N_17649,N_17664);
nand U17811 (N_17811,N_17605,N_17732);
nor U17812 (N_17812,N_17681,N_17672);
and U17813 (N_17813,N_17665,N_17715);
nand U17814 (N_17814,N_17641,N_17702);
or U17815 (N_17815,N_17633,N_17764);
or U17816 (N_17816,N_17720,N_17671);
nor U17817 (N_17817,N_17698,N_17708);
xnor U17818 (N_17818,N_17668,N_17789);
or U17819 (N_17819,N_17763,N_17609);
nor U17820 (N_17820,N_17712,N_17745);
or U17821 (N_17821,N_17622,N_17771);
or U17822 (N_17822,N_17663,N_17760);
and U17823 (N_17823,N_17647,N_17709);
or U17824 (N_17824,N_17770,N_17774);
xor U17825 (N_17825,N_17791,N_17604);
nor U17826 (N_17826,N_17645,N_17768);
nand U17827 (N_17827,N_17784,N_17694);
nand U17828 (N_17828,N_17619,N_17703);
nand U17829 (N_17829,N_17637,N_17635);
nand U17830 (N_17830,N_17723,N_17689);
xor U17831 (N_17831,N_17602,N_17747);
nor U17832 (N_17832,N_17728,N_17677);
xnor U17833 (N_17833,N_17614,N_17741);
or U17834 (N_17834,N_17790,N_17678);
or U17835 (N_17835,N_17690,N_17621);
xnor U17836 (N_17836,N_17717,N_17666);
xor U17837 (N_17837,N_17607,N_17610);
xnor U17838 (N_17838,N_17624,N_17786);
and U17839 (N_17839,N_17754,N_17767);
nand U17840 (N_17840,N_17603,N_17683);
and U17841 (N_17841,N_17631,N_17659);
xnor U17842 (N_17842,N_17776,N_17796);
or U17843 (N_17843,N_17697,N_17655);
and U17844 (N_17844,N_17730,N_17696);
or U17845 (N_17845,N_17656,N_17799);
nor U17846 (N_17846,N_17727,N_17795);
and U17847 (N_17847,N_17700,N_17615);
and U17848 (N_17848,N_17661,N_17669);
xor U17849 (N_17849,N_17731,N_17612);
or U17850 (N_17850,N_17687,N_17724);
or U17851 (N_17851,N_17618,N_17748);
xor U17852 (N_17852,N_17705,N_17743);
xor U17853 (N_17853,N_17788,N_17758);
nand U17854 (N_17854,N_17787,N_17766);
xor U17855 (N_17855,N_17657,N_17682);
xor U17856 (N_17856,N_17695,N_17667);
nand U17857 (N_17857,N_17777,N_17755);
xor U17858 (N_17858,N_17674,N_17740);
xor U17859 (N_17859,N_17749,N_17710);
nand U17860 (N_17860,N_17797,N_17693);
or U17861 (N_17861,N_17601,N_17620);
nor U17862 (N_17862,N_17744,N_17735);
or U17863 (N_17863,N_17630,N_17634);
or U17864 (N_17864,N_17746,N_17642);
or U17865 (N_17865,N_17648,N_17685);
nand U17866 (N_17866,N_17686,N_17707);
or U17867 (N_17867,N_17716,N_17736);
and U17868 (N_17868,N_17782,N_17636);
xor U17869 (N_17869,N_17785,N_17757);
or U17870 (N_17870,N_17765,N_17739);
nor U17871 (N_17871,N_17711,N_17751);
nor U17872 (N_17872,N_17778,N_17753);
or U17873 (N_17873,N_17646,N_17644);
nand U17874 (N_17874,N_17653,N_17652);
nand U17875 (N_17875,N_17651,N_17680);
and U17876 (N_17876,N_17606,N_17726);
and U17877 (N_17877,N_17779,N_17679);
nand U17878 (N_17878,N_17628,N_17660);
or U17879 (N_17879,N_17792,N_17608);
or U17880 (N_17880,N_17725,N_17617);
nand U17881 (N_17881,N_17654,N_17773);
nor U17882 (N_17882,N_17734,N_17638);
xnor U17883 (N_17883,N_17639,N_17675);
nor U17884 (N_17884,N_17704,N_17718);
or U17885 (N_17885,N_17762,N_17780);
nor U17886 (N_17886,N_17688,N_17713);
nor U17887 (N_17887,N_17623,N_17662);
nor U17888 (N_17888,N_17719,N_17714);
and U17889 (N_17889,N_17627,N_17742);
and U17890 (N_17890,N_17692,N_17643);
nor U17891 (N_17891,N_17613,N_17699);
xnor U17892 (N_17892,N_17759,N_17722);
or U17893 (N_17893,N_17632,N_17729);
nand U17894 (N_17894,N_17752,N_17629);
and U17895 (N_17895,N_17794,N_17670);
xnor U17896 (N_17896,N_17769,N_17676);
nor U17897 (N_17897,N_17616,N_17798);
xnor U17898 (N_17898,N_17738,N_17781);
nor U17899 (N_17899,N_17701,N_17737);
xnor U17900 (N_17900,N_17753,N_17643);
nand U17901 (N_17901,N_17619,N_17786);
xor U17902 (N_17902,N_17669,N_17732);
or U17903 (N_17903,N_17792,N_17770);
and U17904 (N_17904,N_17741,N_17727);
nand U17905 (N_17905,N_17601,N_17769);
or U17906 (N_17906,N_17620,N_17775);
or U17907 (N_17907,N_17722,N_17773);
nand U17908 (N_17908,N_17695,N_17778);
xnor U17909 (N_17909,N_17769,N_17664);
nor U17910 (N_17910,N_17769,N_17705);
or U17911 (N_17911,N_17791,N_17645);
and U17912 (N_17912,N_17739,N_17655);
nand U17913 (N_17913,N_17785,N_17608);
xnor U17914 (N_17914,N_17770,N_17722);
or U17915 (N_17915,N_17659,N_17707);
or U17916 (N_17916,N_17775,N_17790);
or U17917 (N_17917,N_17789,N_17782);
and U17918 (N_17918,N_17713,N_17641);
xor U17919 (N_17919,N_17685,N_17783);
or U17920 (N_17920,N_17641,N_17721);
or U17921 (N_17921,N_17608,N_17684);
xnor U17922 (N_17922,N_17600,N_17679);
or U17923 (N_17923,N_17662,N_17656);
xnor U17924 (N_17924,N_17710,N_17692);
nor U17925 (N_17925,N_17676,N_17740);
or U17926 (N_17926,N_17624,N_17796);
xor U17927 (N_17927,N_17605,N_17795);
and U17928 (N_17928,N_17779,N_17677);
or U17929 (N_17929,N_17653,N_17681);
nor U17930 (N_17930,N_17783,N_17713);
nor U17931 (N_17931,N_17641,N_17714);
nor U17932 (N_17932,N_17760,N_17706);
nor U17933 (N_17933,N_17658,N_17719);
nor U17934 (N_17934,N_17745,N_17620);
nor U17935 (N_17935,N_17784,N_17695);
xnor U17936 (N_17936,N_17659,N_17783);
xor U17937 (N_17937,N_17728,N_17725);
nand U17938 (N_17938,N_17783,N_17695);
xnor U17939 (N_17939,N_17641,N_17656);
or U17940 (N_17940,N_17647,N_17724);
and U17941 (N_17941,N_17725,N_17609);
and U17942 (N_17942,N_17686,N_17615);
and U17943 (N_17943,N_17770,N_17642);
nand U17944 (N_17944,N_17785,N_17697);
nand U17945 (N_17945,N_17636,N_17674);
and U17946 (N_17946,N_17664,N_17740);
and U17947 (N_17947,N_17680,N_17684);
or U17948 (N_17948,N_17695,N_17698);
or U17949 (N_17949,N_17692,N_17707);
nor U17950 (N_17950,N_17731,N_17687);
xor U17951 (N_17951,N_17778,N_17686);
and U17952 (N_17952,N_17736,N_17620);
or U17953 (N_17953,N_17735,N_17636);
or U17954 (N_17954,N_17778,N_17644);
and U17955 (N_17955,N_17631,N_17798);
and U17956 (N_17956,N_17799,N_17755);
or U17957 (N_17957,N_17649,N_17686);
or U17958 (N_17958,N_17621,N_17785);
nand U17959 (N_17959,N_17770,N_17641);
or U17960 (N_17960,N_17672,N_17659);
or U17961 (N_17961,N_17750,N_17614);
and U17962 (N_17962,N_17668,N_17677);
and U17963 (N_17963,N_17740,N_17739);
and U17964 (N_17964,N_17678,N_17653);
or U17965 (N_17965,N_17607,N_17602);
or U17966 (N_17966,N_17660,N_17746);
or U17967 (N_17967,N_17627,N_17661);
xnor U17968 (N_17968,N_17693,N_17636);
nor U17969 (N_17969,N_17772,N_17777);
nor U17970 (N_17970,N_17695,N_17681);
and U17971 (N_17971,N_17628,N_17751);
xnor U17972 (N_17972,N_17716,N_17601);
nand U17973 (N_17973,N_17764,N_17678);
and U17974 (N_17974,N_17764,N_17762);
or U17975 (N_17975,N_17698,N_17789);
or U17976 (N_17976,N_17669,N_17610);
nand U17977 (N_17977,N_17621,N_17680);
and U17978 (N_17978,N_17797,N_17603);
xor U17979 (N_17979,N_17767,N_17638);
or U17980 (N_17980,N_17770,N_17779);
nand U17981 (N_17981,N_17772,N_17750);
xor U17982 (N_17982,N_17781,N_17756);
nand U17983 (N_17983,N_17657,N_17609);
nor U17984 (N_17984,N_17762,N_17646);
and U17985 (N_17985,N_17630,N_17619);
nand U17986 (N_17986,N_17620,N_17694);
nor U17987 (N_17987,N_17626,N_17714);
xor U17988 (N_17988,N_17631,N_17743);
or U17989 (N_17989,N_17747,N_17635);
xnor U17990 (N_17990,N_17758,N_17787);
and U17991 (N_17991,N_17678,N_17613);
or U17992 (N_17992,N_17661,N_17743);
or U17993 (N_17993,N_17610,N_17718);
xnor U17994 (N_17994,N_17780,N_17745);
and U17995 (N_17995,N_17787,N_17625);
or U17996 (N_17996,N_17772,N_17789);
nor U17997 (N_17997,N_17625,N_17649);
nand U17998 (N_17998,N_17746,N_17636);
or U17999 (N_17999,N_17728,N_17789);
nand U18000 (N_18000,N_17805,N_17960);
and U18001 (N_18001,N_17800,N_17840);
nor U18002 (N_18002,N_17809,N_17869);
or U18003 (N_18003,N_17835,N_17989);
xor U18004 (N_18004,N_17900,N_17877);
xor U18005 (N_18005,N_17820,N_17910);
or U18006 (N_18006,N_17932,N_17911);
nand U18007 (N_18007,N_17996,N_17917);
nand U18008 (N_18008,N_17857,N_17811);
nand U18009 (N_18009,N_17824,N_17944);
or U18010 (N_18010,N_17838,N_17897);
and U18011 (N_18011,N_17872,N_17982);
nor U18012 (N_18012,N_17969,N_17926);
or U18013 (N_18013,N_17889,N_17974);
nor U18014 (N_18014,N_17898,N_17846);
xor U18015 (N_18015,N_17916,N_17810);
nand U18016 (N_18016,N_17803,N_17892);
nand U18017 (N_18017,N_17918,N_17876);
nand U18018 (N_18018,N_17972,N_17853);
nor U18019 (N_18019,N_17962,N_17906);
nor U18020 (N_18020,N_17886,N_17887);
and U18021 (N_18021,N_17814,N_17881);
nand U18022 (N_18022,N_17885,N_17823);
nand U18023 (N_18023,N_17826,N_17848);
or U18024 (N_18024,N_17977,N_17939);
or U18025 (N_18025,N_17935,N_17883);
and U18026 (N_18026,N_17981,N_17808);
and U18027 (N_18027,N_17818,N_17984);
nor U18028 (N_18028,N_17806,N_17965);
nor U18029 (N_18029,N_17976,N_17888);
or U18030 (N_18030,N_17951,N_17925);
or U18031 (N_18031,N_17968,N_17955);
nand U18032 (N_18032,N_17832,N_17943);
nor U18033 (N_18033,N_17891,N_17850);
and U18034 (N_18034,N_17836,N_17860);
nor U18035 (N_18035,N_17913,N_17904);
xor U18036 (N_18036,N_17844,N_17933);
and U18037 (N_18037,N_17952,N_17953);
and U18038 (N_18038,N_17866,N_17862);
nand U18039 (N_18039,N_17954,N_17940);
and U18040 (N_18040,N_17902,N_17946);
nor U18041 (N_18041,N_17864,N_17971);
nand U18042 (N_18042,N_17845,N_17807);
or U18043 (N_18043,N_17880,N_17992);
and U18044 (N_18044,N_17947,N_17870);
nand U18045 (N_18045,N_17804,N_17979);
nand U18046 (N_18046,N_17914,N_17997);
nor U18047 (N_18047,N_17978,N_17819);
or U18048 (N_18048,N_17959,N_17868);
and U18049 (N_18049,N_17936,N_17929);
nand U18050 (N_18050,N_17874,N_17957);
nand U18051 (N_18051,N_17890,N_17871);
nand U18052 (N_18052,N_17958,N_17967);
nor U18053 (N_18053,N_17834,N_17995);
nor U18054 (N_18054,N_17829,N_17990);
and U18055 (N_18055,N_17937,N_17945);
and U18056 (N_18056,N_17988,N_17884);
nor U18057 (N_18057,N_17948,N_17921);
xor U18058 (N_18058,N_17994,N_17812);
or U18059 (N_18059,N_17816,N_17923);
xor U18060 (N_18060,N_17882,N_17828);
xnor U18061 (N_18061,N_17856,N_17894);
xnor U18062 (N_18062,N_17956,N_17815);
nand U18063 (N_18063,N_17985,N_17863);
nand U18064 (N_18064,N_17841,N_17987);
and U18065 (N_18065,N_17802,N_17896);
nor U18066 (N_18066,N_17973,N_17942);
xnor U18067 (N_18067,N_17905,N_17999);
or U18068 (N_18068,N_17919,N_17915);
or U18069 (N_18069,N_17843,N_17813);
xnor U18070 (N_18070,N_17920,N_17878);
and U18071 (N_18071,N_17938,N_17963);
and U18072 (N_18072,N_17822,N_17852);
nand U18073 (N_18073,N_17817,N_17851);
nor U18074 (N_18074,N_17961,N_17901);
xor U18075 (N_18075,N_17859,N_17833);
nor U18076 (N_18076,N_17927,N_17930);
nand U18077 (N_18077,N_17875,N_17993);
nand U18078 (N_18078,N_17931,N_17909);
nor U18079 (N_18079,N_17941,N_17861);
nor U18080 (N_18080,N_17998,N_17975);
nand U18081 (N_18081,N_17825,N_17855);
and U18082 (N_18082,N_17949,N_17950);
nand U18083 (N_18083,N_17986,N_17922);
or U18084 (N_18084,N_17847,N_17879);
or U18085 (N_18085,N_17839,N_17980);
and U18086 (N_18086,N_17849,N_17837);
and U18087 (N_18087,N_17970,N_17991);
and U18088 (N_18088,N_17895,N_17842);
nand U18089 (N_18089,N_17966,N_17873);
nand U18090 (N_18090,N_17903,N_17964);
or U18091 (N_18091,N_17830,N_17899);
nor U18092 (N_18092,N_17867,N_17924);
xor U18093 (N_18093,N_17831,N_17893);
nand U18094 (N_18094,N_17801,N_17827);
nand U18095 (N_18095,N_17983,N_17854);
nand U18096 (N_18096,N_17934,N_17907);
or U18097 (N_18097,N_17908,N_17865);
nand U18098 (N_18098,N_17928,N_17858);
or U18099 (N_18099,N_17821,N_17912);
and U18100 (N_18100,N_17943,N_17936);
or U18101 (N_18101,N_17939,N_17832);
or U18102 (N_18102,N_17985,N_17841);
nor U18103 (N_18103,N_17972,N_17895);
xnor U18104 (N_18104,N_17825,N_17878);
xnor U18105 (N_18105,N_17869,N_17967);
or U18106 (N_18106,N_17879,N_17849);
nand U18107 (N_18107,N_17801,N_17963);
nor U18108 (N_18108,N_17884,N_17905);
nor U18109 (N_18109,N_17918,N_17986);
or U18110 (N_18110,N_17906,N_17917);
nand U18111 (N_18111,N_17912,N_17824);
nand U18112 (N_18112,N_17919,N_17982);
and U18113 (N_18113,N_17800,N_17843);
xor U18114 (N_18114,N_17900,N_17894);
nand U18115 (N_18115,N_17992,N_17809);
nand U18116 (N_18116,N_17892,N_17898);
nand U18117 (N_18117,N_17828,N_17935);
xnor U18118 (N_18118,N_17998,N_17895);
nor U18119 (N_18119,N_17991,N_17939);
and U18120 (N_18120,N_17952,N_17845);
and U18121 (N_18121,N_17906,N_17972);
nand U18122 (N_18122,N_17889,N_17872);
or U18123 (N_18123,N_17916,N_17983);
nor U18124 (N_18124,N_17892,N_17841);
or U18125 (N_18125,N_17844,N_17901);
or U18126 (N_18126,N_17954,N_17810);
nor U18127 (N_18127,N_17866,N_17871);
and U18128 (N_18128,N_17887,N_17810);
nand U18129 (N_18129,N_17982,N_17913);
xnor U18130 (N_18130,N_17877,N_17830);
nor U18131 (N_18131,N_17873,N_17926);
xor U18132 (N_18132,N_17910,N_17861);
and U18133 (N_18133,N_17942,N_17967);
nand U18134 (N_18134,N_17829,N_17983);
or U18135 (N_18135,N_17969,N_17955);
and U18136 (N_18136,N_17885,N_17883);
or U18137 (N_18137,N_17876,N_17970);
xnor U18138 (N_18138,N_17801,N_17852);
nor U18139 (N_18139,N_17817,N_17876);
or U18140 (N_18140,N_17913,N_17965);
xor U18141 (N_18141,N_17924,N_17959);
nand U18142 (N_18142,N_17925,N_17965);
and U18143 (N_18143,N_17951,N_17999);
nor U18144 (N_18144,N_17832,N_17811);
or U18145 (N_18145,N_17940,N_17887);
nor U18146 (N_18146,N_17808,N_17836);
nand U18147 (N_18147,N_17946,N_17964);
or U18148 (N_18148,N_17990,N_17986);
and U18149 (N_18149,N_17984,N_17829);
nand U18150 (N_18150,N_17828,N_17857);
or U18151 (N_18151,N_17895,N_17994);
or U18152 (N_18152,N_17958,N_17984);
and U18153 (N_18153,N_17974,N_17859);
nand U18154 (N_18154,N_17930,N_17857);
and U18155 (N_18155,N_17958,N_17965);
or U18156 (N_18156,N_17845,N_17971);
or U18157 (N_18157,N_17903,N_17801);
nand U18158 (N_18158,N_17921,N_17934);
nand U18159 (N_18159,N_17988,N_17993);
xor U18160 (N_18160,N_17847,N_17811);
nor U18161 (N_18161,N_17960,N_17951);
nand U18162 (N_18162,N_17916,N_17848);
xnor U18163 (N_18163,N_17849,N_17871);
xnor U18164 (N_18164,N_17913,N_17812);
nor U18165 (N_18165,N_17994,N_17945);
xnor U18166 (N_18166,N_17973,N_17928);
nor U18167 (N_18167,N_17817,N_17945);
xnor U18168 (N_18168,N_17992,N_17998);
nor U18169 (N_18169,N_17897,N_17934);
xor U18170 (N_18170,N_17962,N_17813);
nor U18171 (N_18171,N_17973,N_17964);
xor U18172 (N_18172,N_17843,N_17812);
nor U18173 (N_18173,N_17899,N_17878);
nor U18174 (N_18174,N_17850,N_17988);
xnor U18175 (N_18175,N_17917,N_17971);
and U18176 (N_18176,N_17863,N_17826);
or U18177 (N_18177,N_17941,N_17967);
nor U18178 (N_18178,N_17957,N_17809);
and U18179 (N_18179,N_17849,N_17860);
nand U18180 (N_18180,N_17874,N_17944);
xor U18181 (N_18181,N_17969,N_17865);
and U18182 (N_18182,N_17939,N_17830);
or U18183 (N_18183,N_17912,N_17812);
nor U18184 (N_18184,N_17869,N_17962);
or U18185 (N_18185,N_17870,N_17975);
or U18186 (N_18186,N_17989,N_17871);
nand U18187 (N_18187,N_17999,N_17863);
xnor U18188 (N_18188,N_17967,N_17814);
and U18189 (N_18189,N_17830,N_17903);
and U18190 (N_18190,N_17989,N_17847);
nand U18191 (N_18191,N_17851,N_17922);
or U18192 (N_18192,N_17988,N_17889);
nand U18193 (N_18193,N_17847,N_17947);
xnor U18194 (N_18194,N_17853,N_17970);
nand U18195 (N_18195,N_17915,N_17936);
xor U18196 (N_18196,N_17986,N_17809);
nor U18197 (N_18197,N_17973,N_17828);
and U18198 (N_18198,N_17905,N_17845);
nor U18199 (N_18199,N_17944,N_17857);
nand U18200 (N_18200,N_18027,N_18114);
nor U18201 (N_18201,N_18192,N_18096);
and U18202 (N_18202,N_18159,N_18031);
and U18203 (N_18203,N_18152,N_18092);
nor U18204 (N_18204,N_18182,N_18128);
or U18205 (N_18205,N_18148,N_18003);
or U18206 (N_18206,N_18095,N_18013);
xnor U18207 (N_18207,N_18017,N_18066);
or U18208 (N_18208,N_18195,N_18084);
nor U18209 (N_18209,N_18113,N_18072);
and U18210 (N_18210,N_18076,N_18083);
and U18211 (N_18211,N_18150,N_18140);
nand U18212 (N_18212,N_18030,N_18020);
nor U18213 (N_18213,N_18002,N_18011);
or U18214 (N_18214,N_18161,N_18044);
nand U18215 (N_18215,N_18025,N_18042);
nand U18216 (N_18216,N_18187,N_18109);
or U18217 (N_18217,N_18009,N_18121);
or U18218 (N_18218,N_18060,N_18028);
or U18219 (N_18219,N_18024,N_18055);
nand U18220 (N_18220,N_18110,N_18081);
nand U18221 (N_18221,N_18078,N_18093);
xnor U18222 (N_18222,N_18132,N_18149);
or U18223 (N_18223,N_18177,N_18087);
nand U18224 (N_18224,N_18143,N_18063);
and U18225 (N_18225,N_18054,N_18176);
and U18226 (N_18226,N_18033,N_18018);
xnor U18227 (N_18227,N_18100,N_18080);
xnor U18228 (N_18228,N_18133,N_18144);
or U18229 (N_18229,N_18035,N_18116);
nor U18230 (N_18230,N_18029,N_18154);
xor U18231 (N_18231,N_18034,N_18036);
and U18232 (N_18232,N_18122,N_18174);
or U18233 (N_18233,N_18146,N_18090);
and U18234 (N_18234,N_18099,N_18094);
nand U18235 (N_18235,N_18186,N_18022);
nor U18236 (N_18236,N_18155,N_18131);
and U18237 (N_18237,N_18198,N_18037);
xnor U18238 (N_18238,N_18086,N_18138);
or U18239 (N_18239,N_18021,N_18126);
or U18240 (N_18240,N_18091,N_18059);
nor U18241 (N_18241,N_18194,N_18048);
nor U18242 (N_18242,N_18000,N_18179);
nor U18243 (N_18243,N_18073,N_18160);
and U18244 (N_18244,N_18165,N_18075);
and U18245 (N_18245,N_18124,N_18163);
xor U18246 (N_18246,N_18164,N_18047);
nor U18247 (N_18247,N_18147,N_18015);
nand U18248 (N_18248,N_18130,N_18052);
nor U18249 (N_18249,N_18134,N_18079);
nor U18250 (N_18250,N_18115,N_18162);
or U18251 (N_18251,N_18064,N_18057);
nand U18252 (N_18252,N_18172,N_18097);
xnor U18253 (N_18253,N_18171,N_18180);
xor U18254 (N_18254,N_18061,N_18136);
nor U18255 (N_18255,N_18107,N_18105);
or U18256 (N_18256,N_18008,N_18101);
nand U18257 (N_18257,N_18039,N_18151);
xor U18258 (N_18258,N_18181,N_18199);
or U18259 (N_18259,N_18188,N_18169);
or U18260 (N_18260,N_18108,N_18197);
or U18261 (N_18261,N_18046,N_18127);
or U18262 (N_18262,N_18045,N_18167);
and U18263 (N_18263,N_18053,N_18049);
nand U18264 (N_18264,N_18118,N_18117);
nor U18265 (N_18265,N_18189,N_18129);
and U18266 (N_18266,N_18178,N_18156);
nand U18267 (N_18267,N_18191,N_18023);
and U18268 (N_18268,N_18185,N_18014);
nor U18269 (N_18269,N_18001,N_18119);
and U18270 (N_18270,N_18065,N_18157);
or U18271 (N_18271,N_18196,N_18102);
nor U18272 (N_18272,N_18089,N_18016);
nor U18273 (N_18273,N_18175,N_18032);
and U18274 (N_18274,N_18184,N_18103);
or U18275 (N_18275,N_18058,N_18193);
xor U18276 (N_18276,N_18043,N_18019);
nand U18277 (N_18277,N_18137,N_18088);
and U18278 (N_18278,N_18026,N_18038);
or U18279 (N_18279,N_18145,N_18006);
xnor U18280 (N_18280,N_18141,N_18085);
xnor U18281 (N_18281,N_18125,N_18170);
or U18282 (N_18282,N_18183,N_18153);
and U18283 (N_18283,N_18067,N_18166);
nor U18284 (N_18284,N_18041,N_18158);
or U18285 (N_18285,N_18050,N_18062);
nor U18286 (N_18286,N_18077,N_18012);
or U18287 (N_18287,N_18173,N_18106);
and U18288 (N_18288,N_18004,N_18082);
nand U18289 (N_18289,N_18190,N_18120);
nor U18290 (N_18290,N_18111,N_18112);
and U18291 (N_18291,N_18010,N_18142);
and U18292 (N_18292,N_18071,N_18168);
nand U18293 (N_18293,N_18007,N_18068);
and U18294 (N_18294,N_18056,N_18135);
and U18295 (N_18295,N_18070,N_18074);
and U18296 (N_18296,N_18123,N_18051);
and U18297 (N_18297,N_18098,N_18069);
or U18298 (N_18298,N_18040,N_18005);
and U18299 (N_18299,N_18104,N_18139);
or U18300 (N_18300,N_18166,N_18036);
and U18301 (N_18301,N_18012,N_18022);
xnor U18302 (N_18302,N_18035,N_18151);
nor U18303 (N_18303,N_18149,N_18143);
or U18304 (N_18304,N_18112,N_18192);
and U18305 (N_18305,N_18160,N_18195);
nand U18306 (N_18306,N_18077,N_18050);
xnor U18307 (N_18307,N_18174,N_18047);
or U18308 (N_18308,N_18062,N_18052);
nor U18309 (N_18309,N_18136,N_18028);
nand U18310 (N_18310,N_18166,N_18099);
and U18311 (N_18311,N_18121,N_18073);
xor U18312 (N_18312,N_18017,N_18172);
and U18313 (N_18313,N_18194,N_18102);
or U18314 (N_18314,N_18104,N_18092);
nor U18315 (N_18315,N_18125,N_18098);
nor U18316 (N_18316,N_18146,N_18143);
nor U18317 (N_18317,N_18127,N_18064);
nor U18318 (N_18318,N_18130,N_18092);
xor U18319 (N_18319,N_18117,N_18115);
xnor U18320 (N_18320,N_18065,N_18170);
or U18321 (N_18321,N_18051,N_18089);
and U18322 (N_18322,N_18131,N_18034);
nor U18323 (N_18323,N_18168,N_18070);
xnor U18324 (N_18324,N_18163,N_18048);
or U18325 (N_18325,N_18109,N_18065);
nand U18326 (N_18326,N_18078,N_18018);
and U18327 (N_18327,N_18062,N_18089);
nand U18328 (N_18328,N_18097,N_18028);
nand U18329 (N_18329,N_18152,N_18055);
nor U18330 (N_18330,N_18160,N_18139);
xor U18331 (N_18331,N_18111,N_18020);
nor U18332 (N_18332,N_18044,N_18097);
nand U18333 (N_18333,N_18157,N_18116);
or U18334 (N_18334,N_18160,N_18106);
nor U18335 (N_18335,N_18172,N_18170);
and U18336 (N_18336,N_18048,N_18010);
xor U18337 (N_18337,N_18171,N_18176);
nor U18338 (N_18338,N_18127,N_18119);
nor U18339 (N_18339,N_18159,N_18162);
nand U18340 (N_18340,N_18178,N_18182);
and U18341 (N_18341,N_18049,N_18123);
and U18342 (N_18342,N_18022,N_18054);
xor U18343 (N_18343,N_18167,N_18175);
and U18344 (N_18344,N_18196,N_18153);
nand U18345 (N_18345,N_18103,N_18113);
xnor U18346 (N_18346,N_18068,N_18047);
xnor U18347 (N_18347,N_18088,N_18036);
nor U18348 (N_18348,N_18007,N_18180);
nand U18349 (N_18349,N_18174,N_18068);
or U18350 (N_18350,N_18168,N_18104);
and U18351 (N_18351,N_18070,N_18067);
or U18352 (N_18352,N_18078,N_18016);
nor U18353 (N_18353,N_18081,N_18153);
nor U18354 (N_18354,N_18070,N_18090);
nor U18355 (N_18355,N_18100,N_18058);
nor U18356 (N_18356,N_18095,N_18165);
or U18357 (N_18357,N_18017,N_18060);
xnor U18358 (N_18358,N_18020,N_18025);
or U18359 (N_18359,N_18050,N_18179);
xnor U18360 (N_18360,N_18068,N_18104);
nand U18361 (N_18361,N_18180,N_18144);
or U18362 (N_18362,N_18175,N_18086);
or U18363 (N_18363,N_18083,N_18172);
nor U18364 (N_18364,N_18135,N_18187);
nand U18365 (N_18365,N_18175,N_18154);
xnor U18366 (N_18366,N_18098,N_18048);
nor U18367 (N_18367,N_18153,N_18123);
xnor U18368 (N_18368,N_18181,N_18180);
and U18369 (N_18369,N_18125,N_18099);
nand U18370 (N_18370,N_18062,N_18131);
nand U18371 (N_18371,N_18032,N_18185);
nor U18372 (N_18372,N_18149,N_18163);
and U18373 (N_18373,N_18049,N_18171);
xor U18374 (N_18374,N_18041,N_18169);
nand U18375 (N_18375,N_18197,N_18182);
nor U18376 (N_18376,N_18066,N_18088);
xor U18377 (N_18377,N_18123,N_18021);
xor U18378 (N_18378,N_18095,N_18084);
xnor U18379 (N_18379,N_18170,N_18141);
nor U18380 (N_18380,N_18102,N_18005);
nand U18381 (N_18381,N_18096,N_18084);
nand U18382 (N_18382,N_18121,N_18155);
and U18383 (N_18383,N_18091,N_18090);
nor U18384 (N_18384,N_18155,N_18091);
nor U18385 (N_18385,N_18106,N_18039);
nand U18386 (N_18386,N_18195,N_18181);
xnor U18387 (N_18387,N_18110,N_18152);
xor U18388 (N_18388,N_18025,N_18093);
and U18389 (N_18389,N_18177,N_18103);
nor U18390 (N_18390,N_18028,N_18165);
nor U18391 (N_18391,N_18098,N_18127);
nand U18392 (N_18392,N_18078,N_18086);
and U18393 (N_18393,N_18140,N_18154);
xnor U18394 (N_18394,N_18105,N_18184);
nand U18395 (N_18395,N_18014,N_18103);
or U18396 (N_18396,N_18038,N_18022);
nand U18397 (N_18397,N_18118,N_18073);
xnor U18398 (N_18398,N_18081,N_18187);
and U18399 (N_18399,N_18137,N_18033);
and U18400 (N_18400,N_18319,N_18304);
and U18401 (N_18401,N_18334,N_18276);
and U18402 (N_18402,N_18355,N_18284);
xnor U18403 (N_18403,N_18349,N_18314);
or U18404 (N_18404,N_18331,N_18200);
or U18405 (N_18405,N_18384,N_18392);
nand U18406 (N_18406,N_18260,N_18263);
nand U18407 (N_18407,N_18214,N_18318);
and U18408 (N_18408,N_18267,N_18369);
nor U18409 (N_18409,N_18381,N_18273);
and U18410 (N_18410,N_18330,N_18307);
or U18411 (N_18411,N_18213,N_18327);
nor U18412 (N_18412,N_18306,N_18219);
nand U18413 (N_18413,N_18382,N_18370);
nand U18414 (N_18414,N_18309,N_18275);
xor U18415 (N_18415,N_18385,N_18301);
nor U18416 (N_18416,N_18253,N_18345);
and U18417 (N_18417,N_18338,N_18238);
nor U18418 (N_18418,N_18336,N_18278);
or U18419 (N_18419,N_18320,N_18230);
xnor U18420 (N_18420,N_18302,N_18371);
and U18421 (N_18421,N_18212,N_18285);
or U18422 (N_18422,N_18347,N_18256);
and U18423 (N_18423,N_18298,N_18364);
nor U18424 (N_18424,N_18265,N_18358);
xnor U18425 (N_18425,N_18311,N_18246);
xnor U18426 (N_18426,N_18234,N_18356);
or U18427 (N_18427,N_18373,N_18380);
nor U18428 (N_18428,N_18288,N_18249);
nand U18429 (N_18429,N_18360,N_18341);
xnor U18430 (N_18430,N_18289,N_18317);
or U18431 (N_18431,N_18243,N_18312);
and U18432 (N_18432,N_18296,N_18223);
xnor U18433 (N_18433,N_18261,N_18332);
or U18434 (N_18434,N_18375,N_18272);
xor U18435 (N_18435,N_18368,N_18376);
or U18436 (N_18436,N_18286,N_18335);
xnor U18437 (N_18437,N_18300,N_18205);
and U18438 (N_18438,N_18344,N_18269);
xor U18439 (N_18439,N_18348,N_18248);
or U18440 (N_18440,N_18351,N_18325);
nor U18441 (N_18441,N_18244,N_18342);
nand U18442 (N_18442,N_18383,N_18262);
or U18443 (N_18443,N_18291,N_18329);
nor U18444 (N_18444,N_18220,N_18268);
xor U18445 (N_18445,N_18316,N_18391);
nand U18446 (N_18446,N_18207,N_18353);
and U18447 (N_18447,N_18233,N_18390);
xnor U18448 (N_18448,N_18326,N_18237);
xor U18449 (N_18449,N_18204,N_18362);
nor U18450 (N_18450,N_18216,N_18203);
nor U18451 (N_18451,N_18290,N_18374);
and U18452 (N_18452,N_18366,N_18283);
nor U18453 (N_18453,N_18395,N_18202);
or U18454 (N_18454,N_18271,N_18310);
nand U18455 (N_18455,N_18240,N_18270);
and U18456 (N_18456,N_18379,N_18232);
xor U18457 (N_18457,N_18264,N_18337);
nand U18458 (N_18458,N_18287,N_18250);
nand U18459 (N_18459,N_18235,N_18357);
nand U18460 (N_18460,N_18363,N_18313);
nand U18461 (N_18461,N_18252,N_18201);
nor U18462 (N_18462,N_18305,N_18333);
xnor U18463 (N_18463,N_18292,N_18293);
or U18464 (N_18464,N_18394,N_18239);
nand U18465 (N_18465,N_18321,N_18322);
nor U18466 (N_18466,N_18258,N_18211);
nor U18467 (N_18467,N_18227,N_18282);
xnor U18468 (N_18468,N_18294,N_18388);
nor U18469 (N_18469,N_18225,N_18323);
or U18470 (N_18470,N_18352,N_18297);
nor U18471 (N_18471,N_18277,N_18372);
xnor U18472 (N_18472,N_18257,N_18209);
xor U18473 (N_18473,N_18361,N_18339);
xnor U18474 (N_18474,N_18308,N_18254);
or U18475 (N_18475,N_18245,N_18346);
nand U18476 (N_18476,N_18222,N_18350);
nand U18477 (N_18477,N_18295,N_18266);
nor U18478 (N_18478,N_18354,N_18241);
nand U18479 (N_18479,N_18226,N_18359);
or U18480 (N_18480,N_18324,N_18208);
xor U18481 (N_18481,N_18377,N_18228);
xnor U18482 (N_18482,N_18315,N_18218);
xor U18483 (N_18483,N_18398,N_18217);
or U18484 (N_18484,N_18328,N_18231);
or U18485 (N_18485,N_18386,N_18251);
nor U18486 (N_18486,N_18299,N_18206);
and U18487 (N_18487,N_18397,N_18279);
nor U18488 (N_18488,N_18399,N_18210);
nand U18489 (N_18489,N_18303,N_18259);
or U18490 (N_18490,N_18236,N_18340);
nor U18491 (N_18491,N_18221,N_18247);
xnor U18492 (N_18492,N_18365,N_18281);
nor U18493 (N_18493,N_18387,N_18229);
and U18494 (N_18494,N_18389,N_18224);
or U18495 (N_18495,N_18396,N_18393);
nand U18496 (N_18496,N_18274,N_18242);
xor U18497 (N_18497,N_18378,N_18280);
nor U18498 (N_18498,N_18215,N_18343);
nand U18499 (N_18499,N_18367,N_18255);
nor U18500 (N_18500,N_18268,N_18256);
xnor U18501 (N_18501,N_18372,N_18242);
and U18502 (N_18502,N_18204,N_18258);
or U18503 (N_18503,N_18231,N_18250);
or U18504 (N_18504,N_18330,N_18255);
xor U18505 (N_18505,N_18209,N_18292);
or U18506 (N_18506,N_18298,N_18353);
xnor U18507 (N_18507,N_18303,N_18267);
nor U18508 (N_18508,N_18279,N_18326);
nor U18509 (N_18509,N_18357,N_18253);
nor U18510 (N_18510,N_18274,N_18357);
xor U18511 (N_18511,N_18353,N_18326);
and U18512 (N_18512,N_18334,N_18347);
or U18513 (N_18513,N_18275,N_18208);
nor U18514 (N_18514,N_18254,N_18235);
and U18515 (N_18515,N_18384,N_18311);
xor U18516 (N_18516,N_18259,N_18314);
nor U18517 (N_18517,N_18310,N_18369);
nand U18518 (N_18518,N_18274,N_18374);
nand U18519 (N_18519,N_18348,N_18306);
xnor U18520 (N_18520,N_18297,N_18320);
and U18521 (N_18521,N_18233,N_18301);
nand U18522 (N_18522,N_18212,N_18395);
or U18523 (N_18523,N_18334,N_18232);
xnor U18524 (N_18524,N_18259,N_18313);
and U18525 (N_18525,N_18315,N_18237);
or U18526 (N_18526,N_18356,N_18316);
nor U18527 (N_18527,N_18328,N_18235);
xnor U18528 (N_18528,N_18294,N_18276);
or U18529 (N_18529,N_18339,N_18245);
nor U18530 (N_18530,N_18229,N_18313);
or U18531 (N_18531,N_18285,N_18242);
nor U18532 (N_18532,N_18261,N_18298);
xnor U18533 (N_18533,N_18362,N_18260);
nand U18534 (N_18534,N_18389,N_18346);
nand U18535 (N_18535,N_18348,N_18282);
nand U18536 (N_18536,N_18227,N_18207);
nand U18537 (N_18537,N_18225,N_18379);
nand U18538 (N_18538,N_18206,N_18254);
nor U18539 (N_18539,N_18252,N_18215);
or U18540 (N_18540,N_18212,N_18256);
and U18541 (N_18541,N_18329,N_18342);
nor U18542 (N_18542,N_18248,N_18281);
and U18543 (N_18543,N_18253,N_18278);
nor U18544 (N_18544,N_18294,N_18364);
xnor U18545 (N_18545,N_18374,N_18331);
nand U18546 (N_18546,N_18305,N_18267);
and U18547 (N_18547,N_18227,N_18299);
nand U18548 (N_18548,N_18352,N_18308);
or U18549 (N_18549,N_18389,N_18329);
xor U18550 (N_18550,N_18344,N_18316);
and U18551 (N_18551,N_18207,N_18311);
and U18552 (N_18552,N_18224,N_18319);
nand U18553 (N_18553,N_18393,N_18230);
xor U18554 (N_18554,N_18394,N_18336);
nand U18555 (N_18555,N_18244,N_18395);
xnor U18556 (N_18556,N_18355,N_18314);
nand U18557 (N_18557,N_18306,N_18254);
and U18558 (N_18558,N_18231,N_18237);
xnor U18559 (N_18559,N_18298,N_18241);
or U18560 (N_18560,N_18303,N_18230);
nor U18561 (N_18561,N_18309,N_18374);
or U18562 (N_18562,N_18281,N_18289);
xor U18563 (N_18563,N_18205,N_18254);
xor U18564 (N_18564,N_18287,N_18223);
nand U18565 (N_18565,N_18294,N_18226);
xor U18566 (N_18566,N_18323,N_18342);
or U18567 (N_18567,N_18287,N_18215);
nor U18568 (N_18568,N_18356,N_18204);
nor U18569 (N_18569,N_18380,N_18331);
or U18570 (N_18570,N_18395,N_18330);
nand U18571 (N_18571,N_18281,N_18241);
xor U18572 (N_18572,N_18239,N_18242);
xnor U18573 (N_18573,N_18251,N_18215);
and U18574 (N_18574,N_18265,N_18219);
or U18575 (N_18575,N_18235,N_18301);
xnor U18576 (N_18576,N_18273,N_18356);
and U18577 (N_18577,N_18249,N_18234);
nor U18578 (N_18578,N_18329,N_18209);
nand U18579 (N_18579,N_18325,N_18355);
and U18580 (N_18580,N_18331,N_18296);
and U18581 (N_18581,N_18294,N_18292);
and U18582 (N_18582,N_18385,N_18263);
and U18583 (N_18583,N_18225,N_18328);
xor U18584 (N_18584,N_18383,N_18358);
xnor U18585 (N_18585,N_18243,N_18245);
nand U18586 (N_18586,N_18200,N_18247);
and U18587 (N_18587,N_18390,N_18282);
or U18588 (N_18588,N_18246,N_18389);
nand U18589 (N_18589,N_18294,N_18242);
or U18590 (N_18590,N_18349,N_18259);
nand U18591 (N_18591,N_18237,N_18238);
nand U18592 (N_18592,N_18347,N_18307);
nand U18593 (N_18593,N_18221,N_18388);
nor U18594 (N_18594,N_18249,N_18348);
xor U18595 (N_18595,N_18224,N_18253);
nor U18596 (N_18596,N_18263,N_18350);
xnor U18597 (N_18597,N_18350,N_18329);
xor U18598 (N_18598,N_18357,N_18273);
or U18599 (N_18599,N_18234,N_18292);
nor U18600 (N_18600,N_18536,N_18514);
nand U18601 (N_18601,N_18517,N_18416);
or U18602 (N_18602,N_18581,N_18574);
and U18603 (N_18603,N_18501,N_18493);
and U18604 (N_18604,N_18473,N_18489);
or U18605 (N_18605,N_18445,N_18556);
nor U18606 (N_18606,N_18408,N_18504);
nand U18607 (N_18607,N_18502,N_18437);
nor U18608 (N_18608,N_18503,N_18465);
nand U18609 (N_18609,N_18446,N_18407);
and U18610 (N_18610,N_18469,N_18464);
or U18611 (N_18611,N_18568,N_18570);
nor U18612 (N_18612,N_18543,N_18566);
xnor U18613 (N_18613,N_18577,N_18494);
xnor U18614 (N_18614,N_18497,N_18561);
nor U18615 (N_18615,N_18554,N_18506);
or U18616 (N_18616,N_18591,N_18460);
or U18617 (N_18617,N_18576,N_18491);
and U18618 (N_18618,N_18466,N_18401);
nand U18619 (N_18619,N_18511,N_18414);
or U18620 (N_18620,N_18425,N_18563);
and U18621 (N_18621,N_18426,N_18589);
nand U18622 (N_18622,N_18528,N_18512);
xnor U18623 (N_18623,N_18569,N_18524);
nand U18624 (N_18624,N_18499,N_18546);
or U18625 (N_18625,N_18564,N_18553);
nor U18626 (N_18626,N_18427,N_18451);
or U18627 (N_18627,N_18418,N_18537);
nand U18628 (N_18628,N_18551,N_18450);
xnor U18629 (N_18629,N_18478,N_18540);
xor U18630 (N_18630,N_18498,N_18444);
xor U18631 (N_18631,N_18583,N_18412);
or U18632 (N_18632,N_18548,N_18484);
and U18633 (N_18633,N_18420,N_18482);
or U18634 (N_18634,N_18441,N_18458);
nand U18635 (N_18635,N_18526,N_18505);
xnor U18636 (N_18636,N_18456,N_18559);
nor U18637 (N_18637,N_18558,N_18532);
nand U18638 (N_18638,N_18409,N_18495);
and U18639 (N_18639,N_18402,N_18455);
nor U18640 (N_18640,N_18541,N_18463);
and U18641 (N_18641,N_18599,N_18405);
or U18642 (N_18642,N_18474,N_18417);
nand U18643 (N_18643,N_18421,N_18529);
xor U18644 (N_18644,N_18467,N_18587);
or U18645 (N_18645,N_18555,N_18567);
xnor U18646 (N_18646,N_18457,N_18406);
xnor U18647 (N_18647,N_18435,N_18507);
or U18648 (N_18648,N_18578,N_18513);
and U18649 (N_18649,N_18552,N_18462);
nor U18650 (N_18650,N_18492,N_18515);
nor U18651 (N_18651,N_18485,N_18522);
nand U18652 (N_18652,N_18580,N_18510);
nand U18653 (N_18653,N_18475,N_18550);
or U18654 (N_18654,N_18448,N_18443);
or U18655 (N_18655,N_18440,N_18411);
or U18656 (N_18656,N_18423,N_18545);
or U18657 (N_18657,N_18508,N_18571);
or U18658 (N_18658,N_18410,N_18477);
xor U18659 (N_18659,N_18500,N_18403);
nand U18660 (N_18660,N_18509,N_18594);
nor U18661 (N_18661,N_18582,N_18527);
and U18662 (N_18662,N_18496,N_18480);
xor U18663 (N_18663,N_18472,N_18415);
xor U18664 (N_18664,N_18481,N_18468);
or U18665 (N_18665,N_18442,N_18454);
and U18666 (N_18666,N_18471,N_18530);
xnor U18667 (N_18667,N_18584,N_18518);
xor U18668 (N_18668,N_18521,N_18596);
and U18669 (N_18669,N_18486,N_18470);
and U18670 (N_18670,N_18424,N_18519);
xor U18671 (N_18671,N_18557,N_18565);
nand U18672 (N_18672,N_18431,N_18516);
nor U18673 (N_18673,N_18588,N_18479);
nor U18674 (N_18674,N_18447,N_18573);
xnor U18675 (N_18675,N_18535,N_18597);
and U18676 (N_18676,N_18429,N_18487);
nand U18677 (N_18677,N_18523,N_18572);
xnor U18678 (N_18678,N_18534,N_18593);
and U18679 (N_18679,N_18542,N_18449);
and U18680 (N_18680,N_18560,N_18439);
xor U18681 (N_18681,N_18476,N_18531);
and U18682 (N_18682,N_18452,N_18598);
or U18683 (N_18683,N_18422,N_18438);
nand U18684 (N_18684,N_18490,N_18538);
or U18685 (N_18685,N_18525,N_18433);
or U18686 (N_18686,N_18547,N_18434);
xor U18687 (N_18687,N_18428,N_18539);
xnor U18688 (N_18688,N_18579,N_18585);
nand U18689 (N_18689,N_18488,N_18544);
xor U18690 (N_18690,N_18520,N_18590);
nand U18691 (N_18691,N_18400,N_18575);
and U18692 (N_18692,N_18586,N_18533);
xor U18693 (N_18693,N_18436,N_18430);
nand U18694 (N_18694,N_18592,N_18562);
and U18695 (N_18695,N_18453,N_18595);
and U18696 (N_18696,N_18419,N_18549);
xnor U18697 (N_18697,N_18461,N_18404);
xor U18698 (N_18698,N_18432,N_18483);
or U18699 (N_18699,N_18459,N_18413);
or U18700 (N_18700,N_18542,N_18562);
xor U18701 (N_18701,N_18551,N_18556);
or U18702 (N_18702,N_18455,N_18517);
and U18703 (N_18703,N_18545,N_18582);
and U18704 (N_18704,N_18557,N_18544);
or U18705 (N_18705,N_18434,N_18403);
xnor U18706 (N_18706,N_18417,N_18578);
nor U18707 (N_18707,N_18579,N_18505);
xnor U18708 (N_18708,N_18494,N_18530);
or U18709 (N_18709,N_18577,N_18451);
nor U18710 (N_18710,N_18510,N_18489);
nor U18711 (N_18711,N_18534,N_18510);
nor U18712 (N_18712,N_18446,N_18460);
nand U18713 (N_18713,N_18479,N_18500);
nor U18714 (N_18714,N_18576,N_18408);
xor U18715 (N_18715,N_18552,N_18548);
nor U18716 (N_18716,N_18425,N_18502);
or U18717 (N_18717,N_18566,N_18472);
nor U18718 (N_18718,N_18559,N_18413);
nor U18719 (N_18719,N_18404,N_18422);
nor U18720 (N_18720,N_18483,N_18529);
and U18721 (N_18721,N_18479,N_18563);
and U18722 (N_18722,N_18528,N_18538);
nand U18723 (N_18723,N_18493,N_18440);
nand U18724 (N_18724,N_18571,N_18587);
nand U18725 (N_18725,N_18556,N_18558);
nor U18726 (N_18726,N_18461,N_18589);
and U18727 (N_18727,N_18572,N_18529);
nand U18728 (N_18728,N_18553,N_18554);
or U18729 (N_18729,N_18524,N_18578);
or U18730 (N_18730,N_18403,N_18527);
xnor U18731 (N_18731,N_18538,N_18417);
nor U18732 (N_18732,N_18543,N_18522);
nand U18733 (N_18733,N_18536,N_18555);
nand U18734 (N_18734,N_18425,N_18455);
nor U18735 (N_18735,N_18570,N_18489);
and U18736 (N_18736,N_18595,N_18597);
or U18737 (N_18737,N_18512,N_18567);
and U18738 (N_18738,N_18546,N_18463);
nor U18739 (N_18739,N_18486,N_18580);
or U18740 (N_18740,N_18468,N_18527);
nor U18741 (N_18741,N_18524,N_18520);
nor U18742 (N_18742,N_18460,N_18568);
and U18743 (N_18743,N_18437,N_18409);
xor U18744 (N_18744,N_18578,N_18505);
and U18745 (N_18745,N_18560,N_18573);
and U18746 (N_18746,N_18567,N_18486);
nand U18747 (N_18747,N_18563,N_18464);
xor U18748 (N_18748,N_18405,N_18550);
nor U18749 (N_18749,N_18479,N_18531);
xor U18750 (N_18750,N_18410,N_18560);
xor U18751 (N_18751,N_18446,N_18428);
and U18752 (N_18752,N_18570,N_18581);
nand U18753 (N_18753,N_18435,N_18486);
or U18754 (N_18754,N_18522,N_18489);
nand U18755 (N_18755,N_18584,N_18408);
xor U18756 (N_18756,N_18590,N_18492);
or U18757 (N_18757,N_18566,N_18597);
and U18758 (N_18758,N_18442,N_18554);
and U18759 (N_18759,N_18560,N_18443);
or U18760 (N_18760,N_18458,N_18598);
and U18761 (N_18761,N_18559,N_18410);
nand U18762 (N_18762,N_18468,N_18436);
nor U18763 (N_18763,N_18436,N_18425);
nand U18764 (N_18764,N_18574,N_18538);
xnor U18765 (N_18765,N_18569,N_18561);
nand U18766 (N_18766,N_18411,N_18516);
or U18767 (N_18767,N_18542,N_18593);
xor U18768 (N_18768,N_18501,N_18410);
or U18769 (N_18769,N_18489,N_18526);
xnor U18770 (N_18770,N_18542,N_18439);
xnor U18771 (N_18771,N_18527,N_18452);
xnor U18772 (N_18772,N_18553,N_18484);
or U18773 (N_18773,N_18406,N_18410);
and U18774 (N_18774,N_18514,N_18560);
xnor U18775 (N_18775,N_18520,N_18440);
and U18776 (N_18776,N_18492,N_18522);
xor U18777 (N_18777,N_18509,N_18419);
nand U18778 (N_18778,N_18546,N_18466);
and U18779 (N_18779,N_18440,N_18427);
xnor U18780 (N_18780,N_18448,N_18504);
nor U18781 (N_18781,N_18538,N_18595);
and U18782 (N_18782,N_18583,N_18571);
or U18783 (N_18783,N_18448,N_18545);
nor U18784 (N_18784,N_18563,N_18514);
or U18785 (N_18785,N_18439,N_18533);
xnor U18786 (N_18786,N_18546,N_18464);
nand U18787 (N_18787,N_18488,N_18452);
and U18788 (N_18788,N_18408,N_18445);
and U18789 (N_18789,N_18450,N_18557);
nor U18790 (N_18790,N_18495,N_18578);
xnor U18791 (N_18791,N_18497,N_18477);
nor U18792 (N_18792,N_18480,N_18414);
nand U18793 (N_18793,N_18522,N_18439);
xor U18794 (N_18794,N_18414,N_18592);
xnor U18795 (N_18795,N_18538,N_18599);
or U18796 (N_18796,N_18552,N_18500);
nand U18797 (N_18797,N_18440,N_18446);
nand U18798 (N_18798,N_18504,N_18554);
nor U18799 (N_18799,N_18559,N_18412);
xor U18800 (N_18800,N_18789,N_18763);
and U18801 (N_18801,N_18724,N_18625);
and U18802 (N_18802,N_18755,N_18691);
nand U18803 (N_18803,N_18657,N_18608);
and U18804 (N_18804,N_18642,N_18716);
and U18805 (N_18805,N_18651,N_18614);
nor U18806 (N_18806,N_18797,N_18692);
nand U18807 (N_18807,N_18680,N_18672);
nand U18808 (N_18808,N_18606,N_18664);
or U18809 (N_18809,N_18654,N_18784);
and U18810 (N_18810,N_18718,N_18698);
xnor U18811 (N_18811,N_18669,N_18773);
or U18812 (N_18812,N_18686,N_18757);
and U18813 (N_18813,N_18613,N_18634);
nor U18814 (N_18814,N_18780,N_18701);
and U18815 (N_18815,N_18626,N_18772);
and U18816 (N_18816,N_18779,N_18618);
nor U18817 (N_18817,N_18725,N_18603);
or U18818 (N_18818,N_18743,N_18783);
xnor U18819 (N_18819,N_18735,N_18611);
nand U18820 (N_18820,N_18717,N_18726);
nor U18821 (N_18821,N_18629,N_18781);
nor U18822 (N_18822,N_18689,N_18786);
xor U18823 (N_18823,N_18697,N_18631);
nor U18824 (N_18824,N_18700,N_18675);
xnor U18825 (N_18825,N_18742,N_18794);
nand U18826 (N_18826,N_18740,N_18759);
nand U18827 (N_18827,N_18741,N_18760);
and U18828 (N_18828,N_18776,N_18667);
nand U18829 (N_18829,N_18696,N_18695);
xor U18830 (N_18830,N_18721,N_18727);
or U18831 (N_18831,N_18720,N_18640);
nand U18832 (N_18832,N_18652,N_18636);
xor U18833 (N_18833,N_18604,N_18681);
xor U18834 (N_18834,N_18655,N_18676);
or U18835 (N_18835,N_18702,N_18771);
nand U18836 (N_18836,N_18737,N_18762);
and U18837 (N_18837,N_18775,N_18621);
and U18838 (N_18838,N_18798,N_18661);
and U18839 (N_18839,N_18766,N_18738);
and U18840 (N_18840,N_18601,N_18615);
xnor U18841 (N_18841,N_18602,N_18722);
nor U18842 (N_18842,N_18677,N_18715);
nor U18843 (N_18843,N_18778,N_18699);
nand U18844 (N_18844,N_18739,N_18728);
nand U18845 (N_18845,N_18768,N_18649);
xor U18846 (N_18846,N_18777,N_18714);
and U18847 (N_18847,N_18612,N_18656);
or U18848 (N_18848,N_18782,N_18765);
xnor U18849 (N_18849,N_18616,N_18736);
nor U18850 (N_18850,N_18650,N_18796);
nand U18851 (N_18851,N_18619,N_18648);
and U18852 (N_18852,N_18756,N_18761);
nand U18853 (N_18853,N_18638,N_18704);
and U18854 (N_18854,N_18785,N_18635);
nor U18855 (N_18855,N_18693,N_18643);
nor U18856 (N_18856,N_18745,N_18607);
nor U18857 (N_18857,N_18733,N_18788);
or U18858 (N_18858,N_18787,N_18666);
or U18859 (N_18859,N_18709,N_18690);
nand U18860 (N_18860,N_18644,N_18665);
xor U18861 (N_18861,N_18605,N_18639);
nand U18862 (N_18862,N_18734,N_18630);
or U18863 (N_18863,N_18645,N_18632);
or U18864 (N_18864,N_18617,N_18791);
and U18865 (N_18865,N_18694,N_18749);
xor U18866 (N_18866,N_18711,N_18622);
and U18867 (N_18867,N_18679,N_18712);
xnor U18868 (N_18868,N_18770,N_18663);
xnor U18869 (N_18869,N_18747,N_18752);
and U18870 (N_18870,N_18793,N_18729);
nor U18871 (N_18871,N_18646,N_18731);
nand U18872 (N_18872,N_18637,N_18792);
xor U18873 (N_18873,N_18688,N_18730);
or U18874 (N_18874,N_18662,N_18758);
or U18875 (N_18875,N_18620,N_18678);
and U18876 (N_18876,N_18609,N_18703);
xnor U18877 (N_18877,N_18732,N_18627);
xnor U18878 (N_18878,N_18683,N_18795);
nor U18879 (N_18879,N_18653,N_18799);
xor U18880 (N_18880,N_18713,N_18658);
xnor U18881 (N_18881,N_18706,N_18790);
or U18882 (N_18882,N_18660,N_18624);
nor U18883 (N_18883,N_18668,N_18764);
and U18884 (N_18884,N_18769,N_18641);
and U18885 (N_18885,N_18751,N_18600);
nand U18886 (N_18886,N_18708,N_18674);
nor U18887 (N_18887,N_18671,N_18767);
and U18888 (N_18888,N_18687,N_18719);
nand U18889 (N_18889,N_18684,N_18633);
nor U18890 (N_18890,N_18753,N_18659);
or U18891 (N_18891,N_18744,N_18682);
nand U18892 (N_18892,N_18628,N_18754);
nand U18893 (N_18893,N_18610,N_18705);
xnor U18894 (N_18894,N_18647,N_18685);
nand U18895 (N_18895,N_18750,N_18746);
or U18896 (N_18896,N_18710,N_18670);
xnor U18897 (N_18897,N_18748,N_18774);
or U18898 (N_18898,N_18623,N_18723);
and U18899 (N_18899,N_18673,N_18707);
xnor U18900 (N_18900,N_18667,N_18653);
xor U18901 (N_18901,N_18724,N_18609);
or U18902 (N_18902,N_18603,N_18756);
or U18903 (N_18903,N_18760,N_18768);
nand U18904 (N_18904,N_18727,N_18665);
nand U18905 (N_18905,N_18792,N_18714);
and U18906 (N_18906,N_18709,N_18738);
and U18907 (N_18907,N_18702,N_18604);
or U18908 (N_18908,N_18642,N_18720);
xnor U18909 (N_18909,N_18654,N_18780);
nand U18910 (N_18910,N_18737,N_18609);
nand U18911 (N_18911,N_18705,N_18617);
and U18912 (N_18912,N_18793,N_18767);
or U18913 (N_18913,N_18669,N_18632);
or U18914 (N_18914,N_18724,N_18729);
nor U18915 (N_18915,N_18773,N_18696);
xor U18916 (N_18916,N_18751,N_18754);
nor U18917 (N_18917,N_18610,N_18673);
and U18918 (N_18918,N_18631,N_18634);
xor U18919 (N_18919,N_18768,N_18701);
and U18920 (N_18920,N_18648,N_18625);
nand U18921 (N_18921,N_18762,N_18712);
xnor U18922 (N_18922,N_18769,N_18732);
nor U18923 (N_18923,N_18784,N_18689);
and U18924 (N_18924,N_18790,N_18608);
or U18925 (N_18925,N_18627,N_18679);
xnor U18926 (N_18926,N_18675,N_18642);
or U18927 (N_18927,N_18756,N_18659);
and U18928 (N_18928,N_18748,N_18784);
or U18929 (N_18929,N_18760,N_18747);
and U18930 (N_18930,N_18776,N_18699);
nand U18931 (N_18931,N_18726,N_18700);
nand U18932 (N_18932,N_18741,N_18680);
nor U18933 (N_18933,N_18743,N_18606);
and U18934 (N_18934,N_18729,N_18626);
nor U18935 (N_18935,N_18741,N_18776);
or U18936 (N_18936,N_18751,N_18693);
xor U18937 (N_18937,N_18643,N_18745);
xnor U18938 (N_18938,N_18676,N_18692);
and U18939 (N_18939,N_18792,N_18633);
xor U18940 (N_18940,N_18631,N_18726);
or U18941 (N_18941,N_18677,N_18744);
nor U18942 (N_18942,N_18691,N_18798);
or U18943 (N_18943,N_18718,N_18621);
nand U18944 (N_18944,N_18749,N_18742);
nor U18945 (N_18945,N_18670,N_18734);
xor U18946 (N_18946,N_18779,N_18778);
nand U18947 (N_18947,N_18613,N_18672);
xor U18948 (N_18948,N_18784,N_18788);
nand U18949 (N_18949,N_18769,N_18692);
nand U18950 (N_18950,N_18756,N_18652);
nand U18951 (N_18951,N_18647,N_18699);
and U18952 (N_18952,N_18673,N_18620);
or U18953 (N_18953,N_18617,N_18743);
xor U18954 (N_18954,N_18773,N_18694);
or U18955 (N_18955,N_18662,N_18729);
or U18956 (N_18956,N_18625,N_18654);
nand U18957 (N_18957,N_18707,N_18731);
xor U18958 (N_18958,N_18794,N_18758);
xor U18959 (N_18959,N_18726,N_18640);
nand U18960 (N_18960,N_18643,N_18733);
nand U18961 (N_18961,N_18726,N_18769);
nand U18962 (N_18962,N_18654,N_18709);
nor U18963 (N_18963,N_18629,N_18754);
xnor U18964 (N_18964,N_18668,N_18763);
nand U18965 (N_18965,N_18732,N_18755);
or U18966 (N_18966,N_18642,N_18696);
xnor U18967 (N_18967,N_18748,N_18765);
and U18968 (N_18968,N_18657,N_18769);
nor U18969 (N_18969,N_18691,N_18686);
xor U18970 (N_18970,N_18619,N_18686);
and U18971 (N_18971,N_18714,N_18700);
nor U18972 (N_18972,N_18668,N_18687);
xor U18973 (N_18973,N_18672,N_18754);
nor U18974 (N_18974,N_18711,N_18651);
or U18975 (N_18975,N_18714,N_18723);
xnor U18976 (N_18976,N_18777,N_18799);
or U18977 (N_18977,N_18721,N_18723);
or U18978 (N_18978,N_18748,N_18657);
nand U18979 (N_18979,N_18786,N_18746);
xor U18980 (N_18980,N_18754,N_18723);
or U18981 (N_18981,N_18739,N_18688);
or U18982 (N_18982,N_18708,N_18772);
nor U18983 (N_18983,N_18786,N_18656);
xnor U18984 (N_18984,N_18772,N_18749);
xor U18985 (N_18985,N_18649,N_18658);
or U18986 (N_18986,N_18734,N_18672);
xnor U18987 (N_18987,N_18747,N_18679);
or U18988 (N_18988,N_18793,N_18740);
or U18989 (N_18989,N_18661,N_18648);
nand U18990 (N_18990,N_18603,N_18738);
or U18991 (N_18991,N_18663,N_18660);
nor U18992 (N_18992,N_18685,N_18759);
nand U18993 (N_18993,N_18723,N_18720);
and U18994 (N_18994,N_18693,N_18781);
nand U18995 (N_18995,N_18673,N_18647);
nand U18996 (N_18996,N_18704,N_18764);
or U18997 (N_18997,N_18651,N_18792);
and U18998 (N_18998,N_18608,N_18713);
and U18999 (N_18999,N_18731,N_18673);
nor U19000 (N_19000,N_18962,N_18864);
xor U19001 (N_19001,N_18880,N_18909);
nand U19002 (N_19002,N_18941,N_18885);
xor U19003 (N_19003,N_18971,N_18802);
or U19004 (N_19004,N_18946,N_18968);
nand U19005 (N_19005,N_18993,N_18922);
or U19006 (N_19006,N_18845,N_18969);
or U19007 (N_19007,N_18811,N_18850);
or U19008 (N_19008,N_18840,N_18870);
nor U19009 (N_19009,N_18872,N_18925);
nand U19010 (N_19010,N_18826,N_18890);
or U19011 (N_19011,N_18945,N_18851);
nand U19012 (N_19012,N_18810,N_18895);
nand U19013 (N_19013,N_18956,N_18858);
and U19014 (N_19014,N_18806,N_18988);
and U19015 (N_19015,N_18915,N_18821);
nor U19016 (N_19016,N_18817,N_18947);
nand U19017 (N_19017,N_18861,N_18839);
xnor U19018 (N_19018,N_18914,N_18856);
nor U19019 (N_19019,N_18996,N_18819);
nand U19020 (N_19020,N_18935,N_18884);
and U19021 (N_19021,N_18854,N_18959);
nor U19022 (N_19022,N_18828,N_18906);
nor U19023 (N_19023,N_18877,N_18844);
and U19024 (N_19024,N_18957,N_18897);
xor U19025 (N_19025,N_18836,N_18995);
or U19026 (N_19026,N_18830,N_18837);
or U19027 (N_19027,N_18936,N_18980);
nand U19028 (N_19028,N_18847,N_18938);
nand U19029 (N_19029,N_18902,N_18904);
nand U19030 (N_19030,N_18813,N_18822);
xor U19031 (N_19031,N_18990,N_18905);
xor U19032 (N_19032,N_18888,N_18917);
or U19033 (N_19033,N_18866,N_18863);
nor U19034 (N_19034,N_18991,N_18886);
xnor U19035 (N_19035,N_18984,N_18874);
nor U19036 (N_19036,N_18910,N_18809);
or U19037 (N_19037,N_18841,N_18934);
or U19038 (N_19038,N_18825,N_18808);
nand U19039 (N_19039,N_18901,N_18940);
nand U19040 (N_19040,N_18961,N_18986);
nor U19041 (N_19041,N_18801,N_18949);
or U19042 (N_19042,N_18992,N_18865);
nor U19043 (N_19043,N_18816,N_18882);
xnor U19044 (N_19044,N_18893,N_18989);
nor U19045 (N_19045,N_18939,N_18903);
or U19046 (N_19046,N_18800,N_18804);
nor U19047 (N_19047,N_18849,N_18964);
or U19048 (N_19048,N_18918,N_18951);
or U19049 (N_19049,N_18827,N_18948);
nor U19050 (N_19050,N_18852,N_18912);
and U19051 (N_19051,N_18921,N_18927);
nand U19052 (N_19052,N_18883,N_18873);
nand U19053 (N_19053,N_18965,N_18944);
and U19054 (N_19054,N_18973,N_18871);
nand U19055 (N_19055,N_18955,N_18994);
nand U19056 (N_19056,N_18878,N_18982);
and U19057 (N_19057,N_18920,N_18977);
nand U19058 (N_19058,N_18815,N_18860);
and U19059 (N_19059,N_18943,N_18967);
and U19060 (N_19060,N_18853,N_18997);
nor U19061 (N_19061,N_18950,N_18859);
or U19062 (N_19062,N_18919,N_18881);
and U19063 (N_19063,N_18876,N_18879);
or U19064 (N_19064,N_18981,N_18892);
nor U19065 (N_19065,N_18975,N_18823);
xor U19066 (N_19066,N_18829,N_18924);
nor U19067 (N_19067,N_18926,N_18831);
nand U19068 (N_19068,N_18807,N_18834);
and U19069 (N_19069,N_18985,N_18954);
xor U19070 (N_19070,N_18929,N_18966);
or U19071 (N_19071,N_18999,N_18931);
or U19072 (N_19072,N_18896,N_18930);
xor U19073 (N_19073,N_18953,N_18987);
xnor U19074 (N_19074,N_18867,N_18818);
xnor U19075 (N_19075,N_18887,N_18838);
nand U19076 (N_19076,N_18916,N_18891);
and U19077 (N_19077,N_18846,N_18970);
xor U19078 (N_19078,N_18843,N_18869);
and U19079 (N_19079,N_18978,N_18842);
xor U19080 (N_19080,N_18911,N_18960);
nor U19081 (N_19081,N_18857,N_18900);
nor U19082 (N_19082,N_18998,N_18972);
nor U19083 (N_19083,N_18899,N_18894);
or U19084 (N_19084,N_18923,N_18983);
and U19085 (N_19085,N_18976,N_18868);
xor U19086 (N_19086,N_18979,N_18952);
nand U19087 (N_19087,N_18824,N_18805);
and U19088 (N_19088,N_18942,N_18848);
and U19089 (N_19089,N_18958,N_18862);
nor U19090 (N_19090,N_18875,N_18832);
and U19091 (N_19091,N_18833,N_18855);
or U19092 (N_19092,N_18803,N_18907);
nor U19093 (N_19093,N_18812,N_18937);
nor U19094 (N_19094,N_18933,N_18908);
nand U19095 (N_19095,N_18820,N_18898);
nor U19096 (N_19096,N_18932,N_18928);
and U19097 (N_19097,N_18974,N_18835);
nand U19098 (N_19098,N_18913,N_18814);
or U19099 (N_19099,N_18889,N_18963);
or U19100 (N_19100,N_18810,N_18983);
and U19101 (N_19101,N_18960,N_18804);
or U19102 (N_19102,N_18809,N_18901);
xor U19103 (N_19103,N_18811,N_18810);
xnor U19104 (N_19104,N_18819,N_18925);
xnor U19105 (N_19105,N_18812,N_18828);
xor U19106 (N_19106,N_18832,N_18930);
nand U19107 (N_19107,N_18892,N_18963);
nor U19108 (N_19108,N_18957,N_18919);
xor U19109 (N_19109,N_18908,N_18973);
nand U19110 (N_19110,N_18964,N_18843);
or U19111 (N_19111,N_18880,N_18927);
and U19112 (N_19112,N_18907,N_18887);
and U19113 (N_19113,N_18855,N_18805);
nand U19114 (N_19114,N_18900,N_18820);
xnor U19115 (N_19115,N_18871,N_18809);
nand U19116 (N_19116,N_18906,N_18888);
or U19117 (N_19117,N_18909,N_18864);
and U19118 (N_19118,N_18910,N_18898);
xnor U19119 (N_19119,N_18971,N_18947);
or U19120 (N_19120,N_18813,N_18843);
or U19121 (N_19121,N_18816,N_18887);
or U19122 (N_19122,N_18982,N_18826);
xor U19123 (N_19123,N_18906,N_18959);
and U19124 (N_19124,N_18953,N_18922);
xor U19125 (N_19125,N_18803,N_18954);
and U19126 (N_19126,N_18833,N_18888);
or U19127 (N_19127,N_18837,N_18953);
nand U19128 (N_19128,N_18892,N_18856);
xnor U19129 (N_19129,N_18995,N_18878);
and U19130 (N_19130,N_18940,N_18801);
xor U19131 (N_19131,N_18915,N_18962);
and U19132 (N_19132,N_18810,N_18861);
and U19133 (N_19133,N_18824,N_18954);
xor U19134 (N_19134,N_18808,N_18878);
or U19135 (N_19135,N_18823,N_18896);
and U19136 (N_19136,N_18910,N_18860);
xor U19137 (N_19137,N_18963,N_18926);
nand U19138 (N_19138,N_18980,N_18907);
xnor U19139 (N_19139,N_18929,N_18998);
nor U19140 (N_19140,N_18986,N_18894);
nand U19141 (N_19141,N_18923,N_18820);
nand U19142 (N_19142,N_18915,N_18889);
nor U19143 (N_19143,N_18807,N_18851);
or U19144 (N_19144,N_18898,N_18819);
nand U19145 (N_19145,N_18904,N_18943);
xnor U19146 (N_19146,N_18890,N_18829);
or U19147 (N_19147,N_18858,N_18968);
and U19148 (N_19148,N_18853,N_18977);
nand U19149 (N_19149,N_18819,N_18858);
or U19150 (N_19150,N_18890,N_18966);
nor U19151 (N_19151,N_18907,N_18900);
xor U19152 (N_19152,N_18887,N_18934);
and U19153 (N_19153,N_18824,N_18952);
xor U19154 (N_19154,N_18991,N_18947);
xor U19155 (N_19155,N_18892,N_18844);
xor U19156 (N_19156,N_18905,N_18940);
xnor U19157 (N_19157,N_18844,N_18867);
nand U19158 (N_19158,N_18834,N_18829);
nand U19159 (N_19159,N_18800,N_18918);
nand U19160 (N_19160,N_18842,N_18909);
and U19161 (N_19161,N_18903,N_18865);
nor U19162 (N_19162,N_18985,N_18825);
or U19163 (N_19163,N_18802,N_18989);
nand U19164 (N_19164,N_18939,N_18983);
or U19165 (N_19165,N_18965,N_18893);
xnor U19166 (N_19166,N_18812,N_18930);
and U19167 (N_19167,N_18891,N_18800);
nor U19168 (N_19168,N_18848,N_18964);
xor U19169 (N_19169,N_18830,N_18838);
xnor U19170 (N_19170,N_18955,N_18976);
xnor U19171 (N_19171,N_18998,N_18928);
and U19172 (N_19172,N_18903,N_18982);
nand U19173 (N_19173,N_18839,N_18862);
or U19174 (N_19174,N_18869,N_18802);
nand U19175 (N_19175,N_18864,N_18983);
and U19176 (N_19176,N_18954,N_18952);
nor U19177 (N_19177,N_18855,N_18906);
and U19178 (N_19178,N_18813,N_18867);
nand U19179 (N_19179,N_18977,N_18845);
nor U19180 (N_19180,N_18971,N_18975);
xnor U19181 (N_19181,N_18825,N_18861);
xnor U19182 (N_19182,N_18993,N_18900);
and U19183 (N_19183,N_18884,N_18919);
or U19184 (N_19184,N_18997,N_18925);
or U19185 (N_19185,N_18848,N_18921);
or U19186 (N_19186,N_18871,N_18834);
or U19187 (N_19187,N_18907,N_18831);
and U19188 (N_19188,N_18879,N_18888);
xnor U19189 (N_19189,N_18908,N_18878);
and U19190 (N_19190,N_18986,N_18837);
or U19191 (N_19191,N_18917,N_18873);
xor U19192 (N_19192,N_18850,N_18876);
nor U19193 (N_19193,N_18970,N_18897);
nand U19194 (N_19194,N_18877,N_18803);
and U19195 (N_19195,N_18891,N_18877);
nand U19196 (N_19196,N_18833,N_18813);
or U19197 (N_19197,N_18892,N_18814);
nor U19198 (N_19198,N_18951,N_18809);
and U19199 (N_19199,N_18902,N_18822);
or U19200 (N_19200,N_19142,N_19151);
nand U19201 (N_19201,N_19141,N_19023);
xnor U19202 (N_19202,N_19196,N_19183);
and U19203 (N_19203,N_19044,N_19077);
xnor U19204 (N_19204,N_19029,N_19128);
nor U19205 (N_19205,N_19006,N_19106);
nand U19206 (N_19206,N_19157,N_19099);
and U19207 (N_19207,N_19081,N_19059);
and U19208 (N_19208,N_19042,N_19010);
nand U19209 (N_19209,N_19007,N_19137);
and U19210 (N_19210,N_19066,N_19055);
and U19211 (N_19211,N_19039,N_19037);
or U19212 (N_19212,N_19114,N_19086);
xor U19213 (N_19213,N_19144,N_19145);
nand U19214 (N_19214,N_19062,N_19028);
xor U19215 (N_19215,N_19111,N_19171);
nor U19216 (N_19216,N_19045,N_19074);
nand U19217 (N_19217,N_19064,N_19150);
or U19218 (N_19218,N_19002,N_19052);
nand U19219 (N_19219,N_19125,N_19143);
and U19220 (N_19220,N_19087,N_19000);
or U19221 (N_19221,N_19152,N_19119);
and U19222 (N_19222,N_19097,N_19192);
xor U19223 (N_19223,N_19149,N_19176);
nor U19224 (N_19224,N_19001,N_19065);
nand U19225 (N_19225,N_19167,N_19168);
nand U19226 (N_19226,N_19035,N_19079);
nand U19227 (N_19227,N_19108,N_19186);
nand U19228 (N_19228,N_19138,N_19069);
and U19229 (N_19229,N_19158,N_19173);
or U19230 (N_19230,N_19027,N_19004);
nor U19231 (N_19231,N_19082,N_19139);
xnor U19232 (N_19232,N_19022,N_19172);
xor U19233 (N_19233,N_19085,N_19191);
nor U19234 (N_19234,N_19067,N_19076);
and U19235 (N_19235,N_19102,N_19032);
xnor U19236 (N_19236,N_19003,N_19090);
or U19237 (N_19237,N_19084,N_19041);
xor U19238 (N_19238,N_19043,N_19104);
nor U19239 (N_19239,N_19073,N_19020);
nor U19240 (N_19240,N_19019,N_19146);
or U19241 (N_19241,N_19190,N_19013);
or U19242 (N_19242,N_19034,N_19091);
nand U19243 (N_19243,N_19133,N_19130);
nor U19244 (N_19244,N_19060,N_19101);
nor U19245 (N_19245,N_19197,N_19100);
or U19246 (N_19246,N_19193,N_19054);
or U19247 (N_19247,N_19170,N_19040);
and U19248 (N_19248,N_19018,N_19058);
nand U19249 (N_19249,N_19134,N_19036);
nor U19250 (N_19250,N_19123,N_19198);
nand U19251 (N_19251,N_19163,N_19147);
xor U19252 (N_19252,N_19153,N_19113);
nor U19253 (N_19253,N_19159,N_19175);
nand U19254 (N_19254,N_19031,N_19120);
or U19255 (N_19255,N_19103,N_19072);
and U19256 (N_19256,N_19135,N_19030);
xnor U19257 (N_19257,N_19051,N_19188);
xnor U19258 (N_19258,N_19169,N_19187);
nand U19259 (N_19259,N_19110,N_19046);
xor U19260 (N_19260,N_19122,N_19057);
and U19261 (N_19261,N_19180,N_19083);
nor U19262 (N_19262,N_19050,N_19199);
and U19263 (N_19263,N_19154,N_19017);
nand U19264 (N_19264,N_19012,N_19092);
xor U19265 (N_19265,N_19025,N_19179);
nand U19266 (N_19266,N_19165,N_19021);
nand U19267 (N_19267,N_19112,N_19089);
nand U19268 (N_19268,N_19162,N_19116);
and U19269 (N_19269,N_19178,N_19068);
xnor U19270 (N_19270,N_19185,N_19063);
nor U19271 (N_19271,N_19105,N_19174);
nor U19272 (N_19272,N_19109,N_19016);
or U19273 (N_19273,N_19155,N_19009);
nand U19274 (N_19274,N_19107,N_19075);
nand U19275 (N_19275,N_19088,N_19049);
xnor U19276 (N_19276,N_19184,N_19166);
nor U19277 (N_19277,N_19124,N_19195);
nor U19278 (N_19278,N_19177,N_19160);
xor U19279 (N_19279,N_19131,N_19015);
nand U19280 (N_19280,N_19156,N_19011);
and U19281 (N_19281,N_19117,N_19038);
nand U19282 (N_19282,N_19136,N_19070);
and U19283 (N_19283,N_19048,N_19078);
nand U19284 (N_19284,N_19056,N_19161);
xor U19285 (N_19285,N_19194,N_19033);
nor U19286 (N_19286,N_19118,N_19014);
and U19287 (N_19287,N_19140,N_19053);
xnor U19288 (N_19288,N_19094,N_19164);
or U19289 (N_19289,N_19127,N_19148);
nand U19290 (N_19290,N_19098,N_19024);
nand U19291 (N_19291,N_19189,N_19095);
xnor U19292 (N_19292,N_19061,N_19005);
nor U19293 (N_19293,N_19008,N_19181);
or U19294 (N_19294,N_19182,N_19071);
or U19295 (N_19295,N_19126,N_19080);
and U19296 (N_19296,N_19115,N_19096);
and U19297 (N_19297,N_19132,N_19129);
nand U19298 (N_19298,N_19047,N_19093);
nand U19299 (N_19299,N_19026,N_19121);
nand U19300 (N_19300,N_19102,N_19190);
or U19301 (N_19301,N_19175,N_19079);
nand U19302 (N_19302,N_19082,N_19017);
xor U19303 (N_19303,N_19165,N_19057);
xor U19304 (N_19304,N_19120,N_19037);
nor U19305 (N_19305,N_19146,N_19090);
or U19306 (N_19306,N_19091,N_19022);
and U19307 (N_19307,N_19146,N_19147);
nand U19308 (N_19308,N_19177,N_19084);
or U19309 (N_19309,N_19001,N_19169);
nand U19310 (N_19310,N_19134,N_19135);
nand U19311 (N_19311,N_19180,N_19056);
nand U19312 (N_19312,N_19080,N_19160);
nand U19313 (N_19313,N_19196,N_19190);
or U19314 (N_19314,N_19043,N_19098);
xor U19315 (N_19315,N_19084,N_19019);
or U19316 (N_19316,N_19166,N_19027);
or U19317 (N_19317,N_19165,N_19093);
nor U19318 (N_19318,N_19075,N_19184);
nor U19319 (N_19319,N_19124,N_19122);
nand U19320 (N_19320,N_19104,N_19154);
xnor U19321 (N_19321,N_19145,N_19021);
and U19322 (N_19322,N_19036,N_19006);
nor U19323 (N_19323,N_19082,N_19006);
nand U19324 (N_19324,N_19009,N_19086);
nor U19325 (N_19325,N_19184,N_19173);
xnor U19326 (N_19326,N_19029,N_19073);
or U19327 (N_19327,N_19028,N_19057);
nor U19328 (N_19328,N_19146,N_19076);
nor U19329 (N_19329,N_19054,N_19138);
xor U19330 (N_19330,N_19132,N_19138);
nand U19331 (N_19331,N_19002,N_19050);
or U19332 (N_19332,N_19120,N_19020);
xnor U19333 (N_19333,N_19179,N_19004);
xnor U19334 (N_19334,N_19161,N_19083);
xor U19335 (N_19335,N_19023,N_19194);
or U19336 (N_19336,N_19199,N_19156);
or U19337 (N_19337,N_19068,N_19030);
xnor U19338 (N_19338,N_19005,N_19031);
xnor U19339 (N_19339,N_19165,N_19187);
nor U19340 (N_19340,N_19190,N_19095);
nor U19341 (N_19341,N_19181,N_19031);
nand U19342 (N_19342,N_19135,N_19141);
and U19343 (N_19343,N_19144,N_19130);
nor U19344 (N_19344,N_19121,N_19142);
nor U19345 (N_19345,N_19186,N_19099);
or U19346 (N_19346,N_19033,N_19129);
and U19347 (N_19347,N_19113,N_19129);
or U19348 (N_19348,N_19014,N_19003);
nand U19349 (N_19349,N_19004,N_19021);
nand U19350 (N_19350,N_19044,N_19171);
and U19351 (N_19351,N_19152,N_19108);
and U19352 (N_19352,N_19099,N_19058);
and U19353 (N_19353,N_19194,N_19100);
or U19354 (N_19354,N_19115,N_19134);
nor U19355 (N_19355,N_19190,N_19118);
nor U19356 (N_19356,N_19070,N_19088);
or U19357 (N_19357,N_19166,N_19042);
nor U19358 (N_19358,N_19041,N_19050);
nor U19359 (N_19359,N_19188,N_19077);
xnor U19360 (N_19360,N_19058,N_19139);
xor U19361 (N_19361,N_19121,N_19048);
and U19362 (N_19362,N_19182,N_19080);
xnor U19363 (N_19363,N_19122,N_19101);
and U19364 (N_19364,N_19136,N_19155);
nor U19365 (N_19365,N_19113,N_19114);
and U19366 (N_19366,N_19039,N_19082);
xnor U19367 (N_19367,N_19060,N_19133);
xor U19368 (N_19368,N_19001,N_19127);
nand U19369 (N_19369,N_19064,N_19170);
and U19370 (N_19370,N_19079,N_19112);
nand U19371 (N_19371,N_19105,N_19173);
nor U19372 (N_19372,N_19056,N_19084);
and U19373 (N_19373,N_19175,N_19046);
and U19374 (N_19374,N_19071,N_19020);
nand U19375 (N_19375,N_19014,N_19049);
nand U19376 (N_19376,N_19150,N_19169);
xor U19377 (N_19377,N_19044,N_19011);
xor U19378 (N_19378,N_19050,N_19044);
nand U19379 (N_19379,N_19181,N_19175);
or U19380 (N_19380,N_19097,N_19029);
or U19381 (N_19381,N_19156,N_19129);
nand U19382 (N_19382,N_19064,N_19060);
or U19383 (N_19383,N_19052,N_19014);
and U19384 (N_19384,N_19176,N_19171);
and U19385 (N_19385,N_19007,N_19194);
or U19386 (N_19386,N_19109,N_19095);
or U19387 (N_19387,N_19177,N_19192);
or U19388 (N_19388,N_19118,N_19128);
or U19389 (N_19389,N_19043,N_19055);
nand U19390 (N_19390,N_19147,N_19020);
nand U19391 (N_19391,N_19075,N_19046);
and U19392 (N_19392,N_19059,N_19175);
nand U19393 (N_19393,N_19104,N_19139);
xnor U19394 (N_19394,N_19101,N_19190);
nand U19395 (N_19395,N_19174,N_19193);
xnor U19396 (N_19396,N_19087,N_19005);
xor U19397 (N_19397,N_19127,N_19019);
nand U19398 (N_19398,N_19160,N_19156);
nor U19399 (N_19399,N_19080,N_19120);
nor U19400 (N_19400,N_19288,N_19277);
and U19401 (N_19401,N_19394,N_19267);
or U19402 (N_19402,N_19321,N_19206);
or U19403 (N_19403,N_19323,N_19265);
xor U19404 (N_19404,N_19378,N_19366);
nand U19405 (N_19405,N_19281,N_19319);
nor U19406 (N_19406,N_19270,N_19228);
nand U19407 (N_19407,N_19343,N_19363);
nand U19408 (N_19408,N_19210,N_19226);
nand U19409 (N_19409,N_19316,N_19306);
nand U19410 (N_19410,N_19374,N_19360);
nor U19411 (N_19411,N_19268,N_19386);
nand U19412 (N_19412,N_19370,N_19275);
xnor U19413 (N_19413,N_19215,N_19318);
xor U19414 (N_19414,N_19391,N_19263);
and U19415 (N_19415,N_19398,N_19242);
and U19416 (N_19416,N_19326,N_19264);
and U19417 (N_19417,N_19369,N_19346);
xnor U19418 (N_19418,N_19376,N_19325);
nor U19419 (N_19419,N_19335,N_19303);
nand U19420 (N_19420,N_19322,N_19236);
or U19421 (N_19421,N_19393,N_19225);
nand U19422 (N_19422,N_19241,N_19254);
or U19423 (N_19423,N_19240,N_19348);
nor U19424 (N_19424,N_19276,N_19310);
xor U19425 (N_19425,N_19273,N_19257);
nor U19426 (N_19426,N_19201,N_19307);
xnor U19427 (N_19427,N_19332,N_19269);
or U19428 (N_19428,N_19249,N_19350);
nor U19429 (N_19429,N_19308,N_19336);
nand U19430 (N_19430,N_19320,N_19364);
nor U19431 (N_19431,N_19224,N_19246);
nor U19432 (N_19432,N_19373,N_19218);
and U19433 (N_19433,N_19255,N_19205);
nand U19434 (N_19434,N_19304,N_19289);
or U19435 (N_19435,N_19368,N_19227);
or U19436 (N_19436,N_19208,N_19247);
nand U19437 (N_19437,N_19293,N_19358);
and U19438 (N_19438,N_19204,N_19251);
nand U19439 (N_19439,N_19200,N_19399);
nand U19440 (N_19440,N_19230,N_19383);
and U19441 (N_19441,N_19287,N_19235);
and U19442 (N_19442,N_19342,N_19387);
xnor U19443 (N_19443,N_19291,N_19232);
or U19444 (N_19444,N_19219,N_19280);
and U19445 (N_19445,N_19233,N_19274);
nand U19446 (N_19446,N_19207,N_19334);
xor U19447 (N_19447,N_19272,N_19300);
or U19448 (N_19448,N_19248,N_19282);
nor U19449 (N_19449,N_19329,N_19216);
nand U19450 (N_19450,N_19330,N_19349);
xor U19451 (N_19451,N_19375,N_19253);
or U19452 (N_19452,N_19365,N_19250);
nand U19453 (N_19453,N_19299,N_19292);
and U19454 (N_19454,N_19295,N_19222);
or U19455 (N_19455,N_19237,N_19256);
and U19456 (N_19456,N_19362,N_19261);
or U19457 (N_19457,N_19359,N_19259);
nand U19458 (N_19458,N_19361,N_19353);
xnor U19459 (N_19459,N_19377,N_19214);
nand U19460 (N_19460,N_19345,N_19301);
xnor U19461 (N_19461,N_19238,N_19324);
and U19462 (N_19462,N_19396,N_19351);
nor U19463 (N_19463,N_19389,N_19313);
and U19464 (N_19464,N_19296,N_19285);
nand U19465 (N_19465,N_19340,N_19258);
or U19466 (N_19466,N_19355,N_19229);
and U19467 (N_19467,N_19209,N_19212);
nand U19468 (N_19468,N_19262,N_19244);
nand U19469 (N_19469,N_19356,N_19385);
or U19470 (N_19470,N_19290,N_19211);
nand U19471 (N_19471,N_19221,N_19309);
xnor U19472 (N_19472,N_19314,N_19317);
nor U19473 (N_19473,N_19311,N_19203);
xnor U19474 (N_19474,N_19327,N_19302);
nand U19475 (N_19475,N_19352,N_19202);
nand U19476 (N_19476,N_19305,N_19341);
xnor U19477 (N_19477,N_19297,N_19245);
nand U19478 (N_19478,N_19371,N_19271);
nor U19479 (N_19479,N_19357,N_19388);
nand U19480 (N_19480,N_19260,N_19315);
xor U19481 (N_19481,N_19284,N_19397);
or U19482 (N_19482,N_19217,N_19278);
and U19483 (N_19483,N_19286,N_19333);
and U19484 (N_19484,N_19298,N_19382);
nand U19485 (N_19485,N_19395,N_19312);
nor U19486 (N_19486,N_19372,N_19338);
nor U19487 (N_19487,N_19223,N_19294);
and U19488 (N_19488,N_19392,N_19347);
xnor U19489 (N_19489,N_19354,N_19279);
or U19490 (N_19490,N_19266,N_19283);
nor U19491 (N_19491,N_19213,N_19390);
and U19492 (N_19492,N_19331,N_19384);
nor U19493 (N_19493,N_19243,N_19337);
xor U19494 (N_19494,N_19252,N_19234);
nor U19495 (N_19495,N_19239,N_19367);
nand U19496 (N_19496,N_19381,N_19344);
nor U19497 (N_19497,N_19379,N_19380);
nand U19498 (N_19498,N_19220,N_19231);
or U19499 (N_19499,N_19339,N_19328);
nor U19500 (N_19500,N_19391,N_19343);
nor U19501 (N_19501,N_19322,N_19323);
nand U19502 (N_19502,N_19305,N_19230);
or U19503 (N_19503,N_19387,N_19231);
nor U19504 (N_19504,N_19380,N_19305);
xor U19505 (N_19505,N_19213,N_19218);
nor U19506 (N_19506,N_19388,N_19316);
or U19507 (N_19507,N_19267,N_19350);
nor U19508 (N_19508,N_19205,N_19376);
nor U19509 (N_19509,N_19282,N_19397);
or U19510 (N_19510,N_19365,N_19202);
nand U19511 (N_19511,N_19229,N_19251);
xor U19512 (N_19512,N_19279,N_19286);
nand U19513 (N_19513,N_19341,N_19291);
nor U19514 (N_19514,N_19398,N_19303);
xor U19515 (N_19515,N_19253,N_19236);
and U19516 (N_19516,N_19389,N_19300);
nor U19517 (N_19517,N_19318,N_19366);
and U19518 (N_19518,N_19368,N_19365);
nor U19519 (N_19519,N_19359,N_19317);
nand U19520 (N_19520,N_19313,N_19332);
and U19521 (N_19521,N_19369,N_19358);
xor U19522 (N_19522,N_19235,N_19274);
xor U19523 (N_19523,N_19396,N_19271);
xnor U19524 (N_19524,N_19279,N_19272);
or U19525 (N_19525,N_19396,N_19239);
xor U19526 (N_19526,N_19328,N_19301);
xnor U19527 (N_19527,N_19247,N_19393);
xnor U19528 (N_19528,N_19219,N_19379);
or U19529 (N_19529,N_19272,N_19382);
nor U19530 (N_19530,N_19217,N_19310);
nand U19531 (N_19531,N_19312,N_19331);
xnor U19532 (N_19532,N_19272,N_19328);
nand U19533 (N_19533,N_19215,N_19213);
nand U19534 (N_19534,N_19368,N_19297);
nor U19535 (N_19535,N_19311,N_19221);
nand U19536 (N_19536,N_19254,N_19208);
xnor U19537 (N_19537,N_19357,N_19396);
nor U19538 (N_19538,N_19316,N_19207);
or U19539 (N_19539,N_19265,N_19281);
and U19540 (N_19540,N_19216,N_19332);
nor U19541 (N_19541,N_19366,N_19260);
or U19542 (N_19542,N_19380,N_19334);
nor U19543 (N_19543,N_19309,N_19327);
xor U19544 (N_19544,N_19379,N_19345);
nor U19545 (N_19545,N_19293,N_19266);
or U19546 (N_19546,N_19388,N_19306);
nand U19547 (N_19547,N_19262,N_19368);
or U19548 (N_19548,N_19218,N_19377);
and U19549 (N_19549,N_19257,N_19376);
xor U19550 (N_19550,N_19357,N_19300);
nand U19551 (N_19551,N_19398,N_19339);
nand U19552 (N_19552,N_19340,N_19379);
and U19553 (N_19553,N_19325,N_19229);
or U19554 (N_19554,N_19371,N_19256);
nor U19555 (N_19555,N_19304,N_19334);
nand U19556 (N_19556,N_19315,N_19318);
xnor U19557 (N_19557,N_19334,N_19222);
nor U19558 (N_19558,N_19360,N_19381);
nor U19559 (N_19559,N_19339,N_19272);
or U19560 (N_19560,N_19207,N_19264);
xnor U19561 (N_19561,N_19376,N_19353);
nand U19562 (N_19562,N_19244,N_19329);
xnor U19563 (N_19563,N_19350,N_19298);
xor U19564 (N_19564,N_19344,N_19221);
and U19565 (N_19565,N_19243,N_19308);
xor U19566 (N_19566,N_19349,N_19264);
nor U19567 (N_19567,N_19256,N_19399);
or U19568 (N_19568,N_19205,N_19244);
or U19569 (N_19569,N_19297,N_19379);
nor U19570 (N_19570,N_19302,N_19307);
nor U19571 (N_19571,N_19334,N_19283);
nor U19572 (N_19572,N_19372,N_19341);
and U19573 (N_19573,N_19398,N_19305);
and U19574 (N_19574,N_19352,N_19341);
and U19575 (N_19575,N_19201,N_19375);
and U19576 (N_19576,N_19200,N_19304);
or U19577 (N_19577,N_19201,N_19283);
xnor U19578 (N_19578,N_19210,N_19224);
and U19579 (N_19579,N_19285,N_19314);
xor U19580 (N_19580,N_19294,N_19296);
nand U19581 (N_19581,N_19284,N_19253);
nor U19582 (N_19582,N_19209,N_19214);
or U19583 (N_19583,N_19299,N_19305);
nor U19584 (N_19584,N_19296,N_19251);
and U19585 (N_19585,N_19254,N_19356);
xnor U19586 (N_19586,N_19346,N_19364);
or U19587 (N_19587,N_19235,N_19324);
and U19588 (N_19588,N_19207,N_19345);
nand U19589 (N_19589,N_19358,N_19277);
xor U19590 (N_19590,N_19344,N_19340);
or U19591 (N_19591,N_19213,N_19313);
xnor U19592 (N_19592,N_19389,N_19228);
or U19593 (N_19593,N_19317,N_19262);
or U19594 (N_19594,N_19271,N_19380);
nand U19595 (N_19595,N_19291,N_19393);
nand U19596 (N_19596,N_19215,N_19237);
and U19597 (N_19597,N_19249,N_19254);
and U19598 (N_19598,N_19346,N_19231);
nor U19599 (N_19599,N_19365,N_19264);
nand U19600 (N_19600,N_19445,N_19455);
and U19601 (N_19601,N_19571,N_19557);
and U19602 (N_19602,N_19566,N_19404);
nor U19603 (N_19603,N_19567,N_19518);
nand U19604 (N_19604,N_19401,N_19575);
nand U19605 (N_19605,N_19466,N_19539);
nand U19606 (N_19606,N_19416,N_19548);
nor U19607 (N_19607,N_19424,N_19436);
xnor U19608 (N_19608,N_19570,N_19407);
nor U19609 (N_19609,N_19594,N_19593);
nand U19610 (N_19610,N_19415,N_19426);
or U19611 (N_19611,N_19574,N_19408);
nand U19612 (N_19612,N_19454,N_19446);
xnor U19613 (N_19613,N_19521,N_19579);
and U19614 (N_19614,N_19498,N_19460);
nor U19615 (N_19615,N_19591,N_19471);
nor U19616 (N_19616,N_19470,N_19502);
xor U19617 (N_19617,N_19427,N_19540);
or U19618 (N_19618,N_19458,N_19501);
xor U19619 (N_19619,N_19546,N_19556);
nand U19620 (N_19620,N_19505,N_19417);
or U19621 (N_19621,N_19480,N_19526);
xnor U19622 (N_19622,N_19550,N_19434);
nor U19623 (N_19623,N_19409,N_19462);
xor U19624 (N_19624,N_19541,N_19595);
nand U19625 (N_19625,N_19523,N_19512);
xnor U19626 (N_19626,N_19584,N_19587);
and U19627 (N_19627,N_19536,N_19422);
xor U19628 (N_19628,N_19485,N_19479);
and U19629 (N_19629,N_19545,N_19547);
or U19630 (N_19630,N_19464,N_19474);
xor U19631 (N_19631,N_19459,N_19520);
xor U19632 (N_19632,N_19484,N_19497);
or U19633 (N_19633,N_19563,N_19469);
nand U19634 (N_19634,N_19421,N_19544);
xor U19635 (N_19635,N_19439,N_19510);
or U19636 (N_19636,N_19585,N_19553);
nand U19637 (N_19637,N_19565,N_19527);
or U19638 (N_19638,N_19465,N_19431);
or U19639 (N_19639,N_19598,N_19405);
xor U19640 (N_19640,N_19572,N_19449);
or U19641 (N_19641,N_19443,N_19487);
nor U19642 (N_19642,N_19514,N_19419);
and U19643 (N_19643,N_19496,N_19414);
or U19644 (N_19644,N_19413,N_19451);
nand U19645 (N_19645,N_19590,N_19423);
nand U19646 (N_19646,N_19583,N_19542);
nor U19647 (N_19647,N_19519,N_19482);
nor U19648 (N_19648,N_19428,N_19491);
or U19649 (N_19649,N_19499,N_19429);
xor U19650 (N_19650,N_19400,N_19435);
xnor U19651 (N_19651,N_19444,N_19433);
and U19652 (N_19652,N_19525,N_19531);
xnor U19653 (N_19653,N_19508,N_19492);
xnor U19654 (N_19654,N_19534,N_19577);
or U19655 (N_19655,N_19549,N_19437);
xnor U19656 (N_19656,N_19442,N_19582);
and U19657 (N_19657,N_19438,N_19513);
xnor U19658 (N_19658,N_19456,N_19473);
and U19659 (N_19659,N_19410,N_19452);
and U19660 (N_19660,N_19551,N_19552);
nor U19661 (N_19661,N_19578,N_19530);
nand U19662 (N_19662,N_19533,N_19580);
xnor U19663 (N_19663,N_19457,N_19411);
or U19664 (N_19664,N_19569,N_19467);
and U19665 (N_19665,N_19463,N_19558);
xor U19666 (N_19666,N_19418,N_19504);
or U19667 (N_19667,N_19529,N_19588);
nand U19668 (N_19668,N_19586,N_19506);
and U19669 (N_19669,N_19477,N_19441);
and U19670 (N_19670,N_19412,N_19495);
or U19671 (N_19671,N_19489,N_19511);
or U19672 (N_19672,N_19576,N_19453);
and U19673 (N_19673,N_19537,N_19447);
or U19674 (N_19674,N_19554,N_19568);
nand U19675 (N_19675,N_19494,N_19559);
nand U19676 (N_19676,N_19425,N_19483);
nor U19677 (N_19677,N_19468,N_19509);
or U19678 (N_19678,N_19478,N_19481);
or U19679 (N_19679,N_19581,N_19528);
or U19680 (N_19680,N_19532,N_19538);
and U19681 (N_19681,N_19461,N_19450);
nor U19682 (N_19682,N_19599,N_19472);
xnor U19683 (N_19683,N_19555,N_19490);
nand U19684 (N_19684,N_19515,N_19516);
nand U19685 (N_19685,N_19517,N_19440);
nand U19686 (N_19686,N_19432,N_19476);
or U19687 (N_19687,N_19561,N_19475);
nand U19688 (N_19688,N_19507,N_19522);
or U19689 (N_19689,N_19564,N_19488);
or U19690 (N_19690,N_19535,N_19596);
nor U19691 (N_19691,N_19589,N_19448);
xor U19692 (N_19692,N_19402,N_19592);
or U19693 (N_19693,N_19486,N_19493);
and U19694 (N_19694,N_19597,N_19562);
nand U19695 (N_19695,N_19503,N_19420);
and U19696 (N_19696,N_19560,N_19403);
or U19697 (N_19697,N_19524,N_19573);
xor U19698 (N_19698,N_19406,N_19500);
or U19699 (N_19699,N_19543,N_19430);
xor U19700 (N_19700,N_19530,N_19565);
xor U19701 (N_19701,N_19411,N_19410);
nor U19702 (N_19702,N_19580,N_19487);
or U19703 (N_19703,N_19500,N_19559);
nor U19704 (N_19704,N_19488,N_19450);
nand U19705 (N_19705,N_19403,N_19423);
xnor U19706 (N_19706,N_19512,N_19445);
and U19707 (N_19707,N_19491,N_19541);
nor U19708 (N_19708,N_19429,N_19478);
nor U19709 (N_19709,N_19525,N_19454);
and U19710 (N_19710,N_19556,N_19402);
nand U19711 (N_19711,N_19416,N_19494);
nor U19712 (N_19712,N_19478,N_19493);
or U19713 (N_19713,N_19465,N_19541);
and U19714 (N_19714,N_19440,N_19402);
and U19715 (N_19715,N_19472,N_19514);
nor U19716 (N_19716,N_19452,N_19456);
nand U19717 (N_19717,N_19594,N_19404);
or U19718 (N_19718,N_19502,N_19428);
nand U19719 (N_19719,N_19567,N_19421);
nor U19720 (N_19720,N_19436,N_19477);
xnor U19721 (N_19721,N_19443,N_19583);
or U19722 (N_19722,N_19577,N_19483);
nand U19723 (N_19723,N_19402,N_19406);
and U19724 (N_19724,N_19401,N_19469);
or U19725 (N_19725,N_19580,N_19438);
xnor U19726 (N_19726,N_19449,N_19567);
and U19727 (N_19727,N_19491,N_19580);
nand U19728 (N_19728,N_19455,N_19565);
nor U19729 (N_19729,N_19583,N_19403);
xnor U19730 (N_19730,N_19491,N_19445);
xnor U19731 (N_19731,N_19414,N_19598);
xor U19732 (N_19732,N_19520,N_19587);
or U19733 (N_19733,N_19482,N_19559);
nand U19734 (N_19734,N_19564,N_19417);
nand U19735 (N_19735,N_19495,N_19567);
nor U19736 (N_19736,N_19499,N_19411);
nand U19737 (N_19737,N_19559,N_19446);
nand U19738 (N_19738,N_19465,N_19517);
xnor U19739 (N_19739,N_19499,N_19584);
nor U19740 (N_19740,N_19554,N_19598);
or U19741 (N_19741,N_19410,N_19565);
nor U19742 (N_19742,N_19575,N_19544);
nor U19743 (N_19743,N_19517,N_19420);
or U19744 (N_19744,N_19572,N_19593);
and U19745 (N_19745,N_19448,N_19413);
nor U19746 (N_19746,N_19431,N_19473);
nand U19747 (N_19747,N_19459,N_19550);
xor U19748 (N_19748,N_19544,N_19560);
and U19749 (N_19749,N_19477,N_19456);
xor U19750 (N_19750,N_19444,N_19403);
and U19751 (N_19751,N_19576,N_19454);
or U19752 (N_19752,N_19591,N_19555);
xnor U19753 (N_19753,N_19438,N_19508);
and U19754 (N_19754,N_19515,N_19425);
or U19755 (N_19755,N_19542,N_19485);
and U19756 (N_19756,N_19480,N_19402);
nand U19757 (N_19757,N_19560,N_19517);
xor U19758 (N_19758,N_19596,N_19530);
nor U19759 (N_19759,N_19581,N_19582);
nand U19760 (N_19760,N_19571,N_19400);
nand U19761 (N_19761,N_19446,N_19407);
and U19762 (N_19762,N_19598,N_19496);
and U19763 (N_19763,N_19433,N_19598);
and U19764 (N_19764,N_19478,N_19518);
or U19765 (N_19765,N_19453,N_19553);
and U19766 (N_19766,N_19464,N_19571);
xnor U19767 (N_19767,N_19479,N_19410);
and U19768 (N_19768,N_19576,N_19567);
or U19769 (N_19769,N_19466,N_19406);
nand U19770 (N_19770,N_19422,N_19586);
or U19771 (N_19771,N_19577,N_19553);
xnor U19772 (N_19772,N_19435,N_19467);
and U19773 (N_19773,N_19471,N_19569);
and U19774 (N_19774,N_19433,N_19472);
nand U19775 (N_19775,N_19562,N_19510);
xnor U19776 (N_19776,N_19516,N_19463);
nand U19777 (N_19777,N_19445,N_19416);
xor U19778 (N_19778,N_19592,N_19424);
nor U19779 (N_19779,N_19419,N_19423);
nand U19780 (N_19780,N_19452,N_19403);
nor U19781 (N_19781,N_19480,N_19412);
nand U19782 (N_19782,N_19441,N_19532);
and U19783 (N_19783,N_19476,N_19415);
nor U19784 (N_19784,N_19429,N_19417);
xor U19785 (N_19785,N_19564,N_19548);
and U19786 (N_19786,N_19551,N_19588);
and U19787 (N_19787,N_19506,N_19407);
nand U19788 (N_19788,N_19514,N_19411);
or U19789 (N_19789,N_19557,N_19539);
nand U19790 (N_19790,N_19579,N_19541);
nor U19791 (N_19791,N_19470,N_19562);
nor U19792 (N_19792,N_19520,N_19551);
nand U19793 (N_19793,N_19476,N_19407);
nor U19794 (N_19794,N_19436,N_19427);
and U19795 (N_19795,N_19587,N_19490);
and U19796 (N_19796,N_19590,N_19570);
nor U19797 (N_19797,N_19421,N_19526);
nand U19798 (N_19798,N_19514,N_19538);
nand U19799 (N_19799,N_19542,N_19572);
xnor U19800 (N_19800,N_19703,N_19795);
or U19801 (N_19801,N_19611,N_19735);
or U19802 (N_19802,N_19684,N_19711);
nor U19803 (N_19803,N_19690,N_19772);
xnor U19804 (N_19804,N_19730,N_19645);
or U19805 (N_19805,N_19693,N_19783);
nand U19806 (N_19806,N_19759,N_19784);
nor U19807 (N_19807,N_19686,N_19746);
or U19808 (N_19808,N_19752,N_19757);
xnor U19809 (N_19809,N_19643,N_19640);
nand U19810 (N_19810,N_19716,N_19774);
xnor U19811 (N_19811,N_19766,N_19639);
xor U19812 (N_19812,N_19767,N_19647);
or U19813 (N_19813,N_19669,N_19790);
xnor U19814 (N_19814,N_19680,N_19677);
xor U19815 (N_19815,N_19729,N_19756);
nor U19816 (N_19816,N_19602,N_19707);
or U19817 (N_19817,N_19732,N_19792);
xor U19818 (N_19818,N_19672,N_19739);
xor U19819 (N_19819,N_19644,N_19664);
nand U19820 (N_19820,N_19666,N_19721);
and U19821 (N_19821,N_19715,N_19787);
nand U19822 (N_19822,N_19788,N_19796);
or U19823 (N_19823,N_19712,N_19731);
nand U19824 (N_19824,N_19610,N_19765);
or U19825 (N_19825,N_19673,N_19709);
nand U19826 (N_19826,N_19654,N_19619);
nor U19827 (N_19827,N_19679,N_19606);
or U19828 (N_19828,N_19681,N_19773);
or U19829 (N_19829,N_19754,N_19725);
and U19830 (N_19830,N_19696,N_19762);
or U19831 (N_19831,N_19785,N_19704);
or U19832 (N_19832,N_19658,N_19710);
xnor U19833 (N_19833,N_19713,N_19662);
xor U19834 (N_19834,N_19612,N_19789);
xor U19835 (N_19835,N_19688,N_19651);
nand U19836 (N_19836,N_19698,N_19764);
or U19837 (N_19837,N_19791,N_19675);
xnor U19838 (N_19838,N_19608,N_19755);
nor U19839 (N_19839,N_19616,N_19699);
and U19840 (N_19840,N_19678,N_19659);
xnor U19841 (N_19841,N_19687,N_19682);
or U19842 (N_19842,N_19742,N_19601);
or U19843 (N_19843,N_19768,N_19617);
and U19844 (N_19844,N_19748,N_19660);
or U19845 (N_19845,N_19702,N_19634);
xnor U19846 (N_19846,N_19727,N_19652);
nor U19847 (N_19847,N_19717,N_19797);
nor U19848 (N_19848,N_19718,N_19719);
and U19849 (N_19849,N_19668,N_19649);
nand U19850 (N_19850,N_19670,N_19769);
nand U19851 (N_19851,N_19760,N_19629);
xor U19852 (N_19852,N_19604,N_19665);
nor U19853 (N_19853,N_19633,N_19741);
or U19854 (N_19854,N_19685,N_19663);
xnor U19855 (N_19855,N_19621,N_19605);
nor U19856 (N_19856,N_19761,N_19655);
and U19857 (N_19857,N_19744,N_19750);
and U19858 (N_19858,N_19671,N_19650);
nand U19859 (N_19859,N_19776,N_19734);
and U19860 (N_19860,N_19623,N_19642);
xnor U19861 (N_19861,N_19620,N_19700);
and U19862 (N_19862,N_19745,N_19692);
and U19863 (N_19863,N_19618,N_19694);
nor U19864 (N_19864,N_19758,N_19724);
and U19865 (N_19865,N_19701,N_19722);
and U19866 (N_19866,N_19674,N_19793);
xor U19867 (N_19867,N_19743,N_19798);
nor U19868 (N_19868,N_19600,N_19656);
or U19869 (N_19869,N_19638,N_19614);
xnor U19870 (N_19870,N_19622,N_19632);
or U19871 (N_19871,N_19630,N_19763);
and U19872 (N_19872,N_19609,N_19706);
or U19873 (N_19873,N_19770,N_19782);
or U19874 (N_19874,N_19708,N_19603);
or U19875 (N_19875,N_19799,N_19794);
nand U19876 (N_19876,N_19613,N_19777);
or U19877 (N_19877,N_19697,N_19667);
nor U19878 (N_19878,N_19705,N_19648);
or U19879 (N_19879,N_19780,N_19683);
nand U19880 (N_19880,N_19615,N_19736);
nor U19881 (N_19881,N_19627,N_19740);
nor U19882 (N_19882,N_19726,N_19626);
xor U19883 (N_19883,N_19781,N_19753);
or U19884 (N_19884,N_19786,N_19607);
and U19885 (N_19885,N_19695,N_19624);
and U19886 (N_19886,N_19636,N_19747);
nand U19887 (N_19887,N_19628,N_19749);
nand U19888 (N_19888,N_19771,N_19720);
xnor U19889 (N_19889,N_19641,N_19657);
nand U19890 (N_19890,N_19751,N_19661);
nand U19891 (N_19891,N_19779,N_19625);
nand U19892 (N_19892,N_19775,N_19778);
and U19893 (N_19893,N_19733,N_19637);
nand U19894 (N_19894,N_19737,N_19738);
or U19895 (N_19895,N_19689,N_19728);
nor U19896 (N_19896,N_19635,N_19714);
or U19897 (N_19897,N_19691,N_19723);
nor U19898 (N_19898,N_19676,N_19653);
or U19899 (N_19899,N_19631,N_19646);
and U19900 (N_19900,N_19769,N_19696);
xor U19901 (N_19901,N_19682,N_19773);
xnor U19902 (N_19902,N_19743,N_19754);
xor U19903 (N_19903,N_19724,N_19708);
xnor U19904 (N_19904,N_19704,N_19706);
and U19905 (N_19905,N_19605,N_19686);
nand U19906 (N_19906,N_19680,N_19643);
nand U19907 (N_19907,N_19714,N_19715);
nand U19908 (N_19908,N_19659,N_19673);
or U19909 (N_19909,N_19719,N_19742);
xor U19910 (N_19910,N_19607,N_19736);
xnor U19911 (N_19911,N_19798,N_19637);
or U19912 (N_19912,N_19676,N_19725);
nand U19913 (N_19913,N_19680,N_19637);
and U19914 (N_19914,N_19732,N_19662);
and U19915 (N_19915,N_19621,N_19796);
nor U19916 (N_19916,N_19722,N_19792);
nor U19917 (N_19917,N_19608,N_19796);
nor U19918 (N_19918,N_19701,N_19611);
and U19919 (N_19919,N_19762,N_19617);
or U19920 (N_19920,N_19799,N_19721);
or U19921 (N_19921,N_19763,N_19692);
or U19922 (N_19922,N_19616,N_19608);
or U19923 (N_19923,N_19758,N_19655);
xor U19924 (N_19924,N_19791,N_19744);
or U19925 (N_19925,N_19673,N_19735);
and U19926 (N_19926,N_19668,N_19759);
nand U19927 (N_19927,N_19723,N_19697);
or U19928 (N_19928,N_19702,N_19631);
or U19929 (N_19929,N_19656,N_19751);
xnor U19930 (N_19930,N_19779,N_19659);
or U19931 (N_19931,N_19666,N_19796);
or U19932 (N_19932,N_19695,N_19687);
nand U19933 (N_19933,N_19704,N_19771);
nor U19934 (N_19934,N_19773,N_19781);
xnor U19935 (N_19935,N_19634,N_19760);
and U19936 (N_19936,N_19723,N_19753);
and U19937 (N_19937,N_19729,N_19698);
and U19938 (N_19938,N_19626,N_19638);
and U19939 (N_19939,N_19644,N_19753);
nand U19940 (N_19940,N_19762,N_19639);
xor U19941 (N_19941,N_19606,N_19618);
and U19942 (N_19942,N_19611,N_19617);
and U19943 (N_19943,N_19776,N_19613);
xnor U19944 (N_19944,N_19716,N_19750);
xor U19945 (N_19945,N_19741,N_19688);
or U19946 (N_19946,N_19796,N_19717);
and U19947 (N_19947,N_19788,N_19687);
nand U19948 (N_19948,N_19712,N_19752);
nor U19949 (N_19949,N_19612,N_19737);
nand U19950 (N_19950,N_19766,N_19721);
or U19951 (N_19951,N_19775,N_19628);
xor U19952 (N_19952,N_19648,N_19678);
and U19953 (N_19953,N_19716,N_19673);
nor U19954 (N_19954,N_19661,N_19734);
nand U19955 (N_19955,N_19602,N_19740);
and U19956 (N_19956,N_19792,N_19640);
nor U19957 (N_19957,N_19702,N_19640);
and U19958 (N_19958,N_19643,N_19748);
and U19959 (N_19959,N_19612,N_19704);
xnor U19960 (N_19960,N_19627,N_19786);
and U19961 (N_19961,N_19620,N_19742);
or U19962 (N_19962,N_19743,N_19738);
nor U19963 (N_19963,N_19737,N_19661);
xor U19964 (N_19964,N_19658,N_19764);
nor U19965 (N_19965,N_19612,N_19604);
or U19966 (N_19966,N_19619,N_19791);
nor U19967 (N_19967,N_19758,N_19662);
nor U19968 (N_19968,N_19682,N_19723);
nor U19969 (N_19969,N_19667,N_19636);
and U19970 (N_19970,N_19623,N_19601);
and U19971 (N_19971,N_19792,N_19761);
nand U19972 (N_19972,N_19651,N_19650);
nor U19973 (N_19973,N_19744,N_19623);
nand U19974 (N_19974,N_19650,N_19737);
or U19975 (N_19975,N_19707,N_19672);
and U19976 (N_19976,N_19714,N_19756);
nor U19977 (N_19977,N_19695,N_19794);
nor U19978 (N_19978,N_19785,N_19747);
nand U19979 (N_19979,N_19683,N_19705);
or U19980 (N_19980,N_19716,N_19780);
and U19981 (N_19981,N_19686,N_19642);
or U19982 (N_19982,N_19626,N_19609);
or U19983 (N_19983,N_19717,N_19766);
nand U19984 (N_19984,N_19632,N_19664);
or U19985 (N_19985,N_19766,N_19768);
nor U19986 (N_19986,N_19611,N_19719);
nor U19987 (N_19987,N_19743,N_19735);
nor U19988 (N_19988,N_19704,N_19662);
xor U19989 (N_19989,N_19790,N_19760);
xnor U19990 (N_19990,N_19725,N_19621);
xor U19991 (N_19991,N_19660,N_19755);
or U19992 (N_19992,N_19669,N_19787);
nor U19993 (N_19993,N_19618,N_19743);
nand U19994 (N_19994,N_19703,N_19610);
xor U19995 (N_19995,N_19798,N_19751);
or U19996 (N_19996,N_19722,N_19726);
nor U19997 (N_19997,N_19784,N_19612);
xnor U19998 (N_19998,N_19662,N_19641);
or U19999 (N_19999,N_19731,N_19686);
nand U20000 (N_20000,N_19907,N_19816);
or U20001 (N_20001,N_19857,N_19882);
xor U20002 (N_20002,N_19993,N_19910);
nor U20003 (N_20003,N_19871,N_19976);
and U20004 (N_20004,N_19820,N_19999);
and U20005 (N_20005,N_19988,N_19879);
nand U20006 (N_20006,N_19945,N_19918);
nor U20007 (N_20007,N_19893,N_19962);
nor U20008 (N_20008,N_19883,N_19942);
xor U20009 (N_20009,N_19828,N_19866);
nor U20010 (N_20010,N_19905,N_19824);
nor U20011 (N_20011,N_19951,N_19902);
and U20012 (N_20012,N_19899,N_19880);
nand U20013 (N_20013,N_19920,N_19849);
or U20014 (N_20014,N_19870,N_19914);
nand U20015 (N_20015,N_19888,N_19844);
and U20016 (N_20016,N_19830,N_19854);
nand U20017 (N_20017,N_19843,N_19821);
xor U20018 (N_20018,N_19968,N_19935);
xor U20019 (N_20019,N_19904,N_19929);
nand U20020 (N_20020,N_19877,N_19847);
or U20021 (N_20021,N_19803,N_19874);
xnor U20022 (N_20022,N_19994,N_19878);
and U20023 (N_20023,N_19832,N_19991);
nor U20024 (N_20024,N_19977,N_19833);
nand U20025 (N_20025,N_19919,N_19851);
or U20026 (N_20026,N_19875,N_19979);
nor U20027 (N_20027,N_19971,N_19808);
nand U20028 (N_20028,N_19890,N_19986);
nor U20029 (N_20029,N_19841,N_19804);
xnor U20030 (N_20030,N_19855,N_19826);
and U20031 (N_20031,N_19923,N_19809);
and U20032 (N_20032,N_19838,N_19831);
nor U20033 (N_20033,N_19806,N_19970);
nand U20034 (N_20034,N_19961,N_19944);
or U20035 (N_20035,N_19811,N_19934);
xor U20036 (N_20036,N_19865,N_19925);
nand U20037 (N_20037,N_19872,N_19852);
xor U20038 (N_20038,N_19800,N_19895);
xnor U20039 (N_20039,N_19818,N_19814);
and U20040 (N_20040,N_19949,N_19867);
or U20041 (N_20041,N_19903,N_19959);
or U20042 (N_20042,N_19958,N_19813);
nand U20043 (N_20043,N_19829,N_19954);
or U20044 (N_20044,N_19965,N_19881);
or U20045 (N_20045,N_19996,N_19840);
nand U20046 (N_20046,N_19807,N_19916);
or U20047 (N_20047,N_19887,N_19896);
xnor U20048 (N_20048,N_19969,N_19836);
nand U20049 (N_20049,N_19839,N_19931);
or U20050 (N_20050,N_19897,N_19846);
xnor U20051 (N_20051,N_19964,N_19876);
nor U20052 (N_20052,N_19859,N_19848);
nand U20053 (N_20053,N_19911,N_19805);
nor U20054 (N_20054,N_19909,N_19823);
and U20055 (N_20055,N_19884,N_19952);
and U20056 (N_20056,N_19819,N_19930);
and U20057 (N_20057,N_19898,N_19963);
and U20058 (N_20058,N_19981,N_19978);
nor U20059 (N_20059,N_19984,N_19936);
nand U20060 (N_20060,N_19975,N_19802);
or U20061 (N_20061,N_19869,N_19982);
and U20062 (N_20062,N_19927,N_19926);
nand U20063 (N_20063,N_19815,N_19928);
nand U20064 (N_20064,N_19932,N_19860);
nand U20065 (N_20065,N_19987,N_19983);
and U20066 (N_20066,N_19825,N_19998);
and U20067 (N_20067,N_19992,N_19889);
xor U20068 (N_20068,N_19924,N_19845);
or U20069 (N_20069,N_19853,N_19812);
nand U20070 (N_20070,N_19834,N_19900);
and U20071 (N_20071,N_19915,N_19908);
or U20072 (N_20072,N_19972,N_19950);
nand U20073 (N_20073,N_19891,N_19901);
xnor U20074 (N_20074,N_19973,N_19817);
or U20075 (N_20075,N_19933,N_19985);
or U20076 (N_20076,N_19941,N_19940);
nor U20077 (N_20077,N_19939,N_19921);
or U20078 (N_20078,N_19906,N_19892);
and U20079 (N_20079,N_19912,N_19948);
nand U20080 (N_20080,N_19864,N_19980);
nand U20081 (N_20081,N_19997,N_19863);
and U20082 (N_20082,N_19885,N_19947);
xnor U20083 (N_20083,N_19810,N_19917);
nor U20084 (N_20084,N_19956,N_19827);
nor U20085 (N_20085,N_19967,N_19913);
and U20086 (N_20086,N_19937,N_19966);
nor U20087 (N_20087,N_19955,N_19850);
xnor U20088 (N_20088,N_19873,N_19953);
and U20089 (N_20089,N_19943,N_19960);
or U20090 (N_20090,N_19995,N_19974);
nand U20091 (N_20091,N_19835,N_19922);
nand U20092 (N_20092,N_19990,N_19862);
nor U20093 (N_20093,N_19957,N_19894);
nor U20094 (N_20094,N_19858,N_19856);
xnor U20095 (N_20095,N_19938,N_19861);
nand U20096 (N_20096,N_19886,N_19837);
nand U20097 (N_20097,N_19842,N_19801);
or U20098 (N_20098,N_19822,N_19946);
nor U20099 (N_20099,N_19868,N_19989);
and U20100 (N_20100,N_19815,N_19805);
or U20101 (N_20101,N_19862,N_19857);
xnor U20102 (N_20102,N_19895,N_19954);
nor U20103 (N_20103,N_19807,N_19981);
xnor U20104 (N_20104,N_19820,N_19804);
xnor U20105 (N_20105,N_19914,N_19954);
nor U20106 (N_20106,N_19917,N_19833);
and U20107 (N_20107,N_19855,N_19930);
and U20108 (N_20108,N_19903,N_19873);
xor U20109 (N_20109,N_19825,N_19964);
nor U20110 (N_20110,N_19813,N_19994);
xnor U20111 (N_20111,N_19865,N_19854);
xnor U20112 (N_20112,N_19968,N_19923);
nor U20113 (N_20113,N_19986,N_19848);
xor U20114 (N_20114,N_19804,N_19985);
xor U20115 (N_20115,N_19943,N_19846);
or U20116 (N_20116,N_19997,N_19860);
nor U20117 (N_20117,N_19847,N_19917);
nor U20118 (N_20118,N_19975,N_19973);
and U20119 (N_20119,N_19996,N_19804);
nor U20120 (N_20120,N_19970,N_19987);
nor U20121 (N_20121,N_19979,N_19876);
and U20122 (N_20122,N_19880,N_19836);
nor U20123 (N_20123,N_19928,N_19975);
nand U20124 (N_20124,N_19928,N_19922);
and U20125 (N_20125,N_19842,N_19803);
xor U20126 (N_20126,N_19917,N_19950);
and U20127 (N_20127,N_19935,N_19855);
and U20128 (N_20128,N_19858,N_19974);
and U20129 (N_20129,N_19824,N_19979);
and U20130 (N_20130,N_19830,N_19855);
xnor U20131 (N_20131,N_19949,N_19865);
and U20132 (N_20132,N_19821,N_19834);
and U20133 (N_20133,N_19986,N_19817);
xor U20134 (N_20134,N_19982,N_19898);
or U20135 (N_20135,N_19891,N_19815);
xor U20136 (N_20136,N_19958,N_19876);
xnor U20137 (N_20137,N_19946,N_19986);
nor U20138 (N_20138,N_19980,N_19935);
nand U20139 (N_20139,N_19817,N_19908);
xor U20140 (N_20140,N_19858,N_19829);
or U20141 (N_20141,N_19813,N_19822);
and U20142 (N_20142,N_19853,N_19872);
xor U20143 (N_20143,N_19874,N_19804);
nor U20144 (N_20144,N_19939,N_19801);
xnor U20145 (N_20145,N_19829,N_19876);
nand U20146 (N_20146,N_19956,N_19859);
and U20147 (N_20147,N_19840,N_19866);
nand U20148 (N_20148,N_19891,N_19869);
nand U20149 (N_20149,N_19833,N_19966);
nor U20150 (N_20150,N_19899,N_19920);
nand U20151 (N_20151,N_19922,N_19862);
nand U20152 (N_20152,N_19981,N_19918);
and U20153 (N_20153,N_19853,N_19948);
and U20154 (N_20154,N_19906,N_19809);
and U20155 (N_20155,N_19933,N_19826);
and U20156 (N_20156,N_19840,N_19862);
xor U20157 (N_20157,N_19903,N_19802);
or U20158 (N_20158,N_19846,N_19884);
xor U20159 (N_20159,N_19976,N_19808);
xnor U20160 (N_20160,N_19836,N_19999);
xor U20161 (N_20161,N_19971,N_19868);
nor U20162 (N_20162,N_19970,N_19977);
nand U20163 (N_20163,N_19883,N_19852);
xnor U20164 (N_20164,N_19965,N_19980);
nand U20165 (N_20165,N_19858,N_19836);
and U20166 (N_20166,N_19889,N_19932);
nor U20167 (N_20167,N_19965,N_19897);
nor U20168 (N_20168,N_19944,N_19804);
nor U20169 (N_20169,N_19886,N_19902);
or U20170 (N_20170,N_19865,N_19814);
xor U20171 (N_20171,N_19851,N_19829);
or U20172 (N_20172,N_19901,N_19807);
and U20173 (N_20173,N_19935,N_19880);
xnor U20174 (N_20174,N_19945,N_19806);
nor U20175 (N_20175,N_19969,N_19938);
nand U20176 (N_20176,N_19869,N_19830);
and U20177 (N_20177,N_19944,N_19936);
and U20178 (N_20178,N_19973,N_19824);
nor U20179 (N_20179,N_19982,N_19845);
nor U20180 (N_20180,N_19824,N_19953);
xor U20181 (N_20181,N_19977,N_19972);
nor U20182 (N_20182,N_19976,N_19946);
or U20183 (N_20183,N_19804,N_19819);
xnor U20184 (N_20184,N_19846,N_19847);
or U20185 (N_20185,N_19931,N_19916);
nand U20186 (N_20186,N_19952,N_19916);
and U20187 (N_20187,N_19952,N_19959);
nand U20188 (N_20188,N_19888,N_19980);
xor U20189 (N_20189,N_19994,N_19984);
xnor U20190 (N_20190,N_19956,N_19906);
nor U20191 (N_20191,N_19851,N_19990);
or U20192 (N_20192,N_19821,N_19825);
nor U20193 (N_20193,N_19874,N_19907);
nor U20194 (N_20194,N_19983,N_19818);
nor U20195 (N_20195,N_19888,N_19891);
xor U20196 (N_20196,N_19884,N_19906);
or U20197 (N_20197,N_19976,N_19819);
or U20198 (N_20198,N_19930,N_19926);
or U20199 (N_20199,N_19890,N_19848);
nand U20200 (N_20200,N_20130,N_20084);
and U20201 (N_20201,N_20060,N_20108);
nor U20202 (N_20202,N_20137,N_20182);
or U20203 (N_20203,N_20165,N_20090);
nand U20204 (N_20204,N_20076,N_20194);
or U20205 (N_20205,N_20107,N_20074);
nand U20206 (N_20206,N_20038,N_20007);
nor U20207 (N_20207,N_20135,N_20131);
and U20208 (N_20208,N_20173,N_20013);
and U20209 (N_20209,N_20197,N_20053);
and U20210 (N_20210,N_20061,N_20187);
nor U20211 (N_20211,N_20099,N_20039);
and U20212 (N_20212,N_20155,N_20158);
and U20213 (N_20213,N_20044,N_20123);
or U20214 (N_20214,N_20035,N_20014);
and U20215 (N_20215,N_20188,N_20047);
nor U20216 (N_20216,N_20032,N_20012);
xor U20217 (N_20217,N_20140,N_20078);
or U20218 (N_20218,N_20015,N_20120);
or U20219 (N_20219,N_20069,N_20113);
and U20220 (N_20220,N_20098,N_20095);
nand U20221 (N_20221,N_20093,N_20126);
nand U20222 (N_20222,N_20055,N_20059);
or U20223 (N_20223,N_20091,N_20097);
nor U20224 (N_20224,N_20104,N_20116);
nor U20225 (N_20225,N_20148,N_20161);
and U20226 (N_20226,N_20086,N_20077);
or U20227 (N_20227,N_20021,N_20138);
and U20228 (N_20228,N_20017,N_20178);
nor U20229 (N_20229,N_20167,N_20189);
nor U20230 (N_20230,N_20191,N_20185);
nand U20231 (N_20231,N_20036,N_20141);
nand U20232 (N_20232,N_20081,N_20163);
and U20233 (N_20233,N_20087,N_20043);
and U20234 (N_20234,N_20029,N_20121);
nand U20235 (N_20235,N_20162,N_20005);
and U20236 (N_20236,N_20171,N_20106);
or U20237 (N_20237,N_20070,N_20100);
nand U20238 (N_20238,N_20139,N_20147);
nand U20239 (N_20239,N_20125,N_20124);
xnor U20240 (N_20240,N_20033,N_20159);
and U20241 (N_20241,N_20096,N_20192);
and U20242 (N_20242,N_20050,N_20134);
nor U20243 (N_20243,N_20152,N_20127);
or U20244 (N_20244,N_20048,N_20118);
nor U20245 (N_20245,N_20068,N_20057);
nor U20246 (N_20246,N_20199,N_20198);
xor U20247 (N_20247,N_20105,N_20051);
or U20248 (N_20248,N_20071,N_20008);
or U20249 (N_20249,N_20072,N_20002);
nor U20250 (N_20250,N_20164,N_20063);
nor U20251 (N_20251,N_20018,N_20000);
or U20252 (N_20252,N_20174,N_20157);
and U20253 (N_20253,N_20114,N_20058);
xnor U20254 (N_20254,N_20042,N_20101);
and U20255 (N_20255,N_20085,N_20009);
xor U20256 (N_20256,N_20196,N_20146);
nand U20257 (N_20257,N_20089,N_20031);
nand U20258 (N_20258,N_20102,N_20016);
nand U20259 (N_20259,N_20142,N_20064);
nor U20260 (N_20260,N_20150,N_20103);
and U20261 (N_20261,N_20186,N_20094);
and U20262 (N_20262,N_20169,N_20193);
nor U20263 (N_20263,N_20056,N_20166);
xnor U20264 (N_20264,N_20129,N_20181);
xor U20265 (N_20265,N_20062,N_20082);
or U20266 (N_20266,N_20195,N_20046);
nand U20267 (N_20267,N_20092,N_20179);
and U20268 (N_20268,N_20175,N_20170);
or U20269 (N_20269,N_20168,N_20001);
or U20270 (N_20270,N_20144,N_20119);
or U20271 (N_20271,N_20019,N_20034);
nor U20272 (N_20272,N_20022,N_20011);
nor U20273 (N_20273,N_20075,N_20025);
and U20274 (N_20274,N_20183,N_20024);
nor U20275 (N_20275,N_20117,N_20037);
nand U20276 (N_20276,N_20052,N_20066);
nor U20277 (N_20277,N_20023,N_20111);
nand U20278 (N_20278,N_20045,N_20115);
or U20279 (N_20279,N_20030,N_20020);
xnor U20280 (N_20280,N_20112,N_20176);
and U20281 (N_20281,N_20190,N_20133);
nor U20282 (N_20282,N_20177,N_20128);
or U20283 (N_20283,N_20079,N_20028);
xnor U20284 (N_20284,N_20088,N_20172);
nor U20285 (N_20285,N_20080,N_20083);
nor U20286 (N_20286,N_20004,N_20145);
nand U20287 (N_20287,N_20040,N_20132);
and U20288 (N_20288,N_20026,N_20153);
nand U20289 (N_20289,N_20122,N_20151);
xor U20290 (N_20290,N_20003,N_20109);
and U20291 (N_20291,N_20027,N_20149);
nand U20292 (N_20292,N_20110,N_20067);
xnor U20293 (N_20293,N_20049,N_20143);
nor U20294 (N_20294,N_20154,N_20156);
or U20295 (N_20295,N_20184,N_20065);
nor U20296 (N_20296,N_20054,N_20041);
nor U20297 (N_20297,N_20073,N_20010);
nor U20298 (N_20298,N_20180,N_20136);
nand U20299 (N_20299,N_20160,N_20006);
nor U20300 (N_20300,N_20090,N_20091);
xor U20301 (N_20301,N_20071,N_20110);
and U20302 (N_20302,N_20051,N_20008);
or U20303 (N_20303,N_20011,N_20117);
and U20304 (N_20304,N_20087,N_20105);
xor U20305 (N_20305,N_20186,N_20130);
nor U20306 (N_20306,N_20137,N_20051);
xnor U20307 (N_20307,N_20138,N_20192);
xnor U20308 (N_20308,N_20018,N_20109);
or U20309 (N_20309,N_20180,N_20137);
and U20310 (N_20310,N_20043,N_20106);
nor U20311 (N_20311,N_20024,N_20027);
or U20312 (N_20312,N_20011,N_20163);
nor U20313 (N_20313,N_20188,N_20066);
or U20314 (N_20314,N_20177,N_20032);
nand U20315 (N_20315,N_20002,N_20151);
xnor U20316 (N_20316,N_20023,N_20083);
or U20317 (N_20317,N_20167,N_20186);
nor U20318 (N_20318,N_20099,N_20104);
nor U20319 (N_20319,N_20111,N_20177);
nand U20320 (N_20320,N_20117,N_20102);
and U20321 (N_20321,N_20138,N_20189);
xor U20322 (N_20322,N_20038,N_20148);
nor U20323 (N_20323,N_20078,N_20151);
nand U20324 (N_20324,N_20144,N_20028);
xor U20325 (N_20325,N_20074,N_20094);
xnor U20326 (N_20326,N_20139,N_20122);
or U20327 (N_20327,N_20009,N_20016);
xor U20328 (N_20328,N_20140,N_20014);
and U20329 (N_20329,N_20035,N_20156);
nand U20330 (N_20330,N_20103,N_20174);
and U20331 (N_20331,N_20005,N_20170);
nand U20332 (N_20332,N_20135,N_20150);
nor U20333 (N_20333,N_20095,N_20039);
nand U20334 (N_20334,N_20187,N_20058);
and U20335 (N_20335,N_20065,N_20116);
or U20336 (N_20336,N_20029,N_20179);
or U20337 (N_20337,N_20026,N_20075);
nand U20338 (N_20338,N_20182,N_20149);
xor U20339 (N_20339,N_20027,N_20196);
xor U20340 (N_20340,N_20177,N_20194);
nand U20341 (N_20341,N_20191,N_20120);
nor U20342 (N_20342,N_20039,N_20016);
nand U20343 (N_20343,N_20162,N_20188);
nor U20344 (N_20344,N_20100,N_20161);
nand U20345 (N_20345,N_20002,N_20099);
or U20346 (N_20346,N_20123,N_20197);
nand U20347 (N_20347,N_20044,N_20101);
and U20348 (N_20348,N_20037,N_20047);
xor U20349 (N_20349,N_20110,N_20163);
xor U20350 (N_20350,N_20139,N_20150);
nor U20351 (N_20351,N_20074,N_20166);
or U20352 (N_20352,N_20035,N_20095);
nor U20353 (N_20353,N_20099,N_20161);
xor U20354 (N_20354,N_20114,N_20003);
xor U20355 (N_20355,N_20114,N_20175);
or U20356 (N_20356,N_20040,N_20022);
nand U20357 (N_20357,N_20155,N_20080);
and U20358 (N_20358,N_20075,N_20137);
and U20359 (N_20359,N_20090,N_20197);
nor U20360 (N_20360,N_20096,N_20126);
nand U20361 (N_20361,N_20153,N_20067);
and U20362 (N_20362,N_20080,N_20068);
or U20363 (N_20363,N_20085,N_20093);
nor U20364 (N_20364,N_20121,N_20015);
or U20365 (N_20365,N_20005,N_20168);
nor U20366 (N_20366,N_20044,N_20136);
nor U20367 (N_20367,N_20151,N_20071);
and U20368 (N_20368,N_20021,N_20066);
or U20369 (N_20369,N_20044,N_20197);
nor U20370 (N_20370,N_20070,N_20172);
nand U20371 (N_20371,N_20125,N_20156);
or U20372 (N_20372,N_20104,N_20136);
and U20373 (N_20373,N_20124,N_20082);
nand U20374 (N_20374,N_20109,N_20095);
xor U20375 (N_20375,N_20027,N_20056);
nor U20376 (N_20376,N_20077,N_20045);
nand U20377 (N_20377,N_20171,N_20121);
nand U20378 (N_20378,N_20031,N_20088);
and U20379 (N_20379,N_20046,N_20124);
nand U20380 (N_20380,N_20062,N_20096);
and U20381 (N_20381,N_20068,N_20130);
nor U20382 (N_20382,N_20011,N_20080);
nor U20383 (N_20383,N_20152,N_20027);
and U20384 (N_20384,N_20087,N_20086);
nor U20385 (N_20385,N_20083,N_20043);
xor U20386 (N_20386,N_20045,N_20078);
or U20387 (N_20387,N_20048,N_20079);
xnor U20388 (N_20388,N_20139,N_20195);
nor U20389 (N_20389,N_20044,N_20098);
nor U20390 (N_20390,N_20079,N_20042);
nand U20391 (N_20391,N_20020,N_20079);
and U20392 (N_20392,N_20065,N_20132);
or U20393 (N_20393,N_20163,N_20187);
nand U20394 (N_20394,N_20150,N_20093);
xnor U20395 (N_20395,N_20030,N_20101);
nor U20396 (N_20396,N_20084,N_20043);
nor U20397 (N_20397,N_20000,N_20111);
nand U20398 (N_20398,N_20100,N_20113);
and U20399 (N_20399,N_20142,N_20103);
xor U20400 (N_20400,N_20289,N_20387);
nand U20401 (N_20401,N_20276,N_20321);
and U20402 (N_20402,N_20334,N_20281);
nand U20403 (N_20403,N_20298,N_20234);
or U20404 (N_20404,N_20242,N_20355);
nand U20405 (N_20405,N_20279,N_20274);
xnor U20406 (N_20406,N_20288,N_20314);
and U20407 (N_20407,N_20297,N_20383);
or U20408 (N_20408,N_20358,N_20285);
or U20409 (N_20409,N_20398,N_20206);
nor U20410 (N_20410,N_20397,N_20339);
nor U20411 (N_20411,N_20213,N_20301);
xnor U20412 (N_20412,N_20336,N_20230);
and U20413 (N_20413,N_20233,N_20311);
nor U20414 (N_20414,N_20286,N_20280);
nand U20415 (N_20415,N_20265,N_20259);
or U20416 (N_20416,N_20377,N_20203);
nor U20417 (N_20417,N_20248,N_20337);
xor U20418 (N_20418,N_20241,N_20293);
nor U20419 (N_20419,N_20340,N_20344);
nor U20420 (N_20420,N_20369,N_20226);
or U20421 (N_20421,N_20390,N_20367);
nand U20422 (N_20422,N_20375,N_20341);
or U20423 (N_20423,N_20238,N_20331);
nand U20424 (N_20424,N_20356,N_20245);
or U20425 (N_20425,N_20309,N_20345);
nand U20426 (N_20426,N_20218,N_20296);
or U20427 (N_20427,N_20262,N_20216);
xor U20428 (N_20428,N_20389,N_20227);
or U20429 (N_20429,N_20214,N_20335);
nor U20430 (N_20430,N_20256,N_20329);
and U20431 (N_20431,N_20254,N_20243);
and U20432 (N_20432,N_20208,N_20350);
and U20433 (N_20433,N_20332,N_20222);
nor U20434 (N_20434,N_20361,N_20205);
and U20435 (N_20435,N_20394,N_20300);
nor U20436 (N_20436,N_20210,N_20231);
xnor U20437 (N_20437,N_20257,N_20326);
nand U20438 (N_20438,N_20235,N_20362);
nor U20439 (N_20439,N_20322,N_20373);
nand U20440 (N_20440,N_20221,N_20328);
nor U20441 (N_20441,N_20302,N_20215);
xnor U20442 (N_20442,N_20284,N_20273);
nor U20443 (N_20443,N_20207,N_20278);
nand U20444 (N_20444,N_20385,N_20201);
and U20445 (N_20445,N_20323,N_20357);
xnor U20446 (N_20446,N_20379,N_20232);
nand U20447 (N_20447,N_20342,N_20371);
nor U20448 (N_20448,N_20204,N_20384);
xnor U20449 (N_20449,N_20354,N_20224);
and U20450 (N_20450,N_20312,N_20366);
and U20451 (N_20451,N_20212,N_20292);
nand U20452 (N_20452,N_20351,N_20391);
nor U20453 (N_20453,N_20343,N_20318);
and U20454 (N_20454,N_20381,N_20395);
nor U20455 (N_20455,N_20378,N_20277);
or U20456 (N_20456,N_20290,N_20299);
nor U20457 (N_20457,N_20319,N_20347);
nor U20458 (N_20458,N_20255,N_20229);
or U20459 (N_20459,N_20368,N_20223);
or U20460 (N_20460,N_20236,N_20388);
nor U20461 (N_20461,N_20310,N_20399);
or U20462 (N_20462,N_20303,N_20266);
or U20463 (N_20463,N_20209,N_20220);
and U20464 (N_20464,N_20240,N_20264);
nor U20465 (N_20465,N_20225,N_20338);
or U20466 (N_20466,N_20320,N_20386);
or U20467 (N_20467,N_20370,N_20305);
or U20468 (N_20468,N_20268,N_20348);
or U20469 (N_20469,N_20380,N_20315);
nor U20470 (N_20470,N_20237,N_20219);
nor U20471 (N_20471,N_20267,N_20324);
nor U20472 (N_20472,N_20271,N_20396);
and U20473 (N_20473,N_20275,N_20252);
nor U20474 (N_20474,N_20392,N_20202);
nand U20475 (N_20475,N_20250,N_20200);
and U20476 (N_20476,N_20349,N_20333);
xnor U20477 (N_20477,N_20249,N_20247);
xor U20478 (N_20478,N_20294,N_20263);
and U20479 (N_20479,N_20359,N_20270);
nor U20480 (N_20480,N_20327,N_20393);
or U20481 (N_20481,N_20376,N_20295);
nand U20482 (N_20482,N_20346,N_20283);
and U20483 (N_20483,N_20360,N_20306);
nand U20484 (N_20484,N_20282,N_20253);
or U20485 (N_20485,N_20217,N_20304);
nand U20486 (N_20486,N_20269,N_20260);
or U20487 (N_20487,N_20372,N_20251);
and U20488 (N_20488,N_20244,N_20364);
xnor U20489 (N_20489,N_20374,N_20239);
or U20490 (N_20490,N_20308,N_20330);
or U20491 (N_20491,N_20365,N_20352);
and U20492 (N_20492,N_20317,N_20291);
nand U20493 (N_20493,N_20211,N_20313);
xnor U20494 (N_20494,N_20353,N_20316);
and U20495 (N_20495,N_20258,N_20287);
or U20496 (N_20496,N_20382,N_20228);
and U20497 (N_20497,N_20307,N_20325);
or U20498 (N_20498,N_20363,N_20261);
and U20499 (N_20499,N_20246,N_20272);
nor U20500 (N_20500,N_20206,N_20296);
nor U20501 (N_20501,N_20263,N_20392);
xor U20502 (N_20502,N_20262,N_20388);
or U20503 (N_20503,N_20268,N_20282);
nor U20504 (N_20504,N_20393,N_20376);
nor U20505 (N_20505,N_20272,N_20398);
nand U20506 (N_20506,N_20321,N_20217);
or U20507 (N_20507,N_20255,N_20345);
and U20508 (N_20508,N_20276,N_20203);
and U20509 (N_20509,N_20356,N_20386);
nor U20510 (N_20510,N_20249,N_20291);
and U20511 (N_20511,N_20338,N_20208);
or U20512 (N_20512,N_20203,N_20353);
xnor U20513 (N_20513,N_20328,N_20237);
and U20514 (N_20514,N_20263,N_20212);
nor U20515 (N_20515,N_20363,N_20321);
xor U20516 (N_20516,N_20330,N_20275);
nand U20517 (N_20517,N_20373,N_20286);
nor U20518 (N_20518,N_20377,N_20336);
nand U20519 (N_20519,N_20379,N_20380);
nor U20520 (N_20520,N_20243,N_20354);
nand U20521 (N_20521,N_20268,N_20275);
nand U20522 (N_20522,N_20348,N_20308);
xnor U20523 (N_20523,N_20325,N_20227);
nor U20524 (N_20524,N_20375,N_20378);
xor U20525 (N_20525,N_20362,N_20365);
or U20526 (N_20526,N_20380,N_20287);
nor U20527 (N_20527,N_20213,N_20285);
nor U20528 (N_20528,N_20395,N_20287);
xor U20529 (N_20529,N_20366,N_20300);
nor U20530 (N_20530,N_20225,N_20295);
and U20531 (N_20531,N_20235,N_20221);
and U20532 (N_20532,N_20287,N_20307);
xor U20533 (N_20533,N_20265,N_20209);
xor U20534 (N_20534,N_20203,N_20242);
nand U20535 (N_20535,N_20287,N_20232);
xor U20536 (N_20536,N_20306,N_20357);
xnor U20537 (N_20537,N_20394,N_20208);
or U20538 (N_20538,N_20227,N_20321);
nor U20539 (N_20539,N_20364,N_20311);
nand U20540 (N_20540,N_20352,N_20341);
or U20541 (N_20541,N_20293,N_20371);
nor U20542 (N_20542,N_20276,N_20274);
xnor U20543 (N_20543,N_20270,N_20282);
and U20544 (N_20544,N_20368,N_20208);
nand U20545 (N_20545,N_20352,N_20362);
xor U20546 (N_20546,N_20300,N_20281);
or U20547 (N_20547,N_20211,N_20212);
xnor U20548 (N_20548,N_20387,N_20332);
and U20549 (N_20549,N_20389,N_20378);
nand U20550 (N_20550,N_20244,N_20351);
xor U20551 (N_20551,N_20254,N_20287);
nor U20552 (N_20552,N_20393,N_20273);
nand U20553 (N_20553,N_20302,N_20243);
or U20554 (N_20554,N_20306,N_20230);
xor U20555 (N_20555,N_20263,N_20282);
and U20556 (N_20556,N_20333,N_20202);
and U20557 (N_20557,N_20205,N_20359);
xnor U20558 (N_20558,N_20270,N_20219);
nor U20559 (N_20559,N_20308,N_20214);
xor U20560 (N_20560,N_20301,N_20256);
nor U20561 (N_20561,N_20337,N_20300);
xnor U20562 (N_20562,N_20313,N_20236);
nand U20563 (N_20563,N_20303,N_20383);
nand U20564 (N_20564,N_20396,N_20373);
nand U20565 (N_20565,N_20257,N_20378);
xnor U20566 (N_20566,N_20312,N_20219);
xor U20567 (N_20567,N_20332,N_20361);
xor U20568 (N_20568,N_20296,N_20318);
nand U20569 (N_20569,N_20325,N_20372);
and U20570 (N_20570,N_20292,N_20203);
xnor U20571 (N_20571,N_20303,N_20364);
or U20572 (N_20572,N_20293,N_20286);
nor U20573 (N_20573,N_20310,N_20215);
or U20574 (N_20574,N_20287,N_20387);
or U20575 (N_20575,N_20398,N_20302);
or U20576 (N_20576,N_20260,N_20279);
nand U20577 (N_20577,N_20233,N_20399);
nor U20578 (N_20578,N_20230,N_20255);
nor U20579 (N_20579,N_20233,N_20345);
or U20580 (N_20580,N_20242,N_20267);
nor U20581 (N_20581,N_20252,N_20295);
nor U20582 (N_20582,N_20383,N_20277);
or U20583 (N_20583,N_20250,N_20317);
nand U20584 (N_20584,N_20211,N_20319);
and U20585 (N_20585,N_20244,N_20324);
xnor U20586 (N_20586,N_20343,N_20333);
and U20587 (N_20587,N_20270,N_20231);
nand U20588 (N_20588,N_20237,N_20379);
nor U20589 (N_20589,N_20263,N_20235);
nor U20590 (N_20590,N_20303,N_20290);
nand U20591 (N_20591,N_20385,N_20316);
xor U20592 (N_20592,N_20255,N_20304);
nand U20593 (N_20593,N_20380,N_20290);
xnor U20594 (N_20594,N_20355,N_20276);
or U20595 (N_20595,N_20363,N_20380);
xnor U20596 (N_20596,N_20393,N_20231);
nor U20597 (N_20597,N_20255,N_20338);
or U20598 (N_20598,N_20240,N_20226);
nor U20599 (N_20599,N_20341,N_20357);
and U20600 (N_20600,N_20430,N_20400);
xnor U20601 (N_20601,N_20482,N_20544);
xor U20602 (N_20602,N_20407,N_20418);
nor U20603 (N_20603,N_20467,N_20556);
nand U20604 (N_20604,N_20554,N_20420);
and U20605 (N_20605,N_20582,N_20589);
nor U20606 (N_20606,N_20532,N_20486);
or U20607 (N_20607,N_20452,N_20475);
nor U20608 (N_20608,N_20523,N_20565);
nand U20609 (N_20609,N_20503,N_20599);
or U20610 (N_20610,N_20485,N_20542);
nand U20611 (N_20611,N_20562,N_20449);
nor U20612 (N_20612,N_20598,N_20447);
nor U20613 (N_20613,N_20591,N_20442);
nor U20614 (N_20614,N_20538,N_20581);
or U20615 (N_20615,N_20553,N_20497);
nand U20616 (N_20616,N_20507,N_20463);
xnor U20617 (N_20617,N_20477,N_20585);
or U20618 (N_20618,N_20517,N_20576);
or U20619 (N_20619,N_20437,N_20483);
nor U20620 (N_20620,N_20406,N_20525);
or U20621 (N_20621,N_20559,N_20519);
and U20622 (N_20622,N_20469,N_20533);
nand U20623 (N_20623,N_20550,N_20416);
nor U20624 (N_20624,N_20411,N_20560);
or U20625 (N_20625,N_20530,N_20410);
nor U20626 (N_20626,N_20403,N_20462);
nor U20627 (N_20627,N_20505,N_20439);
nor U20628 (N_20628,N_20425,N_20487);
nand U20629 (N_20629,N_20458,N_20588);
or U20630 (N_20630,N_20408,N_20541);
and U20631 (N_20631,N_20595,N_20453);
nor U20632 (N_20632,N_20522,N_20568);
or U20633 (N_20633,N_20584,N_20432);
nor U20634 (N_20634,N_20413,N_20521);
nand U20635 (N_20635,N_20501,N_20441);
and U20636 (N_20636,N_20490,N_20514);
nor U20637 (N_20637,N_20428,N_20566);
or U20638 (N_20638,N_20529,N_20421);
or U20639 (N_20639,N_20578,N_20459);
and U20640 (N_20640,N_20548,N_20540);
nand U20641 (N_20641,N_20417,N_20551);
or U20642 (N_20642,N_20579,N_20510);
and U20643 (N_20643,N_20431,N_20474);
and U20644 (N_20644,N_20572,N_20440);
or U20645 (N_20645,N_20434,N_20549);
nand U20646 (N_20646,N_20488,N_20456);
xnor U20647 (N_20647,N_20423,N_20518);
nand U20648 (N_20648,N_20546,N_20583);
xor U20649 (N_20649,N_20448,N_20569);
nand U20650 (N_20650,N_20481,N_20586);
xnor U20651 (N_20651,N_20573,N_20444);
nor U20652 (N_20652,N_20552,N_20446);
xor U20653 (N_20653,N_20470,N_20593);
nand U20654 (N_20654,N_20401,N_20454);
nor U20655 (N_20655,N_20433,N_20405);
nor U20656 (N_20656,N_20478,N_20587);
nor U20657 (N_20657,N_20493,N_20502);
xor U20658 (N_20658,N_20412,N_20457);
xnor U20659 (N_20659,N_20535,N_20415);
and U20660 (N_20660,N_20466,N_20409);
and U20661 (N_20661,N_20506,N_20547);
nor U20662 (N_20662,N_20592,N_20480);
nor U20663 (N_20663,N_20574,N_20515);
nor U20664 (N_20664,N_20536,N_20594);
xnor U20665 (N_20665,N_20516,N_20512);
and U20666 (N_20666,N_20557,N_20476);
and U20667 (N_20667,N_20473,N_20537);
or U20668 (N_20668,N_20464,N_20404);
nand U20669 (N_20669,N_20526,N_20513);
or U20670 (N_20670,N_20527,N_20531);
or U20671 (N_20671,N_20511,N_20509);
nor U20672 (N_20672,N_20419,N_20500);
or U20673 (N_20673,N_20580,N_20504);
xnor U20674 (N_20674,N_20494,N_20471);
or U20675 (N_20675,N_20524,N_20491);
or U20676 (N_20676,N_20429,N_20495);
nand U20677 (N_20677,N_20499,N_20590);
and U20678 (N_20678,N_20451,N_20461);
nor U20679 (N_20679,N_20435,N_20414);
xor U20680 (N_20680,N_20520,N_20561);
or U20681 (N_20681,N_20571,N_20577);
or U20682 (N_20682,N_20436,N_20528);
xor U20683 (N_20683,N_20424,N_20596);
nand U20684 (N_20684,N_20498,N_20508);
nor U20685 (N_20685,N_20438,N_20555);
or U20686 (N_20686,N_20450,N_20534);
nor U20687 (N_20687,N_20402,N_20496);
and U20688 (N_20688,N_20558,N_20597);
nor U20689 (N_20689,N_20445,N_20468);
nor U20690 (N_20690,N_20479,N_20472);
nand U20691 (N_20691,N_20484,N_20426);
and U20692 (N_20692,N_20567,N_20539);
nand U20693 (N_20693,N_20492,N_20563);
xor U20694 (N_20694,N_20564,N_20443);
nand U20695 (N_20695,N_20422,N_20545);
and U20696 (N_20696,N_20455,N_20570);
and U20697 (N_20697,N_20575,N_20489);
nand U20698 (N_20698,N_20460,N_20427);
or U20699 (N_20699,N_20465,N_20543);
nand U20700 (N_20700,N_20572,N_20461);
and U20701 (N_20701,N_20503,N_20521);
xor U20702 (N_20702,N_20401,N_20476);
xor U20703 (N_20703,N_20479,N_20463);
or U20704 (N_20704,N_20422,N_20598);
xor U20705 (N_20705,N_20590,N_20459);
or U20706 (N_20706,N_20560,N_20528);
and U20707 (N_20707,N_20595,N_20409);
xor U20708 (N_20708,N_20416,N_20477);
and U20709 (N_20709,N_20564,N_20466);
nor U20710 (N_20710,N_20497,N_20429);
nor U20711 (N_20711,N_20573,N_20478);
and U20712 (N_20712,N_20592,N_20436);
nor U20713 (N_20713,N_20564,N_20469);
and U20714 (N_20714,N_20465,N_20523);
xnor U20715 (N_20715,N_20539,N_20464);
nor U20716 (N_20716,N_20477,N_20499);
nand U20717 (N_20717,N_20536,N_20599);
nor U20718 (N_20718,N_20486,N_20490);
and U20719 (N_20719,N_20592,N_20520);
nand U20720 (N_20720,N_20569,N_20409);
and U20721 (N_20721,N_20431,N_20460);
nor U20722 (N_20722,N_20435,N_20442);
nand U20723 (N_20723,N_20471,N_20500);
xor U20724 (N_20724,N_20422,N_20507);
nor U20725 (N_20725,N_20449,N_20511);
or U20726 (N_20726,N_20541,N_20400);
or U20727 (N_20727,N_20492,N_20465);
and U20728 (N_20728,N_20520,N_20494);
xnor U20729 (N_20729,N_20477,N_20520);
nor U20730 (N_20730,N_20551,N_20527);
nand U20731 (N_20731,N_20410,N_20498);
nor U20732 (N_20732,N_20414,N_20524);
and U20733 (N_20733,N_20509,N_20469);
nor U20734 (N_20734,N_20411,N_20512);
nor U20735 (N_20735,N_20451,N_20492);
xnor U20736 (N_20736,N_20510,N_20444);
and U20737 (N_20737,N_20439,N_20595);
nor U20738 (N_20738,N_20590,N_20427);
and U20739 (N_20739,N_20571,N_20507);
nor U20740 (N_20740,N_20589,N_20449);
nor U20741 (N_20741,N_20554,N_20408);
or U20742 (N_20742,N_20558,N_20413);
and U20743 (N_20743,N_20469,N_20528);
or U20744 (N_20744,N_20407,N_20475);
nand U20745 (N_20745,N_20481,N_20457);
nand U20746 (N_20746,N_20491,N_20469);
and U20747 (N_20747,N_20475,N_20583);
or U20748 (N_20748,N_20413,N_20473);
and U20749 (N_20749,N_20529,N_20486);
nor U20750 (N_20750,N_20428,N_20556);
nand U20751 (N_20751,N_20447,N_20460);
xor U20752 (N_20752,N_20440,N_20515);
or U20753 (N_20753,N_20588,N_20519);
and U20754 (N_20754,N_20528,N_20420);
xor U20755 (N_20755,N_20529,N_20478);
and U20756 (N_20756,N_20545,N_20497);
or U20757 (N_20757,N_20548,N_20535);
nor U20758 (N_20758,N_20522,N_20473);
xor U20759 (N_20759,N_20439,N_20417);
or U20760 (N_20760,N_20427,N_20457);
nand U20761 (N_20761,N_20549,N_20496);
nor U20762 (N_20762,N_20455,N_20443);
nor U20763 (N_20763,N_20594,N_20446);
and U20764 (N_20764,N_20435,N_20595);
xnor U20765 (N_20765,N_20406,N_20425);
nand U20766 (N_20766,N_20503,N_20547);
and U20767 (N_20767,N_20534,N_20490);
nor U20768 (N_20768,N_20470,N_20515);
and U20769 (N_20769,N_20553,N_20532);
xor U20770 (N_20770,N_20478,N_20566);
xnor U20771 (N_20771,N_20517,N_20492);
nand U20772 (N_20772,N_20496,N_20426);
xor U20773 (N_20773,N_20516,N_20493);
nor U20774 (N_20774,N_20422,N_20474);
nand U20775 (N_20775,N_20592,N_20441);
and U20776 (N_20776,N_20550,N_20485);
xor U20777 (N_20777,N_20442,N_20456);
xnor U20778 (N_20778,N_20490,N_20557);
xnor U20779 (N_20779,N_20526,N_20448);
and U20780 (N_20780,N_20573,N_20591);
or U20781 (N_20781,N_20506,N_20441);
nor U20782 (N_20782,N_20420,N_20532);
nor U20783 (N_20783,N_20462,N_20433);
nor U20784 (N_20784,N_20467,N_20531);
nor U20785 (N_20785,N_20550,N_20527);
or U20786 (N_20786,N_20556,N_20548);
xor U20787 (N_20787,N_20429,N_20412);
xnor U20788 (N_20788,N_20491,N_20439);
or U20789 (N_20789,N_20430,N_20529);
nand U20790 (N_20790,N_20417,N_20564);
nand U20791 (N_20791,N_20551,N_20459);
or U20792 (N_20792,N_20520,N_20441);
or U20793 (N_20793,N_20594,N_20458);
xor U20794 (N_20794,N_20596,N_20444);
nand U20795 (N_20795,N_20534,N_20522);
nor U20796 (N_20796,N_20476,N_20584);
nor U20797 (N_20797,N_20491,N_20519);
and U20798 (N_20798,N_20581,N_20433);
xor U20799 (N_20799,N_20417,N_20557);
nor U20800 (N_20800,N_20692,N_20626);
or U20801 (N_20801,N_20727,N_20663);
or U20802 (N_20802,N_20781,N_20694);
xor U20803 (N_20803,N_20655,N_20620);
nand U20804 (N_20804,N_20678,N_20754);
nor U20805 (N_20805,N_20799,N_20774);
or U20806 (N_20806,N_20758,N_20632);
and U20807 (N_20807,N_20648,N_20734);
nand U20808 (N_20808,N_20710,N_20798);
or U20809 (N_20809,N_20725,N_20689);
xnor U20810 (N_20810,N_20757,N_20625);
xor U20811 (N_20811,N_20677,N_20664);
and U20812 (N_20812,N_20613,N_20768);
and U20813 (N_20813,N_20797,N_20631);
and U20814 (N_20814,N_20776,N_20662);
nand U20815 (N_20815,N_20687,N_20607);
or U20816 (N_20816,N_20759,N_20769);
nor U20817 (N_20817,N_20735,N_20646);
or U20818 (N_20818,N_20762,N_20704);
nand U20819 (N_20819,N_20638,N_20621);
nand U20820 (N_20820,N_20791,N_20745);
nand U20821 (N_20821,N_20610,N_20614);
nand U20822 (N_20822,N_20702,N_20772);
and U20823 (N_20823,N_20658,N_20667);
xnor U20824 (N_20824,N_20688,N_20778);
nand U20825 (N_20825,N_20630,N_20649);
xnor U20826 (N_20826,N_20647,N_20764);
xor U20827 (N_20827,N_20628,N_20756);
or U20828 (N_20828,N_20615,N_20784);
and U20829 (N_20829,N_20656,N_20682);
nand U20830 (N_20830,N_20605,N_20748);
nand U20831 (N_20831,N_20696,N_20695);
nor U20832 (N_20832,N_20653,N_20752);
nor U20833 (N_20833,N_20782,N_20675);
nand U20834 (N_20834,N_20672,N_20718);
nor U20835 (N_20835,N_20603,N_20706);
or U20836 (N_20836,N_20690,N_20627);
xnor U20837 (N_20837,N_20780,N_20766);
nand U20838 (N_20838,N_20760,N_20708);
and U20839 (N_20839,N_20739,N_20779);
nor U20840 (N_20840,N_20701,N_20767);
nor U20841 (N_20841,N_20652,N_20697);
xor U20842 (N_20842,N_20673,N_20716);
xor U20843 (N_20843,N_20777,N_20700);
or U20844 (N_20844,N_20622,N_20732);
nor U20845 (N_20845,N_20792,N_20693);
and U20846 (N_20846,N_20643,N_20733);
xor U20847 (N_20847,N_20711,N_20608);
nand U20848 (N_20848,N_20763,N_20707);
and U20849 (N_20849,N_20602,N_20709);
nand U20850 (N_20850,N_20747,N_20750);
and U20851 (N_20851,N_20761,N_20669);
or U20852 (N_20852,N_20715,N_20660);
and U20853 (N_20853,N_20606,N_20611);
and U20854 (N_20854,N_20641,N_20618);
nand U20855 (N_20855,N_20651,N_20786);
nand U20856 (N_20856,N_20686,N_20736);
xor U20857 (N_20857,N_20666,N_20665);
and U20858 (N_20858,N_20657,N_20729);
nand U20859 (N_20859,N_20601,N_20624);
nor U20860 (N_20860,N_20659,N_20719);
xor U20861 (N_20861,N_20650,N_20717);
nand U20862 (N_20862,N_20728,N_20742);
or U20863 (N_20863,N_20785,N_20788);
nand U20864 (N_20864,N_20644,N_20712);
or U20865 (N_20865,N_20691,N_20753);
xor U20866 (N_20866,N_20671,N_20722);
xor U20867 (N_20867,N_20773,N_20731);
xnor U20868 (N_20868,N_20684,N_20793);
nand U20869 (N_20869,N_20668,N_20744);
xnor U20870 (N_20870,N_20794,N_20683);
xnor U20871 (N_20871,N_20635,N_20680);
or U20872 (N_20872,N_20670,N_20714);
or U20873 (N_20873,N_20787,N_20699);
nand U20874 (N_20874,N_20743,N_20737);
nand U20875 (N_20875,N_20616,N_20789);
or U20876 (N_20876,N_20751,N_20685);
nand U20877 (N_20877,N_20749,N_20770);
nand U20878 (N_20878,N_20617,N_20636);
or U20879 (N_20879,N_20674,N_20726);
nand U20880 (N_20880,N_20738,N_20619);
nor U20881 (N_20881,N_20720,N_20703);
nand U20882 (N_20882,N_20746,N_20740);
or U20883 (N_20883,N_20713,N_20724);
nor U20884 (N_20884,N_20790,N_20723);
or U20885 (N_20885,N_20609,N_20645);
and U20886 (N_20886,N_20698,N_20730);
and U20887 (N_20887,N_20676,N_20741);
and U20888 (N_20888,N_20796,N_20681);
nor U20889 (N_20889,N_20795,N_20755);
and U20890 (N_20890,N_20639,N_20640);
nand U20891 (N_20891,N_20642,N_20637);
and U20892 (N_20892,N_20634,N_20765);
nor U20893 (N_20893,N_20679,N_20633);
or U20894 (N_20894,N_20661,N_20721);
xor U20895 (N_20895,N_20705,N_20654);
or U20896 (N_20896,N_20783,N_20612);
nand U20897 (N_20897,N_20629,N_20600);
nor U20898 (N_20898,N_20623,N_20775);
or U20899 (N_20899,N_20604,N_20771);
nand U20900 (N_20900,N_20733,N_20787);
xor U20901 (N_20901,N_20710,N_20729);
and U20902 (N_20902,N_20635,N_20692);
xnor U20903 (N_20903,N_20794,N_20632);
nor U20904 (N_20904,N_20646,N_20792);
and U20905 (N_20905,N_20795,N_20662);
xor U20906 (N_20906,N_20743,N_20679);
nand U20907 (N_20907,N_20765,N_20769);
and U20908 (N_20908,N_20632,N_20796);
nor U20909 (N_20909,N_20685,N_20766);
nand U20910 (N_20910,N_20760,N_20703);
xnor U20911 (N_20911,N_20752,N_20768);
nand U20912 (N_20912,N_20720,N_20622);
nor U20913 (N_20913,N_20619,N_20686);
xor U20914 (N_20914,N_20673,N_20600);
and U20915 (N_20915,N_20757,N_20746);
or U20916 (N_20916,N_20606,N_20631);
nor U20917 (N_20917,N_20745,N_20680);
and U20918 (N_20918,N_20687,N_20604);
xnor U20919 (N_20919,N_20708,N_20794);
nor U20920 (N_20920,N_20773,N_20635);
and U20921 (N_20921,N_20758,N_20686);
xnor U20922 (N_20922,N_20674,N_20683);
or U20923 (N_20923,N_20778,N_20716);
nand U20924 (N_20924,N_20675,N_20650);
nor U20925 (N_20925,N_20778,N_20770);
nand U20926 (N_20926,N_20636,N_20715);
or U20927 (N_20927,N_20727,N_20771);
nor U20928 (N_20928,N_20764,N_20680);
xor U20929 (N_20929,N_20726,N_20624);
or U20930 (N_20930,N_20798,N_20711);
xnor U20931 (N_20931,N_20742,N_20719);
nand U20932 (N_20932,N_20762,N_20692);
xnor U20933 (N_20933,N_20659,N_20635);
nand U20934 (N_20934,N_20791,N_20728);
or U20935 (N_20935,N_20623,N_20681);
nor U20936 (N_20936,N_20650,N_20750);
nand U20937 (N_20937,N_20678,N_20606);
or U20938 (N_20938,N_20769,N_20624);
nand U20939 (N_20939,N_20624,N_20654);
xor U20940 (N_20940,N_20749,N_20689);
nor U20941 (N_20941,N_20662,N_20626);
xor U20942 (N_20942,N_20762,N_20651);
and U20943 (N_20943,N_20665,N_20756);
xor U20944 (N_20944,N_20703,N_20766);
or U20945 (N_20945,N_20632,N_20750);
nand U20946 (N_20946,N_20782,N_20766);
nand U20947 (N_20947,N_20615,N_20606);
xor U20948 (N_20948,N_20766,N_20681);
nor U20949 (N_20949,N_20770,N_20753);
nand U20950 (N_20950,N_20637,N_20766);
nand U20951 (N_20951,N_20714,N_20794);
nor U20952 (N_20952,N_20662,N_20774);
nand U20953 (N_20953,N_20741,N_20736);
or U20954 (N_20954,N_20758,N_20607);
or U20955 (N_20955,N_20635,N_20622);
nand U20956 (N_20956,N_20791,N_20776);
nor U20957 (N_20957,N_20661,N_20719);
and U20958 (N_20958,N_20674,N_20629);
nand U20959 (N_20959,N_20789,N_20687);
and U20960 (N_20960,N_20662,N_20792);
or U20961 (N_20961,N_20720,N_20604);
nand U20962 (N_20962,N_20608,N_20676);
or U20963 (N_20963,N_20738,N_20687);
xor U20964 (N_20964,N_20664,N_20758);
or U20965 (N_20965,N_20773,N_20794);
nor U20966 (N_20966,N_20776,N_20640);
nor U20967 (N_20967,N_20635,N_20771);
nor U20968 (N_20968,N_20717,N_20657);
or U20969 (N_20969,N_20688,N_20731);
and U20970 (N_20970,N_20605,N_20680);
nor U20971 (N_20971,N_20720,N_20723);
and U20972 (N_20972,N_20618,N_20635);
or U20973 (N_20973,N_20713,N_20686);
and U20974 (N_20974,N_20739,N_20758);
or U20975 (N_20975,N_20743,N_20683);
and U20976 (N_20976,N_20752,N_20622);
nor U20977 (N_20977,N_20748,N_20747);
xor U20978 (N_20978,N_20711,N_20796);
or U20979 (N_20979,N_20635,N_20663);
or U20980 (N_20980,N_20734,N_20766);
xnor U20981 (N_20981,N_20635,N_20706);
nor U20982 (N_20982,N_20755,N_20626);
nand U20983 (N_20983,N_20638,N_20615);
xor U20984 (N_20984,N_20786,N_20639);
nand U20985 (N_20985,N_20612,N_20635);
nor U20986 (N_20986,N_20645,N_20795);
or U20987 (N_20987,N_20742,N_20611);
nand U20988 (N_20988,N_20675,N_20714);
xor U20989 (N_20989,N_20743,N_20730);
and U20990 (N_20990,N_20670,N_20763);
nand U20991 (N_20991,N_20688,N_20783);
and U20992 (N_20992,N_20726,N_20791);
xnor U20993 (N_20993,N_20693,N_20626);
or U20994 (N_20994,N_20658,N_20796);
xor U20995 (N_20995,N_20744,N_20645);
or U20996 (N_20996,N_20707,N_20671);
xnor U20997 (N_20997,N_20630,N_20629);
and U20998 (N_20998,N_20768,N_20631);
nor U20999 (N_20999,N_20756,N_20623);
or U21000 (N_21000,N_20822,N_20818);
and U21001 (N_21001,N_20902,N_20827);
or U21002 (N_21002,N_20973,N_20922);
or U21003 (N_21003,N_20881,N_20976);
nand U21004 (N_21004,N_20999,N_20950);
or U21005 (N_21005,N_20908,N_20966);
xor U21006 (N_21006,N_20808,N_20895);
nand U21007 (N_21007,N_20916,N_20880);
or U21008 (N_21008,N_20944,N_20947);
or U21009 (N_21009,N_20876,N_20939);
xor U21010 (N_21010,N_20833,N_20938);
or U21011 (N_21011,N_20959,N_20982);
xor U21012 (N_21012,N_20933,N_20905);
or U21013 (N_21013,N_20963,N_20830);
nand U21014 (N_21014,N_20893,N_20987);
and U21015 (N_21015,N_20865,N_20824);
and U21016 (N_21016,N_20864,N_20952);
nor U21017 (N_21017,N_20906,N_20968);
nand U21018 (N_21018,N_20937,N_20898);
and U21019 (N_21019,N_20981,N_20883);
nand U21020 (N_21020,N_20839,N_20979);
and U21021 (N_21021,N_20921,N_20857);
and U21022 (N_21022,N_20866,N_20985);
nand U21023 (N_21023,N_20826,N_20888);
and U21024 (N_21024,N_20832,N_20819);
nor U21025 (N_21025,N_20951,N_20925);
or U21026 (N_21026,N_20961,N_20945);
and U21027 (N_21027,N_20934,N_20810);
nor U21028 (N_21028,N_20941,N_20917);
nor U21029 (N_21029,N_20860,N_20804);
nand U21030 (N_21030,N_20802,N_20991);
xnor U21031 (N_21031,N_20854,N_20929);
xor U21032 (N_21032,N_20875,N_20807);
and U21033 (N_21033,N_20867,N_20840);
xor U21034 (N_21034,N_20958,N_20960);
nor U21035 (N_21035,N_20871,N_20978);
nor U21036 (N_21036,N_20800,N_20836);
and U21037 (N_21037,N_20862,N_20835);
nand U21038 (N_21038,N_20964,N_20954);
or U21039 (N_21039,N_20879,N_20899);
xnor U21040 (N_21040,N_20986,N_20998);
and U21041 (N_21041,N_20816,N_20889);
or U21042 (N_21042,N_20930,N_20900);
or U21043 (N_21043,N_20913,N_20825);
and U21044 (N_21044,N_20843,N_20988);
or U21045 (N_21045,N_20926,N_20817);
nand U21046 (N_21046,N_20859,N_20855);
and U21047 (N_21047,N_20896,N_20853);
xor U21048 (N_21048,N_20993,N_20990);
and U21049 (N_21049,N_20831,N_20872);
and U21050 (N_21050,N_20918,N_20935);
nor U21051 (N_21051,N_20995,N_20953);
or U21052 (N_21052,N_20983,N_20809);
nand U21053 (N_21053,N_20920,N_20837);
or U21054 (N_21054,N_20845,N_20844);
or U21055 (N_21055,N_20972,N_20834);
or U21056 (N_21056,N_20901,N_20936);
nand U21057 (N_21057,N_20984,N_20891);
nand U21058 (N_21058,N_20910,N_20823);
and U21059 (N_21059,N_20940,N_20914);
nand U21060 (N_21060,N_20828,N_20887);
and U21061 (N_21061,N_20992,N_20846);
or U21062 (N_21062,N_20868,N_20838);
or U21063 (N_21063,N_20892,N_20863);
nor U21064 (N_21064,N_20969,N_20870);
nor U21065 (N_21065,N_20849,N_20803);
or U21066 (N_21066,N_20932,N_20814);
nand U21067 (N_21067,N_20965,N_20850);
xnor U21068 (N_21068,N_20931,N_20873);
nand U21069 (N_21069,N_20980,N_20856);
and U21070 (N_21070,N_20847,N_20805);
or U21071 (N_21071,N_20903,N_20848);
and U21072 (N_21072,N_20897,N_20907);
xor U21073 (N_21073,N_20919,N_20877);
or U21074 (N_21074,N_20924,N_20975);
nand U21075 (N_21075,N_20801,N_20861);
and U21076 (N_21076,N_20815,N_20894);
nor U21077 (N_21077,N_20943,N_20909);
and U21078 (N_21078,N_20852,N_20904);
nand U21079 (N_21079,N_20946,N_20915);
xnor U21080 (N_21080,N_20994,N_20949);
and U21081 (N_21081,N_20874,N_20971);
xnor U21082 (N_21082,N_20885,N_20812);
and U21083 (N_21083,N_20806,N_20997);
and U21084 (N_21084,N_20948,N_20912);
nor U21085 (N_21085,N_20928,N_20923);
and U21086 (N_21086,N_20977,N_20996);
or U21087 (N_21087,N_20886,N_20858);
xnor U21088 (N_21088,N_20882,N_20957);
xnor U21089 (N_21089,N_20842,N_20890);
nand U21090 (N_21090,N_20962,N_20956);
or U21091 (N_21091,N_20869,N_20927);
xor U21092 (N_21092,N_20989,N_20911);
xnor U21093 (N_21093,N_20851,N_20820);
xor U21094 (N_21094,N_20955,N_20821);
nand U21095 (N_21095,N_20811,N_20970);
xnor U21096 (N_21096,N_20967,N_20813);
or U21097 (N_21097,N_20841,N_20878);
and U21098 (N_21098,N_20942,N_20829);
nor U21099 (N_21099,N_20884,N_20974);
or U21100 (N_21100,N_20916,N_20947);
or U21101 (N_21101,N_20837,N_20866);
nor U21102 (N_21102,N_20815,N_20969);
nand U21103 (N_21103,N_20850,N_20994);
nand U21104 (N_21104,N_20861,N_20856);
nor U21105 (N_21105,N_20887,N_20842);
or U21106 (N_21106,N_20988,N_20899);
xnor U21107 (N_21107,N_20962,N_20888);
nor U21108 (N_21108,N_20861,N_20800);
nor U21109 (N_21109,N_20901,N_20820);
and U21110 (N_21110,N_20938,N_20821);
xor U21111 (N_21111,N_20970,N_20962);
nand U21112 (N_21112,N_20948,N_20817);
and U21113 (N_21113,N_20810,N_20813);
nand U21114 (N_21114,N_20895,N_20967);
nor U21115 (N_21115,N_20815,N_20835);
and U21116 (N_21116,N_20824,N_20931);
and U21117 (N_21117,N_20878,N_20872);
or U21118 (N_21118,N_20850,N_20915);
and U21119 (N_21119,N_20935,N_20924);
or U21120 (N_21120,N_20935,N_20966);
nand U21121 (N_21121,N_20973,N_20960);
nand U21122 (N_21122,N_20903,N_20998);
and U21123 (N_21123,N_20865,N_20850);
nor U21124 (N_21124,N_20950,N_20896);
xnor U21125 (N_21125,N_20990,N_20913);
or U21126 (N_21126,N_20936,N_20849);
nor U21127 (N_21127,N_20866,N_20886);
nor U21128 (N_21128,N_20884,N_20995);
or U21129 (N_21129,N_20979,N_20817);
xor U21130 (N_21130,N_20962,N_20811);
nor U21131 (N_21131,N_20874,N_20999);
nand U21132 (N_21132,N_20830,N_20865);
and U21133 (N_21133,N_20815,N_20831);
or U21134 (N_21134,N_20850,N_20851);
or U21135 (N_21135,N_20953,N_20990);
or U21136 (N_21136,N_20935,N_20945);
or U21137 (N_21137,N_20812,N_20820);
and U21138 (N_21138,N_20993,N_20871);
nand U21139 (N_21139,N_20840,N_20826);
xnor U21140 (N_21140,N_20911,N_20893);
and U21141 (N_21141,N_20989,N_20843);
and U21142 (N_21142,N_20887,N_20939);
nand U21143 (N_21143,N_20800,N_20819);
or U21144 (N_21144,N_20984,N_20901);
xor U21145 (N_21145,N_20878,N_20882);
xnor U21146 (N_21146,N_20992,N_20982);
and U21147 (N_21147,N_20947,N_20837);
and U21148 (N_21148,N_20803,N_20836);
or U21149 (N_21149,N_20949,N_20929);
xor U21150 (N_21150,N_20813,N_20952);
and U21151 (N_21151,N_20847,N_20986);
and U21152 (N_21152,N_20945,N_20885);
xnor U21153 (N_21153,N_20883,N_20815);
xor U21154 (N_21154,N_20991,N_20876);
or U21155 (N_21155,N_20958,N_20863);
and U21156 (N_21156,N_20925,N_20859);
xor U21157 (N_21157,N_20896,N_20980);
nand U21158 (N_21158,N_20831,N_20802);
or U21159 (N_21159,N_20966,N_20851);
or U21160 (N_21160,N_20851,N_20919);
xnor U21161 (N_21161,N_20997,N_20942);
xor U21162 (N_21162,N_20986,N_20903);
nor U21163 (N_21163,N_20833,N_20876);
or U21164 (N_21164,N_20973,N_20837);
and U21165 (N_21165,N_20827,N_20997);
nor U21166 (N_21166,N_20903,N_20881);
nand U21167 (N_21167,N_20951,N_20826);
nand U21168 (N_21168,N_20992,N_20957);
nand U21169 (N_21169,N_20935,N_20952);
nand U21170 (N_21170,N_20956,N_20811);
and U21171 (N_21171,N_20886,N_20905);
xor U21172 (N_21172,N_20867,N_20994);
and U21173 (N_21173,N_20919,N_20899);
nor U21174 (N_21174,N_20990,N_20935);
or U21175 (N_21175,N_20923,N_20996);
nand U21176 (N_21176,N_20951,N_20845);
or U21177 (N_21177,N_20894,N_20902);
and U21178 (N_21178,N_20853,N_20906);
xnor U21179 (N_21179,N_20883,N_20920);
nor U21180 (N_21180,N_20928,N_20987);
xnor U21181 (N_21181,N_20857,N_20801);
nand U21182 (N_21182,N_20957,N_20999);
nor U21183 (N_21183,N_20938,N_20829);
nor U21184 (N_21184,N_20925,N_20962);
and U21185 (N_21185,N_20941,N_20909);
xor U21186 (N_21186,N_20952,N_20861);
and U21187 (N_21187,N_20801,N_20983);
or U21188 (N_21188,N_20927,N_20993);
and U21189 (N_21189,N_20947,N_20899);
and U21190 (N_21190,N_20981,N_20993);
xor U21191 (N_21191,N_20963,N_20833);
nand U21192 (N_21192,N_20985,N_20881);
nand U21193 (N_21193,N_20907,N_20946);
or U21194 (N_21194,N_20898,N_20934);
nand U21195 (N_21195,N_20800,N_20899);
and U21196 (N_21196,N_20881,N_20818);
nor U21197 (N_21197,N_20811,N_20986);
and U21198 (N_21198,N_20871,N_20980);
nor U21199 (N_21199,N_20924,N_20828);
nor U21200 (N_21200,N_21138,N_21037);
xnor U21201 (N_21201,N_21185,N_21099);
xor U21202 (N_21202,N_21007,N_21126);
xnor U21203 (N_21203,N_21114,N_21090);
and U21204 (N_21204,N_21022,N_21174);
nand U21205 (N_21205,N_21014,N_21080);
nand U21206 (N_21206,N_21113,N_21074);
and U21207 (N_21207,N_21192,N_21193);
nand U21208 (N_21208,N_21121,N_21155);
and U21209 (N_21209,N_21048,N_21131);
nand U21210 (N_21210,N_21195,N_21015);
and U21211 (N_21211,N_21191,N_21179);
nand U21212 (N_21212,N_21095,N_21046);
nor U21213 (N_21213,N_21045,N_21120);
nor U21214 (N_21214,N_21033,N_21103);
nand U21215 (N_21215,N_21137,N_21072);
nor U21216 (N_21216,N_21133,N_21110);
or U21217 (N_21217,N_21160,N_21055);
nand U21218 (N_21218,N_21097,N_21198);
nor U21219 (N_21219,N_21165,N_21188);
nand U21220 (N_21220,N_21018,N_21151);
and U21221 (N_21221,N_21023,N_21184);
nor U21222 (N_21222,N_21082,N_21020);
or U21223 (N_21223,N_21163,N_21100);
or U21224 (N_21224,N_21087,N_21056);
and U21225 (N_21225,N_21159,N_21035);
or U21226 (N_21226,N_21065,N_21006);
or U21227 (N_21227,N_21010,N_21096);
nor U21228 (N_21228,N_21132,N_21059);
nor U21229 (N_21229,N_21050,N_21027);
nor U21230 (N_21230,N_21034,N_21102);
nor U21231 (N_21231,N_21101,N_21169);
nor U21232 (N_21232,N_21086,N_21047);
xor U21233 (N_21233,N_21156,N_21153);
nor U21234 (N_21234,N_21017,N_21008);
or U21235 (N_21235,N_21032,N_21058);
and U21236 (N_21236,N_21145,N_21013);
nor U21237 (N_21237,N_21130,N_21190);
xnor U21238 (N_21238,N_21009,N_21049);
or U21239 (N_21239,N_21134,N_21175);
and U21240 (N_21240,N_21173,N_21125);
nand U21241 (N_21241,N_21146,N_21019);
nand U21242 (N_21242,N_21044,N_21129);
and U21243 (N_21243,N_21136,N_21003);
nor U21244 (N_21244,N_21186,N_21119);
nand U21245 (N_21245,N_21147,N_21182);
nand U21246 (N_21246,N_21177,N_21052);
xnor U21247 (N_21247,N_21029,N_21043);
xor U21248 (N_21248,N_21063,N_21053);
nor U21249 (N_21249,N_21005,N_21092);
xor U21250 (N_21250,N_21161,N_21077);
and U21251 (N_21251,N_21158,N_21122);
nor U21252 (N_21252,N_21139,N_21143);
xnor U21253 (N_21253,N_21016,N_21197);
nand U21254 (N_21254,N_21109,N_21026);
and U21255 (N_21255,N_21199,N_21094);
xor U21256 (N_21256,N_21093,N_21166);
xor U21257 (N_21257,N_21112,N_21106);
and U21258 (N_21258,N_21030,N_21061);
or U21259 (N_21259,N_21181,N_21001);
nor U21260 (N_21260,N_21062,N_21039);
nor U21261 (N_21261,N_21168,N_21031);
xor U21262 (N_21262,N_21128,N_21091);
and U21263 (N_21263,N_21117,N_21081);
or U21264 (N_21264,N_21083,N_21124);
nand U21265 (N_21265,N_21028,N_21150);
nor U21266 (N_21266,N_21069,N_21021);
nor U21267 (N_21267,N_21054,N_21012);
nor U21268 (N_21268,N_21183,N_21152);
and U21269 (N_21269,N_21076,N_21075);
and U21270 (N_21270,N_21170,N_21194);
and U21271 (N_21271,N_21157,N_21067);
and U21272 (N_21272,N_21068,N_21141);
xnor U21273 (N_21273,N_21088,N_21024);
nor U21274 (N_21274,N_21036,N_21040);
nor U21275 (N_21275,N_21084,N_21079);
nand U21276 (N_21276,N_21098,N_21135);
xnor U21277 (N_21277,N_21104,N_21042);
nand U21278 (N_21278,N_21038,N_21071);
xor U21279 (N_21279,N_21025,N_21123);
or U21280 (N_21280,N_21164,N_21180);
nor U21281 (N_21281,N_21078,N_21011);
nand U21282 (N_21282,N_21189,N_21144);
or U21283 (N_21283,N_21000,N_21089);
nor U21284 (N_21284,N_21002,N_21172);
xnor U21285 (N_21285,N_21187,N_21111);
nand U21286 (N_21286,N_21149,N_21176);
or U21287 (N_21287,N_21085,N_21066);
or U21288 (N_21288,N_21140,N_21118);
and U21289 (N_21289,N_21196,N_21064);
or U21290 (N_21290,N_21041,N_21162);
or U21291 (N_21291,N_21115,N_21051);
or U21292 (N_21292,N_21148,N_21167);
or U21293 (N_21293,N_21154,N_21105);
or U21294 (N_21294,N_21127,N_21116);
and U21295 (N_21295,N_21108,N_21060);
and U21296 (N_21296,N_21171,N_21142);
nor U21297 (N_21297,N_21107,N_21070);
nor U21298 (N_21298,N_21178,N_21073);
xor U21299 (N_21299,N_21004,N_21057);
and U21300 (N_21300,N_21023,N_21126);
xnor U21301 (N_21301,N_21181,N_21082);
or U21302 (N_21302,N_21017,N_21020);
nor U21303 (N_21303,N_21176,N_21171);
or U21304 (N_21304,N_21130,N_21060);
or U21305 (N_21305,N_21057,N_21029);
or U21306 (N_21306,N_21180,N_21099);
or U21307 (N_21307,N_21073,N_21064);
nand U21308 (N_21308,N_21091,N_21040);
and U21309 (N_21309,N_21054,N_21037);
and U21310 (N_21310,N_21072,N_21086);
nor U21311 (N_21311,N_21172,N_21054);
xnor U21312 (N_21312,N_21131,N_21159);
nor U21313 (N_21313,N_21118,N_21054);
or U21314 (N_21314,N_21121,N_21181);
nor U21315 (N_21315,N_21185,N_21026);
xnor U21316 (N_21316,N_21167,N_21080);
and U21317 (N_21317,N_21117,N_21184);
or U21318 (N_21318,N_21124,N_21102);
and U21319 (N_21319,N_21187,N_21019);
or U21320 (N_21320,N_21058,N_21137);
or U21321 (N_21321,N_21149,N_21022);
and U21322 (N_21322,N_21016,N_21181);
nor U21323 (N_21323,N_21052,N_21100);
xor U21324 (N_21324,N_21173,N_21051);
nand U21325 (N_21325,N_21153,N_21131);
nand U21326 (N_21326,N_21190,N_21069);
or U21327 (N_21327,N_21148,N_21023);
nor U21328 (N_21328,N_21187,N_21193);
and U21329 (N_21329,N_21143,N_21070);
nor U21330 (N_21330,N_21057,N_21068);
and U21331 (N_21331,N_21061,N_21133);
nand U21332 (N_21332,N_21110,N_21047);
xor U21333 (N_21333,N_21179,N_21122);
xnor U21334 (N_21334,N_21024,N_21031);
and U21335 (N_21335,N_21197,N_21083);
nand U21336 (N_21336,N_21031,N_21055);
nand U21337 (N_21337,N_21044,N_21157);
nand U21338 (N_21338,N_21125,N_21181);
nor U21339 (N_21339,N_21164,N_21051);
xnor U21340 (N_21340,N_21117,N_21042);
nor U21341 (N_21341,N_21170,N_21023);
nor U21342 (N_21342,N_21109,N_21084);
and U21343 (N_21343,N_21181,N_21139);
or U21344 (N_21344,N_21148,N_21194);
and U21345 (N_21345,N_21156,N_21038);
nand U21346 (N_21346,N_21175,N_21160);
or U21347 (N_21347,N_21188,N_21144);
and U21348 (N_21348,N_21149,N_21190);
or U21349 (N_21349,N_21019,N_21060);
or U21350 (N_21350,N_21060,N_21180);
nand U21351 (N_21351,N_21144,N_21054);
nand U21352 (N_21352,N_21025,N_21172);
nor U21353 (N_21353,N_21173,N_21148);
nor U21354 (N_21354,N_21092,N_21192);
and U21355 (N_21355,N_21130,N_21036);
and U21356 (N_21356,N_21025,N_21193);
and U21357 (N_21357,N_21082,N_21178);
xor U21358 (N_21358,N_21058,N_21070);
xor U21359 (N_21359,N_21139,N_21048);
nor U21360 (N_21360,N_21111,N_21091);
nand U21361 (N_21361,N_21066,N_21069);
nand U21362 (N_21362,N_21153,N_21187);
or U21363 (N_21363,N_21085,N_21180);
or U21364 (N_21364,N_21163,N_21071);
or U21365 (N_21365,N_21138,N_21079);
and U21366 (N_21366,N_21159,N_21092);
nor U21367 (N_21367,N_21030,N_21018);
xor U21368 (N_21368,N_21020,N_21044);
nor U21369 (N_21369,N_21070,N_21052);
nor U21370 (N_21370,N_21047,N_21162);
nor U21371 (N_21371,N_21192,N_21088);
xnor U21372 (N_21372,N_21085,N_21134);
nor U21373 (N_21373,N_21196,N_21033);
or U21374 (N_21374,N_21015,N_21083);
xnor U21375 (N_21375,N_21182,N_21014);
nor U21376 (N_21376,N_21074,N_21066);
nor U21377 (N_21377,N_21132,N_21199);
or U21378 (N_21378,N_21111,N_21199);
and U21379 (N_21379,N_21037,N_21161);
nand U21380 (N_21380,N_21118,N_21078);
or U21381 (N_21381,N_21018,N_21166);
nor U21382 (N_21382,N_21057,N_21115);
or U21383 (N_21383,N_21182,N_21137);
xnor U21384 (N_21384,N_21046,N_21134);
and U21385 (N_21385,N_21180,N_21134);
xor U21386 (N_21386,N_21108,N_21062);
nand U21387 (N_21387,N_21123,N_21003);
xnor U21388 (N_21388,N_21162,N_21006);
or U21389 (N_21389,N_21165,N_21066);
nor U21390 (N_21390,N_21059,N_21161);
and U21391 (N_21391,N_21066,N_21140);
nand U21392 (N_21392,N_21002,N_21165);
nor U21393 (N_21393,N_21062,N_21199);
or U21394 (N_21394,N_21011,N_21056);
and U21395 (N_21395,N_21104,N_21194);
nor U21396 (N_21396,N_21158,N_21120);
nand U21397 (N_21397,N_21041,N_21078);
nand U21398 (N_21398,N_21174,N_21013);
nand U21399 (N_21399,N_21195,N_21132);
nor U21400 (N_21400,N_21318,N_21373);
xor U21401 (N_21401,N_21282,N_21330);
nor U21402 (N_21402,N_21207,N_21249);
nor U21403 (N_21403,N_21382,N_21385);
and U21404 (N_21404,N_21320,N_21348);
xor U21405 (N_21405,N_21384,N_21323);
or U21406 (N_21406,N_21327,N_21204);
xnor U21407 (N_21407,N_21391,N_21266);
nand U21408 (N_21408,N_21233,N_21220);
and U21409 (N_21409,N_21369,N_21309);
and U21410 (N_21410,N_21375,N_21275);
xnor U21411 (N_21411,N_21253,N_21294);
and U21412 (N_21412,N_21231,N_21364);
and U21413 (N_21413,N_21374,N_21290);
and U21414 (N_21414,N_21223,N_21243);
or U21415 (N_21415,N_21350,N_21345);
and U21416 (N_21416,N_21281,N_21315);
and U21417 (N_21417,N_21319,N_21277);
nand U21418 (N_21418,N_21254,N_21239);
and U21419 (N_21419,N_21212,N_21366);
nand U21420 (N_21420,N_21317,N_21390);
or U21421 (N_21421,N_21280,N_21300);
or U21422 (N_21422,N_21200,N_21201);
nand U21423 (N_21423,N_21340,N_21232);
nor U21424 (N_21424,N_21289,N_21214);
nand U21425 (N_21425,N_21376,N_21218);
nand U21426 (N_21426,N_21227,N_21298);
or U21427 (N_21427,N_21341,N_21228);
and U21428 (N_21428,N_21236,N_21326);
xor U21429 (N_21429,N_21324,N_21355);
xor U21430 (N_21430,N_21328,N_21276);
or U21431 (N_21431,N_21274,N_21358);
nand U21432 (N_21432,N_21237,N_21217);
xor U21433 (N_21433,N_21392,N_21325);
or U21434 (N_21434,N_21304,N_21396);
or U21435 (N_21435,N_21271,N_21262);
nor U21436 (N_21436,N_21263,N_21372);
or U21437 (N_21437,N_21339,N_21241);
or U21438 (N_21438,N_21399,N_21338);
nor U21439 (N_21439,N_21205,N_21370);
and U21440 (N_21440,N_21221,N_21208);
nand U21441 (N_21441,N_21367,N_21343);
nand U21442 (N_21442,N_21206,N_21332);
or U21443 (N_21443,N_21305,N_21347);
or U21444 (N_21444,N_21297,N_21256);
and U21445 (N_21445,N_21377,N_21394);
xnor U21446 (N_21446,N_21251,N_21238);
nand U21447 (N_21447,N_21351,N_21291);
nand U21448 (N_21448,N_21329,N_21337);
xor U21449 (N_21449,N_21216,N_21219);
nor U21450 (N_21450,N_21359,N_21273);
and U21451 (N_21451,N_21334,N_21378);
nand U21452 (N_21452,N_21224,N_21397);
xor U21453 (N_21453,N_21259,N_21265);
xnor U21454 (N_21454,N_21283,N_21310);
nor U21455 (N_21455,N_21316,N_21285);
nor U21456 (N_21456,N_21303,N_21244);
or U21457 (N_21457,N_21308,N_21307);
nor U21458 (N_21458,N_21215,N_21296);
nor U21459 (N_21459,N_21362,N_21333);
xor U21460 (N_21460,N_21247,N_21242);
xnor U21461 (N_21461,N_21357,N_21398);
nor U21462 (N_21462,N_21225,N_21250);
nand U21463 (N_21463,N_21299,N_21361);
and U21464 (N_21464,N_21295,N_21349);
or U21465 (N_21465,N_21248,N_21229);
and U21466 (N_21466,N_21383,N_21314);
nor U21467 (N_21467,N_21356,N_21381);
or U21468 (N_21468,N_21269,N_21311);
nand U21469 (N_21469,N_21222,N_21331);
xor U21470 (N_21470,N_21261,N_21258);
nand U21471 (N_21471,N_21246,N_21313);
or U21472 (N_21472,N_21260,N_21240);
and U21473 (N_21473,N_21230,N_21203);
or U21474 (N_21474,N_21267,N_21211);
and U21475 (N_21475,N_21387,N_21252);
nor U21476 (N_21476,N_21302,N_21363);
nor U21477 (N_21477,N_21353,N_21234);
xnor U21478 (N_21478,N_21245,N_21270);
or U21479 (N_21479,N_21388,N_21210);
nor U21480 (N_21480,N_21255,N_21321);
nor U21481 (N_21481,N_21371,N_21380);
xor U21482 (N_21482,N_21360,N_21386);
xor U21483 (N_21483,N_21389,N_21342);
nand U21484 (N_21484,N_21336,N_21346);
xor U21485 (N_21485,N_21335,N_21278);
or U21486 (N_21486,N_21279,N_21287);
nand U21487 (N_21487,N_21354,N_21284);
nand U21488 (N_21488,N_21393,N_21202);
or U21489 (N_21489,N_21272,N_21352);
nand U21490 (N_21490,N_21379,N_21257);
nor U21491 (N_21491,N_21306,N_21344);
nor U21492 (N_21492,N_21226,N_21365);
nor U21493 (N_21493,N_21293,N_21264);
nand U21494 (N_21494,N_21368,N_21286);
nand U21495 (N_21495,N_21312,N_21235);
nand U21496 (N_21496,N_21292,N_21395);
xnor U21497 (N_21497,N_21322,N_21301);
nor U21498 (N_21498,N_21209,N_21288);
or U21499 (N_21499,N_21213,N_21268);
or U21500 (N_21500,N_21391,N_21277);
nor U21501 (N_21501,N_21387,N_21276);
nand U21502 (N_21502,N_21273,N_21348);
xnor U21503 (N_21503,N_21355,N_21216);
xnor U21504 (N_21504,N_21312,N_21250);
nor U21505 (N_21505,N_21312,N_21357);
nand U21506 (N_21506,N_21348,N_21230);
or U21507 (N_21507,N_21214,N_21343);
and U21508 (N_21508,N_21276,N_21380);
and U21509 (N_21509,N_21325,N_21277);
xnor U21510 (N_21510,N_21202,N_21287);
nand U21511 (N_21511,N_21256,N_21338);
or U21512 (N_21512,N_21245,N_21364);
nor U21513 (N_21513,N_21365,N_21333);
nand U21514 (N_21514,N_21240,N_21221);
and U21515 (N_21515,N_21308,N_21205);
nand U21516 (N_21516,N_21325,N_21331);
and U21517 (N_21517,N_21265,N_21329);
or U21518 (N_21518,N_21299,N_21213);
nand U21519 (N_21519,N_21329,N_21346);
xor U21520 (N_21520,N_21273,N_21353);
and U21521 (N_21521,N_21291,N_21223);
or U21522 (N_21522,N_21358,N_21264);
xor U21523 (N_21523,N_21291,N_21315);
xnor U21524 (N_21524,N_21323,N_21237);
or U21525 (N_21525,N_21206,N_21376);
nand U21526 (N_21526,N_21261,N_21377);
and U21527 (N_21527,N_21363,N_21343);
xnor U21528 (N_21528,N_21203,N_21327);
or U21529 (N_21529,N_21357,N_21294);
xor U21530 (N_21530,N_21382,N_21328);
xnor U21531 (N_21531,N_21285,N_21210);
and U21532 (N_21532,N_21389,N_21266);
nand U21533 (N_21533,N_21264,N_21382);
nor U21534 (N_21534,N_21346,N_21375);
nor U21535 (N_21535,N_21257,N_21367);
xor U21536 (N_21536,N_21296,N_21398);
and U21537 (N_21537,N_21338,N_21325);
xnor U21538 (N_21538,N_21288,N_21235);
and U21539 (N_21539,N_21241,N_21386);
nand U21540 (N_21540,N_21376,N_21265);
nor U21541 (N_21541,N_21231,N_21240);
nand U21542 (N_21542,N_21249,N_21399);
nand U21543 (N_21543,N_21286,N_21392);
or U21544 (N_21544,N_21310,N_21315);
nor U21545 (N_21545,N_21278,N_21396);
and U21546 (N_21546,N_21290,N_21359);
or U21547 (N_21547,N_21364,N_21351);
and U21548 (N_21548,N_21200,N_21282);
xnor U21549 (N_21549,N_21334,N_21321);
or U21550 (N_21550,N_21374,N_21317);
and U21551 (N_21551,N_21385,N_21214);
xor U21552 (N_21552,N_21346,N_21252);
xor U21553 (N_21553,N_21257,N_21200);
nand U21554 (N_21554,N_21248,N_21276);
and U21555 (N_21555,N_21229,N_21319);
nand U21556 (N_21556,N_21397,N_21278);
nand U21557 (N_21557,N_21328,N_21244);
nand U21558 (N_21558,N_21293,N_21237);
or U21559 (N_21559,N_21263,N_21225);
or U21560 (N_21560,N_21359,N_21205);
xor U21561 (N_21561,N_21215,N_21213);
or U21562 (N_21562,N_21223,N_21226);
and U21563 (N_21563,N_21377,N_21271);
or U21564 (N_21564,N_21371,N_21200);
nor U21565 (N_21565,N_21234,N_21322);
nor U21566 (N_21566,N_21258,N_21245);
nor U21567 (N_21567,N_21270,N_21259);
nand U21568 (N_21568,N_21370,N_21300);
and U21569 (N_21569,N_21278,N_21375);
nor U21570 (N_21570,N_21284,N_21269);
or U21571 (N_21571,N_21298,N_21395);
or U21572 (N_21572,N_21321,N_21253);
nor U21573 (N_21573,N_21393,N_21254);
nand U21574 (N_21574,N_21375,N_21241);
xor U21575 (N_21575,N_21380,N_21379);
or U21576 (N_21576,N_21345,N_21309);
nand U21577 (N_21577,N_21268,N_21304);
xor U21578 (N_21578,N_21241,N_21271);
nand U21579 (N_21579,N_21221,N_21318);
or U21580 (N_21580,N_21359,N_21231);
xnor U21581 (N_21581,N_21292,N_21224);
xnor U21582 (N_21582,N_21314,N_21242);
nand U21583 (N_21583,N_21389,N_21353);
or U21584 (N_21584,N_21269,N_21344);
and U21585 (N_21585,N_21311,N_21305);
and U21586 (N_21586,N_21294,N_21397);
or U21587 (N_21587,N_21221,N_21356);
and U21588 (N_21588,N_21362,N_21304);
nand U21589 (N_21589,N_21314,N_21265);
or U21590 (N_21590,N_21345,N_21257);
nand U21591 (N_21591,N_21315,N_21303);
nor U21592 (N_21592,N_21264,N_21204);
and U21593 (N_21593,N_21286,N_21328);
xnor U21594 (N_21594,N_21247,N_21209);
nand U21595 (N_21595,N_21206,N_21302);
and U21596 (N_21596,N_21240,N_21378);
or U21597 (N_21597,N_21380,N_21237);
or U21598 (N_21598,N_21324,N_21260);
and U21599 (N_21599,N_21306,N_21244);
nor U21600 (N_21600,N_21402,N_21578);
nand U21601 (N_21601,N_21410,N_21443);
xnor U21602 (N_21602,N_21441,N_21480);
and U21603 (N_21603,N_21486,N_21533);
or U21604 (N_21604,N_21587,N_21432);
nand U21605 (N_21605,N_21564,N_21456);
and U21606 (N_21606,N_21535,N_21401);
xor U21607 (N_21607,N_21433,N_21559);
xor U21608 (N_21608,N_21526,N_21507);
nor U21609 (N_21609,N_21414,N_21588);
and U21610 (N_21610,N_21566,N_21462);
and U21611 (N_21611,N_21453,N_21424);
or U21612 (N_21612,N_21591,N_21419);
xor U21613 (N_21613,N_21552,N_21506);
nand U21614 (N_21614,N_21428,N_21571);
nand U21615 (N_21615,N_21468,N_21455);
xnor U21616 (N_21616,N_21523,N_21412);
nor U21617 (N_21617,N_21517,N_21420);
xnor U21618 (N_21618,N_21452,N_21522);
nor U21619 (N_21619,N_21575,N_21471);
nand U21620 (N_21620,N_21498,N_21444);
and U21621 (N_21621,N_21413,N_21596);
nand U21622 (N_21622,N_21448,N_21421);
xor U21623 (N_21623,N_21423,N_21567);
xor U21624 (N_21624,N_21404,N_21497);
nand U21625 (N_21625,N_21514,N_21585);
or U21626 (N_21626,N_21560,N_21536);
or U21627 (N_21627,N_21426,N_21416);
xor U21628 (N_21628,N_21437,N_21580);
or U21629 (N_21629,N_21574,N_21487);
or U21630 (N_21630,N_21569,N_21593);
nor U21631 (N_21631,N_21520,N_21467);
nor U21632 (N_21632,N_21577,N_21547);
and U21633 (N_21633,N_21430,N_21509);
xor U21634 (N_21634,N_21495,N_21494);
or U21635 (N_21635,N_21508,N_21440);
nand U21636 (N_21636,N_21582,N_21565);
and U21637 (N_21637,N_21563,N_21447);
and U21638 (N_21638,N_21479,N_21406);
and U21639 (N_21639,N_21446,N_21546);
xor U21640 (N_21640,N_21477,N_21597);
or U21641 (N_21641,N_21461,N_21472);
and U21642 (N_21642,N_21484,N_21543);
nor U21643 (N_21643,N_21435,N_21541);
or U21644 (N_21644,N_21449,N_21521);
nor U21645 (N_21645,N_21463,N_21457);
and U21646 (N_21646,N_21465,N_21445);
and U21647 (N_21647,N_21482,N_21553);
nand U21648 (N_21648,N_21519,N_21422);
xor U21649 (N_21649,N_21470,N_21562);
nand U21650 (N_21650,N_21530,N_21451);
xnor U21651 (N_21651,N_21439,N_21550);
nor U21652 (N_21652,N_21476,N_21531);
or U21653 (N_21653,N_21500,N_21594);
xnor U21654 (N_21654,N_21475,N_21570);
or U21655 (N_21655,N_21572,N_21545);
xnor U21656 (N_21656,N_21542,N_21548);
nand U21657 (N_21657,N_21556,N_21474);
nand U21658 (N_21658,N_21425,N_21586);
xor U21659 (N_21659,N_21539,N_21436);
nor U21660 (N_21660,N_21576,N_21431);
and U21661 (N_21661,N_21518,N_21493);
and U21662 (N_21662,N_21459,N_21418);
and U21663 (N_21663,N_21501,N_21434);
or U21664 (N_21664,N_21573,N_21554);
nand U21665 (N_21665,N_21442,N_21551);
nand U21666 (N_21666,N_21488,N_21549);
nand U21667 (N_21667,N_21579,N_21454);
xnor U21668 (N_21668,N_21540,N_21532);
nor U21669 (N_21669,N_21458,N_21528);
xor U21670 (N_21670,N_21534,N_21503);
and U21671 (N_21671,N_21481,N_21464);
nand U21672 (N_21672,N_21513,N_21403);
xor U21673 (N_21673,N_21595,N_21589);
nor U21674 (N_21674,N_21483,N_21415);
and U21675 (N_21675,N_21429,N_21511);
xnor U21676 (N_21676,N_21478,N_21581);
xor U21677 (N_21677,N_21583,N_21400);
or U21678 (N_21678,N_21538,N_21407);
xnor U21679 (N_21679,N_21557,N_21555);
nand U21680 (N_21680,N_21408,N_21405);
nor U21681 (N_21681,N_21466,N_21496);
nor U21682 (N_21682,N_21512,N_21473);
and U21683 (N_21683,N_21505,N_21537);
and U21684 (N_21684,N_21409,N_21489);
xnor U21685 (N_21685,N_21525,N_21510);
or U21686 (N_21686,N_21469,N_21502);
nand U21687 (N_21687,N_21485,N_21558);
and U21688 (N_21688,N_21599,N_21527);
nand U21689 (N_21689,N_21499,N_21515);
nor U21690 (N_21690,N_21450,N_21529);
nor U21691 (N_21691,N_21592,N_21427);
nand U21692 (N_21692,N_21561,N_21524);
nor U21693 (N_21693,N_21491,N_21590);
or U21694 (N_21694,N_21438,N_21411);
or U21695 (N_21695,N_21598,N_21544);
or U21696 (N_21696,N_21568,N_21516);
nand U21697 (N_21697,N_21584,N_21504);
xnor U21698 (N_21698,N_21492,N_21417);
or U21699 (N_21699,N_21460,N_21490);
nand U21700 (N_21700,N_21427,N_21591);
or U21701 (N_21701,N_21406,N_21548);
nor U21702 (N_21702,N_21508,N_21565);
nand U21703 (N_21703,N_21484,N_21416);
nor U21704 (N_21704,N_21497,N_21554);
and U21705 (N_21705,N_21460,N_21539);
or U21706 (N_21706,N_21400,N_21526);
xnor U21707 (N_21707,N_21407,N_21411);
xor U21708 (N_21708,N_21455,N_21512);
nand U21709 (N_21709,N_21477,N_21523);
and U21710 (N_21710,N_21595,N_21402);
and U21711 (N_21711,N_21597,N_21486);
xor U21712 (N_21712,N_21450,N_21456);
nand U21713 (N_21713,N_21485,N_21515);
nor U21714 (N_21714,N_21489,N_21505);
xor U21715 (N_21715,N_21495,N_21535);
or U21716 (N_21716,N_21529,N_21476);
nand U21717 (N_21717,N_21482,N_21427);
nand U21718 (N_21718,N_21537,N_21596);
nor U21719 (N_21719,N_21452,N_21551);
and U21720 (N_21720,N_21441,N_21559);
or U21721 (N_21721,N_21594,N_21561);
xnor U21722 (N_21722,N_21436,N_21536);
nor U21723 (N_21723,N_21550,N_21427);
nand U21724 (N_21724,N_21537,N_21567);
and U21725 (N_21725,N_21478,N_21445);
nor U21726 (N_21726,N_21429,N_21562);
xor U21727 (N_21727,N_21582,N_21587);
or U21728 (N_21728,N_21497,N_21527);
xor U21729 (N_21729,N_21541,N_21475);
nand U21730 (N_21730,N_21506,N_21457);
xnor U21731 (N_21731,N_21564,N_21525);
nor U21732 (N_21732,N_21415,N_21487);
xnor U21733 (N_21733,N_21425,N_21506);
and U21734 (N_21734,N_21540,N_21546);
xor U21735 (N_21735,N_21427,N_21437);
nand U21736 (N_21736,N_21539,N_21529);
nor U21737 (N_21737,N_21559,N_21444);
nor U21738 (N_21738,N_21410,N_21425);
nor U21739 (N_21739,N_21596,N_21487);
nand U21740 (N_21740,N_21486,N_21459);
or U21741 (N_21741,N_21409,N_21463);
and U21742 (N_21742,N_21485,N_21568);
or U21743 (N_21743,N_21589,N_21472);
nor U21744 (N_21744,N_21403,N_21453);
xnor U21745 (N_21745,N_21559,N_21586);
xnor U21746 (N_21746,N_21554,N_21402);
xnor U21747 (N_21747,N_21503,N_21401);
or U21748 (N_21748,N_21564,N_21463);
xor U21749 (N_21749,N_21449,N_21589);
nor U21750 (N_21750,N_21537,N_21539);
xnor U21751 (N_21751,N_21546,N_21407);
nor U21752 (N_21752,N_21592,N_21472);
nor U21753 (N_21753,N_21510,N_21537);
nor U21754 (N_21754,N_21507,N_21501);
nand U21755 (N_21755,N_21532,N_21416);
or U21756 (N_21756,N_21429,N_21464);
nand U21757 (N_21757,N_21502,N_21470);
xnor U21758 (N_21758,N_21455,N_21501);
nor U21759 (N_21759,N_21465,N_21527);
or U21760 (N_21760,N_21532,N_21536);
nand U21761 (N_21761,N_21464,N_21577);
and U21762 (N_21762,N_21440,N_21444);
nor U21763 (N_21763,N_21465,N_21418);
nor U21764 (N_21764,N_21589,N_21430);
nor U21765 (N_21765,N_21445,N_21508);
nand U21766 (N_21766,N_21588,N_21543);
nand U21767 (N_21767,N_21470,N_21525);
nor U21768 (N_21768,N_21556,N_21521);
nor U21769 (N_21769,N_21582,N_21585);
nand U21770 (N_21770,N_21542,N_21471);
xor U21771 (N_21771,N_21432,N_21457);
or U21772 (N_21772,N_21578,N_21536);
or U21773 (N_21773,N_21463,N_21554);
nand U21774 (N_21774,N_21501,N_21493);
and U21775 (N_21775,N_21473,N_21548);
and U21776 (N_21776,N_21405,N_21415);
or U21777 (N_21777,N_21540,N_21424);
nand U21778 (N_21778,N_21505,N_21450);
nor U21779 (N_21779,N_21516,N_21485);
and U21780 (N_21780,N_21437,N_21417);
and U21781 (N_21781,N_21485,N_21570);
nor U21782 (N_21782,N_21587,N_21528);
nand U21783 (N_21783,N_21426,N_21409);
or U21784 (N_21784,N_21456,N_21548);
or U21785 (N_21785,N_21459,N_21475);
xor U21786 (N_21786,N_21590,N_21479);
nor U21787 (N_21787,N_21505,N_21545);
nor U21788 (N_21788,N_21465,N_21459);
and U21789 (N_21789,N_21421,N_21430);
and U21790 (N_21790,N_21489,N_21586);
or U21791 (N_21791,N_21562,N_21548);
nor U21792 (N_21792,N_21456,N_21412);
xor U21793 (N_21793,N_21560,N_21540);
and U21794 (N_21794,N_21447,N_21421);
nand U21795 (N_21795,N_21448,N_21442);
or U21796 (N_21796,N_21427,N_21594);
or U21797 (N_21797,N_21568,N_21558);
nor U21798 (N_21798,N_21573,N_21498);
xor U21799 (N_21799,N_21458,N_21580);
and U21800 (N_21800,N_21706,N_21623);
and U21801 (N_21801,N_21694,N_21691);
nand U21802 (N_21802,N_21617,N_21737);
or U21803 (N_21803,N_21672,N_21656);
nor U21804 (N_21804,N_21682,N_21773);
xor U21805 (N_21805,N_21697,N_21688);
nand U21806 (N_21806,N_21676,N_21727);
nand U21807 (N_21807,N_21792,N_21679);
xor U21808 (N_21808,N_21717,N_21786);
nor U21809 (N_21809,N_21655,N_21742);
or U21810 (N_21810,N_21618,N_21650);
nor U21811 (N_21811,N_21662,N_21739);
or U21812 (N_21812,N_21797,N_21637);
and U21813 (N_21813,N_21761,N_21680);
xnor U21814 (N_21814,N_21675,N_21725);
nor U21815 (N_21815,N_21626,N_21750);
nor U21816 (N_21816,N_21684,N_21602);
and U21817 (N_21817,N_21616,N_21628);
xnor U21818 (N_21818,N_21633,N_21720);
and U21819 (N_21819,N_21765,N_21634);
xnor U21820 (N_21820,N_21639,N_21772);
or U21821 (N_21821,N_21753,N_21659);
nand U21822 (N_21822,N_21619,N_21718);
or U21823 (N_21823,N_21746,N_21651);
and U21824 (N_21824,N_21748,N_21665);
nor U21825 (N_21825,N_21647,N_21741);
nor U21826 (N_21826,N_21621,N_21789);
nand U21827 (N_21827,N_21711,N_21787);
xor U21828 (N_21828,N_21730,N_21778);
and U21829 (N_21829,N_21769,N_21686);
and U21830 (N_21830,N_21632,N_21685);
nand U21831 (N_21831,N_21726,N_21749);
or U21832 (N_21832,N_21704,N_21601);
nand U21833 (N_21833,N_21793,N_21709);
nor U21834 (N_21834,N_21775,N_21640);
and U21835 (N_21835,N_21702,N_21630);
or U21836 (N_21836,N_21710,N_21745);
nor U21837 (N_21837,N_21732,N_21657);
nand U21838 (N_21838,N_21670,N_21707);
xor U21839 (N_21839,N_21603,N_21754);
nor U21840 (N_21840,N_21738,N_21798);
nor U21841 (N_21841,N_21660,N_21692);
xor U21842 (N_21842,N_21620,N_21615);
xor U21843 (N_21843,N_21681,N_21608);
xor U21844 (N_21844,N_21674,N_21690);
or U21845 (N_21845,N_21734,N_21774);
and U21846 (N_21846,N_21794,N_21708);
xnor U21847 (N_21847,N_21767,N_21719);
or U21848 (N_21848,N_21779,N_21715);
nand U21849 (N_21849,N_21678,N_21716);
and U21850 (N_21850,N_21743,N_21612);
or U21851 (N_21851,N_21799,N_21664);
nand U21852 (N_21852,N_21796,N_21714);
and U21853 (N_21853,N_21610,N_21713);
xnor U21854 (N_21854,N_21795,N_21629);
nand U21855 (N_21855,N_21740,N_21784);
and U21856 (N_21856,N_21757,N_21631);
and U21857 (N_21857,N_21782,N_21698);
nand U21858 (N_21858,N_21790,N_21661);
or U21859 (N_21859,N_21723,N_21722);
xnor U21860 (N_21860,N_21671,N_21663);
or U21861 (N_21861,N_21699,N_21763);
or U21862 (N_21862,N_21760,N_21703);
nor U21863 (N_21863,N_21649,N_21600);
nand U21864 (N_21864,N_21747,N_21604);
or U21865 (N_21865,N_21751,N_21728);
nand U21866 (N_21866,N_21770,N_21653);
xnor U21867 (N_21867,N_21712,N_21687);
xnor U21868 (N_21868,N_21622,N_21654);
nor U21869 (N_21869,N_21648,N_21701);
and U21870 (N_21870,N_21669,N_21776);
nand U21871 (N_21871,N_21683,N_21611);
or U21872 (N_21872,N_21666,N_21689);
nor U21873 (N_21873,N_21607,N_21781);
xor U21874 (N_21874,N_21777,N_21744);
and U21875 (N_21875,N_21758,N_21646);
xnor U21876 (N_21876,N_21605,N_21785);
nor U21877 (N_21877,N_21658,N_21693);
or U21878 (N_21878,N_21606,N_21643);
nand U21879 (N_21879,N_21677,N_21766);
or U21880 (N_21880,N_21791,N_21636);
nor U21881 (N_21881,N_21735,N_21695);
and U21882 (N_21882,N_21638,N_21731);
nand U21883 (N_21883,N_21642,N_21673);
and U21884 (N_21884,N_21780,N_21652);
or U21885 (N_21885,N_21705,N_21783);
xnor U21886 (N_21886,N_21667,N_21627);
nor U21887 (N_21887,N_21788,N_21756);
xnor U21888 (N_21888,N_21759,N_21724);
and U21889 (N_21889,N_21768,N_21729);
xor U21890 (N_21890,N_21609,N_21755);
and U21891 (N_21891,N_21624,N_21696);
nand U21892 (N_21892,N_21668,N_21644);
xnor U21893 (N_21893,N_21613,N_21752);
nand U21894 (N_21894,N_21721,N_21625);
nand U21895 (N_21895,N_21771,N_21762);
or U21896 (N_21896,N_21635,N_21700);
xor U21897 (N_21897,N_21733,N_21736);
and U21898 (N_21898,N_21641,N_21645);
and U21899 (N_21899,N_21764,N_21614);
nand U21900 (N_21900,N_21727,N_21642);
and U21901 (N_21901,N_21620,N_21624);
nor U21902 (N_21902,N_21763,N_21609);
or U21903 (N_21903,N_21702,N_21688);
nor U21904 (N_21904,N_21712,N_21679);
nand U21905 (N_21905,N_21644,N_21604);
nand U21906 (N_21906,N_21674,N_21645);
xor U21907 (N_21907,N_21677,N_21774);
nor U21908 (N_21908,N_21625,N_21738);
and U21909 (N_21909,N_21675,N_21611);
xnor U21910 (N_21910,N_21712,N_21722);
or U21911 (N_21911,N_21704,N_21628);
or U21912 (N_21912,N_21635,N_21731);
or U21913 (N_21913,N_21753,N_21685);
nor U21914 (N_21914,N_21652,N_21669);
and U21915 (N_21915,N_21624,N_21751);
nand U21916 (N_21916,N_21686,N_21779);
xnor U21917 (N_21917,N_21764,N_21721);
and U21918 (N_21918,N_21689,N_21662);
and U21919 (N_21919,N_21617,N_21622);
xor U21920 (N_21920,N_21605,N_21601);
or U21921 (N_21921,N_21789,N_21627);
or U21922 (N_21922,N_21642,N_21617);
or U21923 (N_21923,N_21666,N_21706);
xor U21924 (N_21924,N_21614,N_21785);
nor U21925 (N_21925,N_21779,N_21777);
nand U21926 (N_21926,N_21696,N_21726);
nand U21927 (N_21927,N_21701,N_21754);
or U21928 (N_21928,N_21662,N_21668);
or U21929 (N_21929,N_21791,N_21618);
or U21930 (N_21930,N_21719,N_21795);
or U21931 (N_21931,N_21765,N_21661);
and U21932 (N_21932,N_21782,N_21751);
xor U21933 (N_21933,N_21728,N_21646);
and U21934 (N_21934,N_21706,N_21762);
nor U21935 (N_21935,N_21708,N_21742);
and U21936 (N_21936,N_21619,N_21604);
nor U21937 (N_21937,N_21632,N_21600);
xnor U21938 (N_21938,N_21769,N_21795);
nand U21939 (N_21939,N_21620,N_21630);
and U21940 (N_21940,N_21646,N_21676);
nor U21941 (N_21941,N_21664,N_21624);
and U21942 (N_21942,N_21632,N_21690);
nor U21943 (N_21943,N_21688,N_21669);
or U21944 (N_21944,N_21767,N_21788);
nand U21945 (N_21945,N_21759,N_21699);
nor U21946 (N_21946,N_21747,N_21758);
or U21947 (N_21947,N_21789,N_21652);
xnor U21948 (N_21948,N_21777,N_21663);
nand U21949 (N_21949,N_21796,N_21610);
nor U21950 (N_21950,N_21638,N_21668);
and U21951 (N_21951,N_21698,N_21691);
and U21952 (N_21952,N_21640,N_21773);
nand U21953 (N_21953,N_21767,N_21666);
nor U21954 (N_21954,N_21721,N_21681);
or U21955 (N_21955,N_21623,N_21749);
and U21956 (N_21956,N_21771,N_21796);
and U21957 (N_21957,N_21621,N_21749);
xnor U21958 (N_21958,N_21620,N_21676);
xor U21959 (N_21959,N_21780,N_21764);
nor U21960 (N_21960,N_21666,N_21659);
nor U21961 (N_21961,N_21658,N_21757);
nor U21962 (N_21962,N_21713,N_21741);
or U21963 (N_21963,N_21760,N_21610);
nand U21964 (N_21964,N_21763,N_21679);
xor U21965 (N_21965,N_21779,N_21789);
or U21966 (N_21966,N_21622,N_21772);
and U21967 (N_21967,N_21678,N_21734);
xor U21968 (N_21968,N_21746,N_21620);
xnor U21969 (N_21969,N_21734,N_21606);
xor U21970 (N_21970,N_21707,N_21754);
xnor U21971 (N_21971,N_21673,N_21785);
xnor U21972 (N_21972,N_21774,N_21626);
nor U21973 (N_21973,N_21786,N_21736);
and U21974 (N_21974,N_21796,N_21723);
nor U21975 (N_21975,N_21623,N_21707);
nand U21976 (N_21976,N_21614,N_21708);
and U21977 (N_21977,N_21779,N_21642);
or U21978 (N_21978,N_21638,N_21651);
and U21979 (N_21979,N_21635,N_21628);
nand U21980 (N_21980,N_21655,N_21630);
and U21981 (N_21981,N_21695,N_21684);
and U21982 (N_21982,N_21654,N_21643);
and U21983 (N_21983,N_21799,N_21701);
nor U21984 (N_21984,N_21646,N_21617);
nor U21985 (N_21985,N_21631,N_21674);
xor U21986 (N_21986,N_21651,N_21738);
nand U21987 (N_21987,N_21601,N_21655);
nand U21988 (N_21988,N_21766,N_21602);
and U21989 (N_21989,N_21758,N_21661);
nor U21990 (N_21990,N_21750,N_21796);
or U21991 (N_21991,N_21775,N_21659);
nand U21992 (N_21992,N_21660,N_21658);
xor U21993 (N_21993,N_21639,N_21732);
nand U21994 (N_21994,N_21621,N_21730);
nand U21995 (N_21995,N_21643,N_21792);
or U21996 (N_21996,N_21622,N_21729);
nor U21997 (N_21997,N_21730,N_21706);
nor U21998 (N_21998,N_21772,N_21704);
or U21999 (N_21999,N_21733,N_21762);
and U22000 (N_22000,N_21850,N_21954);
and U22001 (N_22001,N_21905,N_21846);
nor U22002 (N_22002,N_21822,N_21899);
xor U22003 (N_22003,N_21889,N_21897);
nand U22004 (N_22004,N_21828,N_21848);
and U22005 (N_22005,N_21935,N_21925);
and U22006 (N_22006,N_21867,N_21912);
xor U22007 (N_22007,N_21808,N_21929);
nor U22008 (N_22008,N_21900,N_21812);
nor U22009 (N_22009,N_21879,N_21964);
xor U22010 (N_22010,N_21920,N_21873);
nor U22011 (N_22011,N_21938,N_21986);
nand U22012 (N_22012,N_21818,N_21934);
nand U22013 (N_22013,N_21815,N_21977);
nand U22014 (N_22014,N_21824,N_21839);
nand U22015 (N_22015,N_21811,N_21999);
or U22016 (N_22016,N_21858,N_21872);
and U22017 (N_22017,N_21886,N_21971);
nor U22018 (N_22018,N_21864,N_21856);
xor U22019 (N_22019,N_21896,N_21805);
xnor U22020 (N_22020,N_21950,N_21882);
nor U22021 (N_22021,N_21926,N_21997);
or U22022 (N_22022,N_21831,N_21957);
xor U22023 (N_22023,N_21817,N_21992);
and U22024 (N_22024,N_21851,N_21809);
xnor U22025 (N_22025,N_21928,N_21940);
or U22026 (N_22026,N_21931,N_21984);
nand U22027 (N_22027,N_21843,N_21861);
and U22028 (N_22028,N_21918,N_21830);
and U22029 (N_22029,N_21901,N_21978);
nand U22030 (N_22030,N_21874,N_21813);
nand U22031 (N_22031,N_21945,N_21814);
and U22032 (N_22032,N_21884,N_21943);
xnor U22033 (N_22033,N_21942,N_21975);
nand U22034 (N_22034,N_21801,N_21859);
nand U22035 (N_22035,N_21883,N_21869);
nor U22036 (N_22036,N_21987,N_21832);
xor U22037 (N_22037,N_21835,N_21800);
xor U22038 (N_22038,N_21909,N_21949);
nand U22039 (N_22039,N_21821,N_21855);
nor U22040 (N_22040,N_21959,N_21904);
nand U22041 (N_22041,N_21870,N_21866);
or U22042 (N_22042,N_21910,N_21941);
nor U22043 (N_22043,N_21985,N_21982);
and U22044 (N_22044,N_21907,N_21952);
and U22045 (N_22045,N_21898,N_21963);
or U22046 (N_22046,N_21979,N_21988);
nand U22047 (N_22047,N_21939,N_21853);
and U22048 (N_22048,N_21823,N_21936);
and U22049 (N_22049,N_21930,N_21967);
nor U22050 (N_22050,N_21902,N_21960);
nand U22051 (N_22051,N_21948,N_21917);
nor U22052 (N_22052,N_21958,N_21807);
nand U22053 (N_22053,N_21955,N_21913);
xor U22054 (N_22054,N_21876,N_21944);
nor U22055 (N_22055,N_21996,N_21819);
nor U22056 (N_22056,N_21890,N_21842);
or U22057 (N_22057,N_21838,N_21933);
and U22058 (N_22058,N_21947,N_21994);
xor U22059 (N_22059,N_21919,N_21892);
or U22060 (N_22060,N_21966,N_21804);
or U22061 (N_22061,N_21860,N_21826);
and U22062 (N_22062,N_21946,N_21998);
nor U22063 (N_22063,N_21922,N_21923);
and U22064 (N_22064,N_21865,N_21837);
and U22065 (N_22065,N_21969,N_21962);
nor U22066 (N_22066,N_21983,N_21916);
xnor U22067 (N_22067,N_21834,N_21976);
or U22068 (N_22068,N_21810,N_21833);
xor U22069 (N_22069,N_21803,N_21915);
nand U22070 (N_22070,N_21951,N_21980);
xor U22071 (N_22071,N_21924,N_21816);
nor U22072 (N_22072,N_21991,N_21970);
nand U22073 (N_22073,N_21965,N_21820);
or U22074 (N_22074,N_21863,N_21868);
and U22075 (N_22075,N_21881,N_21911);
nor U22076 (N_22076,N_21891,N_21802);
nor U22077 (N_22077,N_21852,N_21877);
and U22078 (N_22078,N_21993,N_21906);
or U22079 (N_22079,N_21995,N_21880);
nand U22080 (N_22080,N_21887,N_21847);
or U22081 (N_22081,N_21893,N_21974);
nor U22082 (N_22082,N_21914,N_21968);
or U22083 (N_22083,N_21989,N_21854);
or U22084 (N_22084,N_21937,N_21961);
nand U22085 (N_22085,N_21921,N_21862);
xnor U22086 (N_22086,N_21836,N_21990);
and U22087 (N_22087,N_21840,N_21857);
xnor U22088 (N_22088,N_21829,N_21972);
nor U22089 (N_22089,N_21871,N_21827);
and U22090 (N_22090,N_21878,N_21849);
xnor U22091 (N_22091,N_21825,N_21903);
or U22092 (N_22092,N_21885,N_21875);
xor U22093 (N_22093,N_21973,N_21895);
or U22094 (N_22094,N_21845,N_21844);
nand U22095 (N_22095,N_21927,N_21908);
and U22096 (N_22096,N_21956,N_21841);
and U22097 (N_22097,N_21894,N_21953);
xnor U22098 (N_22098,N_21981,N_21932);
nand U22099 (N_22099,N_21806,N_21888);
nor U22100 (N_22100,N_21851,N_21845);
or U22101 (N_22101,N_21885,N_21972);
nor U22102 (N_22102,N_21822,N_21871);
and U22103 (N_22103,N_21960,N_21953);
nand U22104 (N_22104,N_21856,N_21969);
nor U22105 (N_22105,N_21963,N_21931);
or U22106 (N_22106,N_21848,N_21988);
or U22107 (N_22107,N_21884,N_21933);
nor U22108 (N_22108,N_21994,N_21928);
and U22109 (N_22109,N_21886,N_21978);
and U22110 (N_22110,N_21875,N_21952);
nand U22111 (N_22111,N_21994,N_21831);
nor U22112 (N_22112,N_21963,N_21956);
and U22113 (N_22113,N_21992,N_21872);
nor U22114 (N_22114,N_21945,N_21894);
xnor U22115 (N_22115,N_21989,N_21828);
nor U22116 (N_22116,N_21959,N_21937);
nor U22117 (N_22117,N_21849,N_21918);
nor U22118 (N_22118,N_21894,N_21935);
and U22119 (N_22119,N_21939,N_21975);
nand U22120 (N_22120,N_21993,N_21910);
nand U22121 (N_22121,N_21900,N_21964);
or U22122 (N_22122,N_21843,N_21868);
and U22123 (N_22123,N_21949,N_21814);
xor U22124 (N_22124,N_21939,N_21977);
nor U22125 (N_22125,N_21849,N_21880);
nor U22126 (N_22126,N_21994,N_21822);
nand U22127 (N_22127,N_21929,N_21995);
nor U22128 (N_22128,N_21940,N_21923);
or U22129 (N_22129,N_21891,N_21841);
nand U22130 (N_22130,N_21879,N_21847);
nand U22131 (N_22131,N_21870,N_21860);
xor U22132 (N_22132,N_21941,N_21983);
or U22133 (N_22133,N_21920,N_21883);
or U22134 (N_22134,N_21863,N_21809);
nand U22135 (N_22135,N_21979,N_21895);
or U22136 (N_22136,N_21994,N_21921);
xor U22137 (N_22137,N_21808,N_21974);
nor U22138 (N_22138,N_21955,N_21826);
or U22139 (N_22139,N_21869,N_21800);
and U22140 (N_22140,N_21906,N_21839);
nor U22141 (N_22141,N_21821,N_21980);
xor U22142 (N_22142,N_21841,N_21980);
or U22143 (N_22143,N_21905,N_21977);
nor U22144 (N_22144,N_21961,N_21863);
or U22145 (N_22145,N_21994,N_21866);
xnor U22146 (N_22146,N_21963,N_21921);
or U22147 (N_22147,N_21980,N_21833);
or U22148 (N_22148,N_21937,N_21819);
nor U22149 (N_22149,N_21878,N_21821);
nor U22150 (N_22150,N_21862,N_21983);
nand U22151 (N_22151,N_21962,N_21994);
nand U22152 (N_22152,N_21941,N_21832);
nor U22153 (N_22153,N_21900,N_21897);
xor U22154 (N_22154,N_21945,N_21918);
nor U22155 (N_22155,N_21915,N_21974);
and U22156 (N_22156,N_21822,N_21826);
nand U22157 (N_22157,N_21864,N_21944);
xnor U22158 (N_22158,N_21919,N_21896);
xor U22159 (N_22159,N_21964,N_21934);
nor U22160 (N_22160,N_21868,N_21898);
xnor U22161 (N_22161,N_21940,N_21948);
or U22162 (N_22162,N_21814,N_21996);
nor U22163 (N_22163,N_21818,N_21972);
xor U22164 (N_22164,N_21893,N_21991);
nor U22165 (N_22165,N_21868,N_21884);
and U22166 (N_22166,N_21917,N_21855);
xor U22167 (N_22167,N_21817,N_21883);
and U22168 (N_22168,N_21912,N_21971);
nor U22169 (N_22169,N_21830,N_21997);
and U22170 (N_22170,N_21866,N_21800);
xor U22171 (N_22171,N_21888,N_21964);
or U22172 (N_22172,N_21891,N_21997);
or U22173 (N_22173,N_21884,N_21823);
nand U22174 (N_22174,N_21811,N_21886);
nor U22175 (N_22175,N_21888,N_21855);
xor U22176 (N_22176,N_21979,N_21937);
nor U22177 (N_22177,N_21873,N_21976);
nand U22178 (N_22178,N_21835,N_21911);
nor U22179 (N_22179,N_21856,N_21886);
nand U22180 (N_22180,N_21826,N_21878);
nand U22181 (N_22181,N_21880,N_21811);
nor U22182 (N_22182,N_21920,N_21805);
and U22183 (N_22183,N_21977,N_21963);
xor U22184 (N_22184,N_21893,N_21852);
nor U22185 (N_22185,N_21967,N_21933);
nand U22186 (N_22186,N_21968,N_21913);
or U22187 (N_22187,N_21863,N_21851);
nand U22188 (N_22188,N_21829,N_21811);
nand U22189 (N_22189,N_21824,N_21971);
nor U22190 (N_22190,N_21839,N_21937);
or U22191 (N_22191,N_21884,N_21988);
or U22192 (N_22192,N_21908,N_21803);
xor U22193 (N_22193,N_21824,N_21924);
nor U22194 (N_22194,N_21933,N_21824);
and U22195 (N_22195,N_21937,N_21897);
and U22196 (N_22196,N_21966,N_21889);
nor U22197 (N_22197,N_21839,N_21866);
or U22198 (N_22198,N_21959,N_21842);
and U22199 (N_22199,N_21836,N_21992);
nor U22200 (N_22200,N_22082,N_22129);
or U22201 (N_22201,N_22101,N_22172);
xnor U22202 (N_22202,N_22152,N_22020);
and U22203 (N_22203,N_22125,N_22126);
nor U22204 (N_22204,N_22098,N_22102);
xnor U22205 (N_22205,N_22042,N_22182);
xnor U22206 (N_22206,N_22029,N_22060);
or U22207 (N_22207,N_22096,N_22059);
or U22208 (N_22208,N_22123,N_22167);
xor U22209 (N_22209,N_22108,N_22061);
nand U22210 (N_22210,N_22040,N_22012);
nand U22211 (N_22211,N_22033,N_22157);
nor U22212 (N_22212,N_22124,N_22047);
xor U22213 (N_22213,N_22168,N_22122);
and U22214 (N_22214,N_22189,N_22011);
or U22215 (N_22215,N_22018,N_22155);
or U22216 (N_22216,N_22142,N_22164);
nand U22217 (N_22217,N_22014,N_22071);
and U22218 (N_22218,N_22006,N_22087);
or U22219 (N_22219,N_22095,N_22002);
and U22220 (N_22220,N_22086,N_22174);
xnor U22221 (N_22221,N_22005,N_22092);
and U22222 (N_22222,N_22085,N_22003);
and U22223 (N_22223,N_22181,N_22066);
nand U22224 (N_22224,N_22056,N_22184);
and U22225 (N_22225,N_22022,N_22069);
and U22226 (N_22226,N_22032,N_22074);
xnor U22227 (N_22227,N_22171,N_22045);
xnor U22228 (N_22228,N_22105,N_22008);
xor U22229 (N_22229,N_22179,N_22063);
and U22230 (N_22230,N_22084,N_22013);
xor U22231 (N_22231,N_22099,N_22107);
or U22232 (N_22232,N_22038,N_22148);
xnor U22233 (N_22233,N_22178,N_22049);
nor U22234 (N_22234,N_22026,N_22106);
and U22235 (N_22235,N_22146,N_22076);
nor U22236 (N_22236,N_22068,N_22150);
or U22237 (N_22237,N_22058,N_22153);
xor U22238 (N_22238,N_22021,N_22057);
nand U22239 (N_22239,N_22162,N_22091);
and U22240 (N_22240,N_22139,N_22144);
nand U22241 (N_22241,N_22177,N_22185);
and U22242 (N_22242,N_22036,N_22024);
or U22243 (N_22243,N_22190,N_22134);
and U22244 (N_22244,N_22104,N_22143);
nor U22245 (N_22245,N_22065,N_22183);
and U22246 (N_22246,N_22009,N_22130);
xnor U22247 (N_22247,N_22193,N_22093);
and U22248 (N_22248,N_22050,N_22054);
and U22249 (N_22249,N_22111,N_22023);
or U22250 (N_22250,N_22016,N_22030);
nand U22251 (N_22251,N_22046,N_22180);
nand U22252 (N_22252,N_22132,N_22135);
nor U22253 (N_22253,N_22140,N_22044);
nor U22254 (N_22254,N_22119,N_22037);
xor U22255 (N_22255,N_22112,N_22160);
nor U22256 (N_22256,N_22118,N_22116);
xnor U22257 (N_22257,N_22070,N_22110);
or U22258 (N_22258,N_22034,N_22128);
xor U22259 (N_22259,N_22072,N_22080);
and U22260 (N_22260,N_22062,N_22192);
nor U22261 (N_22261,N_22100,N_22198);
xnor U22262 (N_22262,N_22053,N_22028);
or U22263 (N_22263,N_22141,N_22120);
xor U22264 (N_22264,N_22117,N_22176);
nand U22265 (N_22265,N_22136,N_22035);
xnor U22266 (N_22266,N_22131,N_22186);
nand U22267 (N_22267,N_22115,N_22194);
and U22268 (N_22268,N_22166,N_22170);
and U22269 (N_22269,N_22081,N_22083);
xnor U22270 (N_22270,N_22007,N_22145);
nand U22271 (N_22271,N_22078,N_22159);
or U22272 (N_22272,N_22051,N_22109);
and U22273 (N_22273,N_22048,N_22077);
nor U22274 (N_22274,N_22088,N_22075);
nor U22275 (N_22275,N_22137,N_22173);
nand U22276 (N_22276,N_22191,N_22158);
nand U22277 (N_22277,N_22025,N_22067);
xnor U22278 (N_22278,N_22094,N_22015);
and U22279 (N_22279,N_22175,N_22163);
xnor U22280 (N_22280,N_22103,N_22133);
nor U22281 (N_22281,N_22161,N_22019);
and U22282 (N_22282,N_22052,N_22041);
nor U22283 (N_22283,N_22169,N_22000);
nand U22284 (N_22284,N_22113,N_22127);
nor U22285 (N_22285,N_22154,N_22017);
nor U22286 (N_22286,N_22151,N_22001);
and U22287 (N_22287,N_22188,N_22089);
xnor U22288 (N_22288,N_22196,N_22147);
nand U22289 (N_22289,N_22197,N_22004);
xnor U22290 (N_22290,N_22073,N_22195);
nor U22291 (N_22291,N_22156,N_22043);
nor U22292 (N_22292,N_22097,N_22055);
nand U22293 (N_22293,N_22027,N_22187);
nand U22294 (N_22294,N_22079,N_22039);
or U22295 (N_22295,N_22114,N_22165);
xnor U22296 (N_22296,N_22090,N_22149);
nor U22297 (N_22297,N_22199,N_22031);
or U22298 (N_22298,N_22138,N_22121);
or U22299 (N_22299,N_22064,N_22010);
xor U22300 (N_22300,N_22054,N_22110);
nand U22301 (N_22301,N_22063,N_22188);
and U22302 (N_22302,N_22141,N_22128);
or U22303 (N_22303,N_22043,N_22003);
or U22304 (N_22304,N_22179,N_22170);
or U22305 (N_22305,N_22004,N_22161);
nor U22306 (N_22306,N_22195,N_22017);
nand U22307 (N_22307,N_22025,N_22130);
nand U22308 (N_22308,N_22118,N_22002);
and U22309 (N_22309,N_22057,N_22075);
and U22310 (N_22310,N_22000,N_22155);
or U22311 (N_22311,N_22186,N_22126);
nand U22312 (N_22312,N_22169,N_22053);
xnor U22313 (N_22313,N_22048,N_22181);
and U22314 (N_22314,N_22089,N_22198);
nand U22315 (N_22315,N_22043,N_22187);
or U22316 (N_22316,N_22146,N_22097);
and U22317 (N_22317,N_22062,N_22069);
xor U22318 (N_22318,N_22158,N_22193);
nor U22319 (N_22319,N_22028,N_22091);
xnor U22320 (N_22320,N_22121,N_22060);
or U22321 (N_22321,N_22021,N_22064);
nand U22322 (N_22322,N_22031,N_22066);
nor U22323 (N_22323,N_22104,N_22145);
nand U22324 (N_22324,N_22180,N_22145);
and U22325 (N_22325,N_22030,N_22116);
nor U22326 (N_22326,N_22018,N_22093);
and U22327 (N_22327,N_22036,N_22166);
and U22328 (N_22328,N_22072,N_22037);
and U22329 (N_22329,N_22051,N_22019);
xnor U22330 (N_22330,N_22070,N_22122);
nand U22331 (N_22331,N_22031,N_22189);
or U22332 (N_22332,N_22089,N_22189);
nor U22333 (N_22333,N_22047,N_22162);
xnor U22334 (N_22334,N_22028,N_22132);
xor U22335 (N_22335,N_22184,N_22018);
nor U22336 (N_22336,N_22175,N_22185);
nor U22337 (N_22337,N_22197,N_22122);
xnor U22338 (N_22338,N_22003,N_22160);
nand U22339 (N_22339,N_22065,N_22146);
or U22340 (N_22340,N_22058,N_22021);
or U22341 (N_22341,N_22103,N_22038);
xor U22342 (N_22342,N_22144,N_22156);
nand U22343 (N_22343,N_22122,N_22097);
and U22344 (N_22344,N_22182,N_22053);
xor U22345 (N_22345,N_22183,N_22015);
or U22346 (N_22346,N_22053,N_22146);
or U22347 (N_22347,N_22102,N_22159);
and U22348 (N_22348,N_22073,N_22025);
and U22349 (N_22349,N_22097,N_22113);
nor U22350 (N_22350,N_22156,N_22099);
nand U22351 (N_22351,N_22156,N_22111);
nand U22352 (N_22352,N_22143,N_22017);
or U22353 (N_22353,N_22067,N_22105);
nor U22354 (N_22354,N_22105,N_22029);
xnor U22355 (N_22355,N_22033,N_22069);
and U22356 (N_22356,N_22175,N_22194);
xnor U22357 (N_22357,N_22009,N_22053);
nand U22358 (N_22358,N_22013,N_22041);
nand U22359 (N_22359,N_22005,N_22034);
or U22360 (N_22360,N_22140,N_22117);
and U22361 (N_22361,N_22137,N_22041);
nor U22362 (N_22362,N_22167,N_22142);
nor U22363 (N_22363,N_22135,N_22046);
and U22364 (N_22364,N_22198,N_22036);
nor U22365 (N_22365,N_22158,N_22014);
nand U22366 (N_22366,N_22140,N_22120);
nand U22367 (N_22367,N_22096,N_22043);
nand U22368 (N_22368,N_22031,N_22017);
or U22369 (N_22369,N_22180,N_22194);
and U22370 (N_22370,N_22132,N_22169);
xnor U22371 (N_22371,N_22130,N_22170);
or U22372 (N_22372,N_22174,N_22050);
and U22373 (N_22373,N_22056,N_22136);
and U22374 (N_22374,N_22020,N_22044);
nor U22375 (N_22375,N_22142,N_22103);
xnor U22376 (N_22376,N_22047,N_22084);
nor U22377 (N_22377,N_22188,N_22000);
xnor U22378 (N_22378,N_22117,N_22097);
xor U22379 (N_22379,N_22071,N_22075);
nor U22380 (N_22380,N_22114,N_22091);
xor U22381 (N_22381,N_22060,N_22088);
and U22382 (N_22382,N_22112,N_22186);
and U22383 (N_22383,N_22160,N_22185);
or U22384 (N_22384,N_22043,N_22167);
nor U22385 (N_22385,N_22064,N_22188);
nand U22386 (N_22386,N_22055,N_22017);
nor U22387 (N_22387,N_22113,N_22112);
nor U22388 (N_22388,N_22058,N_22101);
or U22389 (N_22389,N_22115,N_22098);
or U22390 (N_22390,N_22164,N_22090);
or U22391 (N_22391,N_22122,N_22045);
nor U22392 (N_22392,N_22024,N_22101);
xor U22393 (N_22393,N_22188,N_22047);
or U22394 (N_22394,N_22080,N_22094);
or U22395 (N_22395,N_22029,N_22104);
or U22396 (N_22396,N_22107,N_22035);
or U22397 (N_22397,N_22137,N_22171);
xor U22398 (N_22398,N_22077,N_22015);
nand U22399 (N_22399,N_22189,N_22134);
or U22400 (N_22400,N_22283,N_22276);
nor U22401 (N_22401,N_22356,N_22364);
and U22402 (N_22402,N_22312,N_22357);
nor U22403 (N_22403,N_22223,N_22263);
xnor U22404 (N_22404,N_22385,N_22336);
and U22405 (N_22405,N_22320,N_22200);
nor U22406 (N_22406,N_22373,N_22203);
xor U22407 (N_22407,N_22360,N_22341);
and U22408 (N_22408,N_22350,N_22243);
nor U22409 (N_22409,N_22369,N_22308);
or U22410 (N_22410,N_22215,N_22287);
nor U22411 (N_22411,N_22207,N_22240);
xor U22412 (N_22412,N_22296,N_22208);
xor U22413 (N_22413,N_22268,N_22306);
and U22414 (N_22414,N_22251,N_22367);
xor U22415 (N_22415,N_22313,N_22374);
nor U22416 (N_22416,N_22294,N_22222);
xnor U22417 (N_22417,N_22214,N_22379);
nand U22418 (N_22418,N_22376,N_22236);
nand U22419 (N_22419,N_22278,N_22310);
nand U22420 (N_22420,N_22242,N_22372);
nor U22421 (N_22421,N_22212,N_22365);
nand U22422 (N_22422,N_22326,N_22238);
xor U22423 (N_22423,N_22246,N_22255);
and U22424 (N_22424,N_22322,N_22248);
nor U22425 (N_22425,N_22324,N_22217);
xnor U22426 (N_22426,N_22228,N_22247);
xor U22427 (N_22427,N_22388,N_22366);
nor U22428 (N_22428,N_22232,N_22381);
nand U22429 (N_22429,N_22302,N_22275);
nand U22430 (N_22430,N_22216,N_22351);
xnor U22431 (N_22431,N_22288,N_22269);
nor U22432 (N_22432,N_22270,N_22363);
or U22433 (N_22433,N_22397,N_22206);
nand U22434 (N_22434,N_22315,N_22256);
or U22435 (N_22435,N_22390,N_22375);
or U22436 (N_22436,N_22205,N_22301);
nand U22437 (N_22437,N_22224,N_22210);
or U22438 (N_22438,N_22259,N_22384);
xor U22439 (N_22439,N_22330,N_22202);
nand U22440 (N_22440,N_22264,N_22303);
and U22441 (N_22441,N_22359,N_22362);
nand U22442 (N_22442,N_22344,N_22337);
nand U22443 (N_22443,N_22258,N_22386);
or U22444 (N_22444,N_22234,N_22230);
nor U22445 (N_22445,N_22211,N_22305);
or U22446 (N_22446,N_22343,N_22391);
xor U22447 (N_22447,N_22281,N_22393);
or U22448 (N_22448,N_22395,N_22304);
or U22449 (N_22449,N_22358,N_22317);
xor U22450 (N_22450,N_22235,N_22289);
or U22451 (N_22451,N_22282,N_22332);
nor U22452 (N_22452,N_22231,N_22383);
or U22453 (N_22453,N_22273,N_22299);
nor U22454 (N_22454,N_22323,N_22314);
nand U22455 (N_22455,N_22318,N_22220);
nand U22456 (N_22456,N_22227,N_22257);
and U22457 (N_22457,N_22293,N_22345);
and U22458 (N_22458,N_22394,N_22290);
nor U22459 (N_22459,N_22307,N_22377);
xor U22460 (N_22460,N_22319,N_22254);
and U22461 (N_22461,N_22329,N_22298);
xnor U22462 (N_22462,N_22396,N_22285);
nand U22463 (N_22463,N_22219,N_22387);
or U22464 (N_22464,N_22213,N_22327);
and U22465 (N_22465,N_22286,N_22347);
nor U22466 (N_22466,N_22277,N_22368);
or U22467 (N_22467,N_22229,N_22218);
xnor U22468 (N_22468,N_22342,N_22309);
and U22469 (N_22469,N_22253,N_22201);
nor U22470 (N_22470,N_22292,N_22239);
nor U22471 (N_22471,N_22209,N_22295);
nor U22472 (N_22472,N_22245,N_22321);
nand U22473 (N_22473,N_22311,N_22353);
or U22474 (N_22474,N_22316,N_22266);
xor U22475 (N_22475,N_22333,N_22339);
or U22476 (N_22476,N_22280,N_22237);
nor U22477 (N_22477,N_22291,N_22241);
nand U22478 (N_22478,N_22221,N_22279);
nand U22479 (N_22479,N_22233,N_22348);
nor U22480 (N_22480,N_22378,N_22398);
xor U22481 (N_22481,N_22249,N_22328);
nand U22482 (N_22482,N_22297,N_22261);
or U22483 (N_22483,N_22335,N_22252);
and U22484 (N_22484,N_22274,N_22340);
xnor U22485 (N_22485,N_22260,N_22250);
nor U22486 (N_22486,N_22204,N_22399);
nor U22487 (N_22487,N_22334,N_22361);
or U22488 (N_22488,N_22382,N_22272);
nor U22489 (N_22489,N_22346,N_22389);
xor U22490 (N_22490,N_22244,N_22262);
and U22491 (N_22491,N_22352,N_22392);
or U22492 (N_22492,N_22370,N_22225);
nand U22493 (N_22493,N_22325,N_22371);
xnor U22494 (N_22494,N_22349,N_22380);
nand U22495 (N_22495,N_22300,N_22265);
nor U22496 (N_22496,N_22354,N_22267);
and U22497 (N_22497,N_22331,N_22226);
or U22498 (N_22498,N_22338,N_22271);
nand U22499 (N_22499,N_22355,N_22284);
or U22500 (N_22500,N_22329,N_22352);
and U22501 (N_22501,N_22225,N_22362);
and U22502 (N_22502,N_22292,N_22264);
nor U22503 (N_22503,N_22329,N_22291);
or U22504 (N_22504,N_22310,N_22381);
or U22505 (N_22505,N_22357,N_22259);
nor U22506 (N_22506,N_22207,N_22292);
nand U22507 (N_22507,N_22237,N_22340);
nor U22508 (N_22508,N_22232,N_22228);
xor U22509 (N_22509,N_22225,N_22320);
and U22510 (N_22510,N_22313,N_22290);
and U22511 (N_22511,N_22288,N_22247);
and U22512 (N_22512,N_22328,N_22261);
and U22513 (N_22513,N_22288,N_22362);
xnor U22514 (N_22514,N_22328,N_22201);
nand U22515 (N_22515,N_22262,N_22256);
nor U22516 (N_22516,N_22302,N_22240);
and U22517 (N_22517,N_22267,N_22297);
or U22518 (N_22518,N_22271,N_22363);
or U22519 (N_22519,N_22363,N_22372);
nand U22520 (N_22520,N_22330,N_22382);
and U22521 (N_22521,N_22393,N_22320);
xor U22522 (N_22522,N_22262,N_22319);
xor U22523 (N_22523,N_22368,N_22231);
nor U22524 (N_22524,N_22261,N_22249);
nor U22525 (N_22525,N_22321,N_22283);
nor U22526 (N_22526,N_22217,N_22281);
nand U22527 (N_22527,N_22226,N_22362);
nand U22528 (N_22528,N_22384,N_22359);
nor U22529 (N_22529,N_22266,N_22342);
and U22530 (N_22530,N_22388,N_22338);
xor U22531 (N_22531,N_22393,N_22295);
nor U22532 (N_22532,N_22375,N_22202);
or U22533 (N_22533,N_22361,N_22244);
and U22534 (N_22534,N_22231,N_22294);
and U22535 (N_22535,N_22258,N_22374);
nor U22536 (N_22536,N_22395,N_22350);
and U22537 (N_22537,N_22235,N_22270);
or U22538 (N_22538,N_22292,N_22236);
nor U22539 (N_22539,N_22285,N_22351);
xnor U22540 (N_22540,N_22232,N_22336);
xor U22541 (N_22541,N_22260,N_22392);
xnor U22542 (N_22542,N_22361,N_22287);
and U22543 (N_22543,N_22241,N_22362);
and U22544 (N_22544,N_22331,N_22368);
and U22545 (N_22545,N_22215,N_22231);
nand U22546 (N_22546,N_22243,N_22323);
and U22547 (N_22547,N_22346,N_22248);
nor U22548 (N_22548,N_22351,N_22321);
xnor U22549 (N_22549,N_22203,N_22284);
nor U22550 (N_22550,N_22240,N_22349);
nor U22551 (N_22551,N_22253,N_22278);
or U22552 (N_22552,N_22314,N_22237);
nand U22553 (N_22553,N_22236,N_22220);
nor U22554 (N_22554,N_22248,N_22399);
nand U22555 (N_22555,N_22289,N_22231);
or U22556 (N_22556,N_22358,N_22310);
or U22557 (N_22557,N_22246,N_22336);
nand U22558 (N_22558,N_22317,N_22348);
and U22559 (N_22559,N_22326,N_22224);
nor U22560 (N_22560,N_22359,N_22249);
nand U22561 (N_22561,N_22239,N_22316);
and U22562 (N_22562,N_22378,N_22269);
and U22563 (N_22563,N_22291,N_22282);
or U22564 (N_22564,N_22253,N_22250);
or U22565 (N_22565,N_22211,N_22313);
nor U22566 (N_22566,N_22253,N_22226);
and U22567 (N_22567,N_22281,N_22313);
and U22568 (N_22568,N_22370,N_22253);
nor U22569 (N_22569,N_22314,N_22267);
nor U22570 (N_22570,N_22228,N_22278);
nor U22571 (N_22571,N_22268,N_22373);
and U22572 (N_22572,N_22390,N_22204);
nand U22573 (N_22573,N_22272,N_22332);
nor U22574 (N_22574,N_22275,N_22325);
xor U22575 (N_22575,N_22204,N_22278);
nor U22576 (N_22576,N_22203,N_22394);
or U22577 (N_22577,N_22311,N_22386);
or U22578 (N_22578,N_22352,N_22274);
and U22579 (N_22579,N_22253,N_22347);
nor U22580 (N_22580,N_22364,N_22320);
or U22581 (N_22581,N_22296,N_22320);
or U22582 (N_22582,N_22393,N_22366);
xor U22583 (N_22583,N_22213,N_22299);
nor U22584 (N_22584,N_22298,N_22385);
and U22585 (N_22585,N_22311,N_22331);
nor U22586 (N_22586,N_22284,N_22274);
or U22587 (N_22587,N_22367,N_22291);
or U22588 (N_22588,N_22367,N_22372);
and U22589 (N_22589,N_22375,N_22221);
xnor U22590 (N_22590,N_22384,N_22354);
and U22591 (N_22591,N_22265,N_22297);
and U22592 (N_22592,N_22350,N_22237);
xnor U22593 (N_22593,N_22235,N_22390);
and U22594 (N_22594,N_22367,N_22304);
xor U22595 (N_22595,N_22329,N_22305);
nor U22596 (N_22596,N_22237,N_22298);
nor U22597 (N_22597,N_22224,N_22372);
xnor U22598 (N_22598,N_22280,N_22213);
xor U22599 (N_22599,N_22298,N_22327);
xnor U22600 (N_22600,N_22463,N_22581);
nor U22601 (N_22601,N_22579,N_22426);
nor U22602 (N_22602,N_22495,N_22575);
nor U22603 (N_22603,N_22589,N_22492);
nand U22604 (N_22604,N_22455,N_22508);
or U22605 (N_22605,N_22597,N_22442);
or U22606 (N_22606,N_22413,N_22428);
nand U22607 (N_22607,N_22480,N_22474);
nand U22608 (N_22608,N_22444,N_22598);
xor U22609 (N_22609,N_22411,N_22412);
nand U22610 (N_22610,N_22587,N_22502);
nand U22611 (N_22611,N_22530,N_22435);
or U22612 (N_22612,N_22562,N_22491);
nor U22613 (N_22613,N_22592,N_22448);
xnor U22614 (N_22614,N_22402,N_22570);
and U22615 (N_22615,N_22525,N_22542);
xnor U22616 (N_22616,N_22478,N_22445);
nor U22617 (N_22617,N_22487,N_22468);
nor U22618 (N_22618,N_22531,N_22522);
or U22619 (N_22619,N_22432,N_22509);
xnor U22620 (N_22620,N_22452,N_22471);
xor U22621 (N_22621,N_22582,N_22527);
nor U22622 (N_22622,N_22467,N_22573);
and U22623 (N_22623,N_22400,N_22594);
or U22624 (N_22624,N_22517,N_22528);
or U22625 (N_22625,N_22484,N_22519);
xnor U22626 (N_22626,N_22501,N_22585);
nand U22627 (N_22627,N_22456,N_22547);
or U22628 (N_22628,N_22567,N_22459);
or U22629 (N_22629,N_22511,N_22503);
xor U22630 (N_22630,N_22430,N_22533);
or U22631 (N_22631,N_22551,N_22417);
or U22632 (N_22632,N_22588,N_22544);
xor U22633 (N_22633,N_22524,N_22454);
xnor U22634 (N_22634,N_22566,N_22553);
nor U22635 (N_22635,N_22591,N_22541);
or U22636 (N_22636,N_22425,N_22434);
nor U22637 (N_22637,N_22469,N_22540);
and U22638 (N_22638,N_22559,N_22489);
nand U22639 (N_22639,N_22584,N_22496);
nand U22640 (N_22640,N_22409,N_22406);
nor U22641 (N_22641,N_22558,N_22596);
nor U22642 (N_22642,N_22583,N_22565);
nand U22643 (N_22643,N_22407,N_22554);
nor U22644 (N_22644,N_22537,N_22561);
or U22645 (N_22645,N_22479,N_22461);
nand U22646 (N_22646,N_22446,N_22521);
nand U22647 (N_22647,N_22595,N_22518);
nor U22648 (N_22648,N_22490,N_22408);
and U22649 (N_22649,N_22590,N_22534);
and U22650 (N_22650,N_22458,N_22539);
or U22651 (N_22651,N_22416,N_22440);
nand U22652 (N_22652,N_22564,N_22556);
and U22653 (N_22653,N_22488,N_22563);
nor U22654 (N_22654,N_22464,N_22493);
nand U22655 (N_22655,N_22451,N_22443);
and U22656 (N_22656,N_22538,N_22529);
xor U22657 (N_22657,N_22403,N_22462);
or U22658 (N_22658,N_22549,N_22569);
nor U22659 (N_22659,N_22580,N_22431);
or U22660 (N_22660,N_22404,N_22415);
nor U22661 (N_22661,N_22436,N_22470);
and U22662 (N_22662,N_22599,N_22548);
nor U22663 (N_22663,N_22593,N_22473);
nand U22664 (N_22664,N_22449,N_22552);
nor U22665 (N_22665,N_22523,N_22545);
or U22666 (N_22666,N_22405,N_22510);
or U22667 (N_22667,N_22500,N_22465);
nor U22668 (N_22668,N_22433,N_22512);
or U22669 (N_22669,N_22401,N_22577);
xor U22670 (N_22670,N_22520,N_22586);
xor U22671 (N_22671,N_22504,N_22576);
nand U22672 (N_22672,N_22423,N_22505);
or U22673 (N_22673,N_22543,N_22513);
nor U22674 (N_22674,N_22410,N_22472);
nor U22675 (N_22675,N_22421,N_22506);
nand U22676 (N_22676,N_22419,N_22532);
xnor U22677 (N_22677,N_22515,N_22497);
nand U22678 (N_22678,N_22572,N_22453);
or U22679 (N_22679,N_22475,N_22483);
or U22680 (N_22680,N_22526,N_22460);
xnor U22681 (N_22681,N_22574,N_22450);
nor U22682 (N_22682,N_22560,N_22477);
nand U22683 (N_22683,N_22438,N_22546);
and U22684 (N_22684,N_22494,N_22427);
and U22685 (N_22685,N_22420,N_22429);
or U22686 (N_22686,N_22476,N_22457);
nor U22687 (N_22687,N_22466,N_22557);
nor U22688 (N_22688,N_22507,N_22536);
nor U22689 (N_22689,N_22499,N_22555);
nor U22690 (N_22690,N_22578,N_22418);
xor U22691 (N_22691,N_22447,N_22535);
nor U22692 (N_22692,N_22437,N_22498);
nand U22693 (N_22693,N_22568,N_22414);
or U22694 (N_22694,N_22482,N_22439);
and U22695 (N_22695,N_22514,N_22441);
xor U22696 (N_22696,N_22485,N_22571);
nor U22697 (N_22697,N_22424,N_22550);
nand U22698 (N_22698,N_22486,N_22481);
nor U22699 (N_22699,N_22516,N_22422);
nor U22700 (N_22700,N_22475,N_22528);
and U22701 (N_22701,N_22510,N_22464);
or U22702 (N_22702,N_22544,N_22466);
nand U22703 (N_22703,N_22447,N_22470);
nand U22704 (N_22704,N_22595,N_22438);
or U22705 (N_22705,N_22564,N_22463);
nand U22706 (N_22706,N_22446,N_22558);
xor U22707 (N_22707,N_22526,N_22499);
nand U22708 (N_22708,N_22561,N_22571);
or U22709 (N_22709,N_22599,N_22559);
nor U22710 (N_22710,N_22464,N_22590);
or U22711 (N_22711,N_22428,N_22546);
or U22712 (N_22712,N_22471,N_22512);
nor U22713 (N_22713,N_22586,N_22599);
and U22714 (N_22714,N_22415,N_22575);
nor U22715 (N_22715,N_22571,N_22471);
or U22716 (N_22716,N_22486,N_22570);
and U22717 (N_22717,N_22490,N_22423);
nor U22718 (N_22718,N_22409,N_22411);
and U22719 (N_22719,N_22421,N_22449);
xor U22720 (N_22720,N_22478,N_22429);
nor U22721 (N_22721,N_22484,N_22442);
xnor U22722 (N_22722,N_22474,N_22537);
xor U22723 (N_22723,N_22542,N_22426);
or U22724 (N_22724,N_22434,N_22562);
nand U22725 (N_22725,N_22456,N_22513);
xnor U22726 (N_22726,N_22525,N_22527);
or U22727 (N_22727,N_22474,N_22464);
and U22728 (N_22728,N_22553,N_22596);
xor U22729 (N_22729,N_22549,N_22411);
or U22730 (N_22730,N_22481,N_22560);
or U22731 (N_22731,N_22583,N_22458);
nor U22732 (N_22732,N_22496,N_22498);
and U22733 (N_22733,N_22446,N_22564);
and U22734 (N_22734,N_22439,N_22404);
nor U22735 (N_22735,N_22549,N_22423);
and U22736 (N_22736,N_22555,N_22532);
and U22737 (N_22737,N_22497,N_22592);
and U22738 (N_22738,N_22582,N_22515);
and U22739 (N_22739,N_22447,N_22408);
and U22740 (N_22740,N_22550,N_22517);
nand U22741 (N_22741,N_22489,N_22453);
or U22742 (N_22742,N_22438,N_22464);
and U22743 (N_22743,N_22477,N_22406);
xor U22744 (N_22744,N_22463,N_22403);
and U22745 (N_22745,N_22504,N_22595);
nand U22746 (N_22746,N_22583,N_22517);
xor U22747 (N_22747,N_22512,N_22454);
nand U22748 (N_22748,N_22452,N_22451);
and U22749 (N_22749,N_22498,N_22460);
and U22750 (N_22750,N_22552,N_22528);
xnor U22751 (N_22751,N_22458,N_22509);
xor U22752 (N_22752,N_22499,N_22409);
nand U22753 (N_22753,N_22413,N_22493);
nand U22754 (N_22754,N_22566,N_22442);
nand U22755 (N_22755,N_22572,N_22593);
or U22756 (N_22756,N_22444,N_22463);
xor U22757 (N_22757,N_22561,N_22591);
and U22758 (N_22758,N_22526,N_22512);
xnor U22759 (N_22759,N_22428,N_22486);
and U22760 (N_22760,N_22428,N_22455);
nand U22761 (N_22761,N_22409,N_22527);
xor U22762 (N_22762,N_22548,N_22594);
nand U22763 (N_22763,N_22510,N_22475);
xnor U22764 (N_22764,N_22503,N_22462);
nand U22765 (N_22765,N_22449,N_22471);
or U22766 (N_22766,N_22580,N_22559);
xor U22767 (N_22767,N_22568,N_22421);
nor U22768 (N_22768,N_22488,N_22569);
and U22769 (N_22769,N_22537,N_22585);
and U22770 (N_22770,N_22532,N_22516);
xnor U22771 (N_22771,N_22430,N_22543);
and U22772 (N_22772,N_22583,N_22441);
nor U22773 (N_22773,N_22467,N_22594);
or U22774 (N_22774,N_22414,N_22435);
xnor U22775 (N_22775,N_22450,N_22487);
nand U22776 (N_22776,N_22445,N_22451);
nand U22777 (N_22777,N_22452,N_22526);
and U22778 (N_22778,N_22404,N_22588);
or U22779 (N_22779,N_22505,N_22445);
or U22780 (N_22780,N_22414,N_22547);
and U22781 (N_22781,N_22455,N_22405);
and U22782 (N_22782,N_22518,N_22566);
nor U22783 (N_22783,N_22437,N_22442);
and U22784 (N_22784,N_22569,N_22437);
or U22785 (N_22785,N_22594,N_22422);
or U22786 (N_22786,N_22448,N_22586);
xor U22787 (N_22787,N_22487,N_22415);
nand U22788 (N_22788,N_22575,N_22501);
xor U22789 (N_22789,N_22421,N_22518);
or U22790 (N_22790,N_22518,N_22413);
or U22791 (N_22791,N_22480,N_22500);
or U22792 (N_22792,N_22542,N_22547);
or U22793 (N_22793,N_22540,N_22530);
nor U22794 (N_22794,N_22510,N_22555);
nand U22795 (N_22795,N_22519,N_22599);
or U22796 (N_22796,N_22403,N_22511);
nand U22797 (N_22797,N_22514,N_22428);
or U22798 (N_22798,N_22465,N_22468);
nand U22799 (N_22799,N_22455,N_22581);
xor U22800 (N_22800,N_22666,N_22610);
and U22801 (N_22801,N_22646,N_22723);
nor U22802 (N_22802,N_22710,N_22632);
nor U22803 (N_22803,N_22675,N_22604);
nor U22804 (N_22804,N_22640,N_22649);
nand U22805 (N_22805,N_22644,N_22655);
nor U22806 (N_22806,N_22707,N_22794);
and U22807 (N_22807,N_22722,N_22629);
nand U22808 (N_22808,N_22763,N_22661);
nor U22809 (N_22809,N_22663,N_22688);
nor U22810 (N_22810,N_22698,N_22636);
and U22811 (N_22811,N_22695,N_22779);
xnor U22812 (N_22812,N_22713,N_22602);
and U22813 (N_22813,N_22678,N_22738);
and U22814 (N_22814,N_22671,N_22674);
xor U22815 (N_22815,N_22743,N_22765);
nand U22816 (N_22816,N_22751,N_22694);
xor U22817 (N_22817,N_22630,N_22603);
xnor U22818 (N_22818,N_22641,N_22732);
nand U22819 (N_22819,N_22787,N_22623);
xor U22820 (N_22820,N_22783,N_22611);
xnor U22821 (N_22821,N_22731,N_22650);
nand U22822 (N_22822,N_22760,N_22778);
and U22823 (N_22823,N_22672,N_22659);
xnor U22824 (N_22824,N_22724,N_22797);
or U22825 (N_22825,N_22616,N_22648);
xnor U22826 (N_22826,N_22615,N_22761);
and U22827 (N_22827,N_22740,N_22622);
nor U22828 (N_22828,N_22653,N_22711);
or U22829 (N_22829,N_22658,N_22733);
nand U22830 (N_22830,N_22709,N_22749);
nor U22831 (N_22831,N_22638,N_22752);
or U22832 (N_22832,N_22617,N_22756);
xnor U22833 (N_22833,N_22728,N_22725);
nand U22834 (N_22834,N_22795,N_22634);
nand U22835 (N_22835,N_22796,N_22750);
nor U22836 (N_22836,N_22748,N_22645);
nor U22837 (N_22837,N_22764,N_22799);
or U22838 (N_22838,N_22618,N_22777);
and U22839 (N_22839,N_22626,N_22793);
or U22840 (N_22840,N_22770,N_22633);
or U22841 (N_22841,N_22759,N_22716);
xor U22842 (N_22842,N_22746,N_22656);
xnor U22843 (N_22843,N_22687,N_22792);
and U22844 (N_22844,N_22670,N_22775);
nand U22845 (N_22845,N_22665,N_22774);
or U22846 (N_22846,N_22657,N_22766);
or U22847 (N_22847,N_22621,N_22753);
nand U22848 (N_22848,N_22662,N_22668);
or U22849 (N_22849,N_22647,N_22681);
nand U22850 (N_22850,N_22608,N_22721);
nand U22851 (N_22851,N_22789,N_22696);
nand U22852 (N_22852,N_22669,N_22685);
or U22853 (N_22853,N_22736,N_22677);
or U22854 (N_22854,N_22625,N_22673);
xor U22855 (N_22855,N_22734,N_22693);
or U22856 (N_22856,N_22697,N_22742);
nor U22857 (N_22857,N_22691,N_22773);
xnor U22858 (N_22858,N_22660,N_22741);
nand U22859 (N_22859,N_22757,N_22717);
nor U22860 (N_22860,N_22600,N_22624);
and U22861 (N_22861,N_22754,N_22613);
or U22862 (N_22862,N_22790,N_22703);
nor U22863 (N_22863,N_22654,N_22686);
and U22864 (N_22864,N_22784,N_22780);
nand U22865 (N_22865,N_22768,N_22683);
or U22866 (N_22866,N_22719,N_22706);
nor U22867 (N_22867,N_22676,N_22712);
xor U22868 (N_22868,N_22771,N_22781);
nand U22869 (N_22869,N_22607,N_22758);
or U22870 (N_22870,N_22744,N_22680);
nand U22871 (N_22871,N_22619,N_22737);
or U22872 (N_22872,N_22692,N_22729);
nor U22873 (N_22873,N_22628,N_22715);
and U22874 (N_22874,N_22612,N_22652);
and U22875 (N_22875,N_22605,N_22701);
and U22876 (N_22876,N_22679,N_22702);
nand U22877 (N_22877,N_22714,N_22690);
xnor U22878 (N_22878,N_22767,N_22747);
or U22879 (N_22879,N_22772,N_22689);
and U22880 (N_22880,N_22708,N_22620);
nor U22881 (N_22881,N_22798,N_22684);
or U22882 (N_22882,N_22601,N_22664);
nand U22883 (N_22883,N_22762,N_22727);
nand U22884 (N_22884,N_22704,N_22782);
nor U22885 (N_22885,N_22609,N_22631);
and U22886 (N_22886,N_22769,N_22699);
nor U22887 (N_22887,N_22735,N_22720);
nand U22888 (N_22888,N_22776,N_22739);
nand U22889 (N_22889,N_22643,N_22730);
or U22890 (N_22890,N_22700,N_22606);
nand U22891 (N_22891,N_22667,N_22718);
and U22892 (N_22892,N_22785,N_22755);
nand U22893 (N_22893,N_22639,N_22705);
and U22894 (N_22894,N_22726,N_22682);
nand U22895 (N_22895,N_22637,N_22642);
and U22896 (N_22896,N_22791,N_22786);
nand U22897 (N_22897,N_22651,N_22614);
xnor U22898 (N_22898,N_22635,N_22627);
or U22899 (N_22899,N_22788,N_22745);
nand U22900 (N_22900,N_22668,N_22602);
and U22901 (N_22901,N_22657,N_22661);
or U22902 (N_22902,N_22608,N_22694);
and U22903 (N_22903,N_22617,N_22611);
nor U22904 (N_22904,N_22670,N_22660);
and U22905 (N_22905,N_22779,N_22602);
nand U22906 (N_22906,N_22717,N_22726);
nor U22907 (N_22907,N_22785,N_22737);
and U22908 (N_22908,N_22710,N_22601);
or U22909 (N_22909,N_22792,N_22778);
nor U22910 (N_22910,N_22729,N_22682);
and U22911 (N_22911,N_22789,N_22723);
xor U22912 (N_22912,N_22618,N_22766);
xnor U22913 (N_22913,N_22782,N_22787);
nor U22914 (N_22914,N_22620,N_22758);
and U22915 (N_22915,N_22715,N_22723);
or U22916 (N_22916,N_22716,N_22638);
xor U22917 (N_22917,N_22769,N_22793);
xor U22918 (N_22918,N_22683,N_22757);
nand U22919 (N_22919,N_22676,N_22761);
or U22920 (N_22920,N_22691,N_22729);
nor U22921 (N_22921,N_22602,N_22613);
xnor U22922 (N_22922,N_22732,N_22788);
and U22923 (N_22923,N_22691,N_22726);
or U22924 (N_22924,N_22642,N_22748);
or U22925 (N_22925,N_22616,N_22602);
nor U22926 (N_22926,N_22782,N_22726);
xor U22927 (N_22927,N_22725,N_22624);
or U22928 (N_22928,N_22686,N_22645);
nand U22929 (N_22929,N_22625,N_22658);
xor U22930 (N_22930,N_22779,N_22723);
nor U22931 (N_22931,N_22752,N_22748);
or U22932 (N_22932,N_22730,N_22618);
nor U22933 (N_22933,N_22681,N_22791);
or U22934 (N_22934,N_22617,N_22634);
xor U22935 (N_22935,N_22688,N_22774);
nor U22936 (N_22936,N_22600,N_22718);
nand U22937 (N_22937,N_22690,N_22786);
and U22938 (N_22938,N_22727,N_22797);
or U22939 (N_22939,N_22620,N_22756);
nand U22940 (N_22940,N_22770,N_22727);
nand U22941 (N_22941,N_22782,N_22683);
nand U22942 (N_22942,N_22611,N_22684);
xor U22943 (N_22943,N_22726,N_22634);
xor U22944 (N_22944,N_22769,N_22690);
xnor U22945 (N_22945,N_22606,N_22792);
nand U22946 (N_22946,N_22705,N_22607);
or U22947 (N_22947,N_22670,N_22621);
nor U22948 (N_22948,N_22750,N_22714);
or U22949 (N_22949,N_22641,N_22786);
nor U22950 (N_22950,N_22798,N_22736);
nand U22951 (N_22951,N_22780,N_22708);
nor U22952 (N_22952,N_22774,N_22619);
nor U22953 (N_22953,N_22746,N_22760);
nand U22954 (N_22954,N_22697,N_22799);
or U22955 (N_22955,N_22602,N_22672);
or U22956 (N_22956,N_22737,N_22718);
xnor U22957 (N_22957,N_22741,N_22626);
or U22958 (N_22958,N_22722,N_22667);
or U22959 (N_22959,N_22711,N_22671);
nor U22960 (N_22960,N_22753,N_22762);
nand U22961 (N_22961,N_22666,N_22702);
or U22962 (N_22962,N_22782,N_22618);
nand U22963 (N_22963,N_22752,N_22610);
xnor U22964 (N_22964,N_22673,N_22714);
and U22965 (N_22965,N_22729,N_22782);
nor U22966 (N_22966,N_22733,N_22742);
and U22967 (N_22967,N_22743,N_22673);
nor U22968 (N_22968,N_22638,N_22785);
nor U22969 (N_22969,N_22643,N_22661);
xnor U22970 (N_22970,N_22724,N_22785);
nand U22971 (N_22971,N_22650,N_22606);
xor U22972 (N_22972,N_22771,N_22601);
nand U22973 (N_22973,N_22650,N_22601);
and U22974 (N_22974,N_22675,N_22708);
nor U22975 (N_22975,N_22711,N_22714);
xnor U22976 (N_22976,N_22617,N_22664);
xnor U22977 (N_22977,N_22662,N_22612);
xor U22978 (N_22978,N_22684,N_22715);
xnor U22979 (N_22979,N_22744,N_22739);
and U22980 (N_22980,N_22753,N_22693);
nor U22981 (N_22981,N_22632,N_22699);
nor U22982 (N_22982,N_22780,N_22713);
nand U22983 (N_22983,N_22780,N_22660);
nor U22984 (N_22984,N_22786,N_22649);
nor U22985 (N_22985,N_22790,N_22721);
xnor U22986 (N_22986,N_22723,N_22703);
and U22987 (N_22987,N_22758,N_22736);
nor U22988 (N_22988,N_22715,N_22692);
xor U22989 (N_22989,N_22729,N_22762);
nand U22990 (N_22990,N_22645,N_22659);
nor U22991 (N_22991,N_22638,N_22632);
nor U22992 (N_22992,N_22639,N_22632);
and U22993 (N_22993,N_22664,N_22663);
nand U22994 (N_22994,N_22764,N_22717);
nand U22995 (N_22995,N_22714,N_22670);
nor U22996 (N_22996,N_22743,N_22738);
xor U22997 (N_22997,N_22707,N_22710);
nor U22998 (N_22998,N_22640,N_22708);
or U22999 (N_22999,N_22790,N_22651);
nand U23000 (N_23000,N_22901,N_22843);
or U23001 (N_23001,N_22904,N_22871);
nand U23002 (N_23002,N_22846,N_22937);
xnor U23003 (N_23003,N_22854,N_22995);
and U23004 (N_23004,N_22918,N_22897);
or U23005 (N_23005,N_22845,N_22863);
nor U23006 (N_23006,N_22864,N_22900);
and U23007 (N_23007,N_22932,N_22824);
nor U23008 (N_23008,N_22808,N_22917);
nor U23009 (N_23009,N_22923,N_22964);
and U23010 (N_23010,N_22956,N_22892);
or U23011 (N_23011,N_22967,N_22860);
nor U23012 (N_23012,N_22942,N_22936);
nand U23013 (N_23013,N_22998,N_22895);
nor U23014 (N_23014,N_22896,N_22806);
and U23015 (N_23015,N_22838,N_22939);
or U23016 (N_23016,N_22906,N_22934);
nor U23017 (N_23017,N_22841,N_22966);
nand U23018 (N_23018,N_22868,N_22893);
or U23019 (N_23019,N_22850,N_22877);
or U23020 (N_23020,N_22872,N_22993);
nor U23021 (N_23021,N_22980,N_22867);
nand U23022 (N_23022,N_22840,N_22801);
nor U23023 (N_23023,N_22870,N_22800);
nor U23024 (N_23024,N_22990,N_22945);
or U23025 (N_23025,N_22954,N_22855);
or U23026 (N_23026,N_22999,N_22914);
nand U23027 (N_23027,N_22834,N_22813);
nand U23028 (N_23028,N_22852,N_22804);
nor U23029 (N_23029,N_22924,N_22888);
and U23030 (N_23030,N_22989,N_22958);
xnor U23031 (N_23031,N_22984,N_22884);
xnor U23032 (N_23032,N_22886,N_22988);
nor U23033 (N_23033,N_22873,N_22816);
or U23034 (N_23034,N_22920,N_22902);
xnor U23035 (N_23035,N_22817,N_22869);
and U23036 (N_23036,N_22981,N_22927);
xnor U23037 (N_23037,N_22825,N_22851);
or U23038 (N_23038,N_22905,N_22982);
xnor U23039 (N_23039,N_22879,N_22856);
nor U23040 (N_23040,N_22826,N_22944);
or U23041 (N_23041,N_22987,N_22970);
xor U23042 (N_23042,N_22894,N_22887);
nor U23043 (N_23043,N_22857,N_22926);
and U23044 (N_23044,N_22880,N_22885);
nor U23045 (N_23045,N_22922,N_22889);
and U23046 (N_23046,N_22823,N_22890);
xnor U23047 (N_23047,N_22865,N_22968);
nor U23048 (N_23048,N_22812,N_22961);
nand U23049 (N_23049,N_22916,N_22910);
nand U23050 (N_23050,N_22819,N_22952);
or U23051 (N_23051,N_22940,N_22882);
nand U23052 (N_23052,N_22875,N_22960);
and U23053 (N_23053,N_22811,N_22802);
nor U23054 (N_23054,N_22946,N_22947);
and U23055 (N_23055,N_22925,N_22849);
and U23056 (N_23056,N_22977,N_22876);
or U23057 (N_23057,N_22941,N_22909);
nor U23058 (N_23058,N_22949,N_22997);
or U23059 (N_23059,N_22836,N_22818);
and U23060 (N_23060,N_22842,N_22815);
or U23061 (N_23061,N_22837,N_22943);
nor U23062 (N_23062,N_22891,N_22828);
nand U23063 (N_23063,N_22874,N_22844);
and U23064 (N_23064,N_22976,N_22833);
nor U23065 (N_23065,N_22861,N_22907);
or U23066 (N_23066,N_22959,N_22963);
or U23067 (N_23067,N_22994,N_22996);
and U23068 (N_23068,N_22955,N_22809);
nor U23069 (N_23069,N_22950,N_22935);
nor U23070 (N_23070,N_22908,N_22832);
nand U23071 (N_23071,N_22866,N_22911);
and U23072 (N_23072,N_22919,N_22962);
nor U23073 (N_23073,N_22973,N_22830);
nand U23074 (N_23074,N_22829,N_22821);
and U23075 (N_23075,N_22975,N_22931);
and U23076 (N_23076,N_22847,N_22858);
nor U23077 (N_23077,N_22969,N_22898);
xnor U23078 (N_23078,N_22965,N_22848);
nor U23079 (N_23079,N_22915,N_22912);
nor U23080 (N_23080,N_22913,N_22979);
or U23081 (N_23081,N_22807,N_22938);
or U23082 (N_23082,N_22953,N_22862);
or U23083 (N_23083,N_22951,N_22985);
nor U23084 (N_23084,N_22803,N_22948);
nor U23085 (N_23085,N_22859,N_22814);
nor U23086 (N_23086,N_22928,N_22810);
and U23087 (N_23087,N_22957,N_22883);
xor U23088 (N_23088,N_22820,N_22878);
or U23089 (N_23089,N_22853,N_22992);
xor U23090 (N_23090,N_22835,N_22921);
nand U23091 (N_23091,N_22978,N_22933);
nor U23092 (N_23092,N_22881,N_22805);
or U23093 (N_23093,N_22831,N_22974);
nand U23094 (N_23094,N_22971,N_22991);
or U23095 (N_23095,N_22930,N_22827);
nor U23096 (N_23096,N_22983,N_22972);
nor U23097 (N_23097,N_22903,N_22929);
or U23098 (N_23098,N_22822,N_22839);
nand U23099 (N_23099,N_22899,N_22986);
nand U23100 (N_23100,N_22923,N_22849);
xor U23101 (N_23101,N_22909,N_22929);
xor U23102 (N_23102,N_22855,N_22978);
nor U23103 (N_23103,N_22932,N_22853);
nor U23104 (N_23104,N_22832,N_22960);
xor U23105 (N_23105,N_22892,N_22962);
and U23106 (N_23106,N_22852,N_22982);
or U23107 (N_23107,N_22890,N_22985);
nand U23108 (N_23108,N_22907,N_22851);
or U23109 (N_23109,N_22875,N_22928);
nand U23110 (N_23110,N_22885,N_22987);
and U23111 (N_23111,N_22836,N_22908);
or U23112 (N_23112,N_22970,N_22833);
nor U23113 (N_23113,N_22872,N_22850);
and U23114 (N_23114,N_22846,N_22971);
xor U23115 (N_23115,N_22995,N_22809);
nor U23116 (N_23116,N_22881,N_22915);
and U23117 (N_23117,N_22865,N_22991);
nor U23118 (N_23118,N_22944,N_22867);
or U23119 (N_23119,N_22998,N_22942);
or U23120 (N_23120,N_22896,N_22906);
xnor U23121 (N_23121,N_22952,N_22959);
xor U23122 (N_23122,N_22946,N_22994);
and U23123 (N_23123,N_22928,N_22994);
or U23124 (N_23124,N_22881,N_22997);
nand U23125 (N_23125,N_22941,N_22987);
nor U23126 (N_23126,N_22912,N_22997);
and U23127 (N_23127,N_22928,N_22900);
and U23128 (N_23128,N_22989,N_22957);
and U23129 (N_23129,N_22955,N_22835);
nor U23130 (N_23130,N_22822,N_22874);
nor U23131 (N_23131,N_22881,N_22913);
nand U23132 (N_23132,N_22997,N_22988);
or U23133 (N_23133,N_22968,N_22841);
and U23134 (N_23134,N_22915,N_22937);
nor U23135 (N_23135,N_22938,N_22924);
and U23136 (N_23136,N_22894,N_22922);
nor U23137 (N_23137,N_22959,N_22978);
or U23138 (N_23138,N_22832,N_22940);
nand U23139 (N_23139,N_22860,N_22871);
nor U23140 (N_23140,N_22896,N_22853);
and U23141 (N_23141,N_22945,N_22847);
nor U23142 (N_23142,N_22971,N_22858);
nand U23143 (N_23143,N_22975,N_22895);
xnor U23144 (N_23144,N_22924,N_22997);
nor U23145 (N_23145,N_22955,N_22865);
nor U23146 (N_23146,N_22992,N_22815);
nor U23147 (N_23147,N_22885,N_22839);
and U23148 (N_23148,N_22992,N_22956);
or U23149 (N_23149,N_22848,N_22886);
xor U23150 (N_23150,N_22949,N_22833);
and U23151 (N_23151,N_22841,N_22962);
nor U23152 (N_23152,N_22902,N_22960);
or U23153 (N_23153,N_22829,N_22843);
nand U23154 (N_23154,N_22877,N_22833);
xor U23155 (N_23155,N_22967,N_22890);
nand U23156 (N_23156,N_22965,N_22865);
nor U23157 (N_23157,N_22813,N_22892);
nor U23158 (N_23158,N_22802,N_22825);
and U23159 (N_23159,N_22858,N_22871);
and U23160 (N_23160,N_22914,N_22815);
xor U23161 (N_23161,N_22824,N_22979);
or U23162 (N_23162,N_22994,N_22966);
nand U23163 (N_23163,N_22843,N_22880);
nand U23164 (N_23164,N_22870,N_22945);
nor U23165 (N_23165,N_22812,N_22951);
nand U23166 (N_23166,N_22827,N_22854);
nand U23167 (N_23167,N_22983,N_22958);
nand U23168 (N_23168,N_22904,N_22958);
nor U23169 (N_23169,N_22901,N_22902);
and U23170 (N_23170,N_22871,N_22926);
xnor U23171 (N_23171,N_22834,N_22877);
and U23172 (N_23172,N_22894,N_22912);
or U23173 (N_23173,N_22848,N_22972);
or U23174 (N_23174,N_22941,N_22918);
nand U23175 (N_23175,N_22964,N_22808);
xnor U23176 (N_23176,N_22856,N_22904);
or U23177 (N_23177,N_22804,N_22840);
nand U23178 (N_23178,N_22851,N_22858);
nand U23179 (N_23179,N_22816,N_22867);
nor U23180 (N_23180,N_22930,N_22831);
and U23181 (N_23181,N_22901,N_22999);
nand U23182 (N_23182,N_22824,N_22927);
and U23183 (N_23183,N_22826,N_22890);
xor U23184 (N_23184,N_22970,N_22912);
or U23185 (N_23185,N_22991,N_22962);
xnor U23186 (N_23186,N_22841,N_22893);
and U23187 (N_23187,N_22997,N_22873);
and U23188 (N_23188,N_22878,N_22906);
xor U23189 (N_23189,N_22886,N_22981);
and U23190 (N_23190,N_22810,N_22935);
or U23191 (N_23191,N_22822,N_22884);
xor U23192 (N_23192,N_22857,N_22940);
and U23193 (N_23193,N_22900,N_22991);
nand U23194 (N_23194,N_22915,N_22893);
nor U23195 (N_23195,N_22964,N_22810);
nor U23196 (N_23196,N_22984,N_22890);
xnor U23197 (N_23197,N_22861,N_22955);
nor U23198 (N_23198,N_22961,N_22950);
and U23199 (N_23199,N_22871,N_22813);
nand U23200 (N_23200,N_23139,N_23008);
nand U23201 (N_23201,N_23084,N_23050);
xnor U23202 (N_23202,N_23114,N_23130);
nand U23203 (N_23203,N_23106,N_23075);
or U23204 (N_23204,N_23023,N_23198);
and U23205 (N_23205,N_23081,N_23040);
xor U23206 (N_23206,N_23067,N_23027);
nor U23207 (N_23207,N_23115,N_23068);
xnor U23208 (N_23208,N_23090,N_23007);
or U23209 (N_23209,N_23042,N_23053);
and U23210 (N_23210,N_23048,N_23142);
nand U23211 (N_23211,N_23145,N_23051);
nand U23212 (N_23212,N_23095,N_23160);
and U23213 (N_23213,N_23178,N_23055);
xor U23214 (N_23214,N_23118,N_23119);
nor U23215 (N_23215,N_23158,N_23013);
nand U23216 (N_23216,N_23073,N_23127);
xor U23217 (N_23217,N_23021,N_23110);
and U23218 (N_23218,N_23020,N_23086);
nor U23219 (N_23219,N_23098,N_23022);
nand U23220 (N_23220,N_23132,N_23060);
nor U23221 (N_23221,N_23174,N_23025);
and U23222 (N_23222,N_23093,N_23173);
xnor U23223 (N_23223,N_23169,N_23177);
or U23224 (N_23224,N_23011,N_23175);
nand U23225 (N_23225,N_23168,N_23097);
and U23226 (N_23226,N_23144,N_23038);
nor U23227 (N_23227,N_23116,N_23187);
nor U23228 (N_23228,N_23030,N_23165);
nor U23229 (N_23229,N_23141,N_23015);
nand U23230 (N_23230,N_23078,N_23059);
nor U23231 (N_23231,N_23140,N_23171);
xor U23232 (N_23232,N_23049,N_23151);
xnor U23233 (N_23233,N_23157,N_23192);
xor U23234 (N_23234,N_23083,N_23072);
xor U23235 (N_23235,N_23191,N_23080);
nor U23236 (N_23236,N_23052,N_23149);
and U23237 (N_23237,N_23143,N_23193);
xnor U23238 (N_23238,N_23172,N_23071);
or U23239 (N_23239,N_23131,N_23159);
or U23240 (N_23240,N_23056,N_23096);
and U23241 (N_23241,N_23170,N_23146);
xnor U23242 (N_23242,N_23079,N_23010);
or U23243 (N_23243,N_23111,N_23188);
nor U23244 (N_23244,N_23112,N_23091);
xnor U23245 (N_23245,N_23102,N_23100);
nand U23246 (N_23246,N_23189,N_23137);
or U23247 (N_23247,N_23125,N_23005);
nor U23248 (N_23248,N_23087,N_23129);
and U23249 (N_23249,N_23152,N_23164);
and U23250 (N_23250,N_23092,N_23028);
and U23251 (N_23251,N_23155,N_23181);
or U23252 (N_23252,N_23121,N_23122);
xnor U23253 (N_23253,N_23043,N_23004);
xnor U23254 (N_23254,N_23162,N_23179);
nand U23255 (N_23255,N_23085,N_23031);
xnor U23256 (N_23256,N_23006,N_23166);
nor U23257 (N_23257,N_23014,N_23103);
and U23258 (N_23258,N_23065,N_23045);
or U23259 (N_23259,N_23018,N_23182);
or U23260 (N_23260,N_23154,N_23150);
nor U23261 (N_23261,N_23044,N_23126);
or U23262 (N_23262,N_23047,N_23120);
xor U23263 (N_23263,N_23016,N_23077);
nor U23264 (N_23264,N_23058,N_23037);
and U23265 (N_23265,N_23123,N_23147);
xnor U23266 (N_23266,N_23076,N_23185);
nor U23267 (N_23267,N_23190,N_23017);
nor U23268 (N_23268,N_23026,N_23064);
or U23269 (N_23269,N_23046,N_23135);
and U23270 (N_23270,N_23134,N_23066);
or U23271 (N_23271,N_23167,N_23186);
xor U23272 (N_23272,N_23197,N_23032);
xor U23273 (N_23273,N_23196,N_23148);
nand U23274 (N_23274,N_23113,N_23036);
nand U23275 (N_23275,N_23128,N_23104);
and U23276 (N_23276,N_23041,N_23183);
xor U23277 (N_23277,N_23089,N_23199);
nor U23278 (N_23278,N_23109,N_23029);
nor U23279 (N_23279,N_23180,N_23107);
nor U23280 (N_23280,N_23061,N_23156);
or U23281 (N_23281,N_23108,N_23070);
nor U23282 (N_23282,N_23124,N_23133);
or U23283 (N_23283,N_23062,N_23002);
xor U23284 (N_23284,N_23138,N_23099);
or U23285 (N_23285,N_23024,N_23074);
and U23286 (N_23286,N_23057,N_23117);
xnor U23287 (N_23287,N_23034,N_23063);
nand U23288 (N_23288,N_23039,N_23019);
or U23289 (N_23289,N_23088,N_23069);
or U23290 (N_23290,N_23176,N_23054);
nor U23291 (N_23291,N_23094,N_23161);
nor U23292 (N_23292,N_23153,N_23009);
xor U23293 (N_23293,N_23136,N_23035);
xnor U23294 (N_23294,N_23194,N_23000);
and U23295 (N_23295,N_23001,N_23184);
or U23296 (N_23296,N_23033,N_23003);
and U23297 (N_23297,N_23163,N_23195);
nor U23298 (N_23298,N_23105,N_23082);
xor U23299 (N_23299,N_23012,N_23101);
and U23300 (N_23300,N_23014,N_23013);
nand U23301 (N_23301,N_23110,N_23199);
nand U23302 (N_23302,N_23103,N_23016);
xnor U23303 (N_23303,N_23018,N_23187);
and U23304 (N_23304,N_23171,N_23042);
or U23305 (N_23305,N_23086,N_23070);
nor U23306 (N_23306,N_23099,N_23080);
and U23307 (N_23307,N_23043,N_23018);
xnor U23308 (N_23308,N_23195,N_23063);
and U23309 (N_23309,N_23032,N_23072);
and U23310 (N_23310,N_23024,N_23067);
xor U23311 (N_23311,N_23094,N_23157);
xnor U23312 (N_23312,N_23172,N_23047);
nand U23313 (N_23313,N_23048,N_23004);
or U23314 (N_23314,N_23032,N_23056);
and U23315 (N_23315,N_23129,N_23107);
and U23316 (N_23316,N_23130,N_23173);
nor U23317 (N_23317,N_23165,N_23198);
xnor U23318 (N_23318,N_23031,N_23151);
xor U23319 (N_23319,N_23057,N_23089);
nand U23320 (N_23320,N_23148,N_23191);
nand U23321 (N_23321,N_23089,N_23093);
or U23322 (N_23322,N_23056,N_23060);
nand U23323 (N_23323,N_23181,N_23146);
and U23324 (N_23324,N_23149,N_23016);
or U23325 (N_23325,N_23104,N_23072);
nand U23326 (N_23326,N_23119,N_23094);
or U23327 (N_23327,N_23034,N_23097);
xor U23328 (N_23328,N_23025,N_23078);
and U23329 (N_23329,N_23098,N_23017);
xnor U23330 (N_23330,N_23130,N_23132);
and U23331 (N_23331,N_23115,N_23064);
nand U23332 (N_23332,N_23014,N_23197);
nand U23333 (N_23333,N_23085,N_23059);
nor U23334 (N_23334,N_23186,N_23147);
or U23335 (N_23335,N_23158,N_23187);
xor U23336 (N_23336,N_23150,N_23000);
xor U23337 (N_23337,N_23175,N_23187);
xnor U23338 (N_23338,N_23053,N_23124);
xnor U23339 (N_23339,N_23005,N_23016);
nand U23340 (N_23340,N_23137,N_23097);
and U23341 (N_23341,N_23177,N_23122);
or U23342 (N_23342,N_23035,N_23050);
or U23343 (N_23343,N_23071,N_23119);
nor U23344 (N_23344,N_23122,N_23093);
nand U23345 (N_23345,N_23196,N_23123);
nor U23346 (N_23346,N_23121,N_23139);
or U23347 (N_23347,N_23198,N_23195);
and U23348 (N_23348,N_23101,N_23093);
nor U23349 (N_23349,N_23172,N_23074);
and U23350 (N_23350,N_23121,N_23091);
or U23351 (N_23351,N_23189,N_23114);
or U23352 (N_23352,N_23104,N_23199);
and U23353 (N_23353,N_23098,N_23100);
nor U23354 (N_23354,N_23043,N_23072);
nand U23355 (N_23355,N_23107,N_23182);
and U23356 (N_23356,N_23194,N_23133);
or U23357 (N_23357,N_23060,N_23015);
nor U23358 (N_23358,N_23017,N_23040);
and U23359 (N_23359,N_23067,N_23010);
nor U23360 (N_23360,N_23183,N_23129);
and U23361 (N_23361,N_23199,N_23105);
or U23362 (N_23362,N_23190,N_23136);
xor U23363 (N_23363,N_23002,N_23145);
xor U23364 (N_23364,N_23037,N_23014);
nand U23365 (N_23365,N_23177,N_23184);
xnor U23366 (N_23366,N_23018,N_23140);
or U23367 (N_23367,N_23042,N_23070);
and U23368 (N_23368,N_23038,N_23098);
nor U23369 (N_23369,N_23067,N_23022);
and U23370 (N_23370,N_23125,N_23104);
nand U23371 (N_23371,N_23033,N_23062);
nor U23372 (N_23372,N_23195,N_23010);
or U23373 (N_23373,N_23133,N_23183);
or U23374 (N_23374,N_23003,N_23192);
or U23375 (N_23375,N_23114,N_23176);
xnor U23376 (N_23376,N_23067,N_23095);
and U23377 (N_23377,N_23134,N_23033);
and U23378 (N_23378,N_23181,N_23108);
xor U23379 (N_23379,N_23019,N_23114);
or U23380 (N_23380,N_23173,N_23136);
or U23381 (N_23381,N_23077,N_23025);
nor U23382 (N_23382,N_23044,N_23091);
nand U23383 (N_23383,N_23031,N_23120);
or U23384 (N_23384,N_23113,N_23137);
nor U23385 (N_23385,N_23035,N_23081);
and U23386 (N_23386,N_23044,N_23191);
nand U23387 (N_23387,N_23001,N_23161);
and U23388 (N_23388,N_23039,N_23058);
xnor U23389 (N_23389,N_23111,N_23187);
or U23390 (N_23390,N_23138,N_23096);
and U23391 (N_23391,N_23076,N_23173);
and U23392 (N_23392,N_23010,N_23061);
nand U23393 (N_23393,N_23029,N_23180);
nor U23394 (N_23394,N_23125,N_23028);
and U23395 (N_23395,N_23147,N_23143);
xnor U23396 (N_23396,N_23030,N_23197);
nor U23397 (N_23397,N_23010,N_23091);
and U23398 (N_23398,N_23102,N_23158);
xor U23399 (N_23399,N_23064,N_23081);
nand U23400 (N_23400,N_23285,N_23335);
nor U23401 (N_23401,N_23333,N_23374);
xnor U23402 (N_23402,N_23211,N_23379);
or U23403 (N_23403,N_23318,N_23316);
or U23404 (N_23404,N_23219,N_23358);
nand U23405 (N_23405,N_23224,N_23385);
xor U23406 (N_23406,N_23399,N_23209);
nand U23407 (N_23407,N_23249,N_23254);
or U23408 (N_23408,N_23215,N_23227);
xor U23409 (N_23409,N_23206,N_23246);
or U23410 (N_23410,N_23299,N_23326);
or U23411 (N_23411,N_23245,N_23323);
or U23412 (N_23412,N_23300,N_23322);
xor U23413 (N_23413,N_23330,N_23359);
xor U23414 (N_23414,N_23336,N_23252);
and U23415 (N_23415,N_23368,N_23370);
or U23416 (N_23416,N_23353,N_23364);
xnor U23417 (N_23417,N_23208,N_23216);
nand U23418 (N_23418,N_23390,N_23205);
xnor U23419 (N_23419,N_23233,N_23345);
and U23420 (N_23420,N_23306,N_23223);
nand U23421 (N_23421,N_23260,N_23229);
nor U23422 (N_23422,N_23262,N_23239);
nand U23423 (N_23423,N_23220,N_23301);
xnor U23424 (N_23424,N_23349,N_23283);
xnor U23425 (N_23425,N_23331,N_23352);
or U23426 (N_23426,N_23291,N_23253);
nand U23427 (N_23427,N_23392,N_23321);
xnor U23428 (N_23428,N_23210,N_23391);
xnor U23429 (N_23429,N_23338,N_23369);
nor U23430 (N_23430,N_23373,N_23398);
nand U23431 (N_23431,N_23228,N_23313);
or U23432 (N_23432,N_23248,N_23356);
nand U23433 (N_23433,N_23389,N_23367);
nor U23434 (N_23434,N_23222,N_23225);
nand U23435 (N_23435,N_23271,N_23381);
xor U23436 (N_23436,N_23270,N_23341);
nand U23437 (N_23437,N_23231,N_23397);
nor U23438 (N_23438,N_23320,N_23337);
xor U23439 (N_23439,N_23311,N_23268);
nor U23440 (N_23440,N_23278,N_23242);
xor U23441 (N_23441,N_23396,N_23334);
xor U23442 (N_23442,N_23363,N_23376);
and U23443 (N_23443,N_23332,N_23236);
or U23444 (N_23444,N_23212,N_23281);
nor U23445 (N_23445,N_23290,N_23273);
nor U23446 (N_23446,N_23383,N_23366);
nand U23447 (N_23447,N_23380,N_23394);
xor U23448 (N_23448,N_23204,N_23234);
or U23449 (N_23449,N_23258,N_23214);
or U23450 (N_23450,N_23339,N_23276);
and U23451 (N_23451,N_23365,N_23264);
xor U23452 (N_23452,N_23378,N_23267);
nand U23453 (N_23453,N_23296,N_23342);
xor U23454 (N_23454,N_23256,N_23232);
xnor U23455 (N_23455,N_23304,N_23298);
or U23456 (N_23456,N_23388,N_23202);
or U23457 (N_23457,N_23257,N_23360);
nor U23458 (N_23458,N_23293,N_23226);
nor U23459 (N_23459,N_23348,N_23277);
and U23460 (N_23460,N_23375,N_23269);
nor U23461 (N_23461,N_23305,N_23251);
xor U23462 (N_23462,N_23307,N_23286);
nand U23463 (N_23463,N_23218,N_23382);
xnor U23464 (N_23464,N_23325,N_23312);
nand U23465 (N_23465,N_23247,N_23302);
nor U23466 (N_23466,N_23265,N_23310);
nor U23467 (N_23467,N_23272,N_23250);
and U23468 (N_23468,N_23327,N_23279);
and U23469 (N_23469,N_23203,N_23384);
and U23470 (N_23470,N_23395,N_23354);
or U23471 (N_23471,N_23238,N_23207);
nand U23472 (N_23472,N_23213,N_23328);
nand U23473 (N_23473,N_23259,N_23362);
and U23474 (N_23474,N_23237,N_23309);
or U23475 (N_23475,N_23371,N_23372);
xor U23476 (N_23476,N_23340,N_23357);
nor U23477 (N_23477,N_23221,N_23217);
nand U23478 (N_23478,N_23274,N_23355);
xnor U23479 (N_23479,N_23315,N_23263);
or U23480 (N_23480,N_23280,N_23351);
nor U23481 (N_23481,N_23308,N_23387);
or U23482 (N_23482,N_23377,N_23346);
and U23483 (N_23483,N_23317,N_23347);
nor U23484 (N_23484,N_23287,N_23261);
xor U23485 (N_23485,N_23200,N_23329);
and U23486 (N_23486,N_23255,N_23324);
nor U23487 (N_23487,N_23201,N_23393);
nand U23488 (N_23488,N_23275,N_23244);
xnor U23489 (N_23489,N_23295,N_23297);
nor U23490 (N_23490,N_23319,N_23241);
nand U23491 (N_23491,N_23350,N_23284);
or U23492 (N_23492,N_23344,N_23303);
nand U23493 (N_23493,N_23266,N_23230);
nand U23494 (N_23494,N_23243,N_23343);
xor U23495 (N_23495,N_23292,N_23386);
and U23496 (N_23496,N_23294,N_23282);
and U23497 (N_23497,N_23314,N_23235);
or U23498 (N_23498,N_23240,N_23289);
xnor U23499 (N_23499,N_23361,N_23288);
xor U23500 (N_23500,N_23313,N_23369);
xor U23501 (N_23501,N_23240,N_23244);
nand U23502 (N_23502,N_23392,N_23239);
or U23503 (N_23503,N_23323,N_23394);
or U23504 (N_23504,N_23390,N_23353);
nand U23505 (N_23505,N_23268,N_23233);
or U23506 (N_23506,N_23384,N_23270);
nor U23507 (N_23507,N_23281,N_23269);
nor U23508 (N_23508,N_23394,N_23266);
and U23509 (N_23509,N_23291,N_23290);
nor U23510 (N_23510,N_23205,N_23251);
nand U23511 (N_23511,N_23321,N_23347);
and U23512 (N_23512,N_23305,N_23311);
nand U23513 (N_23513,N_23325,N_23226);
nor U23514 (N_23514,N_23325,N_23269);
nor U23515 (N_23515,N_23382,N_23338);
xor U23516 (N_23516,N_23324,N_23223);
xnor U23517 (N_23517,N_23301,N_23336);
and U23518 (N_23518,N_23346,N_23214);
xnor U23519 (N_23519,N_23388,N_23298);
nor U23520 (N_23520,N_23310,N_23273);
nand U23521 (N_23521,N_23328,N_23388);
and U23522 (N_23522,N_23300,N_23216);
xnor U23523 (N_23523,N_23309,N_23376);
and U23524 (N_23524,N_23357,N_23349);
xnor U23525 (N_23525,N_23229,N_23356);
or U23526 (N_23526,N_23299,N_23338);
and U23527 (N_23527,N_23204,N_23212);
nand U23528 (N_23528,N_23305,N_23241);
or U23529 (N_23529,N_23341,N_23280);
and U23530 (N_23530,N_23258,N_23305);
xor U23531 (N_23531,N_23253,N_23219);
or U23532 (N_23532,N_23288,N_23367);
or U23533 (N_23533,N_23294,N_23368);
nand U23534 (N_23534,N_23297,N_23223);
xor U23535 (N_23535,N_23224,N_23326);
nand U23536 (N_23536,N_23332,N_23224);
xnor U23537 (N_23537,N_23260,N_23254);
nor U23538 (N_23538,N_23240,N_23253);
nand U23539 (N_23539,N_23272,N_23323);
and U23540 (N_23540,N_23371,N_23255);
nor U23541 (N_23541,N_23204,N_23299);
xor U23542 (N_23542,N_23372,N_23253);
or U23543 (N_23543,N_23299,N_23276);
nor U23544 (N_23544,N_23277,N_23368);
nand U23545 (N_23545,N_23367,N_23269);
xnor U23546 (N_23546,N_23385,N_23311);
xnor U23547 (N_23547,N_23297,N_23293);
and U23548 (N_23548,N_23252,N_23344);
nand U23549 (N_23549,N_23285,N_23298);
xor U23550 (N_23550,N_23321,N_23268);
xnor U23551 (N_23551,N_23327,N_23208);
or U23552 (N_23552,N_23221,N_23299);
nor U23553 (N_23553,N_23395,N_23257);
xor U23554 (N_23554,N_23239,N_23293);
nand U23555 (N_23555,N_23212,N_23287);
nand U23556 (N_23556,N_23213,N_23207);
or U23557 (N_23557,N_23219,N_23379);
or U23558 (N_23558,N_23317,N_23346);
nor U23559 (N_23559,N_23277,N_23294);
xnor U23560 (N_23560,N_23275,N_23227);
or U23561 (N_23561,N_23204,N_23243);
nor U23562 (N_23562,N_23388,N_23316);
and U23563 (N_23563,N_23269,N_23342);
nand U23564 (N_23564,N_23305,N_23385);
xnor U23565 (N_23565,N_23304,N_23329);
and U23566 (N_23566,N_23258,N_23359);
and U23567 (N_23567,N_23209,N_23396);
and U23568 (N_23568,N_23217,N_23301);
nand U23569 (N_23569,N_23248,N_23290);
nand U23570 (N_23570,N_23206,N_23327);
nand U23571 (N_23571,N_23296,N_23204);
nor U23572 (N_23572,N_23326,N_23281);
xnor U23573 (N_23573,N_23300,N_23278);
and U23574 (N_23574,N_23298,N_23371);
nor U23575 (N_23575,N_23297,N_23268);
and U23576 (N_23576,N_23396,N_23339);
nor U23577 (N_23577,N_23256,N_23328);
and U23578 (N_23578,N_23201,N_23322);
nor U23579 (N_23579,N_23295,N_23242);
nand U23580 (N_23580,N_23378,N_23392);
nand U23581 (N_23581,N_23295,N_23300);
and U23582 (N_23582,N_23330,N_23250);
nor U23583 (N_23583,N_23269,N_23396);
or U23584 (N_23584,N_23245,N_23357);
nand U23585 (N_23585,N_23202,N_23355);
and U23586 (N_23586,N_23215,N_23366);
or U23587 (N_23587,N_23386,N_23351);
xnor U23588 (N_23588,N_23264,N_23296);
and U23589 (N_23589,N_23246,N_23262);
or U23590 (N_23590,N_23211,N_23343);
xor U23591 (N_23591,N_23359,N_23265);
or U23592 (N_23592,N_23248,N_23313);
nand U23593 (N_23593,N_23364,N_23282);
or U23594 (N_23594,N_23391,N_23378);
nor U23595 (N_23595,N_23345,N_23330);
nand U23596 (N_23596,N_23313,N_23214);
xnor U23597 (N_23597,N_23305,N_23247);
and U23598 (N_23598,N_23217,N_23312);
nand U23599 (N_23599,N_23320,N_23310);
nand U23600 (N_23600,N_23435,N_23494);
or U23601 (N_23601,N_23597,N_23577);
nand U23602 (N_23602,N_23485,N_23493);
and U23603 (N_23603,N_23456,N_23587);
or U23604 (N_23604,N_23559,N_23421);
nor U23605 (N_23605,N_23560,N_23512);
nor U23606 (N_23606,N_23442,N_23578);
and U23607 (N_23607,N_23558,N_23572);
xor U23608 (N_23608,N_23490,N_23404);
and U23609 (N_23609,N_23489,N_23424);
nor U23610 (N_23610,N_23486,N_23444);
nor U23611 (N_23611,N_23551,N_23488);
xnor U23612 (N_23612,N_23418,N_23570);
nor U23613 (N_23613,N_23466,N_23415);
nand U23614 (N_23614,N_23440,N_23509);
nand U23615 (N_23615,N_23542,N_23417);
nor U23616 (N_23616,N_23410,N_23580);
nor U23617 (N_23617,N_23487,N_23450);
and U23618 (N_23618,N_23402,N_23514);
and U23619 (N_23619,N_23596,N_23441);
or U23620 (N_23620,N_23430,N_23481);
nand U23621 (N_23621,N_23594,N_23518);
xnor U23622 (N_23622,N_23403,N_23423);
nor U23623 (N_23623,N_23477,N_23476);
or U23624 (N_23624,N_23503,N_23540);
or U23625 (N_23625,N_23567,N_23555);
or U23626 (N_23626,N_23561,N_23407);
xor U23627 (N_23627,N_23523,N_23504);
and U23628 (N_23628,N_23516,N_23508);
and U23629 (N_23629,N_23557,N_23443);
nand U23630 (N_23630,N_23547,N_23491);
and U23631 (N_23631,N_23453,N_23433);
xnor U23632 (N_23632,N_23529,N_23521);
xnor U23633 (N_23633,N_23452,N_23536);
nand U23634 (N_23634,N_23549,N_23499);
nand U23635 (N_23635,N_23590,N_23531);
and U23636 (N_23636,N_23591,N_23544);
nand U23637 (N_23637,N_23585,N_23501);
nand U23638 (N_23638,N_23473,N_23537);
or U23639 (N_23639,N_23552,N_23470);
xnor U23640 (N_23640,N_23538,N_23511);
xnor U23641 (N_23641,N_23575,N_23554);
and U23642 (N_23642,N_23569,N_23405);
or U23643 (N_23643,N_23586,N_23474);
or U23644 (N_23644,N_23520,N_23465);
nand U23645 (N_23645,N_23454,N_23507);
or U23646 (N_23646,N_23460,N_23427);
or U23647 (N_23647,N_23583,N_23513);
nor U23648 (N_23648,N_23522,N_23582);
nor U23649 (N_23649,N_23546,N_23439);
xor U23650 (N_23650,N_23550,N_23445);
nor U23651 (N_23651,N_23406,N_23446);
nor U23652 (N_23652,N_23479,N_23553);
xnor U23653 (N_23653,N_23451,N_23588);
nand U23654 (N_23654,N_23497,N_23595);
nand U23655 (N_23655,N_23478,N_23471);
and U23656 (N_23656,N_23496,N_23419);
xor U23657 (N_23657,N_23416,N_23401);
xnor U23658 (N_23658,N_23498,N_23457);
nand U23659 (N_23659,N_23535,N_23464);
and U23660 (N_23660,N_23431,N_23467);
or U23661 (N_23661,N_23564,N_23425);
and U23662 (N_23662,N_23436,N_23434);
xnor U23663 (N_23663,N_23475,N_23400);
nand U23664 (N_23664,N_23469,N_23472);
or U23665 (N_23665,N_23524,N_23429);
xor U23666 (N_23666,N_23574,N_23432);
nor U23667 (N_23667,N_23562,N_23563);
or U23668 (N_23668,N_23447,N_23539);
and U23669 (N_23669,N_23599,N_23420);
or U23670 (N_23670,N_23571,N_23455);
nor U23671 (N_23671,N_23527,N_23533);
nand U23672 (N_23672,N_23581,N_23573);
or U23673 (N_23673,N_23565,N_23530);
nand U23674 (N_23674,N_23449,N_23480);
nor U23675 (N_23675,N_23426,N_23422);
xnor U23676 (N_23676,N_23506,N_23589);
or U23677 (N_23677,N_23532,N_23468);
nand U23678 (N_23678,N_23438,N_23505);
nand U23679 (N_23679,N_23566,N_23408);
xor U23680 (N_23680,N_23576,N_23579);
and U23681 (N_23681,N_23411,N_23517);
nand U23682 (N_23682,N_23541,N_23495);
and U23683 (N_23683,N_23556,N_23548);
and U23684 (N_23684,N_23500,N_23483);
and U23685 (N_23685,N_23592,N_23545);
and U23686 (N_23686,N_23428,N_23459);
xnor U23687 (N_23687,N_23519,N_23482);
and U23688 (N_23688,N_23593,N_23413);
and U23689 (N_23689,N_23534,N_23409);
nor U23690 (N_23690,N_23515,N_23502);
xnor U23691 (N_23691,N_23526,N_23492);
xor U23692 (N_23692,N_23448,N_23463);
nor U23693 (N_23693,N_23528,N_23543);
or U23694 (N_23694,N_23510,N_23525);
and U23695 (N_23695,N_23598,N_23462);
xor U23696 (N_23696,N_23412,N_23437);
nor U23697 (N_23697,N_23584,N_23458);
and U23698 (N_23698,N_23461,N_23568);
or U23699 (N_23699,N_23484,N_23414);
or U23700 (N_23700,N_23463,N_23507);
xnor U23701 (N_23701,N_23464,N_23525);
nor U23702 (N_23702,N_23505,N_23593);
and U23703 (N_23703,N_23560,N_23551);
nor U23704 (N_23704,N_23490,N_23479);
and U23705 (N_23705,N_23500,N_23405);
nand U23706 (N_23706,N_23450,N_23486);
nand U23707 (N_23707,N_23472,N_23468);
and U23708 (N_23708,N_23555,N_23538);
and U23709 (N_23709,N_23481,N_23500);
and U23710 (N_23710,N_23567,N_23444);
nand U23711 (N_23711,N_23577,N_23464);
nor U23712 (N_23712,N_23592,N_23574);
nand U23713 (N_23713,N_23422,N_23540);
and U23714 (N_23714,N_23432,N_23596);
nor U23715 (N_23715,N_23510,N_23580);
nor U23716 (N_23716,N_23536,N_23448);
or U23717 (N_23717,N_23495,N_23427);
nor U23718 (N_23718,N_23413,N_23420);
and U23719 (N_23719,N_23433,N_23404);
xnor U23720 (N_23720,N_23404,N_23477);
nor U23721 (N_23721,N_23543,N_23479);
or U23722 (N_23722,N_23406,N_23597);
or U23723 (N_23723,N_23523,N_23525);
xor U23724 (N_23724,N_23510,N_23421);
or U23725 (N_23725,N_23414,N_23551);
xor U23726 (N_23726,N_23545,N_23405);
and U23727 (N_23727,N_23536,N_23405);
xor U23728 (N_23728,N_23517,N_23467);
nor U23729 (N_23729,N_23478,N_23441);
nor U23730 (N_23730,N_23552,N_23444);
xor U23731 (N_23731,N_23457,N_23486);
nand U23732 (N_23732,N_23411,N_23591);
and U23733 (N_23733,N_23471,N_23459);
xnor U23734 (N_23734,N_23582,N_23470);
xnor U23735 (N_23735,N_23489,N_23474);
nand U23736 (N_23736,N_23473,N_23574);
nor U23737 (N_23737,N_23496,N_23415);
and U23738 (N_23738,N_23424,N_23482);
or U23739 (N_23739,N_23421,N_23540);
xnor U23740 (N_23740,N_23458,N_23476);
xnor U23741 (N_23741,N_23557,N_23483);
xor U23742 (N_23742,N_23413,N_23405);
xnor U23743 (N_23743,N_23536,N_23413);
and U23744 (N_23744,N_23499,N_23579);
or U23745 (N_23745,N_23478,N_23546);
or U23746 (N_23746,N_23512,N_23486);
or U23747 (N_23747,N_23562,N_23401);
nor U23748 (N_23748,N_23548,N_23413);
or U23749 (N_23749,N_23528,N_23576);
and U23750 (N_23750,N_23491,N_23437);
nor U23751 (N_23751,N_23518,N_23477);
and U23752 (N_23752,N_23545,N_23436);
xnor U23753 (N_23753,N_23572,N_23419);
and U23754 (N_23754,N_23417,N_23484);
or U23755 (N_23755,N_23451,N_23578);
nand U23756 (N_23756,N_23409,N_23446);
nor U23757 (N_23757,N_23442,N_23459);
or U23758 (N_23758,N_23557,N_23572);
nand U23759 (N_23759,N_23502,N_23469);
nor U23760 (N_23760,N_23599,N_23471);
or U23761 (N_23761,N_23479,N_23546);
nor U23762 (N_23762,N_23449,N_23509);
nor U23763 (N_23763,N_23400,N_23531);
xor U23764 (N_23764,N_23449,N_23458);
or U23765 (N_23765,N_23551,N_23463);
and U23766 (N_23766,N_23414,N_23548);
and U23767 (N_23767,N_23529,N_23576);
nor U23768 (N_23768,N_23569,N_23422);
nor U23769 (N_23769,N_23490,N_23538);
nand U23770 (N_23770,N_23423,N_23418);
nand U23771 (N_23771,N_23507,N_23515);
or U23772 (N_23772,N_23414,N_23450);
nand U23773 (N_23773,N_23574,N_23438);
and U23774 (N_23774,N_23478,N_23464);
and U23775 (N_23775,N_23486,N_23432);
xnor U23776 (N_23776,N_23528,N_23508);
xor U23777 (N_23777,N_23428,N_23424);
or U23778 (N_23778,N_23479,N_23489);
xnor U23779 (N_23779,N_23480,N_23484);
or U23780 (N_23780,N_23531,N_23527);
xnor U23781 (N_23781,N_23519,N_23512);
and U23782 (N_23782,N_23575,N_23582);
xor U23783 (N_23783,N_23570,N_23585);
and U23784 (N_23784,N_23503,N_23432);
nand U23785 (N_23785,N_23485,N_23513);
and U23786 (N_23786,N_23536,N_23500);
and U23787 (N_23787,N_23465,N_23572);
nand U23788 (N_23788,N_23592,N_23495);
nand U23789 (N_23789,N_23460,N_23573);
and U23790 (N_23790,N_23548,N_23488);
xor U23791 (N_23791,N_23509,N_23456);
and U23792 (N_23792,N_23553,N_23422);
nand U23793 (N_23793,N_23479,N_23488);
nand U23794 (N_23794,N_23401,N_23465);
xor U23795 (N_23795,N_23528,N_23445);
nor U23796 (N_23796,N_23468,N_23581);
and U23797 (N_23797,N_23527,N_23569);
nand U23798 (N_23798,N_23542,N_23509);
xor U23799 (N_23799,N_23509,N_23469);
and U23800 (N_23800,N_23754,N_23643);
and U23801 (N_23801,N_23794,N_23652);
xor U23802 (N_23802,N_23742,N_23757);
nor U23803 (N_23803,N_23731,N_23610);
xor U23804 (N_23804,N_23620,N_23684);
or U23805 (N_23805,N_23647,N_23673);
xnor U23806 (N_23806,N_23786,N_23772);
nand U23807 (N_23807,N_23792,N_23783);
nor U23808 (N_23808,N_23696,N_23640);
or U23809 (N_23809,N_23709,N_23729);
nor U23810 (N_23810,N_23763,N_23796);
or U23811 (N_23811,N_23769,N_23632);
xor U23812 (N_23812,N_23725,N_23780);
nor U23813 (N_23813,N_23669,N_23750);
nand U23814 (N_23814,N_23623,N_23741);
nand U23815 (N_23815,N_23755,N_23630);
or U23816 (N_23816,N_23723,N_23740);
nor U23817 (N_23817,N_23636,N_23724);
and U23818 (N_23818,N_23722,N_23629);
nand U23819 (N_23819,N_23795,N_23749);
nor U23820 (N_23820,N_23788,N_23716);
or U23821 (N_23821,N_23677,N_23666);
or U23822 (N_23822,N_23770,N_23736);
nand U23823 (N_23823,N_23768,N_23686);
xor U23824 (N_23824,N_23602,N_23762);
xor U23825 (N_23825,N_23656,N_23687);
nand U23826 (N_23826,N_23775,N_23680);
xor U23827 (N_23827,N_23655,N_23789);
nor U23828 (N_23828,N_23700,N_23668);
nor U23829 (N_23829,N_23618,N_23658);
or U23830 (N_23830,N_23714,N_23732);
xnor U23831 (N_23831,N_23627,N_23675);
nor U23832 (N_23832,N_23773,N_23653);
xor U23833 (N_23833,N_23657,N_23699);
nor U23834 (N_23834,N_23682,N_23661);
nor U23835 (N_23835,N_23642,N_23735);
nor U23836 (N_23836,N_23771,N_23764);
or U23837 (N_23837,N_23608,N_23745);
nand U23838 (N_23838,N_23639,N_23782);
and U23839 (N_23839,N_23613,N_23621);
or U23840 (N_23840,N_23738,N_23708);
or U23841 (N_23841,N_23612,N_23759);
or U23842 (N_23842,N_23634,N_23622);
and U23843 (N_23843,N_23798,N_23758);
or U23844 (N_23844,N_23690,N_23785);
nor U23845 (N_23845,N_23633,N_23707);
nand U23846 (N_23846,N_23730,N_23679);
nand U23847 (N_23847,N_23734,N_23779);
xor U23848 (N_23848,N_23781,N_23646);
nand U23849 (N_23849,N_23746,N_23648);
and U23850 (N_23850,N_23774,N_23748);
nor U23851 (N_23851,N_23767,N_23713);
or U23852 (N_23852,N_23739,N_23604);
and U23853 (N_23853,N_23761,N_23665);
xnor U23854 (N_23854,N_23606,N_23737);
or U23855 (N_23855,N_23706,N_23701);
or U23856 (N_23856,N_23719,N_23600);
nand U23857 (N_23857,N_23691,N_23611);
and U23858 (N_23858,N_23791,N_23681);
nor U23859 (N_23859,N_23790,N_23705);
or U23860 (N_23860,N_23635,N_23683);
nor U23861 (N_23861,N_23688,N_23672);
xnor U23862 (N_23862,N_23717,N_23747);
nand U23863 (N_23863,N_23674,N_23631);
or U23864 (N_23864,N_23625,N_23751);
and U23865 (N_23865,N_23628,N_23793);
and U23866 (N_23866,N_23603,N_23784);
nand U23867 (N_23867,N_23711,N_23702);
nor U23868 (N_23868,N_23718,N_23712);
or U23869 (N_23869,N_23644,N_23693);
and U23870 (N_23870,N_23609,N_23671);
or U23871 (N_23871,N_23695,N_23601);
or U23872 (N_23872,N_23703,N_23689);
or U23873 (N_23873,N_23698,N_23694);
nor U23874 (N_23874,N_23663,N_23624);
nor U23875 (N_23875,N_23720,N_23733);
nand U23876 (N_23876,N_23799,N_23776);
and U23877 (N_23877,N_23797,N_23710);
or U23878 (N_23878,N_23721,N_23787);
nor U23879 (N_23879,N_23726,N_23766);
nor U23880 (N_23880,N_23777,N_23619);
or U23881 (N_23881,N_23616,N_23667);
xnor U23882 (N_23882,N_23650,N_23715);
or U23883 (N_23883,N_23637,N_23753);
or U23884 (N_23884,N_23638,N_23697);
nor U23885 (N_23885,N_23645,N_23617);
nor U23886 (N_23886,N_23752,N_23649);
nor U23887 (N_23887,N_23670,N_23660);
xnor U23888 (N_23888,N_23676,N_23778);
or U23889 (N_23889,N_23614,N_23605);
nor U23890 (N_23890,N_23607,N_23692);
or U23891 (N_23891,N_23744,N_23765);
xor U23892 (N_23892,N_23651,N_23727);
xnor U23893 (N_23893,N_23664,N_23615);
and U23894 (N_23894,N_23685,N_23654);
xor U23895 (N_23895,N_23662,N_23728);
xnor U23896 (N_23896,N_23641,N_23743);
nor U23897 (N_23897,N_23760,N_23756);
nand U23898 (N_23898,N_23678,N_23659);
xor U23899 (N_23899,N_23626,N_23704);
nor U23900 (N_23900,N_23793,N_23797);
xor U23901 (N_23901,N_23665,N_23750);
xnor U23902 (N_23902,N_23753,N_23634);
or U23903 (N_23903,N_23780,N_23723);
nor U23904 (N_23904,N_23631,N_23602);
and U23905 (N_23905,N_23724,N_23682);
or U23906 (N_23906,N_23783,N_23679);
nor U23907 (N_23907,N_23700,N_23774);
xnor U23908 (N_23908,N_23673,N_23757);
nand U23909 (N_23909,N_23747,N_23715);
and U23910 (N_23910,N_23700,N_23712);
or U23911 (N_23911,N_23673,N_23725);
nand U23912 (N_23912,N_23732,N_23768);
nand U23913 (N_23913,N_23693,N_23700);
or U23914 (N_23914,N_23655,N_23703);
xnor U23915 (N_23915,N_23605,N_23788);
or U23916 (N_23916,N_23695,N_23732);
and U23917 (N_23917,N_23674,N_23607);
nand U23918 (N_23918,N_23676,N_23652);
and U23919 (N_23919,N_23744,N_23754);
and U23920 (N_23920,N_23635,N_23688);
nor U23921 (N_23921,N_23730,N_23631);
nor U23922 (N_23922,N_23620,N_23707);
xnor U23923 (N_23923,N_23619,N_23667);
xnor U23924 (N_23924,N_23616,N_23759);
or U23925 (N_23925,N_23778,N_23600);
nand U23926 (N_23926,N_23785,N_23695);
or U23927 (N_23927,N_23700,N_23764);
xnor U23928 (N_23928,N_23682,N_23659);
or U23929 (N_23929,N_23613,N_23757);
and U23930 (N_23930,N_23787,N_23770);
nand U23931 (N_23931,N_23760,N_23770);
and U23932 (N_23932,N_23750,N_23736);
nor U23933 (N_23933,N_23631,N_23624);
xnor U23934 (N_23934,N_23783,N_23602);
nor U23935 (N_23935,N_23770,N_23716);
nand U23936 (N_23936,N_23795,N_23766);
nor U23937 (N_23937,N_23702,N_23766);
xor U23938 (N_23938,N_23776,N_23623);
xor U23939 (N_23939,N_23743,N_23631);
or U23940 (N_23940,N_23764,N_23719);
and U23941 (N_23941,N_23773,N_23761);
xnor U23942 (N_23942,N_23626,N_23625);
nand U23943 (N_23943,N_23799,N_23641);
xor U23944 (N_23944,N_23606,N_23700);
or U23945 (N_23945,N_23666,N_23768);
or U23946 (N_23946,N_23747,N_23780);
xnor U23947 (N_23947,N_23799,N_23708);
and U23948 (N_23948,N_23655,N_23716);
nand U23949 (N_23949,N_23720,N_23644);
xor U23950 (N_23950,N_23654,N_23719);
xnor U23951 (N_23951,N_23676,N_23628);
and U23952 (N_23952,N_23647,N_23610);
or U23953 (N_23953,N_23751,N_23724);
nor U23954 (N_23954,N_23788,N_23707);
xnor U23955 (N_23955,N_23614,N_23779);
xor U23956 (N_23956,N_23693,N_23711);
or U23957 (N_23957,N_23683,N_23653);
nand U23958 (N_23958,N_23701,N_23627);
nand U23959 (N_23959,N_23643,N_23714);
and U23960 (N_23960,N_23796,N_23637);
or U23961 (N_23961,N_23608,N_23776);
xor U23962 (N_23962,N_23743,N_23639);
nand U23963 (N_23963,N_23762,N_23685);
xnor U23964 (N_23964,N_23727,N_23721);
and U23965 (N_23965,N_23708,N_23727);
or U23966 (N_23966,N_23767,N_23630);
nor U23967 (N_23967,N_23787,N_23649);
nand U23968 (N_23968,N_23692,N_23788);
nor U23969 (N_23969,N_23650,N_23757);
or U23970 (N_23970,N_23694,N_23642);
or U23971 (N_23971,N_23703,N_23734);
nand U23972 (N_23972,N_23711,N_23729);
or U23973 (N_23973,N_23653,N_23784);
or U23974 (N_23974,N_23602,N_23600);
nor U23975 (N_23975,N_23661,N_23771);
or U23976 (N_23976,N_23617,N_23634);
nor U23977 (N_23977,N_23600,N_23648);
nor U23978 (N_23978,N_23784,N_23651);
nor U23979 (N_23979,N_23726,N_23757);
nor U23980 (N_23980,N_23668,N_23681);
and U23981 (N_23981,N_23703,N_23791);
xor U23982 (N_23982,N_23760,N_23769);
xor U23983 (N_23983,N_23776,N_23751);
or U23984 (N_23984,N_23640,N_23600);
xor U23985 (N_23985,N_23684,N_23638);
nor U23986 (N_23986,N_23721,N_23742);
nor U23987 (N_23987,N_23603,N_23765);
xnor U23988 (N_23988,N_23636,N_23628);
nor U23989 (N_23989,N_23778,N_23650);
and U23990 (N_23990,N_23617,N_23616);
and U23991 (N_23991,N_23604,N_23745);
nand U23992 (N_23992,N_23790,N_23718);
xor U23993 (N_23993,N_23764,N_23773);
or U23994 (N_23994,N_23706,N_23675);
nor U23995 (N_23995,N_23703,N_23726);
xnor U23996 (N_23996,N_23694,N_23782);
nand U23997 (N_23997,N_23683,N_23799);
or U23998 (N_23998,N_23702,N_23683);
and U23999 (N_23999,N_23610,N_23766);
xor U24000 (N_24000,N_23994,N_23975);
or U24001 (N_24001,N_23886,N_23964);
xor U24002 (N_24002,N_23885,N_23913);
or U24003 (N_24003,N_23951,N_23847);
xnor U24004 (N_24004,N_23832,N_23883);
and U24005 (N_24005,N_23826,N_23821);
nor U24006 (N_24006,N_23871,N_23808);
xor U24007 (N_24007,N_23889,N_23955);
and U24008 (N_24008,N_23957,N_23914);
and U24009 (N_24009,N_23859,N_23857);
nor U24010 (N_24010,N_23806,N_23822);
or U24011 (N_24011,N_23846,N_23867);
nor U24012 (N_24012,N_23915,N_23910);
nor U24013 (N_24013,N_23851,N_23980);
or U24014 (N_24014,N_23863,N_23887);
nand U24015 (N_24015,N_23873,N_23929);
nor U24016 (N_24016,N_23986,N_23827);
nand U24017 (N_24017,N_23944,N_23996);
nand U24018 (N_24018,N_23948,N_23833);
nand U24019 (N_24019,N_23958,N_23971);
nand U24020 (N_24020,N_23981,N_23850);
nor U24021 (N_24021,N_23876,N_23999);
nand U24022 (N_24022,N_23942,N_23818);
nor U24023 (N_24023,N_23959,N_23928);
or U24024 (N_24024,N_23860,N_23949);
nor U24025 (N_24025,N_23858,N_23987);
and U24026 (N_24026,N_23834,N_23902);
nand U24027 (N_24027,N_23916,N_23815);
nand U24028 (N_24028,N_23945,N_23920);
or U24029 (N_24029,N_23952,N_23874);
or U24030 (N_24030,N_23954,N_23977);
and U24031 (N_24031,N_23911,N_23922);
and U24032 (N_24032,N_23923,N_23984);
nand U24033 (N_24033,N_23894,N_23807);
nand U24034 (N_24034,N_23809,N_23877);
and U24035 (N_24035,N_23884,N_23879);
and U24036 (N_24036,N_23817,N_23899);
xnor U24037 (N_24037,N_23854,N_23966);
xor U24038 (N_24038,N_23992,N_23925);
nand U24039 (N_24039,N_23901,N_23927);
nor U24040 (N_24040,N_23830,N_23845);
xnor U24041 (N_24041,N_23825,N_23972);
and U24042 (N_24042,N_23880,N_23852);
or U24043 (N_24043,N_23924,N_23893);
xor U24044 (N_24044,N_23993,N_23820);
xnor U24045 (N_24045,N_23848,N_23814);
nand U24046 (N_24046,N_23947,N_23970);
or U24047 (N_24047,N_23819,N_23983);
nor U24048 (N_24048,N_23908,N_23842);
or U24049 (N_24049,N_23982,N_23960);
and U24050 (N_24050,N_23804,N_23962);
and U24051 (N_24051,N_23800,N_23843);
nand U24052 (N_24052,N_23973,N_23805);
nand U24053 (N_24053,N_23813,N_23936);
xor U24054 (N_24054,N_23823,N_23904);
nand U24055 (N_24055,N_23943,N_23935);
nand U24056 (N_24056,N_23941,N_23865);
or U24057 (N_24057,N_23836,N_23837);
nor U24058 (N_24058,N_23892,N_23868);
and U24059 (N_24059,N_23918,N_23991);
nor U24060 (N_24060,N_23898,N_23824);
and U24061 (N_24061,N_23912,N_23988);
xnor U24062 (N_24062,N_23838,N_23866);
nor U24063 (N_24063,N_23919,N_23930);
or U24064 (N_24064,N_23897,N_23881);
or U24065 (N_24065,N_23890,N_23934);
or U24066 (N_24066,N_23976,N_23939);
or U24067 (N_24067,N_23840,N_23844);
xnor U24068 (N_24068,N_23965,N_23940);
xor U24069 (N_24069,N_23906,N_23849);
and U24070 (N_24070,N_23974,N_23907);
xnor U24071 (N_24071,N_23864,N_23926);
nand U24072 (N_24072,N_23896,N_23950);
nor U24073 (N_24073,N_23839,N_23933);
and U24074 (N_24074,N_23855,N_23946);
or U24075 (N_24075,N_23875,N_23998);
or U24076 (N_24076,N_23961,N_23921);
nand U24077 (N_24077,N_23888,N_23990);
and U24078 (N_24078,N_23937,N_23811);
or U24079 (N_24079,N_23872,N_23891);
or U24080 (N_24080,N_23978,N_23900);
xor U24081 (N_24081,N_23979,N_23969);
xnor U24082 (N_24082,N_23870,N_23810);
nor U24083 (N_24083,N_23835,N_23882);
nand U24084 (N_24084,N_23841,N_23997);
nor U24085 (N_24085,N_23968,N_23869);
xnor U24086 (N_24086,N_23828,N_23985);
or U24087 (N_24087,N_23801,N_23903);
nor U24088 (N_24088,N_23816,N_23963);
nand U24089 (N_24089,N_23917,N_23931);
xnor U24090 (N_24090,N_23938,N_23862);
nand U24091 (N_24091,N_23812,N_23803);
xor U24092 (N_24092,N_23932,N_23953);
nor U24093 (N_24093,N_23829,N_23989);
or U24094 (N_24094,N_23856,N_23909);
nand U24095 (N_24095,N_23878,N_23995);
and U24096 (N_24096,N_23905,N_23831);
nand U24097 (N_24097,N_23895,N_23956);
xor U24098 (N_24098,N_23802,N_23861);
nor U24099 (N_24099,N_23967,N_23853);
xor U24100 (N_24100,N_23836,N_23988);
and U24101 (N_24101,N_23885,N_23844);
and U24102 (N_24102,N_23925,N_23995);
xor U24103 (N_24103,N_23873,N_23937);
nand U24104 (N_24104,N_23905,N_23807);
and U24105 (N_24105,N_23850,N_23959);
nand U24106 (N_24106,N_23818,N_23865);
nor U24107 (N_24107,N_23811,N_23943);
nand U24108 (N_24108,N_23850,N_23952);
xnor U24109 (N_24109,N_23933,N_23810);
nand U24110 (N_24110,N_23978,N_23880);
and U24111 (N_24111,N_23941,N_23929);
or U24112 (N_24112,N_23838,N_23924);
nand U24113 (N_24113,N_23956,N_23884);
or U24114 (N_24114,N_23838,N_23967);
nor U24115 (N_24115,N_23821,N_23958);
nand U24116 (N_24116,N_23856,N_23972);
xor U24117 (N_24117,N_23925,N_23834);
nand U24118 (N_24118,N_23998,N_23954);
nand U24119 (N_24119,N_23815,N_23873);
nand U24120 (N_24120,N_23914,N_23894);
or U24121 (N_24121,N_23975,N_23849);
xor U24122 (N_24122,N_23912,N_23880);
xnor U24123 (N_24123,N_23999,N_23936);
nand U24124 (N_24124,N_23992,N_23988);
and U24125 (N_24125,N_23962,N_23966);
xnor U24126 (N_24126,N_23890,N_23867);
and U24127 (N_24127,N_23964,N_23958);
nor U24128 (N_24128,N_23863,N_23819);
xor U24129 (N_24129,N_23995,N_23869);
nand U24130 (N_24130,N_23927,N_23851);
xnor U24131 (N_24131,N_23957,N_23918);
or U24132 (N_24132,N_23915,N_23971);
xnor U24133 (N_24133,N_23857,N_23936);
and U24134 (N_24134,N_23861,N_23879);
nand U24135 (N_24135,N_23994,N_23848);
nor U24136 (N_24136,N_23936,N_23809);
or U24137 (N_24137,N_23806,N_23950);
xor U24138 (N_24138,N_23950,N_23979);
xnor U24139 (N_24139,N_23903,N_23901);
or U24140 (N_24140,N_23837,N_23932);
and U24141 (N_24141,N_23800,N_23922);
nor U24142 (N_24142,N_23972,N_23845);
xor U24143 (N_24143,N_23870,N_23969);
xor U24144 (N_24144,N_23858,N_23830);
and U24145 (N_24145,N_23953,N_23918);
nand U24146 (N_24146,N_23949,N_23973);
or U24147 (N_24147,N_23966,N_23880);
nand U24148 (N_24148,N_23902,N_23928);
nand U24149 (N_24149,N_23841,N_23975);
nor U24150 (N_24150,N_23996,N_23884);
or U24151 (N_24151,N_23813,N_23857);
and U24152 (N_24152,N_23948,N_23972);
or U24153 (N_24153,N_23974,N_23983);
nand U24154 (N_24154,N_23893,N_23821);
nor U24155 (N_24155,N_23867,N_23833);
nor U24156 (N_24156,N_23868,N_23862);
or U24157 (N_24157,N_23994,N_23984);
nor U24158 (N_24158,N_23881,N_23886);
and U24159 (N_24159,N_23981,N_23973);
nand U24160 (N_24160,N_23907,N_23833);
or U24161 (N_24161,N_23936,N_23804);
nor U24162 (N_24162,N_23963,N_23811);
nand U24163 (N_24163,N_23842,N_23968);
xor U24164 (N_24164,N_23946,N_23822);
and U24165 (N_24165,N_23886,N_23972);
and U24166 (N_24166,N_23887,N_23856);
or U24167 (N_24167,N_23854,N_23801);
xnor U24168 (N_24168,N_23985,N_23952);
xnor U24169 (N_24169,N_23908,N_23960);
or U24170 (N_24170,N_23859,N_23880);
xnor U24171 (N_24171,N_23867,N_23983);
and U24172 (N_24172,N_23861,N_23901);
xor U24173 (N_24173,N_23978,N_23893);
and U24174 (N_24174,N_23856,N_23827);
or U24175 (N_24175,N_23973,N_23829);
nand U24176 (N_24176,N_23891,N_23853);
nor U24177 (N_24177,N_23916,N_23913);
xor U24178 (N_24178,N_23928,N_23924);
nor U24179 (N_24179,N_23869,N_23963);
xor U24180 (N_24180,N_23870,N_23800);
xor U24181 (N_24181,N_23801,N_23849);
nand U24182 (N_24182,N_23882,N_23804);
and U24183 (N_24183,N_23999,N_23932);
nand U24184 (N_24184,N_23867,N_23851);
and U24185 (N_24185,N_23920,N_23914);
and U24186 (N_24186,N_23904,N_23801);
nand U24187 (N_24187,N_23911,N_23853);
nand U24188 (N_24188,N_23803,N_23958);
and U24189 (N_24189,N_23840,N_23946);
and U24190 (N_24190,N_23940,N_23882);
nor U24191 (N_24191,N_23873,N_23865);
or U24192 (N_24192,N_23872,N_23802);
nor U24193 (N_24193,N_23938,N_23873);
or U24194 (N_24194,N_23807,N_23946);
xor U24195 (N_24195,N_23819,N_23935);
or U24196 (N_24196,N_23965,N_23993);
or U24197 (N_24197,N_23966,N_23861);
or U24198 (N_24198,N_23983,N_23936);
and U24199 (N_24199,N_23890,N_23971);
and U24200 (N_24200,N_24000,N_24001);
and U24201 (N_24201,N_24187,N_24049);
and U24202 (N_24202,N_24183,N_24038);
nor U24203 (N_24203,N_24150,N_24155);
xor U24204 (N_24204,N_24030,N_24120);
and U24205 (N_24205,N_24088,N_24101);
nand U24206 (N_24206,N_24115,N_24152);
nor U24207 (N_24207,N_24159,N_24141);
xnor U24208 (N_24208,N_24077,N_24035);
nand U24209 (N_24209,N_24067,N_24042);
nand U24210 (N_24210,N_24184,N_24040);
nor U24211 (N_24211,N_24006,N_24161);
xor U24212 (N_24212,N_24068,N_24020);
nand U24213 (N_24213,N_24127,N_24121);
or U24214 (N_24214,N_24104,N_24111);
nor U24215 (N_24215,N_24142,N_24017);
and U24216 (N_24216,N_24128,N_24019);
or U24217 (N_24217,N_24091,N_24158);
nand U24218 (N_24218,N_24056,N_24167);
nor U24219 (N_24219,N_24138,N_24021);
and U24220 (N_24220,N_24177,N_24026);
or U24221 (N_24221,N_24059,N_24083);
nand U24222 (N_24222,N_24163,N_24132);
or U24223 (N_24223,N_24195,N_24018);
xor U24224 (N_24224,N_24078,N_24043);
and U24225 (N_24225,N_24118,N_24129);
nand U24226 (N_24226,N_24060,N_24097);
and U24227 (N_24227,N_24027,N_24005);
and U24228 (N_24228,N_24080,N_24105);
and U24229 (N_24229,N_24063,N_24029);
and U24230 (N_24230,N_24176,N_24034);
xor U24231 (N_24231,N_24076,N_24135);
nor U24232 (N_24232,N_24193,N_24164);
nor U24233 (N_24233,N_24066,N_24082);
or U24234 (N_24234,N_24065,N_24062);
and U24235 (N_24235,N_24174,N_24106);
or U24236 (N_24236,N_24151,N_24079);
nand U24237 (N_24237,N_24188,N_24178);
or U24238 (N_24238,N_24072,N_24089);
nand U24239 (N_24239,N_24037,N_24197);
nor U24240 (N_24240,N_24124,N_24047);
xor U24241 (N_24241,N_24084,N_24094);
and U24242 (N_24242,N_24139,N_24169);
and U24243 (N_24243,N_24173,N_24032);
or U24244 (N_24244,N_24050,N_24051);
xor U24245 (N_24245,N_24190,N_24117);
or U24246 (N_24246,N_24095,N_24045);
nand U24247 (N_24247,N_24055,N_24194);
and U24248 (N_24248,N_24179,N_24033);
and U24249 (N_24249,N_24153,N_24057);
nor U24250 (N_24250,N_24170,N_24146);
nor U24251 (N_24251,N_24149,N_24140);
and U24252 (N_24252,N_24098,N_24073);
nor U24253 (N_24253,N_24100,N_24025);
nor U24254 (N_24254,N_24058,N_24191);
nor U24255 (N_24255,N_24166,N_24192);
or U24256 (N_24256,N_24168,N_24015);
nand U24257 (N_24257,N_24085,N_24012);
xor U24258 (N_24258,N_24157,N_24075);
nand U24259 (N_24259,N_24145,N_24144);
nand U24260 (N_24260,N_24143,N_24010);
or U24261 (N_24261,N_24108,N_24125);
and U24262 (N_24262,N_24130,N_24172);
xor U24263 (N_24263,N_24064,N_24007);
nand U24264 (N_24264,N_24002,N_24013);
and U24265 (N_24265,N_24044,N_24087);
nor U24266 (N_24266,N_24031,N_24014);
and U24267 (N_24267,N_24069,N_24081);
nand U24268 (N_24268,N_24009,N_24103);
or U24269 (N_24269,N_24023,N_24024);
nor U24270 (N_24270,N_24061,N_24148);
nand U24271 (N_24271,N_24028,N_24004);
and U24272 (N_24272,N_24053,N_24054);
or U24273 (N_24273,N_24114,N_24131);
xor U24274 (N_24274,N_24171,N_24136);
and U24275 (N_24275,N_24126,N_24162);
or U24276 (N_24276,N_24165,N_24048);
nor U24277 (N_24277,N_24186,N_24107);
nand U24278 (N_24278,N_24198,N_24016);
nand U24279 (N_24279,N_24011,N_24112);
and U24280 (N_24280,N_24113,N_24160);
nand U24281 (N_24281,N_24154,N_24133);
xnor U24282 (N_24282,N_24102,N_24074);
and U24283 (N_24283,N_24046,N_24199);
xnor U24284 (N_24284,N_24137,N_24134);
xnor U24285 (N_24285,N_24092,N_24109);
and U24286 (N_24286,N_24093,N_24189);
xnor U24287 (N_24287,N_24039,N_24156);
xor U24288 (N_24288,N_24182,N_24022);
or U24289 (N_24289,N_24096,N_24071);
nor U24290 (N_24290,N_24181,N_24086);
and U24291 (N_24291,N_24122,N_24196);
or U24292 (N_24292,N_24041,N_24036);
nand U24293 (N_24293,N_24175,N_24090);
nor U24294 (N_24294,N_24119,N_24052);
nor U24295 (N_24295,N_24070,N_24123);
or U24296 (N_24296,N_24110,N_24180);
nor U24297 (N_24297,N_24147,N_24099);
nor U24298 (N_24298,N_24003,N_24185);
or U24299 (N_24299,N_24008,N_24116);
or U24300 (N_24300,N_24195,N_24094);
and U24301 (N_24301,N_24149,N_24150);
nand U24302 (N_24302,N_24086,N_24196);
and U24303 (N_24303,N_24102,N_24070);
nand U24304 (N_24304,N_24007,N_24143);
or U24305 (N_24305,N_24070,N_24118);
nand U24306 (N_24306,N_24015,N_24113);
or U24307 (N_24307,N_24135,N_24138);
or U24308 (N_24308,N_24046,N_24160);
or U24309 (N_24309,N_24059,N_24116);
nand U24310 (N_24310,N_24072,N_24178);
and U24311 (N_24311,N_24023,N_24099);
xor U24312 (N_24312,N_24046,N_24159);
or U24313 (N_24313,N_24050,N_24100);
xnor U24314 (N_24314,N_24175,N_24073);
and U24315 (N_24315,N_24092,N_24147);
xor U24316 (N_24316,N_24172,N_24095);
nand U24317 (N_24317,N_24028,N_24042);
xor U24318 (N_24318,N_24194,N_24006);
and U24319 (N_24319,N_24186,N_24039);
nor U24320 (N_24320,N_24108,N_24134);
nor U24321 (N_24321,N_24016,N_24155);
nand U24322 (N_24322,N_24131,N_24025);
and U24323 (N_24323,N_24154,N_24045);
and U24324 (N_24324,N_24170,N_24130);
nor U24325 (N_24325,N_24167,N_24091);
nand U24326 (N_24326,N_24198,N_24007);
and U24327 (N_24327,N_24056,N_24067);
nor U24328 (N_24328,N_24134,N_24136);
and U24329 (N_24329,N_24037,N_24193);
nand U24330 (N_24330,N_24137,N_24061);
xor U24331 (N_24331,N_24144,N_24114);
or U24332 (N_24332,N_24172,N_24044);
nand U24333 (N_24333,N_24131,N_24198);
xnor U24334 (N_24334,N_24093,N_24019);
and U24335 (N_24335,N_24178,N_24057);
or U24336 (N_24336,N_24154,N_24135);
nand U24337 (N_24337,N_24194,N_24035);
or U24338 (N_24338,N_24100,N_24067);
xnor U24339 (N_24339,N_24197,N_24187);
or U24340 (N_24340,N_24041,N_24004);
nand U24341 (N_24341,N_24072,N_24085);
nor U24342 (N_24342,N_24189,N_24054);
nor U24343 (N_24343,N_24172,N_24049);
nor U24344 (N_24344,N_24024,N_24022);
or U24345 (N_24345,N_24111,N_24154);
nor U24346 (N_24346,N_24147,N_24107);
or U24347 (N_24347,N_24183,N_24147);
nand U24348 (N_24348,N_24011,N_24017);
or U24349 (N_24349,N_24168,N_24040);
xnor U24350 (N_24350,N_24179,N_24163);
nor U24351 (N_24351,N_24087,N_24101);
nor U24352 (N_24352,N_24052,N_24066);
nor U24353 (N_24353,N_24017,N_24114);
and U24354 (N_24354,N_24162,N_24180);
and U24355 (N_24355,N_24008,N_24180);
and U24356 (N_24356,N_24176,N_24011);
and U24357 (N_24357,N_24137,N_24110);
xor U24358 (N_24358,N_24002,N_24139);
xnor U24359 (N_24359,N_24150,N_24091);
or U24360 (N_24360,N_24169,N_24019);
or U24361 (N_24361,N_24047,N_24115);
and U24362 (N_24362,N_24185,N_24170);
nand U24363 (N_24363,N_24116,N_24087);
and U24364 (N_24364,N_24084,N_24018);
nand U24365 (N_24365,N_24001,N_24126);
nor U24366 (N_24366,N_24104,N_24139);
nor U24367 (N_24367,N_24168,N_24161);
xnor U24368 (N_24368,N_24138,N_24080);
nor U24369 (N_24369,N_24184,N_24028);
and U24370 (N_24370,N_24191,N_24016);
or U24371 (N_24371,N_24089,N_24027);
and U24372 (N_24372,N_24199,N_24173);
or U24373 (N_24373,N_24134,N_24044);
xor U24374 (N_24374,N_24108,N_24095);
nand U24375 (N_24375,N_24123,N_24164);
and U24376 (N_24376,N_24193,N_24138);
and U24377 (N_24377,N_24001,N_24088);
or U24378 (N_24378,N_24134,N_24171);
nand U24379 (N_24379,N_24044,N_24051);
or U24380 (N_24380,N_24038,N_24186);
nor U24381 (N_24381,N_24184,N_24046);
xnor U24382 (N_24382,N_24190,N_24077);
xnor U24383 (N_24383,N_24112,N_24134);
xnor U24384 (N_24384,N_24102,N_24080);
or U24385 (N_24385,N_24138,N_24077);
nand U24386 (N_24386,N_24051,N_24083);
nor U24387 (N_24387,N_24129,N_24176);
or U24388 (N_24388,N_24157,N_24095);
xnor U24389 (N_24389,N_24026,N_24144);
nor U24390 (N_24390,N_24022,N_24045);
nand U24391 (N_24391,N_24192,N_24085);
xnor U24392 (N_24392,N_24080,N_24050);
nor U24393 (N_24393,N_24192,N_24064);
xor U24394 (N_24394,N_24190,N_24071);
and U24395 (N_24395,N_24093,N_24156);
nor U24396 (N_24396,N_24194,N_24140);
nor U24397 (N_24397,N_24092,N_24167);
xnor U24398 (N_24398,N_24198,N_24184);
and U24399 (N_24399,N_24039,N_24185);
and U24400 (N_24400,N_24230,N_24269);
or U24401 (N_24401,N_24370,N_24308);
or U24402 (N_24402,N_24241,N_24254);
xnor U24403 (N_24403,N_24250,N_24376);
or U24404 (N_24404,N_24246,N_24336);
xor U24405 (N_24405,N_24267,N_24390);
or U24406 (N_24406,N_24268,N_24247);
nor U24407 (N_24407,N_24294,N_24212);
or U24408 (N_24408,N_24311,N_24373);
or U24409 (N_24409,N_24392,N_24226);
or U24410 (N_24410,N_24397,N_24209);
nor U24411 (N_24411,N_24204,N_24284);
or U24412 (N_24412,N_24243,N_24380);
xnor U24413 (N_24413,N_24291,N_24389);
xnor U24414 (N_24414,N_24281,N_24235);
and U24415 (N_24415,N_24203,N_24326);
nand U24416 (N_24416,N_24325,N_24200);
xnor U24417 (N_24417,N_24365,N_24224);
nor U24418 (N_24418,N_24378,N_24248);
nand U24419 (N_24419,N_24323,N_24237);
nand U24420 (N_24420,N_24320,N_24331);
nor U24421 (N_24421,N_24322,N_24318);
and U24422 (N_24422,N_24295,N_24290);
nor U24423 (N_24423,N_24345,N_24324);
or U24424 (N_24424,N_24210,N_24251);
xor U24425 (N_24425,N_24381,N_24218);
nor U24426 (N_24426,N_24232,N_24328);
xnor U24427 (N_24427,N_24347,N_24252);
xnor U24428 (N_24428,N_24211,N_24277);
xor U24429 (N_24429,N_24225,N_24259);
or U24430 (N_24430,N_24352,N_24263);
nand U24431 (N_24431,N_24208,N_24223);
xnor U24432 (N_24432,N_24335,N_24272);
or U24433 (N_24433,N_24296,N_24333);
nand U24434 (N_24434,N_24394,N_24302);
or U24435 (N_24435,N_24228,N_24327);
or U24436 (N_24436,N_24292,N_24354);
and U24437 (N_24437,N_24353,N_24286);
and U24438 (N_24438,N_24278,N_24371);
or U24439 (N_24439,N_24242,N_24329);
and U24440 (N_24440,N_24227,N_24202);
and U24441 (N_24441,N_24280,N_24338);
xnor U24442 (N_24442,N_24275,N_24231);
xor U24443 (N_24443,N_24213,N_24360);
or U24444 (N_24444,N_24337,N_24299);
nor U24445 (N_24445,N_24289,N_24382);
or U24446 (N_24446,N_24215,N_24258);
nand U24447 (N_24447,N_24366,N_24355);
xnor U24448 (N_24448,N_24317,N_24361);
nor U24449 (N_24449,N_24349,N_24238);
nand U24450 (N_24450,N_24314,N_24239);
and U24451 (N_24451,N_24298,N_24266);
or U24452 (N_24452,N_24310,N_24393);
or U24453 (N_24453,N_24368,N_24386);
nand U24454 (N_24454,N_24214,N_24396);
nor U24455 (N_24455,N_24244,N_24222);
and U24456 (N_24456,N_24287,N_24303);
nand U24457 (N_24457,N_24274,N_24260);
nor U24458 (N_24458,N_24398,N_24346);
and U24459 (N_24459,N_24315,N_24369);
nor U24460 (N_24460,N_24341,N_24205);
or U24461 (N_24461,N_24344,N_24206);
nand U24462 (N_24462,N_24240,N_24234);
or U24463 (N_24463,N_24316,N_24332);
and U24464 (N_24464,N_24255,N_24334);
and U24465 (N_24465,N_24375,N_24304);
xnor U24466 (N_24466,N_24297,N_24245);
xnor U24467 (N_24467,N_24357,N_24319);
and U24468 (N_24468,N_24293,N_24216);
nor U24469 (N_24469,N_24342,N_24363);
or U24470 (N_24470,N_24273,N_24356);
or U24471 (N_24471,N_24236,N_24201);
nor U24472 (N_24472,N_24276,N_24359);
xnor U24473 (N_24473,N_24364,N_24383);
xnor U24474 (N_24474,N_24388,N_24282);
nand U24475 (N_24475,N_24307,N_24279);
nand U24476 (N_24476,N_24305,N_24262);
nand U24477 (N_24477,N_24256,N_24257);
nand U24478 (N_24478,N_24372,N_24265);
xnor U24479 (N_24479,N_24362,N_24217);
xor U24480 (N_24480,N_24312,N_24229);
nand U24481 (N_24481,N_24321,N_24221);
and U24482 (N_24482,N_24313,N_24233);
or U24483 (N_24483,N_24348,N_24300);
nor U24484 (N_24484,N_24343,N_24220);
nor U24485 (N_24485,N_24330,N_24391);
or U24486 (N_24486,N_24285,N_24358);
and U24487 (N_24487,N_24350,N_24377);
or U24488 (N_24488,N_24270,N_24301);
xnor U24489 (N_24489,N_24249,N_24264);
nand U24490 (N_24490,N_24399,N_24207);
nand U24491 (N_24491,N_24309,N_24261);
or U24492 (N_24492,N_24283,N_24374);
and U24493 (N_24493,N_24339,N_24340);
nand U24494 (N_24494,N_24271,N_24387);
and U24495 (N_24495,N_24288,N_24351);
xor U24496 (N_24496,N_24384,N_24379);
and U24497 (N_24497,N_24219,N_24306);
nand U24498 (N_24498,N_24253,N_24385);
or U24499 (N_24499,N_24395,N_24367);
or U24500 (N_24500,N_24265,N_24387);
and U24501 (N_24501,N_24319,N_24348);
or U24502 (N_24502,N_24283,N_24356);
xor U24503 (N_24503,N_24316,N_24322);
nor U24504 (N_24504,N_24316,N_24259);
and U24505 (N_24505,N_24286,N_24395);
nor U24506 (N_24506,N_24251,N_24255);
or U24507 (N_24507,N_24250,N_24312);
nand U24508 (N_24508,N_24230,N_24224);
and U24509 (N_24509,N_24358,N_24298);
xor U24510 (N_24510,N_24228,N_24242);
and U24511 (N_24511,N_24311,N_24322);
or U24512 (N_24512,N_24213,N_24294);
nor U24513 (N_24513,N_24399,N_24317);
or U24514 (N_24514,N_24258,N_24313);
and U24515 (N_24515,N_24333,N_24359);
nor U24516 (N_24516,N_24229,N_24379);
or U24517 (N_24517,N_24294,N_24315);
xor U24518 (N_24518,N_24238,N_24243);
and U24519 (N_24519,N_24255,N_24266);
or U24520 (N_24520,N_24269,N_24285);
nor U24521 (N_24521,N_24399,N_24254);
nand U24522 (N_24522,N_24370,N_24226);
and U24523 (N_24523,N_24238,N_24220);
and U24524 (N_24524,N_24323,N_24361);
nor U24525 (N_24525,N_24331,N_24304);
nor U24526 (N_24526,N_24274,N_24256);
or U24527 (N_24527,N_24303,N_24257);
or U24528 (N_24528,N_24278,N_24208);
nor U24529 (N_24529,N_24304,N_24311);
nor U24530 (N_24530,N_24312,N_24350);
xor U24531 (N_24531,N_24325,N_24230);
nand U24532 (N_24532,N_24208,N_24366);
nor U24533 (N_24533,N_24261,N_24336);
nand U24534 (N_24534,N_24215,N_24228);
and U24535 (N_24535,N_24382,N_24261);
xor U24536 (N_24536,N_24346,N_24274);
and U24537 (N_24537,N_24261,N_24395);
xnor U24538 (N_24538,N_24255,N_24364);
nor U24539 (N_24539,N_24302,N_24219);
and U24540 (N_24540,N_24383,N_24313);
or U24541 (N_24541,N_24206,N_24387);
and U24542 (N_24542,N_24351,N_24236);
nor U24543 (N_24543,N_24283,N_24323);
and U24544 (N_24544,N_24350,N_24353);
nand U24545 (N_24545,N_24335,N_24284);
or U24546 (N_24546,N_24246,N_24347);
and U24547 (N_24547,N_24239,N_24244);
xor U24548 (N_24548,N_24363,N_24330);
and U24549 (N_24549,N_24313,N_24238);
xnor U24550 (N_24550,N_24239,N_24316);
nor U24551 (N_24551,N_24350,N_24218);
or U24552 (N_24552,N_24394,N_24214);
xnor U24553 (N_24553,N_24352,N_24227);
or U24554 (N_24554,N_24249,N_24385);
nor U24555 (N_24555,N_24231,N_24360);
or U24556 (N_24556,N_24292,N_24258);
xnor U24557 (N_24557,N_24382,N_24349);
nand U24558 (N_24558,N_24259,N_24200);
or U24559 (N_24559,N_24327,N_24379);
or U24560 (N_24560,N_24206,N_24325);
or U24561 (N_24561,N_24215,N_24280);
nand U24562 (N_24562,N_24203,N_24335);
nor U24563 (N_24563,N_24276,N_24398);
xnor U24564 (N_24564,N_24345,N_24318);
xor U24565 (N_24565,N_24340,N_24288);
xnor U24566 (N_24566,N_24385,N_24305);
and U24567 (N_24567,N_24273,N_24380);
xor U24568 (N_24568,N_24356,N_24339);
and U24569 (N_24569,N_24285,N_24267);
and U24570 (N_24570,N_24322,N_24299);
xor U24571 (N_24571,N_24350,N_24324);
nor U24572 (N_24572,N_24311,N_24244);
nand U24573 (N_24573,N_24376,N_24209);
and U24574 (N_24574,N_24313,N_24355);
nor U24575 (N_24575,N_24263,N_24311);
and U24576 (N_24576,N_24339,N_24325);
nand U24577 (N_24577,N_24392,N_24388);
nor U24578 (N_24578,N_24346,N_24324);
nand U24579 (N_24579,N_24277,N_24290);
nand U24580 (N_24580,N_24396,N_24358);
and U24581 (N_24581,N_24349,N_24376);
or U24582 (N_24582,N_24365,N_24295);
or U24583 (N_24583,N_24333,N_24236);
nand U24584 (N_24584,N_24308,N_24310);
or U24585 (N_24585,N_24399,N_24324);
nand U24586 (N_24586,N_24209,N_24234);
nor U24587 (N_24587,N_24281,N_24267);
and U24588 (N_24588,N_24338,N_24248);
xor U24589 (N_24589,N_24323,N_24330);
and U24590 (N_24590,N_24237,N_24393);
nand U24591 (N_24591,N_24227,N_24384);
and U24592 (N_24592,N_24274,N_24352);
and U24593 (N_24593,N_24329,N_24240);
nand U24594 (N_24594,N_24380,N_24302);
nand U24595 (N_24595,N_24291,N_24223);
or U24596 (N_24596,N_24398,N_24284);
xor U24597 (N_24597,N_24265,N_24204);
xnor U24598 (N_24598,N_24278,N_24234);
and U24599 (N_24599,N_24306,N_24250);
nand U24600 (N_24600,N_24598,N_24530);
nor U24601 (N_24601,N_24595,N_24447);
xor U24602 (N_24602,N_24582,N_24492);
nor U24603 (N_24603,N_24585,N_24494);
or U24604 (N_24604,N_24427,N_24451);
or U24605 (N_24605,N_24477,N_24469);
or U24606 (N_24606,N_24566,N_24403);
or U24607 (N_24607,N_24411,N_24545);
nand U24608 (N_24608,N_24572,N_24479);
and U24609 (N_24609,N_24517,N_24467);
nor U24610 (N_24610,N_24504,N_24577);
nor U24611 (N_24611,N_24509,N_24426);
or U24612 (N_24612,N_24575,N_24528);
or U24613 (N_24613,N_24570,N_24516);
or U24614 (N_24614,N_24558,N_24550);
nor U24615 (N_24615,N_24410,N_24519);
and U24616 (N_24616,N_24405,N_24588);
nand U24617 (N_24617,N_24512,N_24465);
and U24618 (N_24618,N_24419,N_24409);
nand U24619 (N_24619,N_24462,N_24526);
xor U24620 (N_24620,N_24597,N_24523);
nor U24621 (N_24621,N_24422,N_24483);
nand U24622 (N_24622,N_24443,N_24536);
nand U24623 (N_24623,N_24448,N_24548);
xor U24624 (N_24624,N_24498,N_24413);
or U24625 (N_24625,N_24440,N_24576);
or U24626 (N_24626,N_24564,N_24420);
or U24627 (N_24627,N_24490,N_24454);
or U24628 (N_24628,N_24476,N_24534);
nor U24629 (N_24629,N_24458,N_24499);
or U24630 (N_24630,N_24445,N_24583);
xnor U24631 (N_24631,N_24402,N_24481);
nor U24632 (N_24632,N_24525,N_24457);
and U24633 (N_24633,N_24537,N_24599);
and U24634 (N_24634,N_24408,N_24450);
xor U24635 (N_24635,N_24417,N_24511);
xnor U24636 (N_24636,N_24508,N_24474);
nor U24637 (N_24637,N_24593,N_24455);
and U24638 (N_24638,N_24518,N_24482);
and U24639 (N_24639,N_24510,N_24425);
nor U24640 (N_24640,N_24429,N_24424);
xnor U24641 (N_24641,N_24501,N_24590);
nor U24642 (N_24642,N_24549,N_24473);
nor U24643 (N_24643,N_24573,N_24546);
and U24644 (N_24644,N_24432,N_24435);
nand U24645 (N_24645,N_24488,N_24529);
nor U24646 (N_24646,N_24506,N_24507);
nor U24647 (N_24647,N_24486,N_24431);
and U24648 (N_24648,N_24553,N_24541);
nand U24649 (N_24649,N_24555,N_24456);
xnor U24650 (N_24650,N_24495,N_24485);
or U24651 (N_24651,N_24491,N_24502);
or U24652 (N_24652,N_24552,N_24452);
nor U24653 (N_24653,N_24542,N_24527);
xnor U24654 (N_24654,N_24478,N_24442);
or U24655 (N_24655,N_24571,N_24586);
nand U24656 (N_24656,N_24580,N_24468);
nand U24657 (N_24657,N_24415,N_24438);
or U24658 (N_24658,N_24406,N_24475);
or U24659 (N_24659,N_24554,N_24500);
nor U24660 (N_24660,N_24416,N_24444);
and U24661 (N_24661,N_24533,N_24493);
and U24662 (N_24662,N_24556,N_24592);
nand U24663 (N_24663,N_24532,N_24531);
nand U24664 (N_24664,N_24515,N_24460);
nand U24665 (N_24665,N_24470,N_24497);
or U24666 (N_24666,N_24407,N_24591);
nor U24667 (N_24667,N_24540,N_24514);
and U24668 (N_24668,N_24459,N_24480);
or U24669 (N_24669,N_24567,N_24579);
and U24670 (N_24670,N_24428,N_24484);
and U24671 (N_24671,N_24505,N_24543);
nand U24672 (N_24672,N_24563,N_24589);
xnor U24673 (N_24673,N_24596,N_24544);
nor U24674 (N_24674,N_24513,N_24559);
xnor U24675 (N_24675,N_24520,N_24565);
xor U24676 (N_24676,N_24496,N_24441);
and U24677 (N_24677,N_24437,N_24569);
or U24678 (N_24678,N_24521,N_24568);
nor U24679 (N_24679,N_24578,N_24461);
or U24680 (N_24680,N_24471,N_24472);
nand U24681 (N_24681,N_24439,N_24587);
xnor U24682 (N_24682,N_24414,N_24538);
or U24683 (N_24683,N_24434,N_24594);
xor U24684 (N_24684,N_24464,N_24449);
nor U24685 (N_24685,N_24418,N_24547);
and U24686 (N_24686,N_24584,N_24400);
or U24687 (N_24687,N_24401,N_24412);
or U24688 (N_24688,N_24433,N_24535);
nor U24689 (N_24689,N_24503,N_24487);
and U24690 (N_24690,N_24560,N_24524);
nand U24691 (N_24691,N_24561,N_24557);
or U24692 (N_24692,N_24489,N_24453);
nand U24693 (N_24693,N_24551,N_24430);
or U24694 (N_24694,N_24423,N_24404);
nor U24695 (N_24695,N_24574,N_24466);
xnor U24696 (N_24696,N_24522,N_24421);
xor U24697 (N_24697,N_24463,N_24436);
and U24698 (N_24698,N_24562,N_24446);
and U24699 (N_24699,N_24581,N_24539);
nor U24700 (N_24700,N_24575,N_24430);
or U24701 (N_24701,N_24510,N_24576);
or U24702 (N_24702,N_24522,N_24468);
nand U24703 (N_24703,N_24565,N_24504);
nor U24704 (N_24704,N_24472,N_24431);
and U24705 (N_24705,N_24528,N_24415);
nor U24706 (N_24706,N_24585,N_24480);
nor U24707 (N_24707,N_24460,N_24418);
or U24708 (N_24708,N_24575,N_24535);
nor U24709 (N_24709,N_24582,N_24479);
or U24710 (N_24710,N_24577,N_24519);
nor U24711 (N_24711,N_24456,N_24450);
and U24712 (N_24712,N_24570,N_24508);
or U24713 (N_24713,N_24594,N_24581);
xor U24714 (N_24714,N_24414,N_24588);
and U24715 (N_24715,N_24486,N_24598);
nor U24716 (N_24716,N_24450,N_24484);
and U24717 (N_24717,N_24544,N_24411);
nor U24718 (N_24718,N_24416,N_24516);
and U24719 (N_24719,N_24436,N_24563);
nand U24720 (N_24720,N_24584,N_24596);
nand U24721 (N_24721,N_24461,N_24411);
and U24722 (N_24722,N_24498,N_24514);
and U24723 (N_24723,N_24487,N_24481);
xor U24724 (N_24724,N_24584,N_24415);
xnor U24725 (N_24725,N_24537,N_24570);
and U24726 (N_24726,N_24501,N_24506);
or U24727 (N_24727,N_24415,N_24563);
xnor U24728 (N_24728,N_24571,N_24484);
nor U24729 (N_24729,N_24406,N_24535);
and U24730 (N_24730,N_24555,N_24546);
and U24731 (N_24731,N_24552,N_24586);
nor U24732 (N_24732,N_24481,N_24411);
xor U24733 (N_24733,N_24429,N_24525);
nor U24734 (N_24734,N_24421,N_24434);
xor U24735 (N_24735,N_24404,N_24514);
nor U24736 (N_24736,N_24579,N_24554);
or U24737 (N_24737,N_24482,N_24547);
nor U24738 (N_24738,N_24442,N_24592);
xnor U24739 (N_24739,N_24404,N_24463);
or U24740 (N_24740,N_24433,N_24452);
and U24741 (N_24741,N_24510,N_24408);
nor U24742 (N_24742,N_24449,N_24438);
or U24743 (N_24743,N_24520,N_24524);
and U24744 (N_24744,N_24534,N_24420);
or U24745 (N_24745,N_24411,N_24561);
or U24746 (N_24746,N_24496,N_24442);
and U24747 (N_24747,N_24451,N_24444);
nand U24748 (N_24748,N_24428,N_24509);
nor U24749 (N_24749,N_24578,N_24566);
nand U24750 (N_24750,N_24583,N_24437);
xnor U24751 (N_24751,N_24515,N_24560);
and U24752 (N_24752,N_24456,N_24510);
or U24753 (N_24753,N_24436,N_24542);
or U24754 (N_24754,N_24429,N_24558);
xor U24755 (N_24755,N_24551,N_24597);
nand U24756 (N_24756,N_24511,N_24520);
and U24757 (N_24757,N_24514,N_24467);
xnor U24758 (N_24758,N_24424,N_24582);
nor U24759 (N_24759,N_24449,N_24567);
xor U24760 (N_24760,N_24528,N_24598);
nor U24761 (N_24761,N_24480,N_24542);
and U24762 (N_24762,N_24543,N_24436);
nor U24763 (N_24763,N_24413,N_24522);
xor U24764 (N_24764,N_24596,N_24565);
nand U24765 (N_24765,N_24582,N_24561);
or U24766 (N_24766,N_24596,N_24462);
and U24767 (N_24767,N_24402,N_24442);
nor U24768 (N_24768,N_24539,N_24483);
nand U24769 (N_24769,N_24461,N_24501);
nor U24770 (N_24770,N_24473,N_24582);
xnor U24771 (N_24771,N_24447,N_24552);
or U24772 (N_24772,N_24554,N_24567);
nor U24773 (N_24773,N_24496,N_24587);
nand U24774 (N_24774,N_24504,N_24508);
xnor U24775 (N_24775,N_24567,N_24461);
nor U24776 (N_24776,N_24506,N_24404);
nor U24777 (N_24777,N_24536,N_24442);
nor U24778 (N_24778,N_24447,N_24414);
nor U24779 (N_24779,N_24444,N_24507);
xnor U24780 (N_24780,N_24524,N_24513);
nand U24781 (N_24781,N_24536,N_24424);
xor U24782 (N_24782,N_24558,N_24417);
nor U24783 (N_24783,N_24440,N_24477);
xor U24784 (N_24784,N_24512,N_24593);
nand U24785 (N_24785,N_24579,N_24584);
and U24786 (N_24786,N_24538,N_24534);
xnor U24787 (N_24787,N_24423,N_24426);
nand U24788 (N_24788,N_24523,N_24517);
nand U24789 (N_24789,N_24524,N_24525);
nand U24790 (N_24790,N_24419,N_24580);
nand U24791 (N_24791,N_24502,N_24548);
nand U24792 (N_24792,N_24578,N_24405);
nor U24793 (N_24793,N_24417,N_24556);
or U24794 (N_24794,N_24418,N_24469);
or U24795 (N_24795,N_24502,N_24473);
and U24796 (N_24796,N_24513,N_24467);
or U24797 (N_24797,N_24594,N_24591);
nor U24798 (N_24798,N_24534,N_24443);
nor U24799 (N_24799,N_24522,N_24429);
xor U24800 (N_24800,N_24657,N_24732);
nor U24801 (N_24801,N_24799,N_24717);
nand U24802 (N_24802,N_24796,N_24630);
nor U24803 (N_24803,N_24793,N_24679);
nor U24804 (N_24804,N_24763,N_24726);
xor U24805 (N_24805,N_24733,N_24741);
nor U24806 (N_24806,N_24696,N_24685);
nand U24807 (N_24807,N_24601,N_24665);
or U24808 (N_24808,N_24683,N_24771);
and U24809 (N_24809,N_24765,N_24634);
and U24810 (N_24810,N_24609,N_24666);
and U24811 (N_24811,N_24739,N_24751);
or U24812 (N_24812,N_24667,N_24690);
nand U24813 (N_24813,N_24721,N_24744);
xnor U24814 (N_24814,N_24714,N_24757);
or U24815 (N_24815,N_24672,N_24737);
xor U24816 (N_24816,N_24627,N_24776);
nand U24817 (N_24817,N_24719,N_24700);
or U24818 (N_24818,N_24727,N_24663);
nor U24819 (N_24819,N_24770,N_24649);
nand U24820 (N_24820,N_24633,N_24754);
nand U24821 (N_24821,N_24798,N_24718);
nand U24822 (N_24822,N_24781,N_24640);
nand U24823 (N_24823,N_24713,N_24661);
nor U24824 (N_24824,N_24703,N_24622);
nor U24825 (N_24825,N_24674,N_24774);
or U24826 (N_24826,N_24606,N_24785);
and U24827 (N_24827,N_24753,N_24682);
nor U24828 (N_24828,N_24600,N_24736);
nand U24829 (N_24829,N_24660,N_24759);
nor U24830 (N_24830,N_24698,N_24791);
nand U24831 (N_24831,N_24687,N_24623);
or U24832 (N_24832,N_24626,N_24694);
or U24833 (N_24833,N_24607,N_24648);
xor U24834 (N_24834,N_24629,N_24605);
xor U24835 (N_24835,N_24693,N_24642);
or U24836 (N_24836,N_24624,N_24653);
and U24837 (N_24837,N_24738,N_24699);
and U24838 (N_24838,N_24631,N_24614);
and U24839 (N_24839,N_24659,N_24706);
nor U24840 (N_24840,N_24745,N_24787);
or U24841 (N_24841,N_24794,N_24767);
nor U24842 (N_24842,N_24777,N_24613);
nor U24843 (N_24843,N_24650,N_24701);
xnor U24844 (N_24844,N_24654,N_24724);
nand U24845 (N_24845,N_24716,N_24681);
nand U24846 (N_24846,N_24638,N_24680);
or U24847 (N_24847,N_24750,N_24628);
and U24848 (N_24848,N_24677,N_24784);
or U24849 (N_24849,N_24782,N_24684);
xnor U24850 (N_24850,N_24612,N_24779);
nand U24851 (N_24851,N_24675,N_24773);
nand U24852 (N_24852,N_24789,N_24655);
or U24853 (N_24853,N_24742,N_24695);
nand U24854 (N_24854,N_24651,N_24720);
xnor U24855 (N_24855,N_24611,N_24615);
and U24856 (N_24856,N_24604,N_24725);
xnor U24857 (N_24857,N_24692,N_24722);
or U24858 (N_24858,N_24748,N_24790);
or U24859 (N_24859,N_24652,N_24710);
or U24860 (N_24860,N_24632,N_24620);
xor U24861 (N_24861,N_24702,N_24641);
and U24862 (N_24862,N_24731,N_24616);
or U24863 (N_24863,N_24755,N_24656);
xnor U24864 (N_24864,N_24617,N_24752);
and U24865 (N_24865,N_24729,N_24610);
nor U24866 (N_24866,N_24673,N_24709);
or U24867 (N_24867,N_24780,N_24715);
nand U24868 (N_24868,N_24669,N_24734);
and U24869 (N_24869,N_24708,N_24768);
xor U24870 (N_24870,N_24761,N_24688);
nand U24871 (N_24871,N_24668,N_24635);
or U24872 (N_24872,N_24728,N_24662);
or U24873 (N_24873,N_24764,N_24792);
and U24874 (N_24874,N_24644,N_24712);
nand U24875 (N_24875,N_24691,N_24772);
nor U24876 (N_24876,N_24797,N_24735);
and U24877 (N_24877,N_24658,N_24670);
and U24878 (N_24878,N_24676,N_24643);
or U24879 (N_24879,N_24678,N_24740);
nand U24880 (N_24880,N_24711,N_24760);
xnor U24881 (N_24881,N_24775,N_24778);
nor U24882 (N_24882,N_24664,N_24697);
xor U24883 (N_24883,N_24621,N_24686);
or U24884 (N_24884,N_24689,N_24758);
nor U24885 (N_24885,N_24769,N_24705);
and U24886 (N_24886,N_24788,N_24645);
nor U24887 (N_24887,N_24762,N_24730);
nor U24888 (N_24888,N_24625,N_24637);
xnor U24889 (N_24889,N_24756,N_24704);
nand U24890 (N_24890,N_24618,N_24619);
xnor U24891 (N_24891,N_24747,N_24749);
xor U24892 (N_24892,N_24707,N_24786);
nand U24893 (N_24893,N_24603,N_24602);
xor U24894 (N_24894,N_24636,N_24795);
or U24895 (N_24895,N_24671,N_24646);
or U24896 (N_24896,N_24766,N_24608);
xnor U24897 (N_24897,N_24723,N_24746);
and U24898 (N_24898,N_24639,N_24743);
and U24899 (N_24899,N_24783,N_24647);
nand U24900 (N_24900,N_24722,N_24639);
and U24901 (N_24901,N_24677,N_24735);
nor U24902 (N_24902,N_24687,N_24791);
nand U24903 (N_24903,N_24644,N_24666);
nand U24904 (N_24904,N_24679,N_24660);
and U24905 (N_24905,N_24624,N_24732);
nor U24906 (N_24906,N_24685,N_24651);
nand U24907 (N_24907,N_24745,N_24622);
and U24908 (N_24908,N_24739,N_24651);
nor U24909 (N_24909,N_24778,N_24622);
xor U24910 (N_24910,N_24688,N_24700);
xor U24911 (N_24911,N_24761,N_24718);
xnor U24912 (N_24912,N_24612,N_24685);
or U24913 (N_24913,N_24684,N_24656);
nor U24914 (N_24914,N_24773,N_24735);
nor U24915 (N_24915,N_24774,N_24692);
nor U24916 (N_24916,N_24607,N_24732);
nand U24917 (N_24917,N_24703,N_24717);
xor U24918 (N_24918,N_24696,N_24601);
xnor U24919 (N_24919,N_24791,N_24679);
and U24920 (N_24920,N_24613,N_24712);
nor U24921 (N_24921,N_24712,N_24719);
nand U24922 (N_24922,N_24730,N_24738);
or U24923 (N_24923,N_24676,N_24651);
and U24924 (N_24924,N_24657,N_24730);
nor U24925 (N_24925,N_24679,N_24663);
nand U24926 (N_24926,N_24693,N_24775);
nand U24927 (N_24927,N_24620,N_24717);
nor U24928 (N_24928,N_24636,N_24670);
nor U24929 (N_24929,N_24781,N_24600);
and U24930 (N_24930,N_24788,N_24707);
nor U24931 (N_24931,N_24705,N_24773);
nor U24932 (N_24932,N_24712,N_24673);
or U24933 (N_24933,N_24640,N_24623);
or U24934 (N_24934,N_24655,N_24758);
or U24935 (N_24935,N_24791,N_24776);
and U24936 (N_24936,N_24784,N_24772);
nor U24937 (N_24937,N_24747,N_24786);
and U24938 (N_24938,N_24607,N_24778);
nor U24939 (N_24939,N_24672,N_24726);
and U24940 (N_24940,N_24618,N_24707);
xnor U24941 (N_24941,N_24785,N_24695);
xor U24942 (N_24942,N_24696,N_24649);
xor U24943 (N_24943,N_24707,N_24757);
xnor U24944 (N_24944,N_24717,N_24607);
nand U24945 (N_24945,N_24646,N_24657);
or U24946 (N_24946,N_24756,N_24665);
or U24947 (N_24947,N_24614,N_24710);
and U24948 (N_24948,N_24675,N_24671);
nor U24949 (N_24949,N_24671,N_24637);
and U24950 (N_24950,N_24660,N_24775);
nand U24951 (N_24951,N_24727,N_24759);
or U24952 (N_24952,N_24616,N_24615);
or U24953 (N_24953,N_24692,N_24715);
or U24954 (N_24954,N_24635,N_24720);
and U24955 (N_24955,N_24775,N_24723);
and U24956 (N_24956,N_24698,N_24676);
nand U24957 (N_24957,N_24779,N_24732);
nor U24958 (N_24958,N_24733,N_24625);
nor U24959 (N_24959,N_24709,N_24722);
nand U24960 (N_24960,N_24718,N_24748);
xnor U24961 (N_24961,N_24638,N_24676);
or U24962 (N_24962,N_24776,N_24681);
nand U24963 (N_24963,N_24718,N_24711);
nor U24964 (N_24964,N_24717,N_24739);
and U24965 (N_24965,N_24627,N_24772);
and U24966 (N_24966,N_24712,N_24788);
and U24967 (N_24967,N_24722,N_24707);
xnor U24968 (N_24968,N_24630,N_24752);
or U24969 (N_24969,N_24749,N_24739);
xor U24970 (N_24970,N_24670,N_24699);
xnor U24971 (N_24971,N_24640,N_24721);
xor U24972 (N_24972,N_24713,N_24762);
xor U24973 (N_24973,N_24790,N_24740);
nor U24974 (N_24974,N_24764,N_24759);
nand U24975 (N_24975,N_24778,N_24709);
or U24976 (N_24976,N_24782,N_24757);
nor U24977 (N_24977,N_24636,N_24657);
or U24978 (N_24978,N_24679,N_24619);
nand U24979 (N_24979,N_24725,N_24745);
nor U24980 (N_24980,N_24772,N_24631);
nor U24981 (N_24981,N_24718,N_24725);
or U24982 (N_24982,N_24688,N_24682);
and U24983 (N_24983,N_24609,N_24724);
nand U24984 (N_24984,N_24749,N_24732);
or U24985 (N_24985,N_24772,N_24693);
nor U24986 (N_24986,N_24746,N_24741);
or U24987 (N_24987,N_24705,N_24655);
nor U24988 (N_24988,N_24693,N_24661);
nor U24989 (N_24989,N_24767,N_24754);
and U24990 (N_24990,N_24773,N_24778);
nand U24991 (N_24991,N_24740,N_24732);
or U24992 (N_24992,N_24785,N_24696);
or U24993 (N_24993,N_24760,N_24620);
nor U24994 (N_24994,N_24715,N_24747);
or U24995 (N_24995,N_24639,N_24770);
nor U24996 (N_24996,N_24604,N_24685);
or U24997 (N_24997,N_24685,N_24752);
and U24998 (N_24998,N_24671,N_24654);
or U24999 (N_24999,N_24615,N_24736);
xnor UO_0 (O_0,N_24815,N_24829);
nand UO_1 (O_1,N_24883,N_24901);
nand UO_2 (O_2,N_24891,N_24861);
xor UO_3 (O_3,N_24852,N_24917);
and UO_4 (O_4,N_24870,N_24949);
nor UO_5 (O_5,N_24988,N_24800);
nor UO_6 (O_6,N_24951,N_24854);
nand UO_7 (O_7,N_24801,N_24804);
nand UO_8 (O_8,N_24997,N_24895);
nor UO_9 (O_9,N_24907,N_24911);
nor UO_10 (O_10,N_24809,N_24953);
nand UO_11 (O_11,N_24814,N_24961);
or UO_12 (O_12,N_24827,N_24900);
or UO_13 (O_13,N_24986,N_24959);
nand UO_14 (O_14,N_24899,N_24926);
and UO_15 (O_15,N_24947,N_24914);
nand UO_16 (O_16,N_24924,N_24821);
or UO_17 (O_17,N_24892,N_24940);
and UO_18 (O_18,N_24882,N_24989);
and UO_19 (O_19,N_24964,N_24972);
nand UO_20 (O_20,N_24876,N_24832);
nor UO_21 (O_21,N_24810,N_24866);
xor UO_22 (O_22,N_24849,N_24839);
nor UO_23 (O_23,N_24845,N_24871);
nor UO_24 (O_24,N_24824,N_24887);
or UO_25 (O_25,N_24803,N_24856);
xor UO_26 (O_26,N_24930,N_24933);
xor UO_27 (O_27,N_24934,N_24807);
or UO_28 (O_28,N_24982,N_24968);
or UO_29 (O_29,N_24987,N_24868);
or UO_30 (O_30,N_24975,N_24913);
nor UO_31 (O_31,N_24909,N_24830);
nand UO_32 (O_32,N_24879,N_24908);
xor UO_33 (O_33,N_24880,N_24978);
or UO_34 (O_34,N_24826,N_24806);
nand UO_35 (O_35,N_24819,N_24939);
or UO_36 (O_36,N_24973,N_24983);
nand UO_37 (O_37,N_24840,N_24812);
and UO_38 (O_38,N_24874,N_24898);
or UO_39 (O_39,N_24817,N_24950);
nor UO_40 (O_40,N_24920,N_24842);
nand UO_41 (O_41,N_24936,N_24831);
or UO_42 (O_42,N_24867,N_24962);
or UO_43 (O_43,N_24935,N_24872);
xor UO_44 (O_44,N_24932,N_24991);
nor UO_45 (O_45,N_24836,N_24881);
xor UO_46 (O_46,N_24999,N_24910);
xnor UO_47 (O_47,N_24890,N_24805);
and UO_48 (O_48,N_24941,N_24837);
or UO_49 (O_49,N_24848,N_24984);
nand UO_50 (O_50,N_24843,N_24902);
xnor UO_51 (O_51,N_24858,N_24860);
xor UO_52 (O_52,N_24931,N_24956);
xor UO_53 (O_53,N_24993,N_24938);
nand UO_54 (O_54,N_24925,N_24969);
nor UO_55 (O_55,N_24808,N_24981);
and UO_56 (O_56,N_24980,N_24893);
and UO_57 (O_57,N_24928,N_24977);
or UO_58 (O_58,N_24967,N_24915);
or UO_59 (O_59,N_24822,N_24853);
xnor UO_60 (O_60,N_24888,N_24954);
and UO_61 (O_61,N_24864,N_24875);
xor UO_62 (O_62,N_24825,N_24841);
nor UO_63 (O_63,N_24922,N_24957);
xor UO_64 (O_64,N_24995,N_24921);
and UO_65 (O_65,N_24990,N_24945);
xor UO_66 (O_66,N_24885,N_24994);
xor UO_67 (O_67,N_24835,N_24912);
nand UO_68 (O_68,N_24966,N_24904);
and UO_69 (O_69,N_24862,N_24865);
or UO_70 (O_70,N_24873,N_24963);
nor UO_71 (O_71,N_24850,N_24919);
nand UO_72 (O_72,N_24823,N_24886);
xor UO_73 (O_73,N_24929,N_24863);
and UO_74 (O_74,N_24958,N_24884);
xor UO_75 (O_75,N_24857,N_24894);
or UO_76 (O_76,N_24844,N_24952);
xnor UO_77 (O_77,N_24802,N_24976);
and UO_78 (O_78,N_24974,N_24897);
nor UO_79 (O_79,N_24979,N_24906);
nand UO_80 (O_80,N_24878,N_24813);
and UO_81 (O_81,N_24903,N_24851);
or UO_82 (O_82,N_24846,N_24985);
xor UO_83 (O_83,N_24955,N_24905);
nand UO_84 (O_84,N_24943,N_24918);
or UO_85 (O_85,N_24818,N_24889);
nor UO_86 (O_86,N_24811,N_24927);
and UO_87 (O_87,N_24847,N_24834);
nor UO_88 (O_88,N_24948,N_24944);
nand UO_89 (O_89,N_24877,N_24946);
xor UO_90 (O_90,N_24923,N_24998);
xnor UO_91 (O_91,N_24960,N_24833);
and UO_92 (O_92,N_24992,N_24916);
or UO_93 (O_93,N_24859,N_24937);
nand UO_94 (O_94,N_24896,N_24970);
and UO_95 (O_95,N_24942,N_24820);
xnor UO_96 (O_96,N_24869,N_24838);
and UO_97 (O_97,N_24965,N_24828);
and UO_98 (O_98,N_24855,N_24816);
xor UO_99 (O_99,N_24971,N_24996);
nand UO_100 (O_100,N_24836,N_24957);
xor UO_101 (O_101,N_24927,N_24837);
and UO_102 (O_102,N_24821,N_24995);
or UO_103 (O_103,N_24909,N_24928);
nand UO_104 (O_104,N_24863,N_24915);
nand UO_105 (O_105,N_24853,N_24856);
nor UO_106 (O_106,N_24879,N_24938);
and UO_107 (O_107,N_24932,N_24844);
nand UO_108 (O_108,N_24946,N_24906);
or UO_109 (O_109,N_24959,N_24899);
nand UO_110 (O_110,N_24878,N_24855);
or UO_111 (O_111,N_24820,N_24928);
xnor UO_112 (O_112,N_24846,N_24915);
nor UO_113 (O_113,N_24993,N_24935);
nor UO_114 (O_114,N_24988,N_24901);
or UO_115 (O_115,N_24995,N_24902);
and UO_116 (O_116,N_24896,N_24930);
nor UO_117 (O_117,N_24896,N_24937);
xnor UO_118 (O_118,N_24890,N_24882);
or UO_119 (O_119,N_24867,N_24827);
nand UO_120 (O_120,N_24948,N_24822);
nor UO_121 (O_121,N_24837,N_24840);
xnor UO_122 (O_122,N_24854,N_24857);
nand UO_123 (O_123,N_24917,N_24899);
xnor UO_124 (O_124,N_24817,N_24913);
xnor UO_125 (O_125,N_24937,N_24802);
nand UO_126 (O_126,N_24971,N_24990);
and UO_127 (O_127,N_24993,N_24945);
and UO_128 (O_128,N_24827,N_24998);
nor UO_129 (O_129,N_24866,N_24826);
xor UO_130 (O_130,N_24976,N_24981);
and UO_131 (O_131,N_24918,N_24871);
or UO_132 (O_132,N_24867,N_24888);
and UO_133 (O_133,N_24921,N_24964);
nand UO_134 (O_134,N_24912,N_24886);
nor UO_135 (O_135,N_24841,N_24804);
xnor UO_136 (O_136,N_24933,N_24995);
and UO_137 (O_137,N_24865,N_24819);
and UO_138 (O_138,N_24841,N_24808);
and UO_139 (O_139,N_24969,N_24886);
xor UO_140 (O_140,N_24828,N_24874);
or UO_141 (O_141,N_24988,N_24893);
nand UO_142 (O_142,N_24949,N_24804);
nor UO_143 (O_143,N_24841,N_24842);
and UO_144 (O_144,N_24829,N_24941);
nand UO_145 (O_145,N_24801,N_24903);
nand UO_146 (O_146,N_24907,N_24848);
and UO_147 (O_147,N_24947,N_24932);
nand UO_148 (O_148,N_24890,N_24816);
nand UO_149 (O_149,N_24938,N_24855);
or UO_150 (O_150,N_24962,N_24986);
nand UO_151 (O_151,N_24889,N_24931);
xnor UO_152 (O_152,N_24978,N_24910);
xor UO_153 (O_153,N_24897,N_24861);
nor UO_154 (O_154,N_24969,N_24944);
and UO_155 (O_155,N_24964,N_24986);
xnor UO_156 (O_156,N_24874,N_24894);
nor UO_157 (O_157,N_24967,N_24881);
xor UO_158 (O_158,N_24856,N_24887);
and UO_159 (O_159,N_24950,N_24917);
or UO_160 (O_160,N_24822,N_24860);
and UO_161 (O_161,N_24975,N_24864);
xor UO_162 (O_162,N_24964,N_24899);
or UO_163 (O_163,N_24858,N_24865);
xor UO_164 (O_164,N_24916,N_24820);
nor UO_165 (O_165,N_24879,N_24865);
xnor UO_166 (O_166,N_24925,N_24872);
nand UO_167 (O_167,N_24993,N_24984);
xor UO_168 (O_168,N_24908,N_24947);
nand UO_169 (O_169,N_24894,N_24923);
or UO_170 (O_170,N_24957,N_24806);
nand UO_171 (O_171,N_24815,N_24847);
nor UO_172 (O_172,N_24847,N_24948);
and UO_173 (O_173,N_24915,N_24848);
and UO_174 (O_174,N_24831,N_24879);
or UO_175 (O_175,N_24927,N_24929);
or UO_176 (O_176,N_24856,N_24967);
nor UO_177 (O_177,N_24862,N_24843);
and UO_178 (O_178,N_24966,N_24938);
nor UO_179 (O_179,N_24991,N_24921);
and UO_180 (O_180,N_24905,N_24834);
or UO_181 (O_181,N_24985,N_24822);
nand UO_182 (O_182,N_24947,N_24912);
nand UO_183 (O_183,N_24871,N_24932);
xnor UO_184 (O_184,N_24978,N_24960);
and UO_185 (O_185,N_24934,N_24919);
nand UO_186 (O_186,N_24822,N_24868);
or UO_187 (O_187,N_24885,N_24803);
xnor UO_188 (O_188,N_24892,N_24861);
and UO_189 (O_189,N_24871,N_24861);
and UO_190 (O_190,N_24916,N_24892);
and UO_191 (O_191,N_24804,N_24962);
or UO_192 (O_192,N_24828,N_24920);
nand UO_193 (O_193,N_24815,N_24823);
nor UO_194 (O_194,N_24934,N_24914);
nor UO_195 (O_195,N_24835,N_24900);
nor UO_196 (O_196,N_24899,N_24834);
and UO_197 (O_197,N_24914,N_24901);
nand UO_198 (O_198,N_24848,N_24971);
or UO_199 (O_199,N_24946,N_24864);
or UO_200 (O_200,N_24989,N_24970);
xnor UO_201 (O_201,N_24946,N_24817);
xor UO_202 (O_202,N_24862,N_24951);
nor UO_203 (O_203,N_24841,N_24800);
or UO_204 (O_204,N_24809,N_24978);
or UO_205 (O_205,N_24877,N_24886);
and UO_206 (O_206,N_24906,N_24891);
xor UO_207 (O_207,N_24815,N_24869);
nor UO_208 (O_208,N_24963,N_24863);
nand UO_209 (O_209,N_24872,N_24937);
xor UO_210 (O_210,N_24880,N_24985);
nor UO_211 (O_211,N_24938,N_24974);
nor UO_212 (O_212,N_24833,N_24930);
and UO_213 (O_213,N_24997,N_24815);
nand UO_214 (O_214,N_24860,N_24980);
xnor UO_215 (O_215,N_24809,N_24946);
or UO_216 (O_216,N_24869,N_24816);
nor UO_217 (O_217,N_24930,N_24959);
xor UO_218 (O_218,N_24879,N_24891);
nand UO_219 (O_219,N_24904,N_24891);
nand UO_220 (O_220,N_24857,N_24828);
xor UO_221 (O_221,N_24908,N_24878);
or UO_222 (O_222,N_24970,N_24996);
or UO_223 (O_223,N_24897,N_24835);
xor UO_224 (O_224,N_24859,N_24895);
nand UO_225 (O_225,N_24934,N_24916);
nor UO_226 (O_226,N_24956,N_24935);
nand UO_227 (O_227,N_24936,N_24927);
xor UO_228 (O_228,N_24833,N_24902);
nand UO_229 (O_229,N_24816,N_24896);
nand UO_230 (O_230,N_24849,N_24989);
nand UO_231 (O_231,N_24805,N_24951);
or UO_232 (O_232,N_24956,N_24859);
or UO_233 (O_233,N_24855,N_24974);
nor UO_234 (O_234,N_24915,N_24904);
nand UO_235 (O_235,N_24843,N_24868);
xor UO_236 (O_236,N_24938,N_24914);
nor UO_237 (O_237,N_24938,N_24880);
nand UO_238 (O_238,N_24963,N_24939);
nand UO_239 (O_239,N_24914,N_24891);
nor UO_240 (O_240,N_24898,N_24988);
nand UO_241 (O_241,N_24834,N_24924);
nand UO_242 (O_242,N_24809,N_24854);
and UO_243 (O_243,N_24924,N_24893);
and UO_244 (O_244,N_24967,N_24943);
or UO_245 (O_245,N_24840,N_24906);
and UO_246 (O_246,N_24981,N_24909);
nor UO_247 (O_247,N_24984,N_24928);
or UO_248 (O_248,N_24966,N_24895);
nor UO_249 (O_249,N_24932,N_24846);
and UO_250 (O_250,N_24857,N_24914);
nand UO_251 (O_251,N_24945,N_24902);
nand UO_252 (O_252,N_24955,N_24942);
or UO_253 (O_253,N_24980,N_24864);
and UO_254 (O_254,N_24828,N_24847);
nor UO_255 (O_255,N_24902,N_24809);
nand UO_256 (O_256,N_24934,N_24909);
nand UO_257 (O_257,N_24998,N_24944);
or UO_258 (O_258,N_24944,N_24845);
nand UO_259 (O_259,N_24810,N_24928);
nand UO_260 (O_260,N_24823,N_24900);
xnor UO_261 (O_261,N_24876,N_24896);
nor UO_262 (O_262,N_24854,N_24910);
and UO_263 (O_263,N_24894,N_24846);
or UO_264 (O_264,N_24875,N_24995);
nand UO_265 (O_265,N_24841,N_24965);
nand UO_266 (O_266,N_24994,N_24884);
or UO_267 (O_267,N_24998,N_24893);
and UO_268 (O_268,N_24828,N_24945);
or UO_269 (O_269,N_24812,N_24855);
nor UO_270 (O_270,N_24804,N_24965);
nand UO_271 (O_271,N_24821,N_24938);
nor UO_272 (O_272,N_24911,N_24968);
xnor UO_273 (O_273,N_24835,N_24823);
xor UO_274 (O_274,N_24896,N_24993);
xor UO_275 (O_275,N_24821,N_24840);
nand UO_276 (O_276,N_24862,N_24999);
nor UO_277 (O_277,N_24976,N_24870);
xnor UO_278 (O_278,N_24800,N_24801);
nor UO_279 (O_279,N_24892,N_24845);
or UO_280 (O_280,N_24953,N_24984);
xor UO_281 (O_281,N_24843,N_24847);
xnor UO_282 (O_282,N_24897,N_24921);
or UO_283 (O_283,N_24951,N_24967);
nand UO_284 (O_284,N_24897,N_24807);
and UO_285 (O_285,N_24890,N_24957);
or UO_286 (O_286,N_24917,N_24952);
xor UO_287 (O_287,N_24908,N_24969);
nand UO_288 (O_288,N_24912,N_24922);
or UO_289 (O_289,N_24952,N_24826);
nand UO_290 (O_290,N_24912,N_24846);
xor UO_291 (O_291,N_24973,N_24972);
xnor UO_292 (O_292,N_24921,N_24944);
xnor UO_293 (O_293,N_24969,N_24870);
nand UO_294 (O_294,N_24929,N_24992);
nand UO_295 (O_295,N_24853,N_24974);
or UO_296 (O_296,N_24853,N_24952);
nand UO_297 (O_297,N_24964,N_24805);
and UO_298 (O_298,N_24969,N_24956);
nand UO_299 (O_299,N_24958,N_24981);
or UO_300 (O_300,N_24870,N_24861);
or UO_301 (O_301,N_24997,N_24931);
nand UO_302 (O_302,N_24838,N_24904);
nor UO_303 (O_303,N_24856,N_24845);
xnor UO_304 (O_304,N_24920,N_24800);
or UO_305 (O_305,N_24802,N_24897);
or UO_306 (O_306,N_24916,N_24910);
and UO_307 (O_307,N_24812,N_24881);
and UO_308 (O_308,N_24947,N_24955);
and UO_309 (O_309,N_24981,N_24926);
xnor UO_310 (O_310,N_24976,N_24986);
nor UO_311 (O_311,N_24933,N_24890);
nor UO_312 (O_312,N_24981,N_24894);
nand UO_313 (O_313,N_24806,N_24945);
and UO_314 (O_314,N_24940,N_24812);
or UO_315 (O_315,N_24805,N_24932);
xor UO_316 (O_316,N_24840,N_24981);
nand UO_317 (O_317,N_24902,N_24903);
nand UO_318 (O_318,N_24914,N_24910);
and UO_319 (O_319,N_24873,N_24894);
xnor UO_320 (O_320,N_24825,N_24818);
or UO_321 (O_321,N_24820,N_24972);
nand UO_322 (O_322,N_24996,N_24868);
xnor UO_323 (O_323,N_24803,N_24807);
and UO_324 (O_324,N_24848,N_24802);
and UO_325 (O_325,N_24941,N_24811);
and UO_326 (O_326,N_24935,N_24885);
or UO_327 (O_327,N_24830,N_24943);
nor UO_328 (O_328,N_24875,N_24924);
nor UO_329 (O_329,N_24843,N_24829);
and UO_330 (O_330,N_24885,N_24829);
or UO_331 (O_331,N_24976,N_24972);
nor UO_332 (O_332,N_24911,N_24878);
or UO_333 (O_333,N_24807,N_24809);
xor UO_334 (O_334,N_24948,N_24919);
nand UO_335 (O_335,N_24830,N_24871);
and UO_336 (O_336,N_24803,N_24835);
or UO_337 (O_337,N_24968,N_24998);
nor UO_338 (O_338,N_24879,N_24887);
xnor UO_339 (O_339,N_24826,N_24813);
nor UO_340 (O_340,N_24991,N_24823);
nor UO_341 (O_341,N_24895,N_24907);
and UO_342 (O_342,N_24924,N_24896);
and UO_343 (O_343,N_24870,N_24971);
or UO_344 (O_344,N_24985,N_24843);
nand UO_345 (O_345,N_24998,N_24890);
xnor UO_346 (O_346,N_24807,N_24922);
xor UO_347 (O_347,N_24820,N_24943);
and UO_348 (O_348,N_24875,N_24918);
nand UO_349 (O_349,N_24902,N_24963);
and UO_350 (O_350,N_24976,N_24823);
and UO_351 (O_351,N_24833,N_24938);
nand UO_352 (O_352,N_24891,N_24852);
or UO_353 (O_353,N_24821,N_24915);
nand UO_354 (O_354,N_24859,N_24874);
nand UO_355 (O_355,N_24830,N_24837);
xor UO_356 (O_356,N_24979,N_24999);
or UO_357 (O_357,N_24888,N_24882);
or UO_358 (O_358,N_24827,N_24886);
and UO_359 (O_359,N_24816,N_24951);
and UO_360 (O_360,N_24849,N_24935);
and UO_361 (O_361,N_24831,N_24902);
and UO_362 (O_362,N_24958,N_24975);
or UO_363 (O_363,N_24862,N_24965);
xor UO_364 (O_364,N_24846,N_24892);
xnor UO_365 (O_365,N_24888,N_24940);
nand UO_366 (O_366,N_24868,N_24960);
nor UO_367 (O_367,N_24890,N_24886);
xor UO_368 (O_368,N_24850,N_24961);
nor UO_369 (O_369,N_24886,N_24818);
nor UO_370 (O_370,N_24905,N_24909);
xor UO_371 (O_371,N_24846,N_24890);
and UO_372 (O_372,N_24806,N_24984);
xnor UO_373 (O_373,N_24885,N_24836);
nand UO_374 (O_374,N_24923,N_24999);
nand UO_375 (O_375,N_24805,N_24876);
and UO_376 (O_376,N_24833,N_24979);
nor UO_377 (O_377,N_24890,N_24953);
nand UO_378 (O_378,N_24919,N_24939);
and UO_379 (O_379,N_24849,N_24955);
or UO_380 (O_380,N_24816,N_24832);
and UO_381 (O_381,N_24917,N_24846);
and UO_382 (O_382,N_24988,N_24891);
and UO_383 (O_383,N_24841,N_24853);
xnor UO_384 (O_384,N_24963,N_24960);
xor UO_385 (O_385,N_24859,N_24949);
nand UO_386 (O_386,N_24876,N_24938);
xor UO_387 (O_387,N_24935,N_24837);
nand UO_388 (O_388,N_24936,N_24813);
nand UO_389 (O_389,N_24885,N_24961);
xor UO_390 (O_390,N_24870,N_24816);
nor UO_391 (O_391,N_24896,N_24992);
nand UO_392 (O_392,N_24928,N_24818);
and UO_393 (O_393,N_24824,N_24934);
nor UO_394 (O_394,N_24958,N_24841);
nor UO_395 (O_395,N_24847,N_24964);
nand UO_396 (O_396,N_24800,N_24812);
nor UO_397 (O_397,N_24927,N_24970);
or UO_398 (O_398,N_24893,N_24967);
and UO_399 (O_399,N_24858,N_24857);
nor UO_400 (O_400,N_24841,N_24935);
nand UO_401 (O_401,N_24926,N_24930);
nor UO_402 (O_402,N_24973,N_24925);
nor UO_403 (O_403,N_24908,N_24948);
nor UO_404 (O_404,N_24967,N_24857);
or UO_405 (O_405,N_24887,N_24815);
nor UO_406 (O_406,N_24812,N_24916);
nor UO_407 (O_407,N_24890,N_24811);
or UO_408 (O_408,N_24827,N_24962);
or UO_409 (O_409,N_24951,N_24847);
or UO_410 (O_410,N_24964,N_24994);
nor UO_411 (O_411,N_24988,N_24832);
nand UO_412 (O_412,N_24869,N_24835);
and UO_413 (O_413,N_24903,N_24931);
xor UO_414 (O_414,N_24816,N_24868);
xnor UO_415 (O_415,N_24829,N_24883);
nand UO_416 (O_416,N_24810,N_24803);
nor UO_417 (O_417,N_24826,N_24855);
and UO_418 (O_418,N_24865,N_24876);
nand UO_419 (O_419,N_24978,N_24931);
or UO_420 (O_420,N_24801,N_24908);
or UO_421 (O_421,N_24821,N_24943);
xor UO_422 (O_422,N_24970,N_24829);
nor UO_423 (O_423,N_24969,N_24867);
nor UO_424 (O_424,N_24973,N_24981);
nor UO_425 (O_425,N_24975,N_24963);
or UO_426 (O_426,N_24938,N_24975);
xor UO_427 (O_427,N_24894,N_24915);
or UO_428 (O_428,N_24995,N_24934);
nor UO_429 (O_429,N_24952,N_24836);
nand UO_430 (O_430,N_24901,N_24842);
nand UO_431 (O_431,N_24891,N_24943);
and UO_432 (O_432,N_24977,N_24875);
xnor UO_433 (O_433,N_24802,N_24891);
or UO_434 (O_434,N_24820,N_24910);
and UO_435 (O_435,N_24867,N_24849);
and UO_436 (O_436,N_24824,N_24801);
or UO_437 (O_437,N_24871,N_24952);
xor UO_438 (O_438,N_24862,N_24815);
and UO_439 (O_439,N_24966,N_24817);
and UO_440 (O_440,N_24804,N_24838);
or UO_441 (O_441,N_24877,N_24970);
xnor UO_442 (O_442,N_24955,N_24896);
or UO_443 (O_443,N_24914,N_24882);
or UO_444 (O_444,N_24894,N_24850);
or UO_445 (O_445,N_24955,N_24930);
or UO_446 (O_446,N_24827,N_24880);
xnor UO_447 (O_447,N_24944,N_24883);
nor UO_448 (O_448,N_24929,N_24813);
xnor UO_449 (O_449,N_24932,N_24850);
or UO_450 (O_450,N_24807,N_24950);
xor UO_451 (O_451,N_24919,N_24932);
or UO_452 (O_452,N_24811,N_24935);
xnor UO_453 (O_453,N_24938,N_24916);
or UO_454 (O_454,N_24890,N_24830);
xor UO_455 (O_455,N_24800,N_24895);
or UO_456 (O_456,N_24868,N_24923);
and UO_457 (O_457,N_24960,N_24844);
xor UO_458 (O_458,N_24999,N_24843);
nor UO_459 (O_459,N_24943,N_24995);
and UO_460 (O_460,N_24801,N_24847);
xnor UO_461 (O_461,N_24961,N_24841);
nor UO_462 (O_462,N_24878,N_24847);
nand UO_463 (O_463,N_24844,N_24826);
or UO_464 (O_464,N_24956,N_24887);
and UO_465 (O_465,N_24862,N_24980);
and UO_466 (O_466,N_24909,N_24923);
or UO_467 (O_467,N_24966,N_24841);
or UO_468 (O_468,N_24866,N_24859);
or UO_469 (O_469,N_24939,N_24946);
nor UO_470 (O_470,N_24918,N_24890);
and UO_471 (O_471,N_24909,N_24860);
and UO_472 (O_472,N_24897,N_24940);
nand UO_473 (O_473,N_24842,N_24880);
and UO_474 (O_474,N_24997,N_24846);
or UO_475 (O_475,N_24899,N_24936);
and UO_476 (O_476,N_24991,N_24803);
xnor UO_477 (O_477,N_24868,N_24976);
or UO_478 (O_478,N_24968,N_24833);
nor UO_479 (O_479,N_24886,N_24838);
and UO_480 (O_480,N_24864,N_24970);
and UO_481 (O_481,N_24840,N_24844);
xnor UO_482 (O_482,N_24994,N_24939);
xnor UO_483 (O_483,N_24998,N_24851);
or UO_484 (O_484,N_24877,N_24823);
xnor UO_485 (O_485,N_24914,N_24945);
and UO_486 (O_486,N_24961,N_24832);
nand UO_487 (O_487,N_24830,N_24950);
or UO_488 (O_488,N_24882,N_24801);
or UO_489 (O_489,N_24872,N_24962);
and UO_490 (O_490,N_24829,N_24918);
nand UO_491 (O_491,N_24905,N_24822);
xor UO_492 (O_492,N_24867,N_24922);
nand UO_493 (O_493,N_24902,N_24856);
nor UO_494 (O_494,N_24816,N_24970);
nand UO_495 (O_495,N_24840,N_24946);
and UO_496 (O_496,N_24813,N_24904);
and UO_497 (O_497,N_24918,N_24886);
and UO_498 (O_498,N_24888,N_24943);
and UO_499 (O_499,N_24886,N_24896);
nand UO_500 (O_500,N_24969,N_24845);
nor UO_501 (O_501,N_24969,N_24855);
nor UO_502 (O_502,N_24929,N_24831);
nand UO_503 (O_503,N_24994,N_24947);
xnor UO_504 (O_504,N_24891,N_24925);
nor UO_505 (O_505,N_24844,N_24831);
xnor UO_506 (O_506,N_24904,N_24840);
nand UO_507 (O_507,N_24888,N_24854);
and UO_508 (O_508,N_24947,N_24855);
xnor UO_509 (O_509,N_24870,N_24894);
or UO_510 (O_510,N_24848,N_24836);
nor UO_511 (O_511,N_24894,N_24886);
nand UO_512 (O_512,N_24953,N_24852);
and UO_513 (O_513,N_24954,N_24913);
xnor UO_514 (O_514,N_24917,N_24996);
nor UO_515 (O_515,N_24833,N_24875);
xnor UO_516 (O_516,N_24933,N_24966);
and UO_517 (O_517,N_24835,N_24849);
nand UO_518 (O_518,N_24946,N_24835);
or UO_519 (O_519,N_24930,N_24882);
nand UO_520 (O_520,N_24891,N_24859);
nor UO_521 (O_521,N_24911,N_24803);
and UO_522 (O_522,N_24957,N_24960);
nand UO_523 (O_523,N_24954,N_24907);
nor UO_524 (O_524,N_24841,N_24836);
nand UO_525 (O_525,N_24986,N_24824);
nor UO_526 (O_526,N_24967,N_24871);
and UO_527 (O_527,N_24960,N_24950);
and UO_528 (O_528,N_24825,N_24877);
and UO_529 (O_529,N_24885,N_24910);
or UO_530 (O_530,N_24923,N_24834);
or UO_531 (O_531,N_24938,N_24800);
nor UO_532 (O_532,N_24841,N_24973);
nor UO_533 (O_533,N_24986,N_24949);
nor UO_534 (O_534,N_24834,N_24814);
or UO_535 (O_535,N_24802,N_24971);
or UO_536 (O_536,N_24804,N_24940);
nor UO_537 (O_537,N_24897,N_24830);
nor UO_538 (O_538,N_24838,N_24806);
nand UO_539 (O_539,N_24838,N_24997);
xnor UO_540 (O_540,N_24866,N_24954);
nor UO_541 (O_541,N_24915,N_24986);
xnor UO_542 (O_542,N_24896,N_24931);
and UO_543 (O_543,N_24935,N_24851);
nand UO_544 (O_544,N_24994,N_24821);
xor UO_545 (O_545,N_24959,N_24964);
nand UO_546 (O_546,N_24944,N_24865);
xor UO_547 (O_547,N_24933,N_24878);
and UO_548 (O_548,N_24929,N_24839);
and UO_549 (O_549,N_24877,N_24822);
and UO_550 (O_550,N_24927,N_24985);
xnor UO_551 (O_551,N_24972,N_24827);
nand UO_552 (O_552,N_24910,N_24880);
xor UO_553 (O_553,N_24823,N_24844);
or UO_554 (O_554,N_24929,N_24864);
or UO_555 (O_555,N_24894,N_24885);
and UO_556 (O_556,N_24849,N_24954);
xor UO_557 (O_557,N_24961,N_24942);
nand UO_558 (O_558,N_24893,N_24913);
nor UO_559 (O_559,N_24818,N_24907);
xnor UO_560 (O_560,N_24962,N_24947);
and UO_561 (O_561,N_24896,N_24947);
nor UO_562 (O_562,N_24852,N_24958);
nand UO_563 (O_563,N_24902,N_24987);
nand UO_564 (O_564,N_24826,N_24994);
or UO_565 (O_565,N_24843,N_24877);
xor UO_566 (O_566,N_24964,N_24940);
nand UO_567 (O_567,N_24860,N_24989);
or UO_568 (O_568,N_24908,N_24835);
nor UO_569 (O_569,N_24800,N_24910);
nor UO_570 (O_570,N_24949,N_24984);
nor UO_571 (O_571,N_24928,N_24877);
xor UO_572 (O_572,N_24907,N_24883);
xnor UO_573 (O_573,N_24959,N_24978);
and UO_574 (O_574,N_24812,N_24801);
or UO_575 (O_575,N_24808,N_24999);
nand UO_576 (O_576,N_24988,N_24948);
or UO_577 (O_577,N_24822,N_24989);
xnor UO_578 (O_578,N_24893,N_24935);
xnor UO_579 (O_579,N_24829,N_24856);
xnor UO_580 (O_580,N_24908,N_24917);
nand UO_581 (O_581,N_24837,N_24801);
or UO_582 (O_582,N_24870,N_24868);
and UO_583 (O_583,N_24842,N_24996);
xnor UO_584 (O_584,N_24800,N_24892);
or UO_585 (O_585,N_24833,N_24887);
and UO_586 (O_586,N_24962,N_24853);
xor UO_587 (O_587,N_24944,N_24997);
and UO_588 (O_588,N_24913,N_24904);
nor UO_589 (O_589,N_24966,N_24860);
or UO_590 (O_590,N_24944,N_24882);
xor UO_591 (O_591,N_24997,N_24893);
nor UO_592 (O_592,N_24918,N_24868);
or UO_593 (O_593,N_24876,N_24869);
and UO_594 (O_594,N_24950,N_24887);
xor UO_595 (O_595,N_24967,N_24823);
nand UO_596 (O_596,N_24822,N_24966);
nor UO_597 (O_597,N_24815,N_24990);
nor UO_598 (O_598,N_24832,N_24933);
xor UO_599 (O_599,N_24911,N_24808);
xor UO_600 (O_600,N_24885,N_24889);
xor UO_601 (O_601,N_24884,N_24961);
nand UO_602 (O_602,N_24868,N_24989);
nand UO_603 (O_603,N_24898,N_24858);
xnor UO_604 (O_604,N_24912,N_24901);
nor UO_605 (O_605,N_24803,N_24964);
and UO_606 (O_606,N_24809,N_24926);
or UO_607 (O_607,N_24867,N_24866);
nor UO_608 (O_608,N_24948,N_24985);
nand UO_609 (O_609,N_24941,N_24942);
nand UO_610 (O_610,N_24967,N_24879);
nor UO_611 (O_611,N_24945,N_24951);
and UO_612 (O_612,N_24844,N_24835);
nand UO_613 (O_613,N_24943,N_24985);
nand UO_614 (O_614,N_24877,N_24820);
and UO_615 (O_615,N_24858,N_24905);
or UO_616 (O_616,N_24972,N_24925);
xor UO_617 (O_617,N_24997,N_24896);
or UO_618 (O_618,N_24932,N_24948);
xor UO_619 (O_619,N_24880,N_24971);
and UO_620 (O_620,N_24974,N_24993);
and UO_621 (O_621,N_24988,N_24887);
or UO_622 (O_622,N_24817,N_24891);
xor UO_623 (O_623,N_24893,N_24851);
xor UO_624 (O_624,N_24936,N_24849);
nand UO_625 (O_625,N_24905,N_24800);
nor UO_626 (O_626,N_24803,N_24864);
nand UO_627 (O_627,N_24919,N_24821);
and UO_628 (O_628,N_24812,N_24997);
xor UO_629 (O_629,N_24871,N_24841);
or UO_630 (O_630,N_24821,N_24918);
nand UO_631 (O_631,N_24951,N_24995);
nor UO_632 (O_632,N_24832,N_24972);
or UO_633 (O_633,N_24983,N_24953);
nor UO_634 (O_634,N_24882,N_24974);
or UO_635 (O_635,N_24958,N_24877);
or UO_636 (O_636,N_24903,N_24811);
and UO_637 (O_637,N_24844,N_24955);
nor UO_638 (O_638,N_24968,N_24816);
nand UO_639 (O_639,N_24830,N_24838);
nand UO_640 (O_640,N_24995,N_24848);
or UO_641 (O_641,N_24836,N_24908);
nand UO_642 (O_642,N_24814,N_24866);
xor UO_643 (O_643,N_24805,N_24908);
xor UO_644 (O_644,N_24968,N_24887);
or UO_645 (O_645,N_24816,N_24830);
or UO_646 (O_646,N_24931,N_24982);
and UO_647 (O_647,N_24915,N_24884);
xnor UO_648 (O_648,N_24961,N_24979);
and UO_649 (O_649,N_24942,N_24917);
and UO_650 (O_650,N_24836,N_24937);
nand UO_651 (O_651,N_24888,N_24837);
and UO_652 (O_652,N_24868,N_24863);
or UO_653 (O_653,N_24984,N_24832);
nand UO_654 (O_654,N_24999,N_24975);
and UO_655 (O_655,N_24886,N_24881);
nand UO_656 (O_656,N_24942,N_24986);
and UO_657 (O_657,N_24890,N_24881);
and UO_658 (O_658,N_24996,N_24814);
nor UO_659 (O_659,N_24902,N_24845);
or UO_660 (O_660,N_24938,N_24847);
xnor UO_661 (O_661,N_24833,N_24921);
or UO_662 (O_662,N_24945,N_24920);
or UO_663 (O_663,N_24874,N_24847);
nor UO_664 (O_664,N_24873,N_24890);
and UO_665 (O_665,N_24969,N_24801);
and UO_666 (O_666,N_24928,N_24845);
and UO_667 (O_667,N_24837,N_24817);
nor UO_668 (O_668,N_24822,N_24969);
xnor UO_669 (O_669,N_24882,N_24942);
nor UO_670 (O_670,N_24849,N_24933);
nand UO_671 (O_671,N_24844,N_24898);
xnor UO_672 (O_672,N_24991,N_24870);
nand UO_673 (O_673,N_24894,N_24960);
and UO_674 (O_674,N_24948,N_24840);
nand UO_675 (O_675,N_24817,N_24874);
nor UO_676 (O_676,N_24816,N_24966);
or UO_677 (O_677,N_24879,N_24939);
xor UO_678 (O_678,N_24947,N_24834);
nor UO_679 (O_679,N_24964,N_24826);
xnor UO_680 (O_680,N_24992,N_24949);
nor UO_681 (O_681,N_24895,N_24845);
nand UO_682 (O_682,N_24955,N_24901);
xor UO_683 (O_683,N_24872,N_24999);
nor UO_684 (O_684,N_24930,N_24851);
and UO_685 (O_685,N_24913,N_24868);
or UO_686 (O_686,N_24979,N_24950);
nor UO_687 (O_687,N_24809,N_24952);
and UO_688 (O_688,N_24958,N_24830);
nor UO_689 (O_689,N_24917,N_24925);
xnor UO_690 (O_690,N_24817,N_24977);
nand UO_691 (O_691,N_24975,N_24970);
nor UO_692 (O_692,N_24891,N_24969);
or UO_693 (O_693,N_24891,N_24942);
and UO_694 (O_694,N_24914,N_24952);
xor UO_695 (O_695,N_24924,N_24888);
and UO_696 (O_696,N_24800,N_24991);
and UO_697 (O_697,N_24907,N_24910);
xor UO_698 (O_698,N_24841,N_24946);
and UO_699 (O_699,N_24813,N_24882);
and UO_700 (O_700,N_24818,N_24936);
nand UO_701 (O_701,N_24992,N_24903);
and UO_702 (O_702,N_24826,N_24835);
and UO_703 (O_703,N_24892,N_24884);
nor UO_704 (O_704,N_24931,N_24838);
and UO_705 (O_705,N_24979,N_24891);
and UO_706 (O_706,N_24844,N_24859);
or UO_707 (O_707,N_24948,N_24949);
nand UO_708 (O_708,N_24904,N_24869);
and UO_709 (O_709,N_24863,N_24805);
xnor UO_710 (O_710,N_24932,N_24879);
or UO_711 (O_711,N_24907,N_24931);
nor UO_712 (O_712,N_24830,N_24846);
nor UO_713 (O_713,N_24862,N_24948);
xnor UO_714 (O_714,N_24911,N_24841);
or UO_715 (O_715,N_24821,N_24917);
nor UO_716 (O_716,N_24833,N_24822);
or UO_717 (O_717,N_24805,N_24847);
nand UO_718 (O_718,N_24835,N_24886);
nor UO_719 (O_719,N_24864,N_24983);
or UO_720 (O_720,N_24893,N_24891);
nand UO_721 (O_721,N_24893,N_24993);
or UO_722 (O_722,N_24965,N_24908);
and UO_723 (O_723,N_24882,N_24983);
nor UO_724 (O_724,N_24871,N_24903);
nand UO_725 (O_725,N_24841,N_24807);
and UO_726 (O_726,N_24964,N_24833);
nor UO_727 (O_727,N_24957,N_24866);
or UO_728 (O_728,N_24825,N_24816);
and UO_729 (O_729,N_24915,N_24951);
or UO_730 (O_730,N_24984,N_24987);
nor UO_731 (O_731,N_24956,N_24992);
and UO_732 (O_732,N_24827,N_24807);
nand UO_733 (O_733,N_24904,N_24907);
xor UO_734 (O_734,N_24993,N_24858);
nor UO_735 (O_735,N_24880,N_24892);
or UO_736 (O_736,N_24906,N_24984);
xnor UO_737 (O_737,N_24995,N_24984);
and UO_738 (O_738,N_24980,N_24873);
or UO_739 (O_739,N_24810,N_24914);
nor UO_740 (O_740,N_24847,N_24990);
nor UO_741 (O_741,N_24866,N_24856);
nand UO_742 (O_742,N_24828,N_24940);
and UO_743 (O_743,N_24918,N_24839);
and UO_744 (O_744,N_24878,N_24999);
xor UO_745 (O_745,N_24954,N_24949);
nor UO_746 (O_746,N_24975,N_24902);
xor UO_747 (O_747,N_24852,N_24803);
nor UO_748 (O_748,N_24859,N_24930);
nand UO_749 (O_749,N_24855,N_24964);
nand UO_750 (O_750,N_24942,N_24878);
or UO_751 (O_751,N_24957,N_24949);
nor UO_752 (O_752,N_24885,N_24979);
and UO_753 (O_753,N_24937,N_24980);
and UO_754 (O_754,N_24891,N_24991);
nor UO_755 (O_755,N_24920,N_24934);
nand UO_756 (O_756,N_24930,N_24886);
or UO_757 (O_757,N_24939,N_24806);
or UO_758 (O_758,N_24943,N_24922);
and UO_759 (O_759,N_24822,N_24932);
xor UO_760 (O_760,N_24803,N_24982);
xor UO_761 (O_761,N_24932,N_24937);
xor UO_762 (O_762,N_24999,N_24866);
or UO_763 (O_763,N_24885,N_24933);
xor UO_764 (O_764,N_24969,N_24901);
nor UO_765 (O_765,N_24869,N_24850);
and UO_766 (O_766,N_24852,N_24820);
and UO_767 (O_767,N_24968,N_24962);
and UO_768 (O_768,N_24853,N_24905);
nand UO_769 (O_769,N_24829,N_24824);
nand UO_770 (O_770,N_24905,N_24839);
xor UO_771 (O_771,N_24813,N_24974);
xor UO_772 (O_772,N_24870,N_24968);
nor UO_773 (O_773,N_24948,N_24838);
xor UO_774 (O_774,N_24886,N_24805);
nand UO_775 (O_775,N_24974,N_24919);
nand UO_776 (O_776,N_24887,N_24899);
nand UO_777 (O_777,N_24867,N_24981);
nand UO_778 (O_778,N_24973,N_24873);
or UO_779 (O_779,N_24819,N_24963);
xor UO_780 (O_780,N_24807,N_24957);
nor UO_781 (O_781,N_24912,N_24810);
nand UO_782 (O_782,N_24992,N_24967);
nand UO_783 (O_783,N_24996,N_24962);
nor UO_784 (O_784,N_24818,N_24829);
nor UO_785 (O_785,N_24934,N_24846);
nor UO_786 (O_786,N_24962,N_24972);
xnor UO_787 (O_787,N_24856,N_24963);
nand UO_788 (O_788,N_24858,N_24953);
or UO_789 (O_789,N_24851,N_24996);
nand UO_790 (O_790,N_24816,N_24820);
xor UO_791 (O_791,N_24866,N_24839);
xor UO_792 (O_792,N_24842,N_24984);
nor UO_793 (O_793,N_24815,N_24875);
xor UO_794 (O_794,N_24980,N_24804);
nor UO_795 (O_795,N_24937,N_24905);
nor UO_796 (O_796,N_24872,N_24838);
nor UO_797 (O_797,N_24978,N_24853);
or UO_798 (O_798,N_24931,N_24977);
xor UO_799 (O_799,N_24837,N_24985);
nor UO_800 (O_800,N_24834,N_24879);
nand UO_801 (O_801,N_24959,N_24916);
xor UO_802 (O_802,N_24990,N_24939);
and UO_803 (O_803,N_24955,N_24851);
and UO_804 (O_804,N_24933,N_24963);
or UO_805 (O_805,N_24993,N_24901);
or UO_806 (O_806,N_24989,N_24960);
nand UO_807 (O_807,N_24834,N_24900);
nand UO_808 (O_808,N_24863,N_24844);
nor UO_809 (O_809,N_24883,N_24919);
and UO_810 (O_810,N_24826,N_24978);
nand UO_811 (O_811,N_24990,N_24873);
xnor UO_812 (O_812,N_24979,N_24892);
xnor UO_813 (O_813,N_24965,N_24889);
or UO_814 (O_814,N_24964,N_24880);
and UO_815 (O_815,N_24978,N_24941);
nand UO_816 (O_816,N_24928,N_24949);
and UO_817 (O_817,N_24902,N_24922);
nor UO_818 (O_818,N_24801,N_24932);
xnor UO_819 (O_819,N_24841,N_24877);
nand UO_820 (O_820,N_24864,N_24812);
nand UO_821 (O_821,N_24930,N_24991);
or UO_822 (O_822,N_24839,N_24837);
nand UO_823 (O_823,N_24905,N_24914);
and UO_824 (O_824,N_24885,N_24862);
or UO_825 (O_825,N_24977,N_24923);
and UO_826 (O_826,N_24853,N_24889);
nor UO_827 (O_827,N_24967,N_24932);
or UO_828 (O_828,N_24909,N_24843);
and UO_829 (O_829,N_24933,N_24801);
and UO_830 (O_830,N_24812,N_24920);
nand UO_831 (O_831,N_24990,N_24868);
and UO_832 (O_832,N_24878,N_24957);
nor UO_833 (O_833,N_24827,N_24800);
xnor UO_834 (O_834,N_24815,N_24813);
nor UO_835 (O_835,N_24874,N_24923);
and UO_836 (O_836,N_24905,N_24989);
xnor UO_837 (O_837,N_24930,N_24905);
nor UO_838 (O_838,N_24997,N_24977);
and UO_839 (O_839,N_24864,N_24914);
and UO_840 (O_840,N_24812,N_24926);
nand UO_841 (O_841,N_24901,N_24854);
and UO_842 (O_842,N_24851,N_24991);
xor UO_843 (O_843,N_24839,N_24803);
and UO_844 (O_844,N_24893,N_24898);
and UO_845 (O_845,N_24816,N_24915);
nor UO_846 (O_846,N_24895,N_24911);
nand UO_847 (O_847,N_24952,N_24996);
and UO_848 (O_848,N_24837,N_24943);
nor UO_849 (O_849,N_24863,N_24823);
or UO_850 (O_850,N_24988,N_24808);
xor UO_851 (O_851,N_24867,N_24874);
or UO_852 (O_852,N_24891,N_24850);
and UO_853 (O_853,N_24980,N_24964);
xnor UO_854 (O_854,N_24950,N_24879);
xnor UO_855 (O_855,N_24912,N_24988);
or UO_856 (O_856,N_24951,N_24860);
nand UO_857 (O_857,N_24944,N_24903);
nor UO_858 (O_858,N_24960,N_24809);
nand UO_859 (O_859,N_24862,N_24975);
nor UO_860 (O_860,N_24900,N_24943);
nand UO_861 (O_861,N_24998,N_24914);
nor UO_862 (O_862,N_24990,N_24974);
and UO_863 (O_863,N_24829,N_24966);
xnor UO_864 (O_864,N_24829,N_24993);
nand UO_865 (O_865,N_24967,N_24959);
or UO_866 (O_866,N_24911,N_24864);
and UO_867 (O_867,N_24992,N_24978);
xor UO_868 (O_868,N_24955,N_24840);
and UO_869 (O_869,N_24852,N_24907);
xnor UO_870 (O_870,N_24828,N_24962);
or UO_871 (O_871,N_24827,N_24988);
nor UO_872 (O_872,N_24949,N_24955);
xnor UO_873 (O_873,N_24906,N_24890);
nand UO_874 (O_874,N_24977,N_24836);
nor UO_875 (O_875,N_24828,N_24931);
xnor UO_876 (O_876,N_24857,N_24992);
and UO_877 (O_877,N_24889,N_24993);
and UO_878 (O_878,N_24807,N_24821);
xor UO_879 (O_879,N_24871,N_24931);
nand UO_880 (O_880,N_24930,N_24970);
nor UO_881 (O_881,N_24983,N_24904);
nand UO_882 (O_882,N_24825,N_24922);
nor UO_883 (O_883,N_24844,N_24816);
nand UO_884 (O_884,N_24925,N_24896);
nor UO_885 (O_885,N_24931,N_24822);
and UO_886 (O_886,N_24876,N_24977);
nor UO_887 (O_887,N_24829,N_24983);
nand UO_888 (O_888,N_24934,N_24981);
and UO_889 (O_889,N_24929,N_24860);
or UO_890 (O_890,N_24979,N_24834);
or UO_891 (O_891,N_24925,N_24869);
nand UO_892 (O_892,N_24828,N_24862);
xnor UO_893 (O_893,N_24844,N_24886);
and UO_894 (O_894,N_24852,N_24914);
nor UO_895 (O_895,N_24805,N_24855);
nand UO_896 (O_896,N_24986,N_24835);
and UO_897 (O_897,N_24883,N_24880);
nor UO_898 (O_898,N_24894,N_24810);
nand UO_899 (O_899,N_24918,N_24982);
nor UO_900 (O_900,N_24877,N_24969);
xnor UO_901 (O_901,N_24803,N_24874);
nand UO_902 (O_902,N_24876,N_24822);
xor UO_903 (O_903,N_24956,N_24970);
nor UO_904 (O_904,N_24874,N_24931);
and UO_905 (O_905,N_24911,N_24897);
or UO_906 (O_906,N_24992,N_24807);
and UO_907 (O_907,N_24965,N_24950);
nor UO_908 (O_908,N_24830,N_24832);
nor UO_909 (O_909,N_24801,N_24836);
nor UO_910 (O_910,N_24976,N_24867);
and UO_911 (O_911,N_24909,N_24877);
and UO_912 (O_912,N_24921,N_24801);
and UO_913 (O_913,N_24866,N_24972);
nor UO_914 (O_914,N_24808,N_24996);
xnor UO_915 (O_915,N_24970,N_24839);
and UO_916 (O_916,N_24833,N_24865);
or UO_917 (O_917,N_24915,N_24866);
and UO_918 (O_918,N_24897,N_24856);
xnor UO_919 (O_919,N_24870,N_24909);
xnor UO_920 (O_920,N_24906,N_24842);
nand UO_921 (O_921,N_24983,N_24945);
nor UO_922 (O_922,N_24986,N_24838);
or UO_923 (O_923,N_24913,N_24885);
and UO_924 (O_924,N_24948,N_24810);
and UO_925 (O_925,N_24810,N_24827);
xor UO_926 (O_926,N_24950,N_24900);
xor UO_927 (O_927,N_24949,N_24993);
xor UO_928 (O_928,N_24880,N_24891);
nand UO_929 (O_929,N_24818,N_24804);
nand UO_930 (O_930,N_24942,N_24880);
and UO_931 (O_931,N_24989,N_24965);
nor UO_932 (O_932,N_24980,N_24955);
xor UO_933 (O_933,N_24932,N_24813);
nor UO_934 (O_934,N_24842,N_24882);
or UO_935 (O_935,N_24991,N_24970);
xor UO_936 (O_936,N_24857,N_24873);
and UO_937 (O_937,N_24893,N_24907);
nand UO_938 (O_938,N_24851,N_24832);
or UO_939 (O_939,N_24943,N_24836);
xnor UO_940 (O_940,N_24919,N_24866);
or UO_941 (O_941,N_24948,N_24857);
and UO_942 (O_942,N_24951,N_24839);
nor UO_943 (O_943,N_24957,N_24906);
or UO_944 (O_944,N_24827,N_24977);
xor UO_945 (O_945,N_24898,N_24911);
nand UO_946 (O_946,N_24866,N_24816);
nand UO_947 (O_947,N_24883,N_24928);
nand UO_948 (O_948,N_24942,N_24822);
nand UO_949 (O_949,N_24862,N_24943);
nor UO_950 (O_950,N_24950,N_24987);
xnor UO_951 (O_951,N_24942,N_24866);
nor UO_952 (O_952,N_24918,N_24898);
xor UO_953 (O_953,N_24858,N_24990);
and UO_954 (O_954,N_24841,N_24943);
nor UO_955 (O_955,N_24829,N_24946);
or UO_956 (O_956,N_24844,N_24991);
and UO_957 (O_957,N_24813,N_24942);
or UO_958 (O_958,N_24942,N_24846);
or UO_959 (O_959,N_24890,N_24919);
or UO_960 (O_960,N_24896,N_24984);
and UO_961 (O_961,N_24829,N_24977);
nand UO_962 (O_962,N_24866,N_24985);
and UO_963 (O_963,N_24868,N_24993);
nor UO_964 (O_964,N_24889,N_24948);
nor UO_965 (O_965,N_24992,N_24913);
xnor UO_966 (O_966,N_24949,N_24904);
or UO_967 (O_967,N_24848,N_24948);
xnor UO_968 (O_968,N_24804,N_24938);
nand UO_969 (O_969,N_24948,N_24911);
nor UO_970 (O_970,N_24850,N_24848);
xnor UO_971 (O_971,N_24956,N_24962);
xor UO_972 (O_972,N_24832,N_24927);
nor UO_973 (O_973,N_24997,N_24869);
xnor UO_974 (O_974,N_24910,N_24867);
nand UO_975 (O_975,N_24873,N_24856);
and UO_976 (O_976,N_24803,N_24846);
nor UO_977 (O_977,N_24971,N_24947);
and UO_978 (O_978,N_24913,N_24826);
xnor UO_979 (O_979,N_24927,N_24926);
and UO_980 (O_980,N_24890,N_24843);
nand UO_981 (O_981,N_24823,N_24826);
or UO_982 (O_982,N_24955,N_24952);
xor UO_983 (O_983,N_24950,N_24892);
xor UO_984 (O_984,N_24901,N_24948);
and UO_985 (O_985,N_24993,N_24854);
nor UO_986 (O_986,N_24944,N_24947);
and UO_987 (O_987,N_24850,N_24943);
nor UO_988 (O_988,N_24929,N_24870);
xor UO_989 (O_989,N_24960,N_24956);
nand UO_990 (O_990,N_24950,N_24840);
and UO_991 (O_991,N_24862,N_24837);
and UO_992 (O_992,N_24845,N_24800);
xor UO_993 (O_993,N_24835,N_24943);
nand UO_994 (O_994,N_24860,N_24866);
or UO_995 (O_995,N_24810,N_24847);
nand UO_996 (O_996,N_24812,N_24903);
nor UO_997 (O_997,N_24845,N_24942);
xnor UO_998 (O_998,N_24969,N_24807);
or UO_999 (O_999,N_24922,N_24915);
xor UO_1000 (O_1000,N_24890,N_24841);
nand UO_1001 (O_1001,N_24874,N_24961);
and UO_1002 (O_1002,N_24870,N_24837);
and UO_1003 (O_1003,N_24848,N_24855);
xnor UO_1004 (O_1004,N_24879,N_24997);
xnor UO_1005 (O_1005,N_24973,N_24956);
nand UO_1006 (O_1006,N_24959,N_24839);
nor UO_1007 (O_1007,N_24935,N_24898);
and UO_1008 (O_1008,N_24823,N_24993);
or UO_1009 (O_1009,N_24929,N_24965);
and UO_1010 (O_1010,N_24956,N_24948);
or UO_1011 (O_1011,N_24939,N_24873);
xor UO_1012 (O_1012,N_24816,N_24804);
or UO_1013 (O_1013,N_24855,N_24918);
and UO_1014 (O_1014,N_24810,N_24886);
or UO_1015 (O_1015,N_24801,N_24910);
xnor UO_1016 (O_1016,N_24826,N_24872);
nor UO_1017 (O_1017,N_24850,N_24815);
and UO_1018 (O_1018,N_24829,N_24942);
xnor UO_1019 (O_1019,N_24954,N_24995);
nand UO_1020 (O_1020,N_24871,N_24873);
nor UO_1021 (O_1021,N_24843,N_24855);
and UO_1022 (O_1022,N_24833,N_24943);
and UO_1023 (O_1023,N_24811,N_24897);
and UO_1024 (O_1024,N_24867,N_24965);
and UO_1025 (O_1025,N_24998,N_24821);
nor UO_1026 (O_1026,N_24864,N_24954);
nand UO_1027 (O_1027,N_24863,N_24819);
and UO_1028 (O_1028,N_24855,N_24932);
nand UO_1029 (O_1029,N_24854,N_24880);
and UO_1030 (O_1030,N_24892,N_24867);
and UO_1031 (O_1031,N_24874,N_24940);
xnor UO_1032 (O_1032,N_24961,N_24890);
or UO_1033 (O_1033,N_24969,N_24874);
nand UO_1034 (O_1034,N_24801,N_24956);
and UO_1035 (O_1035,N_24904,N_24946);
and UO_1036 (O_1036,N_24904,N_24874);
or UO_1037 (O_1037,N_24801,N_24963);
or UO_1038 (O_1038,N_24804,N_24914);
xor UO_1039 (O_1039,N_24858,N_24801);
nor UO_1040 (O_1040,N_24949,N_24997);
nand UO_1041 (O_1041,N_24805,N_24902);
nand UO_1042 (O_1042,N_24996,N_24959);
and UO_1043 (O_1043,N_24980,N_24838);
and UO_1044 (O_1044,N_24963,N_24845);
or UO_1045 (O_1045,N_24983,N_24810);
xnor UO_1046 (O_1046,N_24815,N_24857);
nor UO_1047 (O_1047,N_24804,N_24922);
nor UO_1048 (O_1048,N_24833,N_24937);
and UO_1049 (O_1049,N_24955,N_24913);
nor UO_1050 (O_1050,N_24815,N_24934);
nand UO_1051 (O_1051,N_24813,N_24834);
nor UO_1052 (O_1052,N_24815,N_24832);
or UO_1053 (O_1053,N_24952,N_24804);
xor UO_1054 (O_1054,N_24907,N_24900);
xor UO_1055 (O_1055,N_24828,N_24998);
nor UO_1056 (O_1056,N_24890,N_24972);
and UO_1057 (O_1057,N_24843,N_24889);
or UO_1058 (O_1058,N_24958,N_24913);
nand UO_1059 (O_1059,N_24870,N_24943);
nor UO_1060 (O_1060,N_24806,N_24990);
or UO_1061 (O_1061,N_24881,N_24811);
or UO_1062 (O_1062,N_24835,N_24805);
or UO_1063 (O_1063,N_24836,N_24824);
nand UO_1064 (O_1064,N_24847,N_24906);
nand UO_1065 (O_1065,N_24800,N_24942);
and UO_1066 (O_1066,N_24854,N_24919);
and UO_1067 (O_1067,N_24912,N_24827);
nor UO_1068 (O_1068,N_24996,N_24836);
nor UO_1069 (O_1069,N_24913,N_24875);
and UO_1070 (O_1070,N_24822,N_24834);
xor UO_1071 (O_1071,N_24849,N_24923);
nor UO_1072 (O_1072,N_24875,N_24928);
nor UO_1073 (O_1073,N_24977,N_24848);
nor UO_1074 (O_1074,N_24967,N_24978);
or UO_1075 (O_1075,N_24905,N_24901);
nand UO_1076 (O_1076,N_24830,N_24992);
nand UO_1077 (O_1077,N_24908,N_24821);
nor UO_1078 (O_1078,N_24858,N_24851);
nand UO_1079 (O_1079,N_24958,N_24943);
or UO_1080 (O_1080,N_24949,N_24837);
and UO_1081 (O_1081,N_24906,N_24836);
nor UO_1082 (O_1082,N_24916,N_24862);
nand UO_1083 (O_1083,N_24994,N_24802);
and UO_1084 (O_1084,N_24907,N_24800);
nor UO_1085 (O_1085,N_24845,N_24949);
nand UO_1086 (O_1086,N_24807,N_24981);
or UO_1087 (O_1087,N_24819,N_24981);
and UO_1088 (O_1088,N_24956,N_24929);
xor UO_1089 (O_1089,N_24841,N_24980);
nor UO_1090 (O_1090,N_24838,N_24892);
xnor UO_1091 (O_1091,N_24930,N_24836);
nor UO_1092 (O_1092,N_24925,N_24993);
and UO_1093 (O_1093,N_24970,N_24946);
and UO_1094 (O_1094,N_24993,N_24899);
nor UO_1095 (O_1095,N_24998,N_24889);
nand UO_1096 (O_1096,N_24910,N_24938);
nor UO_1097 (O_1097,N_24964,N_24977);
nor UO_1098 (O_1098,N_24985,N_24912);
and UO_1099 (O_1099,N_24983,N_24920);
nor UO_1100 (O_1100,N_24973,N_24979);
xnor UO_1101 (O_1101,N_24804,N_24848);
nor UO_1102 (O_1102,N_24849,N_24859);
xnor UO_1103 (O_1103,N_24843,N_24990);
and UO_1104 (O_1104,N_24991,N_24843);
nor UO_1105 (O_1105,N_24937,N_24969);
and UO_1106 (O_1106,N_24958,N_24951);
or UO_1107 (O_1107,N_24825,N_24812);
or UO_1108 (O_1108,N_24902,N_24905);
nand UO_1109 (O_1109,N_24877,N_24942);
nand UO_1110 (O_1110,N_24961,N_24951);
nor UO_1111 (O_1111,N_24810,N_24817);
or UO_1112 (O_1112,N_24908,N_24822);
nor UO_1113 (O_1113,N_24943,N_24984);
nand UO_1114 (O_1114,N_24877,N_24809);
or UO_1115 (O_1115,N_24906,N_24944);
nand UO_1116 (O_1116,N_24808,N_24904);
nor UO_1117 (O_1117,N_24822,N_24873);
and UO_1118 (O_1118,N_24880,N_24958);
xor UO_1119 (O_1119,N_24873,N_24968);
nor UO_1120 (O_1120,N_24900,N_24851);
nor UO_1121 (O_1121,N_24915,N_24898);
and UO_1122 (O_1122,N_24820,N_24971);
xor UO_1123 (O_1123,N_24979,N_24872);
xor UO_1124 (O_1124,N_24867,N_24961);
nand UO_1125 (O_1125,N_24909,N_24997);
nand UO_1126 (O_1126,N_24807,N_24843);
or UO_1127 (O_1127,N_24926,N_24997);
and UO_1128 (O_1128,N_24894,N_24897);
and UO_1129 (O_1129,N_24903,N_24897);
or UO_1130 (O_1130,N_24862,N_24891);
nor UO_1131 (O_1131,N_24953,N_24825);
nand UO_1132 (O_1132,N_24907,N_24866);
nand UO_1133 (O_1133,N_24865,N_24994);
xnor UO_1134 (O_1134,N_24815,N_24819);
or UO_1135 (O_1135,N_24980,N_24970);
and UO_1136 (O_1136,N_24968,N_24955);
xor UO_1137 (O_1137,N_24800,N_24930);
nand UO_1138 (O_1138,N_24933,N_24922);
nand UO_1139 (O_1139,N_24800,N_24878);
nor UO_1140 (O_1140,N_24804,N_24941);
nand UO_1141 (O_1141,N_24898,N_24872);
nor UO_1142 (O_1142,N_24910,N_24947);
nand UO_1143 (O_1143,N_24819,N_24807);
or UO_1144 (O_1144,N_24881,N_24876);
or UO_1145 (O_1145,N_24841,N_24884);
xnor UO_1146 (O_1146,N_24989,N_24889);
and UO_1147 (O_1147,N_24879,N_24927);
or UO_1148 (O_1148,N_24873,N_24863);
xnor UO_1149 (O_1149,N_24905,N_24973);
nand UO_1150 (O_1150,N_24873,N_24909);
nor UO_1151 (O_1151,N_24812,N_24897);
and UO_1152 (O_1152,N_24882,N_24932);
nand UO_1153 (O_1153,N_24984,N_24839);
or UO_1154 (O_1154,N_24862,N_24811);
nand UO_1155 (O_1155,N_24812,N_24883);
nand UO_1156 (O_1156,N_24926,N_24911);
or UO_1157 (O_1157,N_24931,N_24972);
and UO_1158 (O_1158,N_24802,N_24902);
and UO_1159 (O_1159,N_24937,N_24862);
nor UO_1160 (O_1160,N_24874,N_24912);
nor UO_1161 (O_1161,N_24869,N_24889);
or UO_1162 (O_1162,N_24846,N_24821);
or UO_1163 (O_1163,N_24853,N_24849);
nand UO_1164 (O_1164,N_24920,N_24834);
xor UO_1165 (O_1165,N_24879,N_24949);
or UO_1166 (O_1166,N_24814,N_24995);
xnor UO_1167 (O_1167,N_24893,N_24856);
nand UO_1168 (O_1168,N_24918,N_24893);
nor UO_1169 (O_1169,N_24993,N_24851);
and UO_1170 (O_1170,N_24936,N_24946);
or UO_1171 (O_1171,N_24851,N_24882);
nand UO_1172 (O_1172,N_24821,N_24950);
or UO_1173 (O_1173,N_24828,N_24843);
xnor UO_1174 (O_1174,N_24970,N_24898);
and UO_1175 (O_1175,N_24879,N_24896);
xor UO_1176 (O_1176,N_24849,N_24851);
nor UO_1177 (O_1177,N_24925,N_24994);
xor UO_1178 (O_1178,N_24892,N_24987);
nand UO_1179 (O_1179,N_24801,N_24813);
and UO_1180 (O_1180,N_24905,N_24868);
and UO_1181 (O_1181,N_24940,N_24867);
and UO_1182 (O_1182,N_24905,N_24835);
nand UO_1183 (O_1183,N_24850,N_24924);
and UO_1184 (O_1184,N_24941,N_24895);
xor UO_1185 (O_1185,N_24972,N_24968);
xnor UO_1186 (O_1186,N_24880,N_24879);
or UO_1187 (O_1187,N_24824,N_24904);
nor UO_1188 (O_1188,N_24880,N_24817);
nand UO_1189 (O_1189,N_24924,N_24897);
nand UO_1190 (O_1190,N_24938,N_24962);
and UO_1191 (O_1191,N_24809,N_24825);
xor UO_1192 (O_1192,N_24861,N_24940);
nand UO_1193 (O_1193,N_24949,N_24963);
nor UO_1194 (O_1194,N_24903,N_24849);
or UO_1195 (O_1195,N_24820,N_24817);
nor UO_1196 (O_1196,N_24840,N_24866);
or UO_1197 (O_1197,N_24985,N_24841);
and UO_1198 (O_1198,N_24888,N_24816);
nand UO_1199 (O_1199,N_24901,N_24870);
and UO_1200 (O_1200,N_24866,N_24929);
and UO_1201 (O_1201,N_24849,N_24982);
nand UO_1202 (O_1202,N_24937,N_24830);
nor UO_1203 (O_1203,N_24959,N_24807);
or UO_1204 (O_1204,N_24879,N_24820);
and UO_1205 (O_1205,N_24818,N_24809);
xnor UO_1206 (O_1206,N_24887,N_24978);
nor UO_1207 (O_1207,N_24966,N_24884);
xnor UO_1208 (O_1208,N_24979,N_24986);
or UO_1209 (O_1209,N_24832,N_24977);
nor UO_1210 (O_1210,N_24847,N_24916);
xor UO_1211 (O_1211,N_24871,N_24896);
nand UO_1212 (O_1212,N_24889,N_24929);
and UO_1213 (O_1213,N_24836,N_24942);
xnor UO_1214 (O_1214,N_24852,N_24915);
and UO_1215 (O_1215,N_24829,N_24921);
and UO_1216 (O_1216,N_24904,N_24934);
and UO_1217 (O_1217,N_24818,N_24967);
or UO_1218 (O_1218,N_24884,N_24912);
xnor UO_1219 (O_1219,N_24865,N_24989);
and UO_1220 (O_1220,N_24871,N_24994);
xor UO_1221 (O_1221,N_24873,N_24833);
and UO_1222 (O_1222,N_24886,N_24897);
and UO_1223 (O_1223,N_24830,N_24997);
or UO_1224 (O_1224,N_24953,N_24874);
and UO_1225 (O_1225,N_24923,N_24964);
and UO_1226 (O_1226,N_24928,N_24972);
xnor UO_1227 (O_1227,N_24967,N_24908);
nor UO_1228 (O_1228,N_24983,N_24975);
or UO_1229 (O_1229,N_24933,N_24839);
xor UO_1230 (O_1230,N_24933,N_24904);
xor UO_1231 (O_1231,N_24861,N_24872);
or UO_1232 (O_1232,N_24914,N_24892);
or UO_1233 (O_1233,N_24822,N_24963);
nand UO_1234 (O_1234,N_24836,N_24948);
nand UO_1235 (O_1235,N_24975,N_24957);
xnor UO_1236 (O_1236,N_24843,N_24952);
nor UO_1237 (O_1237,N_24947,N_24803);
nand UO_1238 (O_1238,N_24977,N_24944);
nand UO_1239 (O_1239,N_24936,N_24970);
xor UO_1240 (O_1240,N_24867,N_24977);
nor UO_1241 (O_1241,N_24974,N_24814);
and UO_1242 (O_1242,N_24870,N_24823);
nand UO_1243 (O_1243,N_24828,N_24810);
xnor UO_1244 (O_1244,N_24842,N_24925);
or UO_1245 (O_1245,N_24949,N_24966);
or UO_1246 (O_1246,N_24958,N_24850);
nor UO_1247 (O_1247,N_24820,N_24933);
xor UO_1248 (O_1248,N_24987,N_24865);
or UO_1249 (O_1249,N_24978,N_24828);
nor UO_1250 (O_1250,N_24917,N_24840);
xor UO_1251 (O_1251,N_24800,N_24953);
nor UO_1252 (O_1252,N_24876,N_24848);
and UO_1253 (O_1253,N_24964,N_24931);
nand UO_1254 (O_1254,N_24915,N_24937);
nor UO_1255 (O_1255,N_24941,N_24959);
and UO_1256 (O_1256,N_24965,N_24870);
nand UO_1257 (O_1257,N_24808,N_24865);
nand UO_1258 (O_1258,N_24931,N_24891);
nor UO_1259 (O_1259,N_24901,N_24857);
xor UO_1260 (O_1260,N_24972,N_24933);
xor UO_1261 (O_1261,N_24839,N_24890);
xor UO_1262 (O_1262,N_24864,N_24891);
and UO_1263 (O_1263,N_24856,N_24950);
or UO_1264 (O_1264,N_24923,N_24856);
xor UO_1265 (O_1265,N_24965,N_24901);
xor UO_1266 (O_1266,N_24807,N_24859);
or UO_1267 (O_1267,N_24808,N_24908);
nand UO_1268 (O_1268,N_24975,N_24810);
xor UO_1269 (O_1269,N_24837,N_24916);
xor UO_1270 (O_1270,N_24853,N_24855);
or UO_1271 (O_1271,N_24857,N_24919);
or UO_1272 (O_1272,N_24931,N_24915);
and UO_1273 (O_1273,N_24959,N_24946);
nor UO_1274 (O_1274,N_24970,N_24972);
or UO_1275 (O_1275,N_24831,N_24911);
or UO_1276 (O_1276,N_24865,N_24920);
xnor UO_1277 (O_1277,N_24897,N_24872);
or UO_1278 (O_1278,N_24822,N_24898);
xnor UO_1279 (O_1279,N_24924,N_24867);
or UO_1280 (O_1280,N_24814,N_24927);
or UO_1281 (O_1281,N_24935,N_24901);
or UO_1282 (O_1282,N_24862,N_24861);
nor UO_1283 (O_1283,N_24929,N_24810);
and UO_1284 (O_1284,N_24931,N_24916);
or UO_1285 (O_1285,N_24850,N_24836);
xnor UO_1286 (O_1286,N_24985,N_24920);
nand UO_1287 (O_1287,N_24921,N_24865);
nor UO_1288 (O_1288,N_24987,N_24852);
nor UO_1289 (O_1289,N_24898,N_24815);
xnor UO_1290 (O_1290,N_24921,N_24869);
xor UO_1291 (O_1291,N_24967,N_24984);
nor UO_1292 (O_1292,N_24836,N_24940);
xor UO_1293 (O_1293,N_24813,N_24886);
and UO_1294 (O_1294,N_24874,N_24956);
nor UO_1295 (O_1295,N_24807,N_24850);
and UO_1296 (O_1296,N_24969,N_24808);
nor UO_1297 (O_1297,N_24828,N_24944);
xnor UO_1298 (O_1298,N_24933,N_24921);
or UO_1299 (O_1299,N_24991,N_24815);
or UO_1300 (O_1300,N_24929,N_24801);
and UO_1301 (O_1301,N_24839,N_24938);
and UO_1302 (O_1302,N_24832,N_24823);
and UO_1303 (O_1303,N_24991,N_24941);
xor UO_1304 (O_1304,N_24854,N_24926);
or UO_1305 (O_1305,N_24802,N_24975);
nand UO_1306 (O_1306,N_24939,N_24962);
and UO_1307 (O_1307,N_24924,N_24899);
or UO_1308 (O_1308,N_24957,N_24886);
nor UO_1309 (O_1309,N_24810,N_24989);
xor UO_1310 (O_1310,N_24802,N_24917);
xor UO_1311 (O_1311,N_24972,N_24899);
nand UO_1312 (O_1312,N_24869,N_24903);
nand UO_1313 (O_1313,N_24802,N_24817);
or UO_1314 (O_1314,N_24968,N_24961);
xnor UO_1315 (O_1315,N_24940,N_24948);
nand UO_1316 (O_1316,N_24861,N_24852);
xnor UO_1317 (O_1317,N_24820,N_24862);
xor UO_1318 (O_1318,N_24889,N_24824);
and UO_1319 (O_1319,N_24871,N_24843);
and UO_1320 (O_1320,N_24904,N_24850);
xor UO_1321 (O_1321,N_24944,N_24989);
and UO_1322 (O_1322,N_24895,N_24829);
or UO_1323 (O_1323,N_24922,N_24857);
nor UO_1324 (O_1324,N_24859,N_24888);
nand UO_1325 (O_1325,N_24961,N_24855);
or UO_1326 (O_1326,N_24849,N_24854);
or UO_1327 (O_1327,N_24901,N_24898);
and UO_1328 (O_1328,N_24850,N_24849);
nor UO_1329 (O_1329,N_24949,N_24812);
nor UO_1330 (O_1330,N_24979,N_24994);
or UO_1331 (O_1331,N_24973,N_24877);
and UO_1332 (O_1332,N_24966,N_24859);
or UO_1333 (O_1333,N_24803,N_24901);
or UO_1334 (O_1334,N_24945,N_24897);
nor UO_1335 (O_1335,N_24868,N_24927);
nand UO_1336 (O_1336,N_24854,N_24879);
and UO_1337 (O_1337,N_24823,N_24960);
nor UO_1338 (O_1338,N_24875,N_24812);
nand UO_1339 (O_1339,N_24954,N_24836);
xor UO_1340 (O_1340,N_24993,N_24977);
nand UO_1341 (O_1341,N_24901,N_24866);
nand UO_1342 (O_1342,N_24902,N_24949);
nor UO_1343 (O_1343,N_24834,N_24811);
xnor UO_1344 (O_1344,N_24806,N_24809);
and UO_1345 (O_1345,N_24868,N_24875);
xnor UO_1346 (O_1346,N_24932,N_24827);
and UO_1347 (O_1347,N_24979,N_24875);
xor UO_1348 (O_1348,N_24847,N_24909);
nor UO_1349 (O_1349,N_24839,N_24869);
or UO_1350 (O_1350,N_24895,N_24855);
nand UO_1351 (O_1351,N_24969,N_24945);
xor UO_1352 (O_1352,N_24805,N_24949);
and UO_1353 (O_1353,N_24819,N_24910);
or UO_1354 (O_1354,N_24942,N_24827);
and UO_1355 (O_1355,N_24871,N_24992);
nand UO_1356 (O_1356,N_24936,N_24869);
xor UO_1357 (O_1357,N_24866,N_24869);
or UO_1358 (O_1358,N_24992,N_24972);
nand UO_1359 (O_1359,N_24888,N_24975);
nand UO_1360 (O_1360,N_24925,N_24919);
nand UO_1361 (O_1361,N_24867,N_24861);
nor UO_1362 (O_1362,N_24804,N_24925);
nand UO_1363 (O_1363,N_24827,N_24936);
nor UO_1364 (O_1364,N_24936,N_24990);
nand UO_1365 (O_1365,N_24958,N_24890);
nand UO_1366 (O_1366,N_24821,N_24961);
nand UO_1367 (O_1367,N_24994,N_24901);
or UO_1368 (O_1368,N_24925,N_24874);
nand UO_1369 (O_1369,N_24949,N_24914);
or UO_1370 (O_1370,N_24896,N_24952);
xor UO_1371 (O_1371,N_24885,N_24997);
nand UO_1372 (O_1372,N_24837,N_24979);
nand UO_1373 (O_1373,N_24903,N_24863);
or UO_1374 (O_1374,N_24853,N_24932);
nor UO_1375 (O_1375,N_24822,N_24832);
xnor UO_1376 (O_1376,N_24954,N_24966);
and UO_1377 (O_1377,N_24863,N_24839);
and UO_1378 (O_1378,N_24932,N_24841);
and UO_1379 (O_1379,N_24875,N_24814);
xnor UO_1380 (O_1380,N_24840,N_24890);
nor UO_1381 (O_1381,N_24942,N_24968);
nor UO_1382 (O_1382,N_24814,N_24952);
nand UO_1383 (O_1383,N_24809,N_24865);
and UO_1384 (O_1384,N_24981,N_24915);
xnor UO_1385 (O_1385,N_24915,N_24818);
or UO_1386 (O_1386,N_24923,N_24906);
nand UO_1387 (O_1387,N_24927,N_24972);
nor UO_1388 (O_1388,N_24885,N_24819);
xor UO_1389 (O_1389,N_24890,N_24851);
and UO_1390 (O_1390,N_24860,N_24961);
nand UO_1391 (O_1391,N_24979,N_24940);
nand UO_1392 (O_1392,N_24864,N_24887);
and UO_1393 (O_1393,N_24973,N_24832);
xor UO_1394 (O_1394,N_24915,N_24812);
or UO_1395 (O_1395,N_24922,N_24994);
xor UO_1396 (O_1396,N_24979,N_24978);
xor UO_1397 (O_1397,N_24812,N_24858);
nand UO_1398 (O_1398,N_24813,N_24916);
nor UO_1399 (O_1399,N_24964,N_24890);
or UO_1400 (O_1400,N_24936,N_24905);
nor UO_1401 (O_1401,N_24833,N_24805);
nand UO_1402 (O_1402,N_24910,N_24832);
or UO_1403 (O_1403,N_24827,N_24963);
nand UO_1404 (O_1404,N_24905,N_24915);
xor UO_1405 (O_1405,N_24804,N_24858);
or UO_1406 (O_1406,N_24803,N_24956);
and UO_1407 (O_1407,N_24957,N_24935);
nand UO_1408 (O_1408,N_24981,N_24890);
or UO_1409 (O_1409,N_24949,N_24882);
xnor UO_1410 (O_1410,N_24947,N_24890);
or UO_1411 (O_1411,N_24827,N_24840);
nor UO_1412 (O_1412,N_24803,N_24853);
or UO_1413 (O_1413,N_24808,N_24926);
xor UO_1414 (O_1414,N_24843,N_24939);
xnor UO_1415 (O_1415,N_24986,N_24848);
or UO_1416 (O_1416,N_24825,N_24868);
or UO_1417 (O_1417,N_24924,N_24975);
xor UO_1418 (O_1418,N_24978,N_24922);
and UO_1419 (O_1419,N_24950,N_24889);
nand UO_1420 (O_1420,N_24931,N_24963);
nor UO_1421 (O_1421,N_24807,N_24857);
nor UO_1422 (O_1422,N_24805,N_24827);
nand UO_1423 (O_1423,N_24909,N_24939);
or UO_1424 (O_1424,N_24925,N_24985);
and UO_1425 (O_1425,N_24961,N_24815);
nor UO_1426 (O_1426,N_24907,N_24918);
nor UO_1427 (O_1427,N_24923,N_24817);
or UO_1428 (O_1428,N_24959,N_24934);
and UO_1429 (O_1429,N_24839,N_24820);
or UO_1430 (O_1430,N_24972,N_24865);
or UO_1431 (O_1431,N_24849,N_24843);
nor UO_1432 (O_1432,N_24924,N_24991);
xor UO_1433 (O_1433,N_24949,N_24885);
or UO_1434 (O_1434,N_24803,N_24957);
nor UO_1435 (O_1435,N_24996,N_24914);
nand UO_1436 (O_1436,N_24983,N_24970);
or UO_1437 (O_1437,N_24937,N_24909);
nor UO_1438 (O_1438,N_24876,N_24945);
or UO_1439 (O_1439,N_24911,N_24890);
nor UO_1440 (O_1440,N_24962,N_24852);
or UO_1441 (O_1441,N_24974,N_24893);
nor UO_1442 (O_1442,N_24966,N_24844);
nor UO_1443 (O_1443,N_24980,N_24907);
or UO_1444 (O_1444,N_24835,N_24985);
nor UO_1445 (O_1445,N_24830,N_24807);
nor UO_1446 (O_1446,N_24954,N_24911);
and UO_1447 (O_1447,N_24941,N_24858);
nor UO_1448 (O_1448,N_24898,N_24892);
xnor UO_1449 (O_1449,N_24956,N_24897);
nand UO_1450 (O_1450,N_24868,N_24949);
nor UO_1451 (O_1451,N_24961,N_24875);
and UO_1452 (O_1452,N_24877,N_24961);
nand UO_1453 (O_1453,N_24909,N_24832);
and UO_1454 (O_1454,N_24961,N_24856);
xor UO_1455 (O_1455,N_24878,N_24839);
or UO_1456 (O_1456,N_24999,N_24877);
and UO_1457 (O_1457,N_24811,N_24808);
or UO_1458 (O_1458,N_24997,N_24938);
xor UO_1459 (O_1459,N_24862,N_24880);
or UO_1460 (O_1460,N_24809,N_24834);
nor UO_1461 (O_1461,N_24924,N_24898);
nor UO_1462 (O_1462,N_24872,N_24810);
nand UO_1463 (O_1463,N_24932,N_24842);
nor UO_1464 (O_1464,N_24945,N_24976);
or UO_1465 (O_1465,N_24852,N_24997);
or UO_1466 (O_1466,N_24947,N_24963);
nand UO_1467 (O_1467,N_24890,N_24922);
and UO_1468 (O_1468,N_24826,N_24981);
and UO_1469 (O_1469,N_24842,N_24941);
and UO_1470 (O_1470,N_24932,N_24812);
nor UO_1471 (O_1471,N_24960,N_24817);
or UO_1472 (O_1472,N_24821,N_24986);
nand UO_1473 (O_1473,N_24995,N_24864);
and UO_1474 (O_1474,N_24816,N_24821);
or UO_1475 (O_1475,N_24830,N_24934);
xnor UO_1476 (O_1476,N_24867,N_24823);
nor UO_1477 (O_1477,N_24876,N_24823);
nor UO_1478 (O_1478,N_24845,N_24878);
or UO_1479 (O_1479,N_24985,N_24980);
and UO_1480 (O_1480,N_24927,N_24928);
nand UO_1481 (O_1481,N_24950,N_24937);
nand UO_1482 (O_1482,N_24958,N_24920);
xnor UO_1483 (O_1483,N_24977,N_24890);
and UO_1484 (O_1484,N_24993,N_24890);
nor UO_1485 (O_1485,N_24997,N_24847);
and UO_1486 (O_1486,N_24807,N_24853);
xor UO_1487 (O_1487,N_24996,N_24827);
nand UO_1488 (O_1488,N_24835,N_24987);
or UO_1489 (O_1489,N_24881,N_24950);
and UO_1490 (O_1490,N_24982,N_24896);
or UO_1491 (O_1491,N_24977,N_24903);
nand UO_1492 (O_1492,N_24974,N_24985);
or UO_1493 (O_1493,N_24807,N_24812);
nand UO_1494 (O_1494,N_24964,N_24908);
or UO_1495 (O_1495,N_24832,N_24890);
or UO_1496 (O_1496,N_24830,N_24917);
nand UO_1497 (O_1497,N_24919,N_24807);
or UO_1498 (O_1498,N_24900,N_24859);
nand UO_1499 (O_1499,N_24859,N_24857);
nor UO_1500 (O_1500,N_24813,N_24828);
or UO_1501 (O_1501,N_24979,N_24846);
nand UO_1502 (O_1502,N_24890,N_24898);
nor UO_1503 (O_1503,N_24949,N_24840);
nor UO_1504 (O_1504,N_24878,N_24866);
and UO_1505 (O_1505,N_24801,N_24844);
nor UO_1506 (O_1506,N_24920,N_24883);
xnor UO_1507 (O_1507,N_24805,N_24871);
or UO_1508 (O_1508,N_24955,N_24814);
xnor UO_1509 (O_1509,N_24957,N_24933);
nor UO_1510 (O_1510,N_24831,N_24834);
or UO_1511 (O_1511,N_24884,N_24990);
and UO_1512 (O_1512,N_24875,N_24835);
nand UO_1513 (O_1513,N_24970,N_24909);
nor UO_1514 (O_1514,N_24981,N_24863);
or UO_1515 (O_1515,N_24951,N_24978);
or UO_1516 (O_1516,N_24980,N_24976);
nand UO_1517 (O_1517,N_24913,N_24963);
or UO_1518 (O_1518,N_24955,N_24808);
nand UO_1519 (O_1519,N_24883,N_24827);
nand UO_1520 (O_1520,N_24819,N_24833);
nor UO_1521 (O_1521,N_24911,N_24922);
nand UO_1522 (O_1522,N_24977,N_24825);
nor UO_1523 (O_1523,N_24947,N_24960);
nand UO_1524 (O_1524,N_24995,N_24927);
nor UO_1525 (O_1525,N_24952,N_24908);
or UO_1526 (O_1526,N_24906,N_24945);
nor UO_1527 (O_1527,N_24960,N_24961);
nor UO_1528 (O_1528,N_24901,N_24836);
nand UO_1529 (O_1529,N_24917,N_24827);
nand UO_1530 (O_1530,N_24966,N_24977);
nand UO_1531 (O_1531,N_24867,N_24978);
nor UO_1532 (O_1532,N_24858,N_24932);
nor UO_1533 (O_1533,N_24878,N_24960);
and UO_1534 (O_1534,N_24994,N_24912);
nand UO_1535 (O_1535,N_24875,N_24870);
and UO_1536 (O_1536,N_24924,N_24927);
nor UO_1537 (O_1537,N_24905,N_24988);
or UO_1538 (O_1538,N_24933,N_24884);
nand UO_1539 (O_1539,N_24870,N_24945);
nor UO_1540 (O_1540,N_24829,N_24975);
xnor UO_1541 (O_1541,N_24959,N_24819);
and UO_1542 (O_1542,N_24878,N_24913);
or UO_1543 (O_1543,N_24869,N_24982);
and UO_1544 (O_1544,N_24816,N_24829);
nor UO_1545 (O_1545,N_24809,N_24992);
or UO_1546 (O_1546,N_24801,N_24842);
or UO_1547 (O_1547,N_24848,N_24954);
nor UO_1548 (O_1548,N_24876,N_24866);
nor UO_1549 (O_1549,N_24900,N_24985);
nor UO_1550 (O_1550,N_24985,N_24898);
xor UO_1551 (O_1551,N_24835,N_24831);
or UO_1552 (O_1552,N_24975,N_24831);
and UO_1553 (O_1553,N_24860,N_24813);
or UO_1554 (O_1554,N_24874,N_24889);
nand UO_1555 (O_1555,N_24819,N_24985);
and UO_1556 (O_1556,N_24952,N_24901);
xor UO_1557 (O_1557,N_24932,N_24980);
and UO_1558 (O_1558,N_24978,N_24907);
nor UO_1559 (O_1559,N_24829,N_24904);
or UO_1560 (O_1560,N_24883,N_24874);
and UO_1561 (O_1561,N_24883,N_24900);
xor UO_1562 (O_1562,N_24831,N_24918);
nor UO_1563 (O_1563,N_24824,N_24811);
nor UO_1564 (O_1564,N_24809,N_24848);
nor UO_1565 (O_1565,N_24877,N_24847);
and UO_1566 (O_1566,N_24962,N_24841);
nand UO_1567 (O_1567,N_24974,N_24981);
and UO_1568 (O_1568,N_24836,N_24985);
nor UO_1569 (O_1569,N_24812,N_24828);
or UO_1570 (O_1570,N_24849,N_24807);
and UO_1571 (O_1571,N_24906,N_24879);
and UO_1572 (O_1572,N_24807,N_24930);
nor UO_1573 (O_1573,N_24928,N_24961);
or UO_1574 (O_1574,N_24926,N_24933);
or UO_1575 (O_1575,N_24812,N_24996);
and UO_1576 (O_1576,N_24899,N_24914);
and UO_1577 (O_1577,N_24975,N_24845);
nor UO_1578 (O_1578,N_24934,N_24800);
and UO_1579 (O_1579,N_24996,N_24927);
and UO_1580 (O_1580,N_24996,N_24997);
xnor UO_1581 (O_1581,N_24850,N_24969);
nor UO_1582 (O_1582,N_24912,N_24811);
and UO_1583 (O_1583,N_24952,N_24801);
and UO_1584 (O_1584,N_24929,N_24805);
nand UO_1585 (O_1585,N_24875,N_24865);
nor UO_1586 (O_1586,N_24947,N_24835);
xor UO_1587 (O_1587,N_24918,N_24828);
xnor UO_1588 (O_1588,N_24962,N_24926);
and UO_1589 (O_1589,N_24906,N_24911);
nand UO_1590 (O_1590,N_24899,N_24828);
nand UO_1591 (O_1591,N_24971,N_24977);
xnor UO_1592 (O_1592,N_24835,N_24891);
and UO_1593 (O_1593,N_24950,N_24925);
or UO_1594 (O_1594,N_24906,N_24959);
nor UO_1595 (O_1595,N_24991,N_24934);
nor UO_1596 (O_1596,N_24916,N_24842);
or UO_1597 (O_1597,N_24863,N_24942);
nand UO_1598 (O_1598,N_24834,N_24808);
nand UO_1599 (O_1599,N_24800,N_24978);
or UO_1600 (O_1600,N_24874,N_24809);
or UO_1601 (O_1601,N_24847,N_24865);
nor UO_1602 (O_1602,N_24895,N_24998);
nand UO_1603 (O_1603,N_24822,N_24946);
or UO_1604 (O_1604,N_24887,N_24947);
or UO_1605 (O_1605,N_24813,N_24949);
xnor UO_1606 (O_1606,N_24897,N_24932);
xnor UO_1607 (O_1607,N_24821,N_24806);
or UO_1608 (O_1608,N_24914,N_24918);
nor UO_1609 (O_1609,N_24847,N_24886);
or UO_1610 (O_1610,N_24903,N_24835);
nor UO_1611 (O_1611,N_24938,N_24951);
nor UO_1612 (O_1612,N_24888,N_24810);
nor UO_1613 (O_1613,N_24801,N_24825);
and UO_1614 (O_1614,N_24807,N_24970);
nor UO_1615 (O_1615,N_24955,N_24830);
nand UO_1616 (O_1616,N_24932,N_24949);
xnor UO_1617 (O_1617,N_24934,N_24994);
nand UO_1618 (O_1618,N_24964,N_24858);
or UO_1619 (O_1619,N_24833,N_24884);
or UO_1620 (O_1620,N_24899,N_24850);
nor UO_1621 (O_1621,N_24928,N_24908);
xor UO_1622 (O_1622,N_24931,N_24942);
and UO_1623 (O_1623,N_24866,N_24899);
xnor UO_1624 (O_1624,N_24960,N_24807);
or UO_1625 (O_1625,N_24802,N_24935);
or UO_1626 (O_1626,N_24918,N_24880);
nor UO_1627 (O_1627,N_24973,N_24887);
nand UO_1628 (O_1628,N_24979,N_24849);
nand UO_1629 (O_1629,N_24804,N_24954);
nand UO_1630 (O_1630,N_24816,N_24897);
nor UO_1631 (O_1631,N_24896,N_24885);
xor UO_1632 (O_1632,N_24911,N_24905);
xnor UO_1633 (O_1633,N_24907,N_24882);
and UO_1634 (O_1634,N_24896,N_24832);
and UO_1635 (O_1635,N_24951,N_24846);
nor UO_1636 (O_1636,N_24950,N_24906);
and UO_1637 (O_1637,N_24849,N_24939);
and UO_1638 (O_1638,N_24912,N_24930);
nand UO_1639 (O_1639,N_24829,N_24929);
xor UO_1640 (O_1640,N_24971,N_24890);
and UO_1641 (O_1641,N_24808,N_24931);
xor UO_1642 (O_1642,N_24836,N_24838);
xnor UO_1643 (O_1643,N_24976,N_24890);
xnor UO_1644 (O_1644,N_24884,N_24971);
nand UO_1645 (O_1645,N_24873,N_24868);
and UO_1646 (O_1646,N_24847,N_24842);
or UO_1647 (O_1647,N_24878,N_24951);
and UO_1648 (O_1648,N_24845,N_24897);
and UO_1649 (O_1649,N_24829,N_24910);
nand UO_1650 (O_1650,N_24871,N_24815);
or UO_1651 (O_1651,N_24838,N_24875);
xor UO_1652 (O_1652,N_24927,N_24914);
and UO_1653 (O_1653,N_24910,N_24966);
and UO_1654 (O_1654,N_24878,N_24868);
nor UO_1655 (O_1655,N_24912,N_24929);
or UO_1656 (O_1656,N_24882,N_24883);
nand UO_1657 (O_1657,N_24894,N_24837);
and UO_1658 (O_1658,N_24898,N_24868);
or UO_1659 (O_1659,N_24883,N_24846);
or UO_1660 (O_1660,N_24923,N_24997);
nand UO_1661 (O_1661,N_24908,N_24810);
xor UO_1662 (O_1662,N_24856,N_24960);
nor UO_1663 (O_1663,N_24874,N_24958);
xnor UO_1664 (O_1664,N_24876,N_24814);
or UO_1665 (O_1665,N_24976,N_24857);
or UO_1666 (O_1666,N_24874,N_24845);
xnor UO_1667 (O_1667,N_24810,N_24926);
or UO_1668 (O_1668,N_24964,N_24942);
nand UO_1669 (O_1669,N_24972,N_24966);
xor UO_1670 (O_1670,N_24998,N_24992);
and UO_1671 (O_1671,N_24978,N_24968);
or UO_1672 (O_1672,N_24809,N_24904);
or UO_1673 (O_1673,N_24826,N_24977);
and UO_1674 (O_1674,N_24901,N_24886);
and UO_1675 (O_1675,N_24995,N_24985);
and UO_1676 (O_1676,N_24804,N_24942);
and UO_1677 (O_1677,N_24817,N_24941);
xor UO_1678 (O_1678,N_24930,N_24936);
or UO_1679 (O_1679,N_24869,N_24829);
xnor UO_1680 (O_1680,N_24976,N_24842);
xnor UO_1681 (O_1681,N_24815,N_24894);
nor UO_1682 (O_1682,N_24944,N_24822);
or UO_1683 (O_1683,N_24816,N_24906);
and UO_1684 (O_1684,N_24801,N_24984);
xor UO_1685 (O_1685,N_24944,N_24843);
or UO_1686 (O_1686,N_24807,N_24833);
xor UO_1687 (O_1687,N_24873,N_24838);
nand UO_1688 (O_1688,N_24886,N_24905);
nor UO_1689 (O_1689,N_24925,N_24823);
xor UO_1690 (O_1690,N_24894,N_24921);
nor UO_1691 (O_1691,N_24945,N_24900);
xnor UO_1692 (O_1692,N_24839,N_24865);
or UO_1693 (O_1693,N_24805,N_24819);
or UO_1694 (O_1694,N_24867,N_24887);
xor UO_1695 (O_1695,N_24987,N_24932);
xor UO_1696 (O_1696,N_24963,N_24818);
or UO_1697 (O_1697,N_24801,N_24909);
xor UO_1698 (O_1698,N_24913,N_24894);
or UO_1699 (O_1699,N_24918,N_24955);
nand UO_1700 (O_1700,N_24986,N_24890);
xnor UO_1701 (O_1701,N_24919,N_24833);
nor UO_1702 (O_1702,N_24972,N_24851);
and UO_1703 (O_1703,N_24887,N_24875);
nand UO_1704 (O_1704,N_24878,N_24956);
or UO_1705 (O_1705,N_24833,N_24975);
and UO_1706 (O_1706,N_24845,N_24901);
nor UO_1707 (O_1707,N_24823,N_24899);
nor UO_1708 (O_1708,N_24832,N_24908);
nor UO_1709 (O_1709,N_24915,N_24913);
nor UO_1710 (O_1710,N_24956,N_24831);
or UO_1711 (O_1711,N_24942,N_24953);
nor UO_1712 (O_1712,N_24955,N_24911);
xor UO_1713 (O_1713,N_24843,N_24945);
or UO_1714 (O_1714,N_24851,N_24995);
and UO_1715 (O_1715,N_24902,N_24861);
nor UO_1716 (O_1716,N_24909,N_24962);
xor UO_1717 (O_1717,N_24820,N_24965);
xor UO_1718 (O_1718,N_24928,N_24819);
nor UO_1719 (O_1719,N_24858,N_24983);
and UO_1720 (O_1720,N_24810,N_24876);
nand UO_1721 (O_1721,N_24886,N_24989);
nor UO_1722 (O_1722,N_24816,N_24924);
or UO_1723 (O_1723,N_24899,N_24861);
or UO_1724 (O_1724,N_24880,N_24943);
or UO_1725 (O_1725,N_24968,N_24868);
xnor UO_1726 (O_1726,N_24922,N_24918);
xor UO_1727 (O_1727,N_24902,N_24884);
nand UO_1728 (O_1728,N_24804,N_24809);
and UO_1729 (O_1729,N_24806,N_24869);
nand UO_1730 (O_1730,N_24804,N_24982);
nor UO_1731 (O_1731,N_24869,N_24875);
xor UO_1732 (O_1732,N_24853,N_24945);
and UO_1733 (O_1733,N_24805,N_24816);
or UO_1734 (O_1734,N_24820,N_24884);
nand UO_1735 (O_1735,N_24946,N_24865);
xnor UO_1736 (O_1736,N_24936,N_24834);
or UO_1737 (O_1737,N_24930,N_24831);
nor UO_1738 (O_1738,N_24867,N_24833);
xor UO_1739 (O_1739,N_24835,N_24968);
nand UO_1740 (O_1740,N_24950,N_24946);
nand UO_1741 (O_1741,N_24997,N_24903);
and UO_1742 (O_1742,N_24939,N_24933);
nand UO_1743 (O_1743,N_24857,N_24981);
or UO_1744 (O_1744,N_24955,N_24824);
nand UO_1745 (O_1745,N_24815,N_24821);
nand UO_1746 (O_1746,N_24886,N_24888);
or UO_1747 (O_1747,N_24902,N_24896);
and UO_1748 (O_1748,N_24994,N_24831);
or UO_1749 (O_1749,N_24996,N_24905);
and UO_1750 (O_1750,N_24850,N_24828);
nor UO_1751 (O_1751,N_24927,N_24908);
nand UO_1752 (O_1752,N_24880,N_24941);
nand UO_1753 (O_1753,N_24886,N_24950);
xor UO_1754 (O_1754,N_24911,N_24987);
xnor UO_1755 (O_1755,N_24875,N_24878);
nor UO_1756 (O_1756,N_24912,N_24992);
and UO_1757 (O_1757,N_24816,N_24873);
xor UO_1758 (O_1758,N_24962,N_24803);
nor UO_1759 (O_1759,N_24879,N_24893);
nor UO_1760 (O_1760,N_24932,N_24821);
xor UO_1761 (O_1761,N_24993,N_24873);
xor UO_1762 (O_1762,N_24944,N_24905);
nor UO_1763 (O_1763,N_24838,N_24912);
or UO_1764 (O_1764,N_24893,N_24823);
xor UO_1765 (O_1765,N_24823,N_24915);
nor UO_1766 (O_1766,N_24848,N_24845);
and UO_1767 (O_1767,N_24930,N_24895);
nand UO_1768 (O_1768,N_24954,N_24927);
and UO_1769 (O_1769,N_24883,N_24886);
xnor UO_1770 (O_1770,N_24980,N_24847);
xnor UO_1771 (O_1771,N_24983,N_24822);
nand UO_1772 (O_1772,N_24956,N_24857);
and UO_1773 (O_1773,N_24903,N_24947);
and UO_1774 (O_1774,N_24839,N_24960);
nor UO_1775 (O_1775,N_24883,N_24817);
and UO_1776 (O_1776,N_24856,N_24857);
nor UO_1777 (O_1777,N_24841,N_24857);
xor UO_1778 (O_1778,N_24994,N_24973);
and UO_1779 (O_1779,N_24930,N_24867);
or UO_1780 (O_1780,N_24863,N_24833);
xnor UO_1781 (O_1781,N_24820,N_24907);
or UO_1782 (O_1782,N_24817,N_24801);
or UO_1783 (O_1783,N_24932,N_24854);
and UO_1784 (O_1784,N_24855,N_24990);
nor UO_1785 (O_1785,N_24806,N_24819);
or UO_1786 (O_1786,N_24815,N_24843);
or UO_1787 (O_1787,N_24948,N_24995);
nand UO_1788 (O_1788,N_24997,N_24950);
and UO_1789 (O_1789,N_24984,N_24804);
or UO_1790 (O_1790,N_24972,N_24844);
or UO_1791 (O_1791,N_24813,N_24924);
xor UO_1792 (O_1792,N_24982,N_24949);
nand UO_1793 (O_1793,N_24968,N_24828);
xor UO_1794 (O_1794,N_24999,N_24836);
or UO_1795 (O_1795,N_24875,N_24843);
and UO_1796 (O_1796,N_24990,N_24908);
or UO_1797 (O_1797,N_24850,N_24832);
and UO_1798 (O_1798,N_24909,N_24927);
xnor UO_1799 (O_1799,N_24854,N_24826);
or UO_1800 (O_1800,N_24965,N_24884);
and UO_1801 (O_1801,N_24940,N_24918);
or UO_1802 (O_1802,N_24843,N_24921);
and UO_1803 (O_1803,N_24843,N_24867);
nand UO_1804 (O_1804,N_24933,N_24843);
nor UO_1805 (O_1805,N_24887,N_24823);
and UO_1806 (O_1806,N_24941,N_24945);
nor UO_1807 (O_1807,N_24914,N_24840);
and UO_1808 (O_1808,N_24969,N_24842);
and UO_1809 (O_1809,N_24918,N_24902);
nand UO_1810 (O_1810,N_24825,N_24960);
nor UO_1811 (O_1811,N_24943,N_24954);
nor UO_1812 (O_1812,N_24859,N_24886);
nand UO_1813 (O_1813,N_24853,N_24951);
nand UO_1814 (O_1814,N_24935,N_24887);
xnor UO_1815 (O_1815,N_24971,N_24909);
or UO_1816 (O_1816,N_24803,N_24844);
xor UO_1817 (O_1817,N_24944,N_24867);
and UO_1818 (O_1818,N_24962,N_24868);
and UO_1819 (O_1819,N_24943,N_24901);
nand UO_1820 (O_1820,N_24835,N_24877);
nor UO_1821 (O_1821,N_24938,N_24929);
xor UO_1822 (O_1822,N_24857,N_24835);
xor UO_1823 (O_1823,N_24827,N_24935);
and UO_1824 (O_1824,N_24950,N_24823);
nand UO_1825 (O_1825,N_24841,N_24858);
or UO_1826 (O_1826,N_24855,N_24983);
nand UO_1827 (O_1827,N_24852,N_24881);
nand UO_1828 (O_1828,N_24988,N_24810);
and UO_1829 (O_1829,N_24865,N_24814);
nor UO_1830 (O_1830,N_24922,N_24949);
nand UO_1831 (O_1831,N_24834,N_24828);
xor UO_1832 (O_1832,N_24968,N_24829);
nor UO_1833 (O_1833,N_24935,N_24814);
nor UO_1834 (O_1834,N_24952,N_24930);
nor UO_1835 (O_1835,N_24806,N_24863);
xor UO_1836 (O_1836,N_24804,N_24937);
or UO_1837 (O_1837,N_24839,N_24940);
xor UO_1838 (O_1838,N_24905,N_24883);
nor UO_1839 (O_1839,N_24963,N_24951);
xnor UO_1840 (O_1840,N_24983,N_24880);
nand UO_1841 (O_1841,N_24868,N_24853);
nand UO_1842 (O_1842,N_24958,N_24839);
nand UO_1843 (O_1843,N_24845,N_24924);
and UO_1844 (O_1844,N_24828,N_24891);
and UO_1845 (O_1845,N_24940,N_24803);
or UO_1846 (O_1846,N_24896,N_24842);
nand UO_1847 (O_1847,N_24940,N_24930);
xnor UO_1848 (O_1848,N_24975,N_24849);
and UO_1849 (O_1849,N_24927,N_24992);
and UO_1850 (O_1850,N_24815,N_24801);
nor UO_1851 (O_1851,N_24851,N_24843);
nor UO_1852 (O_1852,N_24995,N_24937);
nand UO_1853 (O_1853,N_24815,N_24924);
nor UO_1854 (O_1854,N_24821,N_24905);
or UO_1855 (O_1855,N_24910,N_24996);
nor UO_1856 (O_1856,N_24926,N_24877);
and UO_1857 (O_1857,N_24802,N_24842);
nor UO_1858 (O_1858,N_24907,N_24802);
xor UO_1859 (O_1859,N_24967,N_24882);
and UO_1860 (O_1860,N_24828,N_24996);
xnor UO_1861 (O_1861,N_24957,N_24817);
nor UO_1862 (O_1862,N_24939,N_24983);
nor UO_1863 (O_1863,N_24916,N_24875);
and UO_1864 (O_1864,N_24896,N_24942);
xnor UO_1865 (O_1865,N_24891,N_24867);
nand UO_1866 (O_1866,N_24804,N_24814);
nor UO_1867 (O_1867,N_24871,N_24806);
nor UO_1868 (O_1868,N_24808,N_24901);
and UO_1869 (O_1869,N_24984,N_24803);
and UO_1870 (O_1870,N_24951,N_24838);
nand UO_1871 (O_1871,N_24928,N_24851);
nor UO_1872 (O_1872,N_24914,N_24824);
and UO_1873 (O_1873,N_24906,N_24968);
nor UO_1874 (O_1874,N_24953,N_24828);
or UO_1875 (O_1875,N_24823,N_24803);
nor UO_1876 (O_1876,N_24813,N_24961);
and UO_1877 (O_1877,N_24837,N_24860);
xor UO_1878 (O_1878,N_24976,N_24948);
nor UO_1879 (O_1879,N_24816,N_24937);
xnor UO_1880 (O_1880,N_24932,N_24803);
nor UO_1881 (O_1881,N_24847,N_24898);
nand UO_1882 (O_1882,N_24965,N_24886);
or UO_1883 (O_1883,N_24816,N_24849);
xnor UO_1884 (O_1884,N_24907,N_24838);
and UO_1885 (O_1885,N_24915,N_24943);
nor UO_1886 (O_1886,N_24899,N_24805);
or UO_1887 (O_1887,N_24946,N_24879);
and UO_1888 (O_1888,N_24960,N_24846);
and UO_1889 (O_1889,N_24900,N_24839);
xor UO_1890 (O_1890,N_24944,N_24869);
xnor UO_1891 (O_1891,N_24908,N_24932);
and UO_1892 (O_1892,N_24895,N_24831);
xnor UO_1893 (O_1893,N_24846,N_24824);
and UO_1894 (O_1894,N_24962,N_24864);
nand UO_1895 (O_1895,N_24998,N_24942);
nor UO_1896 (O_1896,N_24800,N_24986);
nand UO_1897 (O_1897,N_24813,N_24859);
nand UO_1898 (O_1898,N_24992,N_24827);
or UO_1899 (O_1899,N_24852,N_24819);
xor UO_1900 (O_1900,N_24802,N_24870);
or UO_1901 (O_1901,N_24976,N_24904);
nand UO_1902 (O_1902,N_24806,N_24950);
nor UO_1903 (O_1903,N_24991,N_24872);
or UO_1904 (O_1904,N_24875,N_24848);
nand UO_1905 (O_1905,N_24900,N_24846);
and UO_1906 (O_1906,N_24960,N_24902);
nand UO_1907 (O_1907,N_24842,N_24870);
nand UO_1908 (O_1908,N_24929,N_24922);
xnor UO_1909 (O_1909,N_24816,N_24863);
and UO_1910 (O_1910,N_24819,N_24918);
or UO_1911 (O_1911,N_24875,N_24861);
or UO_1912 (O_1912,N_24991,N_24946);
xor UO_1913 (O_1913,N_24835,N_24846);
nand UO_1914 (O_1914,N_24807,N_24941);
and UO_1915 (O_1915,N_24917,N_24871);
xnor UO_1916 (O_1916,N_24811,N_24829);
xor UO_1917 (O_1917,N_24939,N_24900);
xnor UO_1918 (O_1918,N_24999,N_24858);
nor UO_1919 (O_1919,N_24967,N_24812);
nand UO_1920 (O_1920,N_24809,N_24833);
and UO_1921 (O_1921,N_24864,N_24977);
or UO_1922 (O_1922,N_24820,N_24844);
and UO_1923 (O_1923,N_24877,N_24866);
xor UO_1924 (O_1924,N_24828,N_24948);
and UO_1925 (O_1925,N_24926,N_24896);
and UO_1926 (O_1926,N_24969,N_24910);
or UO_1927 (O_1927,N_24836,N_24800);
nor UO_1928 (O_1928,N_24828,N_24887);
nand UO_1929 (O_1929,N_24954,N_24838);
or UO_1930 (O_1930,N_24838,N_24842);
xnor UO_1931 (O_1931,N_24889,N_24881);
and UO_1932 (O_1932,N_24996,N_24882);
or UO_1933 (O_1933,N_24930,N_24914);
xor UO_1934 (O_1934,N_24973,N_24953);
nand UO_1935 (O_1935,N_24872,N_24941);
or UO_1936 (O_1936,N_24802,N_24861);
or UO_1937 (O_1937,N_24996,N_24909);
and UO_1938 (O_1938,N_24868,N_24844);
xor UO_1939 (O_1939,N_24850,N_24839);
and UO_1940 (O_1940,N_24867,N_24953);
or UO_1941 (O_1941,N_24856,N_24992);
or UO_1942 (O_1942,N_24833,N_24910);
or UO_1943 (O_1943,N_24866,N_24835);
or UO_1944 (O_1944,N_24865,N_24909);
nor UO_1945 (O_1945,N_24969,N_24838);
nand UO_1946 (O_1946,N_24958,N_24995);
or UO_1947 (O_1947,N_24955,N_24978);
nand UO_1948 (O_1948,N_24816,N_24833);
or UO_1949 (O_1949,N_24867,N_24917);
or UO_1950 (O_1950,N_24812,N_24966);
nor UO_1951 (O_1951,N_24817,N_24985);
nor UO_1952 (O_1952,N_24906,N_24904);
or UO_1953 (O_1953,N_24996,N_24861);
xor UO_1954 (O_1954,N_24900,N_24885);
nand UO_1955 (O_1955,N_24939,N_24948);
and UO_1956 (O_1956,N_24890,N_24914);
xnor UO_1957 (O_1957,N_24908,N_24872);
or UO_1958 (O_1958,N_24853,N_24906);
and UO_1959 (O_1959,N_24920,N_24858);
or UO_1960 (O_1960,N_24941,N_24958);
and UO_1961 (O_1961,N_24998,N_24937);
and UO_1962 (O_1962,N_24958,N_24915);
and UO_1963 (O_1963,N_24919,N_24822);
or UO_1964 (O_1964,N_24816,N_24884);
nor UO_1965 (O_1965,N_24916,N_24974);
and UO_1966 (O_1966,N_24920,N_24994);
nor UO_1967 (O_1967,N_24883,N_24996);
nor UO_1968 (O_1968,N_24979,N_24847);
nor UO_1969 (O_1969,N_24864,N_24931);
nor UO_1970 (O_1970,N_24916,N_24846);
or UO_1971 (O_1971,N_24815,N_24904);
and UO_1972 (O_1972,N_24824,N_24928);
and UO_1973 (O_1973,N_24902,N_24936);
and UO_1974 (O_1974,N_24956,N_24920);
or UO_1975 (O_1975,N_24897,N_24996);
nand UO_1976 (O_1976,N_24819,N_24934);
and UO_1977 (O_1977,N_24911,N_24957);
xor UO_1978 (O_1978,N_24945,N_24954);
nand UO_1979 (O_1979,N_24975,N_24896);
or UO_1980 (O_1980,N_24967,N_24803);
xnor UO_1981 (O_1981,N_24974,N_24890);
nor UO_1982 (O_1982,N_24821,N_24964);
and UO_1983 (O_1983,N_24864,N_24999);
nor UO_1984 (O_1984,N_24961,N_24834);
nand UO_1985 (O_1985,N_24930,N_24889);
and UO_1986 (O_1986,N_24853,N_24862);
xnor UO_1987 (O_1987,N_24837,N_24873);
nor UO_1988 (O_1988,N_24803,N_24840);
and UO_1989 (O_1989,N_24875,N_24942);
nand UO_1990 (O_1990,N_24805,N_24831);
xor UO_1991 (O_1991,N_24860,N_24817);
nor UO_1992 (O_1992,N_24924,N_24972);
and UO_1993 (O_1993,N_24913,N_24825);
nand UO_1994 (O_1994,N_24895,N_24839);
nand UO_1995 (O_1995,N_24807,N_24961);
or UO_1996 (O_1996,N_24971,N_24807);
nand UO_1997 (O_1997,N_24884,N_24832);
or UO_1998 (O_1998,N_24823,N_24841);
nor UO_1999 (O_1999,N_24825,N_24921);
and UO_2000 (O_2000,N_24987,N_24883);
xor UO_2001 (O_2001,N_24842,N_24985);
and UO_2002 (O_2002,N_24840,N_24896);
nor UO_2003 (O_2003,N_24937,N_24801);
and UO_2004 (O_2004,N_24827,N_24819);
nand UO_2005 (O_2005,N_24806,N_24962);
or UO_2006 (O_2006,N_24956,N_24959);
nand UO_2007 (O_2007,N_24955,N_24926);
nand UO_2008 (O_2008,N_24933,N_24823);
xor UO_2009 (O_2009,N_24911,N_24949);
and UO_2010 (O_2010,N_24937,N_24851);
nor UO_2011 (O_2011,N_24831,N_24979);
or UO_2012 (O_2012,N_24992,N_24942);
nand UO_2013 (O_2013,N_24953,N_24854);
nor UO_2014 (O_2014,N_24802,N_24920);
and UO_2015 (O_2015,N_24888,N_24971);
nor UO_2016 (O_2016,N_24814,N_24857);
nor UO_2017 (O_2017,N_24836,N_24928);
nor UO_2018 (O_2018,N_24819,N_24891);
and UO_2019 (O_2019,N_24898,N_24843);
nand UO_2020 (O_2020,N_24921,N_24903);
xnor UO_2021 (O_2021,N_24840,N_24868);
nand UO_2022 (O_2022,N_24980,N_24954);
and UO_2023 (O_2023,N_24835,N_24955);
xnor UO_2024 (O_2024,N_24892,N_24886);
or UO_2025 (O_2025,N_24913,N_24859);
nor UO_2026 (O_2026,N_24971,N_24841);
nand UO_2027 (O_2027,N_24876,N_24990);
xnor UO_2028 (O_2028,N_24869,N_24824);
and UO_2029 (O_2029,N_24980,N_24825);
nor UO_2030 (O_2030,N_24991,N_24833);
nor UO_2031 (O_2031,N_24940,N_24984);
nand UO_2032 (O_2032,N_24825,N_24906);
nor UO_2033 (O_2033,N_24809,N_24897);
or UO_2034 (O_2034,N_24935,N_24919);
nand UO_2035 (O_2035,N_24813,N_24950);
nand UO_2036 (O_2036,N_24835,N_24863);
xor UO_2037 (O_2037,N_24811,N_24838);
nor UO_2038 (O_2038,N_24985,N_24861);
or UO_2039 (O_2039,N_24971,N_24939);
nor UO_2040 (O_2040,N_24849,N_24946);
nand UO_2041 (O_2041,N_24813,N_24877);
nand UO_2042 (O_2042,N_24943,N_24840);
and UO_2043 (O_2043,N_24826,N_24834);
nor UO_2044 (O_2044,N_24935,N_24989);
nor UO_2045 (O_2045,N_24903,N_24916);
nor UO_2046 (O_2046,N_24998,N_24938);
and UO_2047 (O_2047,N_24841,N_24809);
nand UO_2048 (O_2048,N_24916,N_24964);
nor UO_2049 (O_2049,N_24975,N_24942);
nor UO_2050 (O_2050,N_24810,N_24833);
and UO_2051 (O_2051,N_24980,N_24801);
or UO_2052 (O_2052,N_24992,N_24907);
xor UO_2053 (O_2053,N_24834,N_24842);
or UO_2054 (O_2054,N_24829,N_24899);
nand UO_2055 (O_2055,N_24888,N_24814);
nor UO_2056 (O_2056,N_24997,N_24860);
nor UO_2057 (O_2057,N_24966,N_24925);
or UO_2058 (O_2058,N_24994,N_24992);
nor UO_2059 (O_2059,N_24855,N_24936);
nor UO_2060 (O_2060,N_24981,N_24977);
xor UO_2061 (O_2061,N_24923,N_24995);
nor UO_2062 (O_2062,N_24869,N_24915);
nor UO_2063 (O_2063,N_24830,N_24829);
nor UO_2064 (O_2064,N_24925,N_24880);
nor UO_2065 (O_2065,N_24987,N_24976);
xor UO_2066 (O_2066,N_24839,N_24873);
xnor UO_2067 (O_2067,N_24844,N_24979);
nor UO_2068 (O_2068,N_24881,N_24893);
or UO_2069 (O_2069,N_24951,N_24970);
or UO_2070 (O_2070,N_24928,N_24892);
or UO_2071 (O_2071,N_24993,N_24973);
or UO_2072 (O_2072,N_24841,N_24818);
xnor UO_2073 (O_2073,N_24888,N_24836);
xnor UO_2074 (O_2074,N_24849,N_24921);
nand UO_2075 (O_2075,N_24988,N_24963);
and UO_2076 (O_2076,N_24838,N_24900);
and UO_2077 (O_2077,N_24959,N_24854);
nand UO_2078 (O_2078,N_24889,N_24922);
xor UO_2079 (O_2079,N_24989,N_24842);
nand UO_2080 (O_2080,N_24965,N_24881);
nor UO_2081 (O_2081,N_24954,N_24803);
xor UO_2082 (O_2082,N_24915,N_24921);
xnor UO_2083 (O_2083,N_24879,N_24925);
xor UO_2084 (O_2084,N_24982,N_24934);
or UO_2085 (O_2085,N_24973,N_24876);
nand UO_2086 (O_2086,N_24864,N_24892);
and UO_2087 (O_2087,N_24870,N_24859);
nor UO_2088 (O_2088,N_24929,N_24811);
or UO_2089 (O_2089,N_24878,N_24852);
and UO_2090 (O_2090,N_24941,N_24863);
nor UO_2091 (O_2091,N_24983,N_24938);
and UO_2092 (O_2092,N_24890,N_24850);
nand UO_2093 (O_2093,N_24988,N_24881);
nand UO_2094 (O_2094,N_24816,N_24867);
xor UO_2095 (O_2095,N_24801,N_24999);
and UO_2096 (O_2096,N_24856,N_24953);
xor UO_2097 (O_2097,N_24822,N_24892);
xor UO_2098 (O_2098,N_24968,N_24945);
xor UO_2099 (O_2099,N_24845,N_24832);
and UO_2100 (O_2100,N_24817,N_24967);
nand UO_2101 (O_2101,N_24971,N_24989);
nor UO_2102 (O_2102,N_24972,N_24860);
nor UO_2103 (O_2103,N_24916,N_24883);
nor UO_2104 (O_2104,N_24890,N_24980);
and UO_2105 (O_2105,N_24991,N_24835);
or UO_2106 (O_2106,N_24979,N_24901);
xor UO_2107 (O_2107,N_24931,N_24934);
nor UO_2108 (O_2108,N_24928,N_24929);
and UO_2109 (O_2109,N_24817,N_24847);
nand UO_2110 (O_2110,N_24962,N_24854);
xnor UO_2111 (O_2111,N_24927,N_24890);
nor UO_2112 (O_2112,N_24941,N_24862);
or UO_2113 (O_2113,N_24987,N_24992);
nor UO_2114 (O_2114,N_24917,N_24945);
xnor UO_2115 (O_2115,N_24978,N_24837);
and UO_2116 (O_2116,N_24809,N_24828);
and UO_2117 (O_2117,N_24988,N_24931);
and UO_2118 (O_2118,N_24958,N_24972);
or UO_2119 (O_2119,N_24900,N_24842);
nor UO_2120 (O_2120,N_24822,N_24889);
xor UO_2121 (O_2121,N_24981,N_24865);
nor UO_2122 (O_2122,N_24933,N_24835);
xor UO_2123 (O_2123,N_24842,N_24855);
xnor UO_2124 (O_2124,N_24961,N_24998);
nand UO_2125 (O_2125,N_24815,N_24848);
xnor UO_2126 (O_2126,N_24921,N_24817);
or UO_2127 (O_2127,N_24934,N_24858);
and UO_2128 (O_2128,N_24881,N_24939);
nor UO_2129 (O_2129,N_24807,N_24986);
nand UO_2130 (O_2130,N_24993,N_24959);
nor UO_2131 (O_2131,N_24985,N_24944);
nor UO_2132 (O_2132,N_24905,N_24819);
and UO_2133 (O_2133,N_24811,N_24921);
xor UO_2134 (O_2134,N_24961,N_24924);
nor UO_2135 (O_2135,N_24931,N_24969);
xnor UO_2136 (O_2136,N_24867,N_24935);
or UO_2137 (O_2137,N_24956,N_24957);
xnor UO_2138 (O_2138,N_24971,N_24896);
or UO_2139 (O_2139,N_24913,N_24827);
nor UO_2140 (O_2140,N_24830,N_24974);
xnor UO_2141 (O_2141,N_24844,N_24852);
nor UO_2142 (O_2142,N_24845,N_24955);
nand UO_2143 (O_2143,N_24804,N_24966);
xnor UO_2144 (O_2144,N_24817,N_24893);
nor UO_2145 (O_2145,N_24802,N_24942);
nor UO_2146 (O_2146,N_24934,N_24953);
nor UO_2147 (O_2147,N_24981,N_24936);
nor UO_2148 (O_2148,N_24919,N_24996);
nor UO_2149 (O_2149,N_24899,N_24849);
and UO_2150 (O_2150,N_24980,N_24962);
nor UO_2151 (O_2151,N_24877,N_24840);
nor UO_2152 (O_2152,N_24896,N_24919);
nand UO_2153 (O_2153,N_24878,N_24939);
nand UO_2154 (O_2154,N_24927,N_24967);
xor UO_2155 (O_2155,N_24805,N_24872);
and UO_2156 (O_2156,N_24912,N_24907);
nand UO_2157 (O_2157,N_24806,N_24940);
and UO_2158 (O_2158,N_24992,N_24884);
xnor UO_2159 (O_2159,N_24892,N_24919);
or UO_2160 (O_2160,N_24800,N_24977);
xnor UO_2161 (O_2161,N_24883,N_24970);
nand UO_2162 (O_2162,N_24956,N_24946);
or UO_2163 (O_2163,N_24868,N_24920);
nor UO_2164 (O_2164,N_24857,N_24931);
or UO_2165 (O_2165,N_24984,N_24904);
nor UO_2166 (O_2166,N_24921,N_24860);
xnor UO_2167 (O_2167,N_24980,N_24806);
nand UO_2168 (O_2168,N_24932,N_24921);
nor UO_2169 (O_2169,N_24910,N_24927);
nand UO_2170 (O_2170,N_24941,N_24902);
nand UO_2171 (O_2171,N_24977,N_24917);
xor UO_2172 (O_2172,N_24955,N_24877);
and UO_2173 (O_2173,N_24992,N_24925);
nor UO_2174 (O_2174,N_24984,N_24890);
or UO_2175 (O_2175,N_24939,N_24997);
and UO_2176 (O_2176,N_24953,N_24826);
xnor UO_2177 (O_2177,N_24980,N_24968);
xnor UO_2178 (O_2178,N_24837,N_24928);
nor UO_2179 (O_2179,N_24921,N_24812);
nand UO_2180 (O_2180,N_24968,N_24919);
xor UO_2181 (O_2181,N_24891,N_24982);
and UO_2182 (O_2182,N_24879,N_24991);
and UO_2183 (O_2183,N_24876,N_24969);
nor UO_2184 (O_2184,N_24941,N_24815);
or UO_2185 (O_2185,N_24806,N_24850);
or UO_2186 (O_2186,N_24968,N_24813);
xnor UO_2187 (O_2187,N_24983,N_24914);
nand UO_2188 (O_2188,N_24836,N_24990);
xor UO_2189 (O_2189,N_24824,N_24827);
or UO_2190 (O_2190,N_24939,N_24805);
nand UO_2191 (O_2191,N_24853,N_24910);
and UO_2192 (O_2192,N_24847,N_24929);
and UO_2193 (O_2193,N_24818,N_24990);
and UO_2194 (O_2194,N_24894,N_24916);
nand UO_2195 (O_2195,N_24853,N_24996);
nor UO_2196 (O_2196,N_24839,N_24877);
or UO_2197 (O_2197,N_24949,N_24952);
nor UO_2198 (O_2198,N_24984,N_24980);
nor UO_2199 (O_2199,N_24913,N_24807);
xnor UO_2200 (O_2200,N_24888,N_24990);
nand UO_2201 (O_2201,N_24853,N_24826);
xnor UO_2202 (O_2202,N_24891,N_24838);
and UO_2203 (O_2203,N_24902,N_24991);
xor UO_2204 (O_2204,N_24933,N_24886);
and UO_2205 (O_2205,N_24907,N_24968);
nor UO_2206 (O_2206,N_24998,N_24910);
and UO_2207 (O_2207,N_24928,N_24978);
or UO_2208 (O_2208,N_24942,N_24970);
xor UO_2209 (O_2209,N_24843,N_24845);
and UO_2210 (O_2210,N_24891,N_24927);
xnor UO_2211 (O_2211,N_24947,N_24941);
or UO_2212 (O_2212,N_24873,N_24919);
and UO_2213 (O_2213,N_24840,N_24851);
and UO_2214 (O_2214,N_24904,N_24823);
or UO_2215 (O_2215,N_24983,N_24900);
or UO_2216 (O_2216,N_24928,N_24890);
xnor UO_2217 (O_2217,N_24865,N_24908);
nor UO_2218 (O_2218,N_24840,N_24876);
nand UO_2219 (O_2219,N_24878,N_24815);
or UO_2220 (O_2220,N_24960,N_24915);
or UO_2221 (O_2221,N_24822,N_24818);
or UO_2222 (O_2222,N_24880,N_24821);
xnor UO_2223 (O_2223,N_24895,N_24821);
nand UO_2224 (O_2224,N_24988,N_24856);
xnor UO_2225 (O_2225,N_24915,N_24803);
nor UO_2226 (O_2226,N_24801,N_24887);
nor UO_2227 (O_2227,N_24889,N_24964);
xor UO_2228 (O_2228,N_24802,N_24801);
nor UO_2229 (O_2229,N_24861,N_24842);
xnor UO_2230 (O_2230,N_24905,N_24867);
or UO_2231 (O_2231,N_24967,N_24854);
xnor UO_2232 (O_2232,N_24872,N_24997);
nand UO_2233 (O_2233,N_24927,N_24888);
xnor UO_2234 (O_2234,N_24834,N_24983);
nand UO_2235 (O_2235,N_24803,N_24849);
and UO_2236 (O_2236,N_24951,N_24848);
xor UO_2237 (O_2237,N_24922,N_24947);
and UO_2238 (O_2238,N_24888,N_24894);
nand UO_2239 (O_2239,N_24832,N_24960);
nor UO_2240 (O_2240,N_24964,N_24841);
xor UO_2241 (O_2241,N_24819,N_24814);
nor UO_2242 (O_2242,N_24879,N_24964);
and UO_2243 (O_2243,N_24884,N_24887);
nand UO_2244 (O_2244,N_24924,N_24856);
or UO_2245 (O_2245,N_24993,N_24846);
or UO_2246 (O_2246,N_24877,N_24974);
or UO_2247 (O_2247,N_24951,N_24845);
nand UO_2248 (O_2248,N_24935,N_24803);
nor UO_2249 (O_2249,N_24950,N_24850);
nor UO_2250 (O_2250,N_24920,N_24826);
or UO_2251 (O_2251,N_24897,N_24805);
nand UO_2252 (O_2252,N_24952,N_24992);
and UO_2253 (O_2253,N_24912,N_24931);
or UO_2254 (O_2254,N_24907,N_24975);
nand UO_2255 (O_2255,N_24999,N_24888);
nor UO_2256 (O_2256,N_24961,N_24881);
nor UO_2257 (O_2257,N_24911,N_24896);
and UO_2258 (O_2258,N_24851,N_24874);
and UO_2259 (O_2259,N_24934,N_24966);
and UO_2260 (O_2260,N_24976,N_24924);
nand UO_2261 (O_2261,N_24856,N_24891);
xnor UO_2262 (O_2262,N_24974,N_24849);
and UO_2263 (O_2263,N_24951,N_24866);
and UO_2264 (O_2264,N_24919,N_24880);
and UO_2265 (O_2265,N_24970,N_24894);
nor UO_2266 (O_2266,N_24961,N_24876);
nand UO_2267 (O_2267,N_24976,N_24830);
nor UO_2268 (O_2268,N_24916,N_24976);
or UO_2269 (O_2269,N_24811,N_24933);
xor UO_2270 (O_2270,N_24826,N_24957);
nor UO_2271 (O_2271,N_24857,N_24866);
nor UO_2272 (O_2272,N_24809,N_24907);
and UO_2273 (O_2273,N_24844,N_24918);
nor UO_2274 (O_2274,N_24939,N_24930);
xnor UO_2275 (O_2275,N_24917,N_24947);
xnor UO_2276 (O_2276,N_24868,N_24854);
or UO_2277 (O_2277,N_24949,N_24989);
xor UO_2278 (O_2278,N_24976,N_24896);
xnor UO_2279 (O_2279,N_24920,N_24905);
xor UO_2280 (O_2280,N_24816,N_24802);
nor UO_2281 (O_2281,N_24891,N_24918);
nand UO_2282 (O_2282,N_24960,N_24838);
and UO_2283 (O_2283,N_24953,N_24892);
nor UO_2284 (O_2284,N_24844,N_24804);
nor UO_2285 (O_2285,N_24968,N_24902);
nor UO_2286 (O_2286,N_24907,N_24971);
nand UO_2287 (O_2287,N_24987,N_24870);
or UO_2288 (O_2288,N_24839,N_24806);
and UO_2289 (O_2289,N_24921,N_24832);
or UO_2290 (O_2290,N_24936,N_24832);
nand UO_2291 (O_2291,N_24956,N_24817);
nor UO_2292 (O_2292,N_24914,N_24970);
or UO_2293 (O_2293,N_24932,N_24978);
nand UO_2294 (O_2294,N_24851,N_24963);
nor UO_2295 (O_2295,N_24828,N_24856);
nor UO_2296 (O_2296,N_24920,N_24900);
or UO_2297 (O_2297,N_24918,N_24859);
or UO_2298 (O_2298,N_24888,N_24843);
xnor UO_2299 (O_2299,N_24813,N_24837);
nor UO_2300 (O_2300,N_24981,N_24999);
nor UO_2301 (O_2301,N_24889,N_24949);
or UO_2302 (O_2302,N_24937,N_24812);
nor UO_2303 (O_2303,N_24928,N_24878);
xor UO_2304 (O_2304,N_24935,N_24889);
nand UO_2305 (O_2305,N_24804,N_24951);
xnor UO_2306 (O_2306,N_24856,N_24911);
and UO_2307 (O_2307,N_24968,N_24931);
nor UO_2308 (O_2308,N_24851,N_24880);
nand UO_2309 (O_2309,N_24877,N_24944);
xnor UO_2310 (O_2310,N_24883,N_24819);
and UO_2311 (O_2311,N_24966,N_24881);
xor UO_2312 (O_2312,N_24859,N_24848);
xnor UO_2313 (O_2313,N_24855,N_24869);
nor UO_2314 (O_2314,N_24854,N_24814);
and UO_2315 (O_2315,N_24964,N_24968);
nor UO_2316 (O_2316,N_24817,N_24988);
and UO_2317 (O_2317,N_24959,N_24852);
xnor UO_2318 (O_2318,N_24917,N_24863);
and UO_2319 (O_2319,N_24843,N_24837);
nor UO_2320 (O_2320,N_24866,N_24946);
or UO_2321 (O_2321,N_24803,N_24848);
xor UO_2322 (O_2322,N_24882,N_24925);
and UO_2323 (O_2323,N_24868,N_24951);
xnor UO_2324 (O_2324,N_24872,N_24982);
and UO_2325 (O_2325,N_24997,N_24894);
nand UO_2326 (O_2326,N_24970,N_24863);
nand UO_2327 (O_2327,N_24890,N_24895);
nor UO_2328 (O_2328,N_24814,N_24899);
or UO_2329 (O_2329,N_24932,N_24996);
or UO_2330 (O_2330,N_24903,N_24979);
and UO_2331 (O_2331,N_24858,N_24909);
or UO_2332 (O_2332,N_24996,N_24924);
and UO_2333 (O_2333,N_24829,N_24813);
and UO_2334 (O_2334,N_24965,N_24847);
nor UO_2335 (O_2335,N_24982,N_24951);
and UO_2336 (O_2336,N_24845,N_24873);
nor UO_2337 (O_2337,N_24951,N_24905);
or UO_2338 (O_2338,N_24936,N_24820);
xnor UO_2339 (O_2339,N_24832,N_24964);
nand UO_2340 (O_2340,N_24920,N_24853);
nor UO_2341 (O_2341,N_24883,N_24843);
nand UO_2342 (O_2342,N_24914,N_24848);
nand UO_2343 (O_2343,N_24972,N_24855);
nor UO_2344 (O_2344,N_24919,N_24800);
or UO_2345 (O_2345,N_24829,N_24948);
nand UO_2346 (O_2346,N_24856,N_24849);
and UO_2347 (O_2347,N_24950,N_24910);
xnor UO_2348 (O_2348,N_24834,N_24894);
nand UO_2349 (O_2349,N_24931,N_24958);
and UO_2350 (O_2350,N_24930,N_24899);
and UO_2351 (O_2351,N_24860,N_24844);
xor UO_2352 (O_2352,N_24949,N_24860);
or UO_2353 (O_2353,N_24959,N_24836);
nand UO_2354 (O_2354,N_24908,N_24891);
and UO_2355 (O_2355,N_24848,N_24868);
nand UO_2356 (O_2356,N_24831,N_24910);
nor UO_2357 (O_2357,N_24963,N_24809);
xnor UO_2358 (O_2358,N_24973,N_24930);
nand UO_2359 (O_2359,N_24937,N_24815);
or UO_2360 (O_2360,N_24841,N_24998);
or UO_2361 (O_2361,N_24834,N_24845);
xor UO_2362 (O_2362,N_24935,N_24916);
or UO_2363 (O_2363,N_24887,N_24926);
or UO_2364 (O_2364,N_24961,N_24837);
xor UO_2365 (O_2365,N_24988,N_24888);
nor UO_2366 (O_2366,N_24800,N_24871);
or UO_2367 (O_2367,N_24908,N_24988);
and UO_2368 (O_2368,N_24945,N_24818);
xor UO_2369 (O_2369,N_24809,N_24977);
nor UO_2370 (O_2370,N_24932,N_24988);
nand UO_2371 (O_2371,N_24901,N_24897);
nor UO_2372 (O_2372,N_24986,N_24974);
xnor UO_2373 (O_2373,N_24980,N_24948);
xnor UO_2374 (O_2374,N_24952,N_24916);
nor UO_2375 (O_2375,N_24839,N_24816);
and UO_2376 (O_2376,N_24950,N_24933);
nor UO_2377 (O_2377,N_24929,N_24871);
nor UO_2378 (O_2378,N_24838,N_24849);
or UO_2379 (O_2379,N_24884,N_24979);
or UO_2380 (O_2380,N_24910,N_24817);
and UO_2381 (O_2381,N_24882,N_24926);
nor UO_2382 (O_2382,N_24819,N_24979);
or UO_2383 (O_2383,N_24920,N_24874);
and UO_2384 (O_2384,N_24909,N_24914);
xor UO_2385 (O_2385,N_24889,N_24901);
nand UO_2386 (O_2386,N_24933,N_24956);
and UO_2387 (O_2387,N_24895,N_24944);
and UO_2388 (O_2388,N_24841,N_24812);
xnor UO_2389 (O_2389,N_24908,N_24841);
xnor UO_2390 (O_2390,N_24991,N_24979);
nor UO_2391 (O_2391,N_24890,N_24807);
nand UO_2392 (O_2392,N_24916,N_24841);
or UO_2393 (O_2393,N_24995,N_24819);
nor UO_2394 (O_2394,N_24809,N_24802);
xor UO_2395 (O_2395,N_24969,N_24816);
nand UO_2396 (O_2396,N_24996,N_24860);
or UO_2397 (O_2397,N_24809,N_24981);
or UO_2398 (O_2398,N_24929,N_24888);
xnor UO_2399 (O_2399,N_24947,N_24816);
and UO_2400 (O_2400,N_24988,N_24945);
and UO_2401 (O_2401,N_24973,N_24843);
nand UO_2402 (O_2402,N_24981,N_24919);
or UO_2403 (O_2403,N_24898,N_24940);
nor UO_2404 (O_2404,N_24959,N_24832);
and UO_2405 (O_2405,N_24828,N_24999);
xnor UO_2406 (O_2406,N_24802,N_24968);
nor UO_2407 (O_2407,N_24979,N_24853);
or UO_2408 (O_2408,N_24960,N_24931);
or UO_2409 (O_2409,N_24826,N_24949);
nor UO_2410 (O_2410,N_24953,N_24974);
nand UO_2411 (O_2411,N_24823,N_24977);
nor UO_2412 (O_2412,N_24805,N_24837);
nor UO_2413 (O_2413,N_24893,N_24848);
nor UO_2414 (O_2414,N_24814,N_24864);
nand UO_2415 (O_2415,N_24905,N_24972);
and UO_2416 (O_2416,N_24870,N_24879);
nor UO_2417 (O_2417,N_24800,N_24923);
or UO_2418 (O_2418,N_24923,N_24826);
nor UO_2419 (O_2419,N_24815,N_24977);
xor UO_2420 (O_2420,N_24873,N_24807);
nand UO_2421 (O_2421,N_24911,N_24930);
nand UO_2422 (O_2422,N_24881,N_24940);
nor UO_2423 (O_2423,N_24982,N_24919);
or UO_2424 (O_2424,N_24938,N_24835);
nand UO_2425 (O_2425,N_24814,N_24926);
or UO_2426 (O_2426,N_24804,N_24969);
or UO_2427 (O_2427,N_24863,N_24999);
nand UO_2428 (O_2428,N_24889,N_24815);
xor UO_2429 (O_2429,N_24806,N_24898);
xor UO_2430 (O_2430,N_24987,N_24952);
xnor UO_2431 (O_2431,N_24939,N_24807);
nor UO_2432 (O_2432,N_24987,N_24841);
and UO_2433 (O_2433,N_24998,N_24896);
xnor UO_2434 (O_2434,N_24871,N_24899);
and UO_2435 (O_2435,N_24925,N_24846);
and UO_2436 (O_2436,N_24853,N_24997);
nand UO_2437 (O_2437,N_24977,N_24865);
xor UO_2438 (O_2438,N_24917,N_24812);
or UO_2439 (O_2439,N_24896,N_24950);
nand UO_2440 (O_2440,N_24972,N_24879);
and UO_2441 (O_2441,N_24932,N_24935);
nor UO_2442 (O_2442,N_24907,N_24934);
nand UO_2443 (O_2443,N_24892,N_24973);
xor UO_2444 (O_2444,N_24920,N_24907);
nor UO_2445 (O_2445,N_24960,N_24995);
nand UO_2446 (O_2446,N_24998,N_24997);
and UO_2447 (O_2447,N_24906,N_24822);
or UO_2448 (O_2448,N_24997,N_24900);
or UO_2449 (O_2449,N_24818,N_24954);
xnor UO_2450 (O_2450,N_24917,N_24969);
and UO_2451 (O_2451,N_24944,N_24972);
or UO_2452 (O_2452,N_24907,N_24843);
nand UO_2453 (O_2453,N_24903,N_24945);
nor UO_2454 (O_2454,N_24888,N_24865);
nor UO_2455 (O_2455,N_24953,N_24837);
nand UO_2456 (O_2456,N_24891,N_24882);
nand UO_2457 (O_2457,N_24897,N_24949);
xnor UO_2458 (O_2458,N_24943,N_24873);
and UO_2459 (O_2459,N_24882,N_24915);
or UO_2460 (O_2460,N_24974,N_24836);
or UO_2461 (O_2461,N_24944,N_24814);
xnor UO_2462 (O_2462,N_24994,N_24895);
nand UO_2463 (O_2463,N_24888,N_24800);
xnor UO_2464 (O_2464,N_24815,N_24846);
nor UO_2465 (O_2465,N_24827,N_24950);
or UO_2466 (O_2466,N_24982,N_24980);
xor UO_2467 (O_2467,N_24802,N_24960);
or UO_2468 (O_2468,N_24870,N_24983);
nor UO_2469 (O_2469,N_24952,N_24813);
nor UO_2470 (O_2470,N_24947,N_24918);
nand UO_2471 (O_2471,N_24910,N_24866);
nand UO_2472 (O_2472,N_24814,N_24818);
or UO_2473 (O_2473,N_24991,N_24857);
nand UO_2474 (O_2474,N_24939,N_24831);
and UO_2475 (O_2475,N_24924,N_24955);
nand UO_2476 (O_2476,N_24930,N_24946);
xnor UO_2477 (O_2477,N_24972,N_24993);
and UO_2478 (O_2478,N_24902,N_24800);
nor UO_2479 (O_2479,N_24923,N_24951);
nor UO_2480 (O_2480,N_24962,N_24813);
and UO_2481 (O_2481,N_24932,N_24916);
nor UO_2482 (O_2482,N_24819,N_24902);
nor UO_2483 (O_2483,N_24934,N_24822);
and UO_2484 (O_2484,N_24882,N_24848);
and UO_2485 (O_2485,N_24929,N_24917);
xor UO_2486 (O_2486,N_24967,N_24966);
and UO_2487 (O_2487,N_24850,N_24872);
or UO_2488 (O_2488,N_24917,N_24995);
nand UO_2489 (O_2489,N_24990,N_24808);
and UO_2490 (O_2490,N_24981,N_24963);
xor UO_2491 (O_2491,N_24941,N_24931);
and UO_2492 (O_2492,N_24916,N_24968);
nand UO_2493 (O_2493,N_24809,N_24852);
or UO_2494 (O_2494,N_24895,N_24909);
nand UO_2495 (O_2495,N_24942,N_24928);
xnor UO_2496 (O_2496,N_24855,N_24948);
xnor UO_2497 (O_2497,N_24824,N_24905);
and UO_2498 (O_2498,N_24914,N_24935);
xnor UO_2499 (O_2499,N_24804,N_24999);
nor UO_2500 (O_2500,N_24976,N_24817);
nor UO_2501 (O_2501,N_24994,N_24838);
or UO_2502 (O_2502,N_24997,N_24955);
nor UO_2503 (O_2503,N_24878,N_24869);
xor UO_2504 (O_2504,N_24964,N_24840);
and UO_2505 (O_2505,N_24977,N_24952);
nor UO_2506 (O_2506,N_24956,N_24939);
nor UO_2507 (O_2507,N_24821,N_24885);
nor UO_2508 (O_2508,N_24915,N_24805);
nor UO_2509 (O_2509,N_24924,N_24902);
xor UO_2510 (O_2510,N_24908,N_24914);
or UO_2511 (O_2511,N_24909,N_24892);
xnor UO_2512 (O_2512,N_24927,N_24853);
or UO_2513 (O_2513,N_24949,N_24875);
nor UO_2514 (O_2514,N_24908,N_24940);
nand UO_2515 (O_2515,N_24955,N_24916);
and UO_2516 (O_2516,N_24985,N_24961);
nor UO_2517 (O_2517,N_24822,N_24839);
and UO_2518 (O_2518,N_24879,N_24821);
nor UO_2519 (O_2519,N_24991,N_24922);
nor UO_2520 (O_2520,N_24823,N_24941);
nand UO_2521 (O_2521,N_24917,N_24909);
xnor UO_2522 (O_2522,N_24891,N_24977);
nor UO_2523 (O_2523,N_24985,N_24965);
xor UO_2524 (O_2524,N_24978,N_24915);
or UO_2525 (O_2525,N_24824,N_24891);
nand UO_2526 (O_2526,N_24890,N_24955);
or UO_2527 (O_2527,N_24830,N_24928);
or UO_2528 (O_2528,N_24815,N_24960);
and UO_2529 (O_2529,N_24878,N_24805);
xor UO_2530 (O_2530,N_24885,N_24837);
and UO_2531 (O_2531,N_24891,N_24946);
or UO_2532 (O_2532,N_24931,N_24839);
xor UO_2533 (O_2533,N_24946,N_24981);
nand UO_2534 (O_2534,N_24919,N_24914);
xor UO_2535 (O_2535,N_24859,N_24873);
xnor UO_2536 (O_2536,N_24881,N_24978);
nor UO_2537 (O_2537,N_24822,N_24829);
xor UO_2538 (O_2538,N_24987,N_24981);
and UO_2539 (O_2539,N_24834,N_24945);
nand UO_2540 (O_2540,N_24940,N_24875);
nor UO_2541 (O_2541,N_24845,N_24824);
or UO_2542 (O_2542,N_24921,N_24974);
nor UO_2543 (O_2543,N_24961,N_24889);
nand UO_2544 (O_2544,N_24895,N_24836);
nand UO_2545 (O_2545,N_24937,N_24842);
nand UO_2546 (O_2546,N_24981,N_24969);
nand UO_2547 (O_2547,N_24864,N_24868);
and UO_2548 (O_2548,N_24974,N_24801);
nand UO_2549 (O_2549,N_24956,N_24974);
nand UO_2550 (O_2550,N_24974,N_24891);
nor UO_2551 (O_2551,N_24832,N_24853);
and UO_2552 (O_2552,N_24960,N_24986);
and UO_2553 (O_2553,N_24861,N_24807);
nand UO_2554 (O_2554,N_24972,N_24811);
nand UO_2555 (O_2555,N_24985,N_24814);
nor UO_2556 (O_2556,N_24868,N_24847);
nor UO_2557 (O_2557,N_24876,N_24940);
nand UO_2558 (O_2558,N_24860,N_24807);
or UO_2559 (O_2559,N_24965,N_24993);
nand UO_2560 (O_2560,N_24879,N_24995);
and UO_2561 (O_2561,N_24953,N_24904);
nor UO_2562 (O_2562,N_24825,N_24807);
and UO_2563 (O_2563,N_24886,N_24973);
xor UO_2564 (O_2564,N_24874,N_24872);
nor UO_2565 (O_2565,N_24951,N_24824);
nand UO_2566 (O_2566,N_24911,N_24875);
or UO_2567 (O_2567,N_24961,N_24892);
and UO_2568 (O_2568,N_24984,N_24988);
nor UO_2569 (O_2569,N_24822,N_24870);
and UO_2570 (O_2570,N_24844,N_24843);
or UO_2571 (O_2571,N_24944,N_24802);
nand UO_2572 (O_2572,N_24892,N_24907);
and UO_2573 (O_2573,N_24851,N_24983);
nor UO_2574 (O_2574,N_24965,N_24944);
nand UO_2575 (O_2575,N_24907,N_24867);
xor UO_2576 (O_2576,N_24882,N_24979);
xor UO_2577 (O_2577,N_24960,N_24914);
nand UO_2578 (O_2578,N_24826,N_24916);
or UO_2579 (O_2579,N_24854,N_24947);
xnor UO_2580 (O_2580,N_24809,N_24868);
nand UO_2581 (O_2581,N_24898,N_24952);
xnor UO_2582 (O_2582,N_24986,N_24957);
nor UO_2583 (O_2583,N_24938,N_24830);
nand UO_2584 (O_2584,N_24953,N_24869);
nand UO_2585 (O_2585,N_24808,N_24833);
or UO_2586 (O_2586,N_24902,N_24858);
nor UO_2587 (O_2587,N_24900,N_24807);
nor UO_2588 (O_2588,N_24867,N_24878);
nor UO_2589 (O_2589,N_24939,N_24945);
xor UO_2590 (O_2590,N_24948,N_24806);
nor UO_2591 (O_2591,N_24869,N_24852);
or UO_2592 (O_2592,N_24830,N_24936);
nand UO_2593 (O_2593,N_24916,N_24884);
or UO_2594 (O_2594,N_24817,N_24855);
or UO_2595 (O_2595,N_24881,N_24885);
nand UO_2596 (O_2596,N_24917,N_24870);
xor UO_2597 (O_2597,N_24803,N_24942);
nor UO_2598 (O_2598,N_24861,N_24939);
and UO_2599 (O_2599,N_24840,N_24863);
nor UO_2600 (O_2600,N_24800,N_24873);
or UO_2601 (O_2601,N_24938,N_24853);
and UO_2602 (O_2602,N_24868,N_24832);
and UO_2603 (O_2603,N_24874,N_24990);
nor UO_2604 (O_2604,N_24952,N_24980);
or UO_2605 (O_2605,N_24805,N_24977);
nand UO_2606 (O_2606,N_24966,N_24924);
and UO_2607 (O_2607,N_24879,N_24867);
nor UO_2608 (O_2608,N_24826,N_24801);
nand UO_2609 (O_2609,N_24993,N_24912);
and UO_2610 (O_2610,N_24910,N_24815);
nor UO_2611 (O_2611,N_24907,N_24803);
nand UO_2612 (O_2612,N_24965,N_24833);
or UO_2613 (O_2613,N_24856,N_24844);
or UO_2614 (O_2614,N_24968,N_24926);
or UO_2615 (O_2615,N_24818,N_24805);
nand UO_2616 (O_2616,N_24957,N_24973);
or UO_2617 (O_2617,N_24853,N_24840);
nor UO_2618 (O_2618,N_24856,N_24822);
nor UO_2619 (O_2619,N_24907,N_24993);
or UO_2620 (O_2620,N_24964,N_24846);
or UO_2621 (O_2621,N_24811,N_24923);
or UO_2622 (O_2622,N_24895,N_24929);
xnor UO_2623 (O_2623,N_24983,N_24972);
nor UO_2624 (O_2624,N_24878,N_24993);
nor UO_2625 (O_2625,N_24941,N_24946);
xor UO_2626 (O_2626,N_24926,N_24886);
nor UO_2627 (O_2627,N_24854,N_24844);
nand UO_2628 (O_2628,N_24973,N_24963);
nor UO_2629 (O_2629,N_24890,N_24952);
nor UO_2630 (O_2630,N_24898,N_24881);
or UO_2631 (O_2631,N_24824,N_24855);
nand UO_2632 (O_2632,N_24915,N_24865);
nand UO_2633 (O_2633,N_24834,N_24922);
or UO_2634 (O_2634,N_24894,N_24904);
nor UO_2635 (O_2635,N_24913,N_24988);
nand UO_2636 (O_2636,N_24951,N_24827);
nor UO_2637 (O_2637,N_24902,N_24827);
nand UO_2638 (O_2638,N_24927,N_24955);
and UO_2639 (O_2639,N_24972,N_24906);
nand UO_2640 (O_2640,N_24958,N_24856);
xor UO_2641 (O_2641,N_24999,N_24854);
nand UO_2642 (O_2642,N_24977,N_24850);
nand UO_2643 (O_2643,N_24955,N_24858);
and UO_2644 (O_2644,N_24945,N_24915);
and UO_2645 (O_2645,N_24977,N_24937);
nand UO_2646 (O_2646,N_24943,N_24957);
or UO_2647 (O_2647,N_24900,N_24937);
nand UO_2648 (O_2648,N_24819,N_24861);
xnor UO_2649 (O_2649,N_24928,N_24869);
or UO_2650 (O_2650,N_24988,N_24966);
nor UO_2651 (O_2651,N_24877,N_24861);
and UO_2652 (O_2652,N_24979,N_24870);
or UO_2653 (O_2653,N_24830,N_24875);
and UO_2654 (O_2654,N_24831,N_24815);
and UO_2655 (O_2655,N_24953,N_24957);
and UO_2656 (O_2656,N_24953,N_24969);
or UO_2657 (O_2657,N_24922,N_24820);
xor UO_2658 (O_2658,N_24847,N_24892);
nand UO_2659 (O_2659,N_24854,N_24933);
xor UO_2660 (O_2660,N_24832,N_24932);
or UO_2661 (O_2661,N_24822,N_24980);
nor UO_2662 (O_2662,N_24902,N_24997);
nand UO_2663 (O_2663,N_24953,N_24901);
or UO_2664 (O_2664,N_24895,N_24963);
or UO_2665 (O_2665,N_24965,N_24845);
and UO_2666 (O_2666,N_24837,N_24988);
nor UO_2667 (O_2667,N_24974,N_24860);
nor UO_2668 (O_2668,N_24927,N_24973);
nor UO_2669 (O_2669,N_24961,N_24802);
and UO_2670 (O_2670,N_24903,N_24847);
nand UO_2671 (O_2671,N_24905,N_24872);
and UO_2672 (O_2672,N_24969,N_24871);
xnor UO_2673 (O_2673,N_24842,N_24954);
and UO_2674 (O_2674,N_24975,N_24882);
xnor UO_2675 (O_2675,N_24872,N_24888);
xnor UO_2676 (O_2676,N_24810,N_24875);
xor UO_2677 (O_2677,N_24970,N_24973);
or UO_2678 (O_2678,N_24985,N_24940);
xnor UO_2679 (O_2679,N_24978,N_24981);
and UO_2680 (O_2680,N_24817,N_24996);
xor UO_2681 (O_2681,N_24849,N_24932);
nand UO_2682 (O_2682,N_24806,N_24955);
xnor UO_2683 (O_2683,N_24804,N_24963);
xnor UO_2684 (O_2684,N_24862,N_24878);
or UO_2685 (O_2685,N_24860,N_24899);
and UO_2686 (O_2686,N_24807,N_24820);
xnor UO_2687 (O_2687,N_24976,N_24855);
or UO_2688 (O_2688,N_24879,N_24863);
xnor UO_2689 (O_2689,N_24835,N_24816);
nor UO_2690 (O_2690,N_24915,N_24924);
or UO_2691 (O_2691,N_24833,N_24926);
nand UO_2692 (O_2692,N_24876,N_24885);
and UO_2693 (O_2693,N_24963,N_24821);
nand UO_2694 (O_2694,N_24884,N_24907);
nor UO_2695 (O_2695,N_24848,N_24806);
or UO_2696 (O_2696,N_24991,N_24913);
and UO_2697 (O_2697,N_24890,N_24825);
nor UO_2698 (O_2698,N_24957,N_24863);
or UO_2699 (O_2699,N_24873,N_24801);
xnor UO_2700 (O_2700,N_24887,N_24920);
or UO_2701 (O_2701,N_24889,N_24812);
and UO_2702 (O_2702,N_24908,N_24830);
xnor UO_2703 (O_2703,N_24811,N_24866);
nand UO_2704 (O_2704,N_24973,N_24820);
and UO_2705 (O_2705,N_24903,N_24830);
xor UO_2706 (O_2706,N_24825,N_24872);
or UO_2707 (O_2707,N_24995,N_24967);
nand UO_2708 (O_2708,N_24954,N_24984);
nor UO_2709 (O_2709,N_24974,N_24835);
xor UO_2710 (O_2710,N_24811,N_24997);
xor UO_2711 (O_2711,N_24870,N_24954);
or UO_2712 (O_2712,N_24976,N_24994);
or UO_2713 (O_2713,N_24968,N_24853);
or UO_2714 (O_2714,N_24846,N_24923);
and UO_2715 (O_2715,N_24982,N_24870);
and UO_2716 (O_2716,N_24982,N_24861);
nor UO_2717 (O_2717,N_24961,N_24938);
and UO_2718 (O_2718,N_24872,N_24824);
xor UO_2719 (O_2719,N_24940,N_24843);
nor UO_2720 (O_2720,N_24833,N_24905);
or UO_2721 (O_2721,N_24946,N_24968);
nand UO_2722 (O_2722,N_24929,N_24872);
xnor UO_2723 (O_2723,N_24903,N_24985);
or UO_2724 (O_2724,N_24939,N_24979);
nand UO_2725 (O_2725,N_24954,N_24965);
or UO_2726 (O_2726,N_24834,N_24967);
and UO_2727 (O_2727,N_24942,N_24936);
nor UO_2728 (O_2728,N_24868,N_24967);
and UO_2729 (O_2729,N_24891,N_24973);
nand UO_2730 (O_2730,N_24870,N_24846);
nand UO_2731 (O_2731,N_24803,N_24987);
xor UO_2732 (O_2732,N_24996,N_24975);
and UO_2733 (O_2733,N_24823,N_24964);
and UO_2734 (O_2734,N_24986,N_24978);
nand UO_2735 (O_2735,N_24826,N_24958);
xnor UO_2736 (O_2736,N_24971,N_24919);
nand UO_2737 (O_2737,N_24903,N_24873);
and UO_2738 (O_2738,N_24884,N_24919);
xor UO_2739 (O_2739,N_24929,N_24988);
and UO_2740 (O_2740,N_24815,N_24842);
nand UO_2741 (O_2741,N_24957,N_24860);
and UO_2742 (O_2742,N_24885,N_24958);
xnor UO_2743 (O_2743,N_24882,N_24872);
nand UO_2744 (O_2744,N_24814,N_24915);
and UO_2745 (O_2745,N_24837,N_24846);
xor UO_2746 (O_2746,N_24859,N_24828);
nor UO_2747 (O_2747,N_24833,N_24959);
or UO_2748 (O_2748,N_24897,N_24976);
nand UO_2749 (O_2749,N_24934,N_24856);
and UO_2750 (O_2750,N_24875,N_24990);
and UO_2751 (O_2751,N_24881,N_24915);
and UO_2752 (O_2752,N_24839,N_24969);
xor UO_2753 (O_2753,N_24903,N_24834);
nand UO_2754 (O_2754,N_24815,N_24916);
nor UO_2755 (O_2755,N_24900,N_24938);
and UO_2756 (O_2756,N_24828,N_24872);
and UO_2757 (O_2757,N_24939,N_24854);
or UO_2758 (O_2758,N_24985,N_24895);
and UO_2759 (O_2759,N_24923,N_24954);
nand UO_2760 (O_2760,N_24811,N_24870);
nor UO_2761 (O_2761,N_24830,N_24825);
nor UO_2762 (O_2762,N_24832,N_24949);
nand UO_2763 (O_2763,N_24923,N_24828);
nor UO_2764 (O_2764,N_24867,N_24945);
xor UO_2765 (O_2765,N_24977,N_24869);
nor UO_2766 (O_2766,N_24812,N_24805);
xnor UO_2767 (O_2767,N_24995,N_24876);
xnor UO_2768 (O_2768,N_24985,N_24999);
nor UO_2769 (O_2769,N_24847,N_24819);
xnor UO_2770 (O_2770,N_24948,N_24842);
or UO_2771 (O_2771,N_24946,N_24852);
and UO_2772 (O_2772,N_24867,N_24993);
and UO_2773 (O_2773,N_24956,N_24863);
xor UO_2774 (O_2774,N_24857,N_24820);
and UO_2775 (O_2775,N_24864,N_24818);
nor UO_2776 (O_2776,N_24804,N_24807);
nor UO_2777 (O_2777,N_24827,N_24945);
nand UO_2778 (O_2778,N_24964,N_24817);
xor UO_2779 (O_2779,N_24993,N_24847);
or UO_2780 (O_2780,N_24903,N_24958);
nor UO_2781 (O_2781,N_24853,N_24851);
nand UO_2782 (O_2782,N_24902,N_24812);
nand UO_2783 (O_2783,N_24876,N_24986);
nand UO_2784 (O_2784,N_24961,N_24930);
nor UO_2785 (O_2785,N_24938,N_24859);
or UO_2786 (O_2786,N_24987,N_24913);
nand UO_2787 (O_2787,N_24980,N_24967);
xor UO_2788 (O_2788,N_24860,N_24863);
nand UO_2789 (O_2789,N_24897,N_24846);
xnor UO_2790 (O_2790,N_24999,N_24889);
and UO_2791 (O_2791,N_24844,N_24999);
nor UO_2792 (O_2792,N_24861,N_24849);
nand UO_2793 (O_2793,N_24895,N_24864);
and UO_2794 (O_2794,N_24946,N_24893);
and UO_2795 (O_2795,N_24928,N_24980);
nand UO_2796 (O_2796,N_24965,N_24953);
nor UO_2797 (O_2797,N_24836,N_24867);
xnor UO_2798 (O_2798,N_24906,N_24899);
nand UO_2799 (O_2799,N_24912,N_24919);
and UO_2800 (O_2800,N_24821,N_24911);
xnor UO_2801 (O_2801,N_24856,N_24831);
and UO_2802 (O_2802,N_24964,N_24830);
xnor UO_2803 (O_2803,N_24809,N_24991);
nand UO_2804 (O_2804,N_24882,N_24972);
or UO_2805 (O_2805,N_24813,N_24835);
xnor UO_2806 (O_2806,N_24845,N_24990);
nor UO_2807 (O_2807,N_24815,N_24983);
and UO_2808 (O_2808,N_24977,N_24814);
or UO_2809 (O_2809,N_24904,N_24817);
or UO_2810 (O_2810,N_24888,N_24842);
and UO_2811 (O_2811,N_24903,N_24810);
or UO_2812 (O_2812,N_24850,N_24814);
xor UO_2813 (O_2813,N_24899,N_24940);
or UO_2814 (O_2814,N_24937,N_24831);
or UO_2815 (O_2815,N_24851,N_24891);
or UO_2816 (O_2816,N_24878,N_24879);
and UO_2817 (O_2817,N_24817,N_24918);
and UO_2818 (O_2818,N_24935,N_24839);
or UO_2819 (O_2819,N_24825,N_24826);
nand UO_2820 (O_2820,N_24842,N_24917);
xor UO_2821 (O_2821,N_24922,N_24886);
or UO_2822 (O_2822,N_24879,N_24928);
nand UO_2823 (O_2823,N_24874,N_24945);
or UO_2824 (O_2824,N_24921,N_24940);
xnor UO_2825 (O_2825,N_24935,N_24974);
xor UO_2826 (O_2826,N_24871,N_24983);
xnor UO_2827 (O_2827,N_24976,N_24907);
nor UO_2828 (O_2828,N_24932,N_24917);
nand UO_2829 (O_2829,N_24911,N_24855);
xnor UO_2830 (O_2830,N_24993,N_24942);
nand UO_2831 (O_2831,N_24827,N_24896);
nor UO_2832 (O_2832,N_24918,N_24865);
nor UO_2833 (O_2833,N_24910,N_24923);
xor UO_2834 (O_2834,N_24991,N_24888);
and UO_2835 (O_2835,N_24859,N_24945);
or UO_2836 (O_2836,N_24813,N_24960);
nand UO_2837 (O_2837,N_24831,N_24801);
or UO_2838 (O_2838,N_24868,N_24973);
nand UO_2839 (O_2839,N_24984,N_24833);
and UO_2840 (O_2840,N_24828,N_24806);
and UO_2841 (O_2841,N_24984,N_24807);
xnor UO_2842 (O_2842,N_24868,N_24826);
xor UO_2843 (O_2843,N_24893,N_24942);
nor UO_2844 (O_2844,N_24823,N_24913);
and UO_2845 (O_2845,N_24821,N_24957);
nand UO_2846 (O_2846,N_24923,N_24841);
xor UO_2847 (O_2847,N_24979,N_24887);
nor UO_2848 (O_2848,N_24855,N_24830);
xor UO_2849 (O_2849,N_24962,N_24991);
and UO_2850 (O_2850,N_24871,N_24872);
xnor UO_2851 (O_2851,N_24834,N_24916);
or UO_2852 (O_2852,N_24829,N_24875);
nor UO_2853 (O_2853,N_24958,N_24887);
or UO_2854 (O_2854,N_24945,N_24936);
or UO_2855 (O_2855,N_24934,N_24868);
nand UO_2856 (O_2856,N_24896,N_24830);
or UO_2857 (O_2857,N_24922,N_24832);
nand UO_2858 (O_2858,N_24929,N_24894);
or UO_2859 (O_2859,N_24821,N_24968);
nor UO_2860 (O_2860,N_24889,N_24972);
nand UO_2861 (O_2861,N_24915,N_24919);
nand UO_2862 (O_2862,N_24851,N_24987);
and UO_2863 (O_2863,N_24806,N_24981);
xor UO_2864 (O_2864,N_24985,N_24830);
and UO_2865 (O_2865,N_24866,N_24940);
xnor UO_2866 (O_2866,N_24849,N_24964);
nor UO_2867 (O_2867,N_24850,N_24953);
nand UO_2868 (O_2868,N_24978,N_24821);
and UO_2869 (O_2869,N_24952,N_24861);
xor UO_2870 (O_2870,N_24972,N_24950);
nand UO_2871 (O_2871,N_24880,N_24814);
nand UO_2872 (O_2872,N_24875,N_24824);
or UO_2873 (O_2873,N_24814,N_24870);
nand UO_2874 (O_2874,N_24951,N_24959);
nor UO_2875 (O_2875,N_24950,N_24962);
and UO_2876 (O_2876,N_24825,N_24880);
and UO_2877 (O_2877,N_24941,N_24921);
and UO_2878 (O_2878,N_24981,N_24955);
xor UO_2879 (O_2879,N_24907,N_24986);
or UO_2880 (O_2880,N_24929,N_24898);
nor UO_2881 (O_2881,N_24901,N_24950);
and UO_2882 (O_2882,N_24854,N_24900);
and UO_2883 (O_2883,N_24867,N_24921);
or UO_2884 (O_2884,N_24857,N_24880);
nor UO_2885 (O_2885,N_24975,N_24856);
xor UO_2886 (O_2886,N_24907,N_24982);
nand UO_2887 (O_2887,N_24917,N_24911);
and UO_2888 (O_2888,N_24971,N_24842);
and UO_2889 (O_2889,N_24994,N_24999);
nor UO_2890 (O_2890,N_24845,N_24997);
and UO_2891 (O_2891,N_24993,N_24869);
xor UO_2892 (O_2892,N_24958,N_24925);
nand UO_2893 (O_2893,N_24811,N_24887);
nor UO_2894 (O_2894,N_24947,N_24845);
or UO_2895 (O_2895,N_24951,N_24948);
nand UO_2896 (O_2896,N_24997,N_24892);
nor UO_2897 (O_2897,N_24914,N_24964);
or UO_2898 (O_2898,N_24847,N_24942);
nand UO_2899 (O_2899,N_24981,N_24829);
nand UO_2900 (O_2900,N_24803,N_24929);
nand UO_2901 (O_2901,N_24860,N_24956);
xnor UO_2902 (O_2902,N_24830,N_24978);
nand UO_2903 (O_2903,N_24866,N_24952);
or UO_2904 (O_2904,N_24938,N_24992);
nand UO_2905 (O_2905,N_24904,N_24875);
xor UO_2906 (O_2906,N_24820,N_24818);
and UO_2907 (O_2907,N_24964,N_24904);
xnor UO_2908 (O_2908,N_24929,N_24876);
xnor UO_2909 (O_2909,N_24829,N_24825);
and UO_2910 (O_2910,N_24868,N_24858);
and UO_2911 (O_2911,N_24804,N_24975);
nor UO_2912 (O_2912,N_24820,N_24811);
xnor UO_2913 (O_2913,N_24896,N_24958);
nor UO_2914 (O_2914,N_24943,N_24991);
nand UO_2915 (O_2915,N_24815,N_24968);
or UO_2916 (O_2916,N_24879,N_24953);
xor UO_2917 (O_2917,N_24969,N_24903);
or UO_2918 (O_2918,N_24859,N_24884);
and UO_2919 (O_2919,N_24960,N_24980);
xor UO_2920 (O_2920,N_24951,N_24922);
xor UO_2921 (O_2921,N_24949,N_24901);
xnor UO_2922 (O_2922,N_24878,N_24977);
or UO_2923 (O_2923,N_24867,N_24850);
nor UO_2924 (O_2924,N_24965,N_24895);
or UO_2925 (O_2925,N_24889,N_24926);
xor UO_2926 (O_2926,N_24968,N_24840);
nand UO_2927 (O_2927,N_24931,N_24984);
xnor UO_2928 (O_2928,N_24969,N_24932);
nand UO_2929 (O_2929,N_24858,N_24886);
xor UO_2930 (O_2930,N_24894,N_24973);
nand UO_2931 (O_2931,N_24857,N_24882);
or UO_2932 (O_2932,N_24835,N_24819);
and UO_2933 (O_2933,N_24807,N_24944);
or UO_2934 (O_2934,N_24871,N_24965);
xor UO_2935 (O_2935,N_24962,N_24897);
and UO_2936 (O_2936,N_24801,N_24901);
nand UO_2937 (O_2937,N_24963,N_24969);
xor UO_2938 (O_2938,N_24884,N_24810);
nand UO_2939 (O_2939,N_24938,N_24953);
xnor UO_2940 (O_2940,N_24991,N_24980);
and UO_2941 (O_2941,N_24922,N_24936);
xor UO_2942 (O_2942,N_24816,N_24892);
and UO_2943 (O_2943,N_24940,N_24894);
xnor UO_2944 (O_2944,N_24905,N_24954);
nand UO_2945 (O_2945,N_24926,N_24824);
nor UO_2946 (O_2946,N_24834,N_24860);
xor UO_2947 (O_2947,N_24936,N_24809);
and UO_2948 (O_2948,N_24985,N_24913);
and UO_2949 (O_2949,N_24947,N_24953);
nor UO_2950 (O_2950,N_24938,N_24809);
nand UO_2951 (O_2951,N_24870,N_24883);
nand UO_2952 (O_2952,N_24834,N_24803);
nor UO_2953 (O_2953,N_24837,N_24914);
and UO_2954 (O_2954,N_24983,N_24868);
nand UO_2955 (O_2955,N_24966,N_24953);
nor UO_2956 (O_2956,N_24982,N_24899);
nand UO_2957 (O_2957,N_24893,N_24865);
or UO_2958 (O_2958,N_24886,N_24801);
or UO_2959 (O_2959,N_24892,N_24869);
nand UO_2960 (O_2960,N_24808,N_24929);
xor UO_2961 (O_2961,N_24848,N_24860);
nor UO_2962 (O_2962,N_24827,N_24898);
or UO_2963 (O_2963,N_24910,N_24992);
nor UO_2964 (O_2964,N_24950,N_24934);
nor UO_2965 (O_2965,N_24962,N_24954);
xor UO_2966 (O_2966,N_24941,N_24868);
nand UO_2967 (O_2967,N_24826,N_24941);
and UO_2968 (O_2968,N_24908,N_24839);
nand UO_2969 (O_2969,N_24857,N_24851);
nand UO_2970 (O_2970,N_24936,N_24890);
or UO_2971 (O_2971,N_24913,N_24820);
or UO_2972 (O_2972,N_24921,N_24842);
or UO_2973 (O_2973,N_24902,N_24895);
or UO_2974 (O_2974,N_24851,N_24881);
or UO_2975 (O_2975,N_24981,N_24910);
xnor UO_2976 (O_2976,N_24992,N_24973);
or UO_2977 (O_2977,N_24964,N_24891);
or UO_2978 (O_2978,N_24877,N_24989);
or UO_2979 (O_2979,N_24971,N_24827);
xor UO_2980 (O_2980,N_24937,N_24850);
or UO_2981 (O_2981,N_24828,N_24926);
xor UO_2982 (O_2982,N_24895,N_24993);
and UO_2983 (O_2983,N_24906,N_24823);
nor UO_2984 (O_2984,N_24863,N_24872);
xnor UO_2985 (O_2985,N_24950,N_24871);
nor UO_2986 (O_2986,N_24847,N_24921);
nand UO_2987 (O_2987,N_24934,N_24806);
or UO_2988 (O_2988,N_24989,N_24827);
xnor UO_2989 (O_2989,N_24925,N_24837);
nand UO_2990 (O_2990,N_24943,N_24937);
and UO_2991 (O_2991,N_24849,N_24919);
and UO_2992 (O_2992,N_24973,N_24829);
xnor UO_2993 (O_2993,N_24837,N_24996);
and UO_2994 (O_2994,N_24939,N_24908);
xor UO_2995 (O_2995,N_24949,N_24950);
or UO_2996 (O_2996,N_24957,N_24929);
and UO_2997 (O_2997,N_24944,N_24900);
nor UO_2998 (O_2998,N_24985,N_24871);
nor UO_2999 (O_2999,N_24920,N_24925);
endmodule