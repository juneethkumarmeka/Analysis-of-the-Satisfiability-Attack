module basic_750_5000_1000_10_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_263,In_39);
nand U1 (N_1,In_139,In_492);
nor U2 (N_2,In_411,In_424);
and U3 (N_3,In_349,In_161);
xnor U4 (N_4,In_650,In_262);
nand U5 (N_5,In_515,In_249);
nand U6 (N_6,In_350,In_446);
nor U7 (N_7,In_380,In_385);
nor U8 (N_8,In_298,In_149);
and U9 (N_9,In_232,In_425);
xnor U10 (N_10,In_593,In_265);
or U11 (N_11,In_10,In_610);
nand U12 (N_12,In_18,In_16);
and U13 (N_13,In_189,In_62);
or U14 (N_14,In_444,In_697);
or U15 (N_15,In_173,In_412);
nand U16 (N_16,In_307,In_266);
nor U17 (N_17,In_540,In_333);
or U18 (N_18,In_735,In_745);
nand U19 (N_19,In_171,In_662);
or U20 (N_20,In_679,In_282);
nand U21 (N_21,In_562,In_337);
nand U22 (N_22,In_530,In_309);
and U23 (N_23,In_212,In_274);
nand U24 (N_24,In_533,In_12);
nand U25 (N_25,In_82,In_643);
and U26 (N_26,In_739,In_299);
or U27 (N_27,In_365,In_579);
xnor U28 (N_28,In_143,In_211);
nor U29 (N_29,In_419,In_4);
nand U30 (N_30,In_33,In_130);
or U31 (N_31,In_112,In_72);
xor U32 (N_32,In_291,In_378);
or U33 (N_33,In_475,In_723);
nor U34 (N_34,In_401,In_382);
and U35 (N_35,In_23,In_582);
or U36 (N_36,In_482,In_302);
or U37 (N_37,In_206,In_501);
or U38 (N_38,In_354,In_660);
nor U39 (N_39,In_158,In_633);
or U40 (N_40,In_221,In_596);
nand U41 (N_41,In_63,In_222);
and U42 (N_42,In_132,In_372);
or U43 (N_43,In_209,In_499);
or U44 (N_44,In_180,In_229);
and U45 (N_45,In_379,In_352);
nand U46 (N_46,In_199,In_243);
and U47 (N_47,In_652,In_67);
nor U48 (N_48,In_676,In_743);
and U49 (N_49,In_241,In_60);
nand U50 (N_50,In_418,In_702);
and U51 (N_51,In_340,In_258);
nand U52 (N_52,In_551,In_273);
or U53 (N_53,In_688,In_127);
nand U54 (N_54,In_603,In_664);
and U55 (N_55,In_584,In_122);
and U56 (N_56,In_50,In_268);
and U57 (N_57,In_54,In_387);
or U58 (N_58,In_100,In_97);
or U59 (N_59,In_430,In_503);
nor U60 (N_60,In_368,In_29);
nor U61 (N_61,In_71,In_493);
and U62 (N_62,In_187,In_434);
and U63 (N_63,In_597,In_172);
and U64 (N_64,In_733,In_137);
nand U65 (N_65,In_732,In_680);
and U66 (N_66,In_724,In_627);
nand U67 (N_67,In_629,In_160);
or U68 (N_68,In_271,In_134);
nor U69 (N_69,In_522,In_469);
xor U70 (N_70,In_518,In_741);
and U71 (N_71,In_369,In_509);
or U72 (N_72,In_543,In_423);
nor U73 (N_73,In_710,In_330);
and U74 (N_74,In_103,In_73);
nor U75 (N_75,In_449,In_635);
and U76 (N_76,In_438,In_384);
and U77 (N_77,In_729,In_92);
or U78 (N_78,In_601,In_686);
nor U79 (N_79,In_26,In_276);
nor U80 (N_80,In_396,In_460);
and U81 (N_81,In_315,In_96);
xnor U82 (N_82,In_539,In_52);
nor U83 (N_83,In_250,In_304);
or U84 (N_84,In_13,In_318);
nor U85 (N_85,In_604,In_175);
and U86 (N_86,In_3,In_389);
or U87 (N_87,In_79,In_140);
or U88 (N_88,In_86,In_57);
xnor U89 (N_89,In_420,In_131);
nor U90 (N_90,In_466,In_133);
and U91 (N_91,In_407,In_358);
and U92 (N_92,In_66,In_479);
nor U93 (N_93,In_14,In_388);
or U94 (N_94,In_485,In_605);
or U95 (N_95,In_145,In_677);
nor U96 (N_96,In_147,In_520);
xor U97 (N_97,In_747,In_740);
nor U98 (N_98,In_481,In_594);
or U99 (N_99,In_69,In_456);
or U100 (N_100,In_692,In_612);
xor U101 (N_101,In_484,In_355);
nand U102 (N_102,In_285,In_620);
and U103 (N_103,In_101,In_653);
nor U104 (N_104,In_671,In_431);
and U105 (N_105,In_667,In_259);
nor U106 (N_106,In_34,In_687);
nor U107 (N_107,In_359,In_181);
nor U108 (N_108,In_336,In_126);
nand U109 (N_109,In_663,In_666);
nand U110 (N_110,In_706,In_400);
and U111 (N_111,In_496,In_570);
nand U112 (N_112,In_617,In_178);
nor U113 (N_113,In_320,In_441);
xor U114 (N_114,In_670,In_526);
nor U115 (N_115,In_716,In_374);
and U116 (N_116,In_628,In_141);
nor U117 (N_117,In_641,In_339);
or U118 (N_118,In_672,In_203);
xor U119 (N_119,In_223,In_168);
or U120 (N_120,In_701,In_427);
nor U121 (N_121,In_87,In_480);
nand U122 (N_122,In_696,In_421);
nand U123 (N_123,In_689,In_47);
nand U124 (N_124,In_725,In_244);
nor U125 (N_125,In_346,In_587);
nor U126 (N_126,In_386,In_544);
and U127 (N_127,In_297,In_106);
xor U128 (N_128,In_397,In_437);
and U129 (N_129,In_529,In_393);
or U130 (N_130,In_452,In_550);
nand U131 (N_131,In_373,In_321);
or U132 (N_132,In_74,In_602);
nand U133 (N_133,In_744,In_528);
xnor U134 (N_134,In_279,In_281);
and U135 (N_135,In_685,In_693);
and U136 (N_136,In_213,In_534);
nor U137 (N_137,In_447,In_746);
xor U138 (N_138,In_415,In_366);
and U139 (N_139,In_476,In_43);
xor U140 (N_140,In_630,In_348);
xnor U141 (N_141,In_478,In_468);
nand U142 (N_142,In_30,In_600);
and U143 (N_143,In_6,In_606);
nor U144 (N_144,In_319,In_721);
or U145 (N_145,In_580,In_219);
nand U146 (N_146,In_714,In_237);
and U147 (N_147,In_704,In_457);
and U148 (N_148,In_519,In_571);
and U149 (N_149,In_516,In_370);
and U150 (N_150,In_264,In_375);
nor U151 (N_151,In_324,In_623);
and U152 (N_152,In_547,In_68);
or U153 (N_153,In_636,In_202);
nor U154 (N_154,In_713,In_477);
nor U155 (N_155,In_155,In_343);
and U156 (N_156,In_508,In_121);
xnor U157 (N_157,In_642,In_215);
and U158 (N_158,In_621,In_293);
nand U159 (N_159,In_150,In_216);
xnor U160 (N_160,In_502,In_208);
xnor U161 (N_161,In_41,In_694);
nor U162 (N_162,In_156,In_311);
nor U163 (N_163,In_225,In_654);
nor U164 (N_164,In_326,In_95);
nand U165 (N_165,In_737,In_59);
nor U166 (N_166,In_634,In_159);
nor U167 (N_167,In_573,In_169);
nand U168 (N_168,In_283,In_749);
nand U169 (N_169,In_125,In_504);
or U170 (N_170,In_583,In_24);
nand U171 (N_171,In_234,In_2);
nor U172 (N_172,In_410,In_360);
nand U173 (N_173,In_555,In_599);
nand U174 (N_174,In_546,In_7);
and U175 (N_175,In_135,In_316);
and U176 (N_176,In_639,In_246);
and U177 (N_177,In_705,In_428);
and U178 (N_178,In_611,In_89);
nor U179 (N_179,In_84,In_607);
or U180 (N_180,In_269,In_616);
nand U181 (N_181,In_231,In_251);
nor U182 (N_182,In_195,In_422);
or U183 (N_183,In_334,In_19);
nand U184 (N_184,In_497,In_413);
and U185 (N_185,In_191,In_45);
nor U186 (N_186,In_586,In_742);
xor U187 (N_187,In_248,In_618);
xor U188 (N_188,In_270,In_700);
xor U189 (N_189,In_645,In_432);
and U190 (N_190,In_613,In_376);
xnor U191 (N_191,In_328,In_718);
or U192 (N_192,In_659,In_294);
nor U193 (N_193,In_395,In_1);
and U194 (N_194,In_748,In_105);
xor U195 (N_195,In_590,In_254);
or U196 (N_196,In_552,In_179);
nor U197 (N_197,In_568,In_585);
or U198 (N_198,In_129,In_655);
nand U199 (N_199,In_9,In_500);
or U200 (N_200,In_405,In_506);
or U201 (N_201,In_278,In_565);
nand U202 (N_202,In_310,In_403);
and U203 (N_203,In_626,In_690);
nor U204 (N_204,In_454,In_392);
xnor U205 (N_205,In_80,In_107);
or U206 (N_206,In_727,In_98);
and U207 (N_207,In_609,In_78);
or U208 (N_208,In_220,In_442);
nand U209 (N_209,In_556,In_572);
and U210 (N_210,In_669,In_55);
or U211 (N_211,In_495,In_102);
nand U212 (N_212,In_292,In_462);
and U213 (N_213,In_182,In_104);
nor U214 (N_214,In_128,In_228);
nand U215 (N_215,In_314,In_286);
nor U216 (N_216,In_467,In_738);
and U217 (N_217,In_404,In_595);
nor U218 (N_218,In_698,In_303);
nand U219 (N_219,In_510,In_557);
and U220 (N_220,In_111,In_32);
nand U221 (N_221,In_699,In_109);
nand U222 (N_222,In_176,In_185);
nand U223 (N_223,In_545,In_461);
nand U224 (N_224,In_563,In_517);
and U225 (N_225,In_58,In_576);
and U226 (N_226,In_589,In_123);
nand U227 (N_227,In_345,In_204);
nor U228 (N_228,In_371,In_720);
or U229 (N_229,In_505,In_36);
xor U230 (N_230,In_536,In_152);
or U231 (N_231,In_524,In_631);
or U232 (N_232,In_527,In_116);
nor U233 (N_233,In_227,In_674);
nor U234 (N_234,In_364,In_614);
xnor U235 (N_235,In_486,In_312);
or U236 (N_236,In_472,In_272);
and U237 (N_237,In_177,In_657);
xor U238 (N_238,In_569,In_151);
nor U239 (N_239,In_170,In_200);
nand U240 (N_240,In_538,In_31);
nor U241 (N_241,In_406,In_465);
nand U242 (N_242,In_305,In_624);
and U243 (N_243,In_327,In_390);
nor U244 (N_244,In_554,In_494);
nor U245 (N_245,In_56,In_542);
or U246 (N_246,In_91,In_632);
and U247 (N_247,In_335,In_290);
xor U248 (N_248,In_196,In_532);
nand U249 (N_249,In_581,In_473);
nand U250 (N_250,In_317,In_113);
or U251 (N_251,In_474,In_429);
xnor U252 (N_252,In_574,In_255);
nand U253 (N_253,In_230,In_11);
nand U254 (N_254,In_445,In_675);
nand U255 (N_255,In_592,In_489);
and U256 (N_256,In_284,In_17);
nor U257 (N_257,In_306,In_194);
or U258 (N_258,In_665,In_491);
xor U259 (N_259,In_553,In_37);
or U260 (N_260,In_118,In_289);
nand U261 (N_261,In_399,In_673);
nand U262 (N_262,In_577,In_598);
and U263 (N_263,In_22,In_351);
and U264 (N_264,In_88,In_439);
nand U265 (N_265,In_453,In_691);
xor U266 (N_266,In_167,In_525);
and U267 (N_267,In_537,In_166);
nor U268 (N_268,In_414,In_470);
and U269 (N_269,In_435,In_575);
xor U270 (N_270,In_153,In_288);
nor U271 (N_271,In_531,In_711);
and U272 (N_272,In_190,In_193);
nor U273 (N_273,In_588,In_275);
nor U274 (N_274,In_448,In_402);
nand U275 (N_275,In_94,In_235);
and U276 (N_276,In_507,In_341);
or U277 (N_277,In_165,In_114);
nand U278 (N_278,In_541,In_394);
or U279 (N_279,In_48,In_511);
and U280 (N_280,In_521,In_426);
or U281 (N_281,In_566,In_325);
or U282 (N_282,In_362,In_322);
and U283 (N_283,In_83,In_300);
and U284 (N_284,In_367,In_146);
and U285 (N_285,In_0,In_347);
and U286 (N_286,In_483,In_715);
and U287 (N_287,In_5,In_238);
nor U288 (N_288,In_267,In_198);
or U289 (N_289,In_164,In_77);
nor U290 (N_290,In_647,In_184);
nand U291 (N_291,In_734,In_381);
nand U292 (N_292,In_443,In_210);
nand U293 (N_293,In_712,In_148);
and U294 (N_294,In_99,In_683);
nand U295 (N_295,In_214,In_120);
nor U296 (N_296,In_640,In_656);
or U297 (N_297,In_490,In_108);
and U298 (N_298,In_648,In_64);
xnor U299 (N_299,In_560,In_61);
or U300 (N_300,In_558,In_564);
or U301 (N_301,In_695,In_391);
and U302 (N_302,In_76,In_93);
xor U303 (N_303,In_15,In_186);
and U304 (N_304,In_70,In_313);
nand U305 (N_305,In_498,In_638);
nand U306 (N_306,In_408,In_726);
and U307 (N_307,In_398,In_296);
nor U308 (N_308,In_523,In_682);
and U309 (N_309,In_357,In_90);
nor U310 (N_310,In_471,In_256);
or U311 (N_311,In_649,In_455);
nor U312 (N_312,In_28,In_644);
or U313 (N_313,In_201,In_450);
nand U314 (N_314,In_27,In_253);
xor U315 (N_315,In_548,In_615);
nor U316 (N_316,In_207,In_512);
nand U317 (N_317,In_409,In_21);
or U318 (N_318,In_295,In_731);
or U319 (N_319,In_464,In_183);
and U320 (N_320,In_332,In_709);
and U321 (N_321,In_363,In_567);
xnor U322 (N_322,In_163,In_416);
nand U323 (N_323,In_329,In_252);
and U324 (N_324,In_717,In_42);
nand U325 (N_325,In_287,In_703);
xor U326 (N_326,In_561,In_417);
or U327 (N_327,In_8,In_323);
xor U328 (N_328,In_240,In_440);
or U329 (N_329,In_383,In_331);
and U330 (N_330,In_226,In_40);
and U331 (N_331,In_433,In_236);
nor U332 (N_332,In_217,In_233);
and U333 (N_333,In_188,In_261);
and U334 (N_334,In_646,In_174);
and U335 (N_335,In_377,In_344);
nor U336 (N_336,In_142,In_678);
nor U337 (N_337,In_708,In_637);
nor U338 (N_338,In_245,In_458);
and U339 (N_339,In_622,In_154);
nor U340 (N_340,In_681,In_49);
nand U341 (N_341,In_81,In_661);
nand U342 (N_342,In_110,In_684);
xnor U343 (N_343,In_25,In_144);
or U344 (N_344,In_119,In_591);
nand U345 (N_345,In_124,In_338);
or U346 (N_346,In_301,In_668);
or U347 (N_347,In_205,In_459);
nand U348 (N_348,In_736,In_658);
nand U349 (N_349,In_115,In_53);
xnor U350 (N_350,In_361,In_549);
nor U351 (N_351,In_707,In_35);
nor U352 (N_352,In_224,In_136);
nand U353 (N_353,In_218,In_535);
nand U354 (N_354,In_625,In_559);
or U355 (N_355,In_451,In_280);
or U356 (N_356,In_247,In_85);
or U357 (N_357,In_46,In_463);
xnor U358 (N_358,In_197,In_578);
nand U359 (N_359,In_719,In_162);
nand U360 (N_360,In_356,In_192);
nor U361 (N_361,In_513,In_242);
xor U362 (N_362,In_75,In_65);
nor U363 (N_363,In_277,In_487);
or U364 (N_364,In_51,In_619);
nor U365 (N_365,In_117,In_436);
and U366 (N_366,In_722,In_730);
nor U367 (N_367,In_728,In_157);
nand U368 (N_368,In_608,In_353);
nand U369 (N_369,In_257,In_239);
nand U370 (N_370,In_651,In_138);
nor U371 (N_371,In_260,In_38);
xor U372 (N_372,In_514,In_20);
nand U373 (N_373,In_488,In_308);
xor U374 (N_374,In_342,In_44);
and U375 (N_375,In_726,In_102);
nor U376 (N_376,In_649,In_330);
nor U377 (N_377,In_368,In_220);
nand U378 (N_378,In_521,In_250);
and U379 (N_379,In_121,In_440);
nand U380 (N_380,In_692,In_258);
or U381 (N_381,In_279,In_716);
and U382 (N_382,In_681,In_404);
or U383 (N_383,In_595,In_598);
nand U384 (N_384,In_33,In_473);
xor U385 (N_385,In_161,In_256);
and U386 (N_386,In_320,In_728);
or U387 (N_387,In_316,In_273);
and U388 (N_388,In_225,In_147);
nor U389 (N_389,In_736,In_508);
xnor U390 (N_390,In_400,In_596);
and U391 (N_391,In_181,In_219);
nand U392 (N_392,In_41,In_679);
xor U393 (N_393,In_102,In_227);
nor U394 (N_394,In_603,In_430);
and U395 (N_395,In_133,In_581);
and U396 (N_396,In_168,In_72);
or U397 (N_397,In_107,In_150);
or U398 (N_398,In_499,In_640);
xnor U399 (N_399,In_747,In_465);
nor U400 (N_400,In_341,In_644);
or U401 (N_401,In_144,In_592);
and U402 (N_402,In_500,In_714);
and U403 (N_403,In_652,In_386);
nor U404 (N_404,In_542,In_526);
or U405 (N_405,In_191,In_588);
or U406 (N_406,In_121,In_318);
and U407 (N_407,In_389,In_257);
or U408 (N_408,In_6,In_99);
nor U409 (N_409,In_69,In_204);
nand U410 (N_410,In_87,In_348);
or U411 (N_411,In_196,In_264);
and U412 (N_412,In_364,In_420);
xnor U413 (N_413,In_436,In_573);
nand U414 (N_414,In_343,In_692);
nand U415 (N_415,In_628,In_492);
nor U416 (N_416,In_457,In_741);
nand U417 (N_417,In_546,In_609);
and U418 (N_418,In_23,In_740);
nor U419 (N_419,In_602,In_685);
and U420 (N_420,In_535,In_329);
and U421 (N_421,In_598,In_187);
nor U422 (N_422,In_12,In_647);
nand U423 (N_423,In_533,In_129);
or U424 (N_424,In_645,In_14);
nor U425 (N_425,In_274,In_449);
xor U426 (N_426,In_342,In_73);
or U427 (N_427,In_687,In_713);
and U428 (N_428,In_176,In_22);
nand U429 (N_429,In_745,In_157);
nor U430 (N_430,In_97,In_442);
or U431 (N_431,In_591,In_585);
nor U432 (N_432,In_676,In_3);
or U433 (N_433,In_660,In_142);
or U434 (N_434,In_60,In_40);
nand U435 (N_435,In_428,In_410);
nand U436 (N_436,In_233,In_76);
nand U437 (N_437,In_4,In_731);
or U438 (N_438,In_285,In_202);
or U439 (N_439,In_339,In_228);
nor U440 (N_440,In_619,In_474);
xor U441 (N_441,In_677,In_352);
nand U442 (N_442,In_641,In_106);
or U443 (N_443,In_71,In_262);
xor U444 (N_444,In_142,In_454);
nand U445 (N_445,In_106,In_584);
nand U446 (N_446,In_218,In_403);
or U447 (N_447,In_389,In_319);
nor U448 (N_448,In_685,In_668);
nand U449 (N_449,In_659,In_262);
and U450 (N_450,In_433,In_692);
or U451 (N_451,In_232,In_415);
or U452 (N_452,In_94,In_489);
nor U453 (N_453,In_397,In_292);
nand U454 (N_454,In_8,In_565);
nand U455 (N_455,In_258,In_26);
nor U456 (N_456,In_212,In_554);
or U457 (N_457,In_270,In_254);
nor U458 (N_458,In_703,In_582);
or U459 (N_459,In_429,In_730);
or U460 (N_460,In_58,In_25);
and U461 (N_461,In_352,In_233);
or U462 (N_462,In_278,In_684);
nand U463 (N_463,In_477,In_223);
nor U464 (N_464,In_414,In_5);
or U465 (N_465,In_389,In_35);
or U466 (N_466,In_510,In_94);
or U467 (N_467,In_350,In_417);
and U468 (N_468,In_600,In_590);
or U469 (N_469,In_221,In_605);
or U470 (N_470,In_539,In_686);
nor U471 (N_471,In_458,In_156);
xnor U472 (N_472,In_409,In_483);
or U473 (N_473,In_739,In_453);
and U474 (N_474,In_259,In_714);
and U475 (N_475,In_426,In_96);
nor U476 (N_476,In_19,In_423);
or U477 (N_477,In_615,In_485);
nor U478 (N_478,In_92,In_373);
or U479 (N_479,In_617,In_739);
xnor U480 (N_480,In_175,In_516);
nand U481 (N_481,In_271,In_584);
and U482 (N_482,In_358,In_580);
nor U483 (N_483,In_606,In_594);
nand U484 (N_484,In_416,In_228);
nor U485 (N_485,In_83,In_533);
or U486 (N_486,In_301,In_360);
nor U487 (N_487,In_263,In_396);
nor U488 (N_488,In_91,In_359);
xor U489 (N_489,In_255,In_128);
nor U490 (N_490,In_213,In_59);
or U491 (N_491,In_22,In_738);
xor U492 (N_492,In_418,In_29);
xnor U493 (N_493,In_518,In_601);
xor U494 (N_494,In_684,In_558);
or U495 (N_495,In_272,In_70);
xnor U496 (N_496,In_307,In_351);
nor U497 (N_497,In_243,In_533);
nor U498 (N_498,In_567,In_43);
and U499 (N_499,In_96,In_335);
nand U500 (N_500,N_189,N_486);
nand U501 (N_501,N_79,N_149);
xor U502 (N_502,N_430,N_160);
or U503 (N_503,N_58,N_217);
nor U504 (N_504,N_454,N_395);
nor U505 (N_505,N_163,N_328);
or U506 (N_506,N_412,N_226);
and U507 (N_507,N_18,N_129);
nand U508 (N_508,N_305,N_262);
nor U509 (N_509,N_230,N_385);
or U510 (N_510,N_358,N_474);
nor U511 (N_511,N_271,N_369);
nor U512 (N_512,N_487,N_153);
or U513 (N_513,N_158,N_447);
or U514 (N_514,N_164,N_199);
and U515 (N_515,N_135,N_240);
nand U516 (N_516,N_118,N_131);
and U517 (N_517,N_427,N_420);
xnor U518 (N_518,N_111,N_177);
and U519 (N_519,N_59,N_359);
or U520 (N_520,N_216,N_42);
or U521 (N_521,N_197,N_494);
or U522 (N_522,N_146,N_170);
nor U523 (N_523,N_437,N_391);
nand U524 (N_524,N_251,N_92);
nor U525 (N_525,N_80,N_416);
or U526 (N_526,N_288,N_147);
or U527 (N_527,N_282,N_370);
nor U528 (N_528,N_259,N_11);
nand U529 (N_529,N_45,N_17);
nand U530 (N_530,N_83,N_389);
nor U531 (N_531,N_329,N_424);
or U532 (N_532,N_220,N_349);
xnor U533 (N_533,N_224,N_200);
nor U534 (N_534,N_33,N_229);
and U535 (N_535,N_352,N_279);
or U536 (N_536,N_206,N_485);
or U537 (N_537,N_139,N_403);
or U538 (N_538,N_308,N_187);
nand U539 (N_539,N_194,N_449);
nand U540 (N_540,N_300,N_141);
nand U541 (N_541,N_142,N_415);
nor U542 (N_542,N_467,N_360);
nor U543 (N_543,N_128,N_169);
and U544 (N_544,N_397,N_376);
and U545 (N_545,N_211,N_323);
or U546 (N_546,N_425,N_237);
nand U547 (N_547,N_294,N_102);
nand U548 (N_548,N_24,N_417);
and U549 (N_549,N_121,N_339);
nor U550 (N_550,N_405,N_234);
xnor U551 (N_551,N_337,N_366);
nand U552 (N_552,N_433,N_176);
nor U553 (N_553,N_204,N_54);
nor U554 (N_554,N_46,N_428);
and U555 (N_555,N_67,N_411);
xnor U556 (N_556,N_171,N_57);
xor U557 (N_557,N_49,N_399);
nand U558 (N_558,N_312,N_275);
nor U559 (N_559,N_446,N_281);
and U560 (N_560,N_66,N_193);
and U561 (N_561,N_65,N_152);
nor U562 (N_562,N_183,N_0);
nand U563 (N_563,N_296,N_482);
or U564 (N_564,N_267,N_287);
and U565 (N_565,N_440,N_466);
and U566 (N_566,N_367,N_322);
or U567 (N_567,N_445,N_413);
nor U568 (N_568,N_292,N_456);
or U569 (N_569,N_253,N_192);
and U570 (N_570,N_112,N_346);
and U571 (N_571,N_340,N_324);
and U572 (N_572,N_117,N_91);
nand U573 (N_573,N_263,N_400);
nand U574 (N_574,N_317,N_51);
or U575 (N_575,N_293,N_331);
or U576 (N_576,N_161,N_471);
or U577 (N_577,N_110,N_410);
or U578 (N_578,N_455,N_404);
nand U579 (N_579,N_137,N_309);
nor U580 (N_580,N_219,N_101);
nand U581 (N_581,N_319,N_261);
xnor U582 (N_582,N_335,N_64);
and U583 (N_583,N_47,N_448);
nand U584 (N_584,N_386,N_130);
or U585 (N_585,N_250,N_377);
nor U586 (N_586,N_38,N_441);
nand U587 (N_587,N_225,N_12);
nand U588 (N_588,N_123,N_257);
xnor U589 (N_589,N_476,N_132);
and U590 (N_590,N_249,N_277);
nand U591 (N_591,N_483,N_236);
nand U592 (N_592,N_231,N_278);
or U593 (N_593,N_207,N_347);
nand U594 (N_594,N_162,N_144);
nand U595 (N_595,N_473,N_212);
nor U596 (N_596,N_157,N_464);
xor U597 (N_597,N_463,N_168);
or U598 (N_598,N_408,N_451);
xnor U599 (N_599,N_436,N_98);
and U600 (N_600,N_70,N_383);
and U601 (N_601,N_497,N_73);
or U602 (N_602,N_260,N_97);
nor U603 (N_603,N_499,N_266);
and U604 (N_604,N_378,N_396);
xor U605 (N_605,N_39,N_478);
and U606 (N_606,N_107,N_422);
or U607 (N_607,N_356,N_315);
and U608 (N_608,N_61,N_361);
nor U609 (N_609,N_14,N_276);
nor U610 (N_610,N_419,N_184);
nand U611 (N_611,N_2,N_459);
and U612 (N_612,N_450,N_357);
or U613 (N_613,N_390,N_426);
and U614 (N_614,N_336,N_421);
or U615 (N_615,N_490,N_274);
and U616 (N_616,N_30,N_255);
nor U617 (N_617,N_342,N_35);
nand U618 (N_618,N_460,N_109);
and U619 (N_619,N_371,N_34);
or U620 (N_620,N_68,N_373);
or U621 (N_621,N_462,N_232);
nand U622 (N_622,N_246,N_133);
and U623 (N_623,N_432,N_330);
nand U624 (N_624,N_3,N_86);
nor U625 (N_625,N_155,N_63);
nand U626 (N_626,N_5,N_9);
and U627 (N_627,N_241,N_76);
nand U628 (N_628,N_6,N_173);
or U629 (N_629,N_365,N_256);
or U630 (N_630,N_179,N_56);
or U631 (N_631,N_96,N_233);
and U632 (N_632,N_488,N_332);
and U633 (N_633,N_318,N_303);
nor U634 (N_634,N_465,N_484);
nand U635 (N_635,N_444,N_50);
nor U636 (N_636,N_136,N_95);
or U637 (N_637,N_205,N_172);
xor U638 (N_638,N_239,N_181);
nand U639 (N_639,N_381,N_227);
nand U640 (N_640,N_119,N_74);
nand U641 (N_641,N_398,N_325);
nor U642 (N_642,N_201,N_8);
xnor U643 (N_643,N_401,N_36);
and U644 (N_644,N_221,N_85);
and U645 (N_645,N_297,N_355);
nand U646 (N_646,N_406,N_414);
and U647 (N_647,N_333,N_338);
or U648 (N_648,N_492,N_20);
nor U649 (N_649,N_321,N_1);
or U650 (N_650,N_457,N_10);
nor U651 (N_651,N_299,N_245);
and U652 (N_652,N_31,N_264);
or U653 (N_653,N_72,N_84);
nor U654 (N_654,N_88,N_124);
nand U655 (N_655,N_311,N_442);
nor U656 (N_656,N_409,N_418);
or U657 (N_657,N_477,N_71);
xnor U658 (N_658,N_40,N_327);
nor U659 (N_659,N_461,N_113);
or U660 (N_660,N_190,N_468);
nand U661 (N_661,N_55,N_140);
nor U662 (N_662,N_174,N_69);
and U663 (N_663,N_286,N_48);
or U664 (N_664,N_393,N_185);
nor U665 (N_665,N_156,N_105);
nand U666 (N_666,N_180,N_148);
nand U667 (N_667,N_41,N_134);
nand U668 (N_668,N_191,N_196);
and U669 (N_669,N_452,N_374);
nor U670 (N_670,N_89,N_402);
xnor U671 (N_671,N_252,N_82);
nor U672 (N_672,N_429,N_154);
nand U673 (N_673,N_301,N_75);
nor U674 (N_674,N_479,N_203);
and U675 (N_675,N_21,N_93);
nor U676 (N_676,N_202,N_182);
xnor U677 (N_677,N_166,N_316);
and U678 (N_678,N_298,N_28);
nand U679 (N_679,N_150,N_125);
and U680 (N_680,N_351,N_159);
nor U681 (N_681,N_248,N_268);
or U682 (N_682,N_475,N_87);
or U683 (N_683,N_210,N_372);
xor U684 (N_684,N_19,N_431);
or U685 (N_685,N_138,N_81);
nor U686 (N_686,N_392,N_363);
or U687 (N_687,N_285,N_60);
and U688 (N_688,N_27,N_407);
xor U689 (N_689,N_423,N_106);
nand U690 (N_690,N_235,N_472);
and U691 (N_691,N_434,N_104);
nand U692 (N_692,N_443,N_165);
nand U693 (N_693,N_380,N_115);
nand U694 (N_694,N_167,N_127);
nor U695 (N_695,N_348,N_495);
and U696 (N_696,N_7,N_394);
and U697 (N_697,N_37,N_222);
nand U698 (N_698,N_313,N_498);
or U699 (N_699,N_44,N_269);
nor U700 (N_700,N_353,N_280);
or U701 (N_701,N_307,N_188);
nor U702 (N_702,N_439,N_94);
nand U703 (N_703,N_22,N_186);
and U704 (N_704,N_62,N_491);
and U705 (N_705,N_114,N_215);
xor U706 (N_706,N_213,N_480);
nor U707 (N_707,N_218,N_103);
or U708 (N_708,N_481,N_238);
xor U709 (N_709,N_496,N_364);
nand U710 (N_710,N_90,N_320);
and U711 (N_711,N_379,N_198);
and U712 (N_712,N_247,N_25);
or U713 (N_713,N_214,N_326);
nand U714 (N_714,N_15,N_295);
nand U715 (N_715,N_470,N_223);
nor U716 (N_716,N_493,N_284);
and U717 (N_717,N_143,N_344);
nor U718 (N_718,N_126,N_100);
or U719 (N_719,N_32,N_384);
xor U720 (N_720,N_209,N_4);
and U721 (N_721,N_78,N_302);
and U722 (N_722,N_291,N_178);
nor U723 (N_723,N_334,N_310);
and U724 (N_724,N_23,N_151);
and U725 (N_725,N_435,N_314);
nor U726 (N_726,N_489,N_29);
nand U727 (N_727,N_43,N_16);
nor U728 (N_728,N_375,N_26);
or U729 (N_729,N_52,N_108);
nand U730 (N_730,N_122,N_368);
and U731 (N_731,N_13,N_175);
xnor U732 (N_732,N_453,N_77);
and U733 (N_733,N_53,N_345);
or U734 (N_734,N_258,N_469);
nand U735 (N_735,N_244,N_387);
and U736 (N_736,N_289,N_458);
and U737 (N_737,N_382,N_350);
xnor U738 (N_738,N_304,N_242);
nor U739 (N_739,N_99,N_195);
nand U740 (N_740,N_145,N_290);
and U741 (N_741,N_116,N_341);
nor U742 (N_742,N_254,N_343);
nand U743 (N_743,N_228,N_306);
and U744 (N_744,N_208,N_283);
or U745 (N_745,N_354,N_362);
xnor U746 (N_746,N_270,N_120);
and U747 (N_747,N_273,N_243);
or U748 (N_748,N_265,N_438);
nor U749 (N_749,N_388,N_272);
or U750 (N_750,N_276,N_187);
and U751 (N_751,N_123,N_66);
or U752 (N_752,N_283,N_489);
and U753 (N_753,N_55,N_446);
nand U754 (N_754,N_150,N_250);
and U755 (N_755,N_1,N_147);
nor U756 (N_756,N_435,N_394);
nand U757 (N_757,N_413,N_196);
and U758 (N_758,N_235,N_453);
nor U759 (N_759,N_151,N_256);
or U760 (N_760,N_239,N_266);
or U761 (N_761,N_162,N_443);
nand U762 (N_762,N_300,N_384);
or U763 (N_763,N_475,N_46);
xor U764 (N_764,N_41,N_46);
and U765 (N_765,N_202,N_244);
nand U766 (N_766,N_442,N_212);
nand U767 (N_767,N_151,N_269);
xnor U768 (N_768,N_5,N_21);
or U769 (N_769,N_359,N_62);
and U770 (N_770,N_217,N_430);
nand U771 (N_771,N_45,N_94);
or U772 (N_772,N_499,N_165);
or U773 (N_773,N_254,N_356);
nor U774 (N_774,N_446,N_168);
nand U775 (N_775,N_462,N_27);
nor U776 (N_776,N_80,N_496);
or U777 (N_777,N_293,N_147);
nand U778 (N_778,N_247,N_296);
or U779 (N_779,N_494,N_47);
nor U780 (N_780,N_479,N_336);
nor U781 (N_781,N_59,N_200);
nor U782 (N_782,N_41,N_322);
nor U783 (N_783,N_46,N_481);
nand U784 (N_784,N_313,N_260);
or U785 (N_785,N_190,N_427);
nand U786 (N_786,N_84,N_498);
or U787 (N_787,N_98,N_53);
nand U788 (N_788,N_116,N_280);
or U789 (N_789,N_40,N_267);
nor U790 (N_790,N_148,N_429);
nor U791 (N_791,N_321,N_132);
or U792 (N_792,N_93,N_429);
xor U793 (N_793,N_385,N_474);
or U794 (N_794,N_204,N_84);
nor U795 (N_795,N_29,N_119);
or U796 (N_796,N_40,N_446);
nand U797 (N_797,N_30,N_286);
nor U798 (N_798,N_397,N_423);
and U799 (N_799,N_409,N_143);
nor U800 (N_800,N_231,N_167);
nand U801 (N_801,N_255,N_352);
nor U802 (N_802,N_7,N_129);
or U803 (N_803,N_393,N_199);
and U804 (N_804,N_119,N_273);
xor U805 (N_805,N_288,N_215);
nor U806 (N_806,N_342,N_449);
and U807 (N_807,N_401,N_17);
nor U808 (N_808,N_204,N_74);
nor U809 (N_809,N_325,N_419);
and U810 (N_810,N_83,N_247);
nor U811 (N_811,N_180,N_53);
nand U812 (N_812,N_1,N_243);
nand U813 (N_813,N_326,N_107);
or U814 (N_814,N_477,N_379);
and U815 (N_815,N_160,N_373);
or U816 (N_816,N_217,N_48);
and U817 (N_817,N_351,N_261);
nand U818 (N_818,N_225,N_204);
or U819 (N_819,N_123,N_394);
nor U820 (N_820,N_388,N_352);
or U821 (N_821,N_290,N_411);
nor U822 (N_822,N_3,N_201);
nand U823 (N_823,N_152,N_265);
xor U824 (N_824,N_257,N_323);
and U825 (N_825,N_368,N_300);
nand U826 (N_826,N_51,N_22);
nand U827 (N_827,N_132,N_33);
nor U828 (N_828,N_197,N_489);
xor U829 (N_829,N_273,N_191);
and U830 (N_830,N_138,N_267);
nand U831 (N_831,N_495,N_269);
and U832 (N_832,N_400,N_244);
and U833 (N_833,N_56,N_83);
nand U834 (N_834,N_481,N_72);
nand U835 (N_835,N_144,N_46);
nor U836 (N_836,N_130,N_383);
or U837 (N_837,N_45,N_397);
and U838 (N_838,N_301,N_103);
or U839 (N_839,N_477,N_288);
and U840 (N_840,N_261,N_96);
or U841 (N_841,N_429,N_73);
xnor U842 (N_842,N_151,N_440);
and U843 (N_843,N_10,N_198);
nor U844 (N_844,N_369,N_381);
xor U845 (N_845,N_257,N_246);
nor U846 (N_846,N_456,N_159);
nand U847 (N_847,N_336,N_485);
nor U848 (N_848,N_389,N_241);
nand U849 (N_849,N_466,N_198);
and U850 (N_850,N_426,N_54);
xor U851 (N_851,N_204,N_247);
or U852 (N_852,N_496,N_251);
xor U853 (N_853,N_258,N_291);
and U854 (N_854,N_250,N_249);
or U855 (N_855,N_244,N_227);
nand U856 (N_856,N_365,N_182);
nand U857 (N_857,N_200,N_348);
nand U858 (N_858,N_283,N_333);
nand U859 (N_859,N_312,N_293);
nor U860 (N_860,N_59,N_335);
and U861 (N_861,N_60,N_137);
nand U862 (N_862,N_446,N_7);
nor U863 (N_863,N_423,N_498);
or U864 (N_864,N_56,N_108);
nor U865 (N_865,N_295,N_23);
and U866 (N_866,N_368,N_105);
nand U867 (N_867,N_432,N_10);
nor U868 (N_868,N_498,N_206);
nor U869 (N_869,N_209,N_138);
nor U870 (N_870,N_239,N_66);
and U871 (N_871,N_52,N_138);
and U872 (N_872,N_272,N_204);
or U873 (N_873,N_471,N_435);
xor U874 (N_874,N_308,N_491);
and U875 (N_875,N_203,N_69);
nand U876 (N_876,N_373,N_169);
nand U877 (N_877,N_51,N_248);
nor U878 (N_878,N_393,N_235);
or U879 (N_879,N_306,N_337);
nand U880 (N_880,N_469,N_245);
or U881 (N_881,N_475,N_389);
nor U882 (N_882,N_280,N_98);
and U883 (N_883,N_412,N_225);
nand U884 (N_884,N_237,N_446);
nand U885 (N_885,N_402,N_481);
or U886 (N_886,N_383,N_407);
nor U887 (N_887,N_449,N_7);
nor U888 (N_888,N_244,N_44);
xnor U889 (N_889,N_262,N_434);
or U890 (N_890,N_476,N_128);
or U891 (N_891,N_362,N_73);
and U892 (N_892,N_278,N_463);
and U893 (N_893,N_298,N_235);
and U894 (N_894,N_42,N_275);
nor U895 (N_895,N_475,N_183);
or U896 (N_896,N_329,N_194);
or U897 (N_897,N_466,N_335);
and U898 (N_898,N_140,N_171);
or U899 (N_899,N_288,N_141);
xor U900 (N_900,N_326,N_126);
and U901 (N_901,N_389,N_9);
nand U902 (N_902,N_271,N_252);
or U903 (N_903,N_319,N_332);
and U904 (N_904,N_253,N_36);
xnor U905 (N_905,N_65,N_256);
nand U906 (N_906,N_291,N_301);
and U907 (N_907,N_370,N_115);
xor U908 (N_908,N_206,N_460);
nand U909 (N_909,N_193,N_15);
and U910 (N_910,N_57,N_336);
and U911 (N_911,N_135,N_344);
or U912 (N_912,N_335,N_239);
nor U913 (N_913,N_479,N_242);
or U914 (N_914,N_350,N_81);
and U915 (N_915,N_156,N_434);
xor U916 (N_916,N_416,N_407);
and U917 (N_917,N_289,N_365);
nor U918 (N_918,N_181,N_463);
nor U919 (N_919,N_320,N_497);
and U920 (N_920,N_284,N_143);
or U921 (N_921,N_339,N_323);
or U922 (N_922,N_68,N_405);
nor U923 (N_923,N_420,N_104);
and U924 (N_924,N_421,N_6);
xnor U925 (N_925,N_35,N_461);
and U926 (N_926,N_275,N_382);
nor U927 (N_927,N_227,N_401);
or U928 (N_928,N_16,N_64);
or U929 (N_929,N_199,N_122);
nor U930 (N_930,N_2,N_29);
or U931 (N_931,N_137,N_486);
or U932 (N_932,N_93,N_158);
and U933 (N_933,N_429,N_345);
nor U934 (N_934,N_248,N_84);
xnor U935 (N_935,N_171,N_165);
and U936 (N_936,N_96,N_83);
and U937 (N_937,N_423,N_53);
and U938 (N_938,N_233,N_412);
and U939 (N_939,N_6,N_449);
nand U940 (N_940,N_237,N_221);
nor U941 (N_941,N_492,N_11);
nor U942 (N_942,N_301,N_346);
and U943 (N_943,N_222,N_116);
xor U944 (N_944,N_163,N_255);
nor U945 (N_945,N_439,N_474);
nor U946 (N_946,N_57,N_395);
and U947 (N_947,N_492,N_111);
and U948 (N_948,N_232,N_46);
and U949 (N_949,N_79,N_374);
nand U950 (N_950,N_248,N_405);
and U951 (N_951,N_394,N_4);
or U952 (N_952,N_453,N_44);
or U953 (N_953,N_453,N_451);
nand U954 (N_954,N_452,N_256);
nand U955 (N_955,N_436,N_2);
nor U956 (N_956,N_124,N_389);
xnor U957 (N_957,N_49,N_388);
and U958 (N_958,N_265,N_255);
xor U959 (N_959,N_242,N_469);
nor U960 (N_960,N_150,N_233);
and U961 (N_961,N_216,N_451);
nor U962 (N_962,N_73,N_46);
nor U963 (N_963,N_299,N_248);
xor U964 (N_964,N_451,N_371);
and U965 (N_965,N_385,N_249);
nor U966 (N_966,N_96,N_410);
nand U967 (N_967,N_352,N_154);
and U968 (N_968,N_225,N_315);
or U969 (N_969,N_427,N_221);
nand U970 (N_970,N_489,N_380);
xnor U971 (N_971,N_177,N_92);
or U972 (N_972,N_447,N_79);
xnor U973 (N_973,N_242,N_64);
or U974 (N_974,N_266,N_395);
and U975 (N_975,N_462,N_388);
nand U976 (N_976,N_237,N_26);
or U977 (N_977,N_271,N_380);
and U978 (N_978,N_484,N_284);
nand U979 (N_979,N_371,N_234);
or U980 (N_980,N_201,N_145);
xor U981 (N_981,N_10,N_219);
xor U982 (N_982,N_8,N_370);
and U983 (N_983,N_205,N_209);
nor U984 (N_984,N_304,N_181);
or U985 (N_985,N_419,N_141);
nor U986 (N_986,N_324,N_302);
nand U987 (N_987,N_78,N_55);
xnor U988 (N_988,N_144,N_198);
nand U989 (N_989,N_254,N_330);
nand U990 (N_990,N_37,N_10);
nand U991 (N_991,N_125,N_435);
nor U992 (N_992,N_215,N_20);
xnor U993 (N_993,N_400,N_383);
nor U994 (N_994,N_174,N_359);
nand U995 (N_995,N_356,N_305);
nand U996 (N_996,N_316,N_163);
and U997 (N_997,N_28,N_7);
nor U998 (N_998,N_36,N_290);
and U999 (N_999,N_256,N_327);
or U1000 (N_1000,N_763,N_782);
nor U1001 (N_1001,N_954,N_828);
or U1002 (N_1002,N_540,N_975);
xor U1003 (N_1003,N_890,N_500);
or U1004 (N_1004,N_674,N_746);
nand U1005 (N_1005,N_899,N_790);
or U1006 (N_1006,N_772,N_884);
nand U1007 (N_1007,N_513,N_821);
xnor U1008 (N_1008,N_817,N_554);
and U1009 (N_1009,N_648,N_517);
or U1010 (N_1010,N_918,N_693);
or U1011 (N_1011,N_725,N_581);
and U1012 (N_1012,N_728,N_642);
and U1013 (N_1013,N_766,N_986);
and U1014 (N_1014,N_593,N_641);
xnor U1015 (N_1015,N_791,N_998);
xor U1016 (N_1016,N_967,N_920);
or U1017 (N_1017,N_754,N_855);
and U1018 (N_1018,N_708,N_863);
nand U1019 (N_1019,N_559,N_701);
and U1020 (N_1020,N_707,N_927);
and U1021 (N_1021,N_943,N_662);
nor U1022 (N_1022,N_952,N_506);
or U1023 (N_1023,N_972,N_950);
and U1024 (N_1024,N_564,N_563);
and U1025 (N_1025,N_711,N_990);
xor U1026 (N_1026,N_953,N_826);
or U1027 (N_1027,N_809,N_980);
nand U1028 (N_1028,N_555,N_751);
nor U1029 (N_1029,N_777,N_514);
or U1030 (N_1030,N_745,N_675);
nand U1031 (N_1031,N_651,N_710);
or U1032 (N_1032,N_601,N_861);
and U1033 (N_1033,N_729,N_549);
and U1034 (N_1034,N_778,N_647);
nor U1035 (N_1035,N_836,N_716);
or U1036 (N_1036,N_628,N_685);
or U1037 (N_1037,N_659,N_550);
or U1038 (N_1038,N_819,N_535);
nor U1039 (N_1039,N_551,N_803);
or U1040 (N_1040,N_650,N_719);
and U1041 (N_1041,N_678,N_590);
and U1042 (N_1042,N_516,N_961);
and U1043 (N_1043,N_605,N_656);
and U1044 (N_1044,N_621,N_893);
or U1045 (N_1045,N_565,N_706);
and U1046 (N_1046,N_912,N_885);
and U1047 (N_1047,N_668,N_985);
nand U1048 (N_1048,N_835,N_850);
nor U1049 (N_1049,N_811,N_797);
and U1050 (N_1050,N_818,N_794);
and U1051 (N_1051,N_569,N_904);
nor U1052 (N_1052,N_970,N_518);
and U1053 (N_1053,N_793,N_977);
nand U1054 (N_1054,N_684,N_865);
nand U1055 (N_1055,N_692,N_853);
xnor U1056 (N_1056,N_805,N_501);
nand U1057 (N_1057,N_841,N_544);
or U1058 (N_1058,N_947,N_646);
and U1059 (N_1059,N_808,N_915);
nand U1060 (N_1060,N_576,N_829);
or U1061 (N_1061,N_857,N_531);
and U1062 (N_1062,N_773,N_832);
nor U1063 (N_1063,N_546,N_680);
or U1064 (N_1064,N_957,N_767);
xnor U1065 (N_1065,N_911,N_981);
nor U1066 (N_1066,N_543,N_966);
xor U1067 (N_1067,N_798,N_880);
or U1068 (N_1068,N_895,N_936);
or U1069 (N_1069,N_524,N_939);
or U1070 (N_1070,N_713,N_688);
or U1071 (N_1071,N_694,N_823);
and U1072 (N_1072,N_552,N_816);
and U1073 (N_1073,N_958,N_871);
or U1074 (N_1074,N_847,N_994);
xnor U1075 (N_1075,N_741,N_788);
nor U1076 (N_1076,N_897,N_515);
nand U1077 (N_1077,N_681,N_886);
xor U1078 (N_1078,N_834,N_807);
and U1079 (N_1079,N_671,N_858);
nor U1080 (N_1080,N_717,N_643);
and U1081 (N_1081,N_724,N_718);
and U1082 (N_1082,N_672,N_887);
nor U1083 (N_1083,N_537,N_851);
nor U1084 (N_1084,N_783,N_534);
or U1085 (N_1085,N_806,N_536);
and U1086 (N_1086,N_820,N_612);
nand U1087 (N_1087,N_844,N_696);
and U1088 (N_1088,N_833,N_747);
or U1089 (N_1089,N_968,N_891);
or U1090 (N_1090,N_868,N_510);
nor U1091 (N_1091,N_928,N_872);
xor U1092 (N_1092,N_557,N_652);
nor U1093 (N_1093,N_677,N_698);
xor U1094 (N_1094,N_703,N_827);
xnor U1095 (N_1095,N_784,N_520);
and U1096 (N_1096,N_578,N_619);
nor U1097 (N_1097,N_606,N_739);
xnor U1098 (N_1098,N_924,N_976);
nand U1099 (N_1099,N_682,N_866);
xor U1100 (N_1100,N_992,N_721);
nor U1101 (N_1101,N_780,N_588);
nor U1102 (N_1102,N_769,N_690);
nor U1103 (N_1103,N_812,N_732);
or U1104 (N_1104,N_775,N_699);
or U1105 (N_1105,N_849,N_720);
or U1106 (N_1106,N_634,N_771);
nor U1107 (N_1107,N_586,N_542);
and U1108 (N_1108,N_509,N_657);
nand U1109 (N_1109,N_687,N_839);
nor U1110 (N_1110,N_770,N_562);
nand U1111 (N_1111,N_925,N_661);
nor U1112 (N_1112,N_978,N_932);
and U1113 (N_1113,N_963,N_539);
and U1114 (N_1114,N_599,N_759);
and U1115 (N_1115,N_528,N_610);
or U1116 (N_1116,N_523,N_756);
and U1117 (N_1117,N_574,N_587);
and U1118 (N_1118,N_743,N_547);
nand U1119 (N_1119,N_787,N_575);
and U1120 (N_1120,N_760,N_566);
or U1121 (N_1121,N_814,N_802);
or U1122 (N_1122,N_622,N_876);
or U1123 (N_1123,N_956,N_636);
and U1124 (N_1124,N_919,N_874);
nor U1125 (N_1125,N_764,N_704);
nor U1126 (N_1126,N_989,N_779);
xnor U1127 (N_1127,N_988,N_974);
nor U1128 (N_1128,N_618,N_894);
or U1129 (N_1129,N_625,N_785);
and U1130 (N_1130,N_914,N_944);
and U1131 (N_1131,N_591,N_709);
and U1132 (N_1132,N_548,N_620);
nand U1133 (N_1133,N_529,N_774);
nand U1134 (N_1134,N_856,N_987);
or U1135 (N_1135,N_735,N_553);
and U1136 (N_1136,N_792,N_623);
nand U1137 (N_1137,N_916,N_683);
and U1138 (N_1138,N_645,N_592);
or U1139 (N_1139,N_627,N_614);
and U1140 (N_1140,N_649,N_942);
nor U1141 (N_1141,N_583,N_736);
or U1142 (N_1142,N_530,N_860);
nor U1143 (N_1143,N_800,N_949);
and U1144 (N_1144,N_840,N_951);
nor U1145 (N_1145,N_532,N_786);
nor U1146 (N_1146,N_908,N_615);
nor U1147 (N_1147,N_589,N_870);
and U1148 (N_1148,N_511,N_603);
nor U1149 (N_1149,N_852,N_600);
nor U1150 (N_1150,N_996,N_755);
nor U1151 (N_1151,N_881,N_519);
xor U1152 (N_1152,N_984,N_705);
or U1153 (N_1153,N_512,N_731);
nand U1154 (N_1154,N_907,N_561);
or U1155 (N_1155,N_873,N_753);
nand U1156 (N_1156,N_663,N_796);
nor U1157 (N_1157,N_862,N_658);
nand U1158 (N_1158,N_776,N_843);
and U1159 (N_1159,N_630,N_525);
nor U1160 (N_1160,N_697,N_505);
nand U1161 (N_1161,N_888,N_585);
nand U1162 (N_1162,N_991,N_637);
nor U1163 (N_1163,N_629,N_626);
or U1164 (N_1164,N_595,N_813);
nand U1165 (N_1165,N_758,N_946);
nor U1166 (N_1166,N_973,N_877);
and U1167 (N_1167,N_567,N_742);
nand U1168 (N_1168,N_664,N_979);
nor U1169 (N_1169,N_882,N_905);
and U1170 (N_1170,N_815,N_744);
nor U1171 (N_1171,N_935,N_631);
and U1172 (N_1172,N_864,N_582);
or U1173 (N_1173,N_971,N_541);
nor U1174 (N_1174,N_660,N_527);
or U1175 (N_1175,N_902,N_962);
and U1176 (N_1176,N_573,N_913);
or U1177 (N_1177,N_635,N_789);
nor U1178 (N_1178,N_995,N_930);
nand U1179 (N_1179,N_969,N_571);
nor U1180 (N_1180,N_982,N_560);
xor U1181 (N_1181,N_923,N_695);
and U1182 (N_1182,N_632,N_526);
and U1183 (N_1183,N_714,N_580);
or U1184 (N_1184,N_700,N_613);
and U1185 (N_1185,N_837,N_673);
nand U1186 (N_1186,N_889,N_558);
or U1187 (N_1187,N_538,N_616);
and U1188 (N_1188,N_568,N_666);
or U1189 (N_1189,N_941,N_702);
nor U1190 (N_1190,N_579,N_508);
or U1191 (N_1191,N_765,N_999);
xor U1192 (N_1192,N_598,N_848);
and U1193 (N_1193,N_584,N_665);
nor U1194 (N_1194,N_609,N_761);
and U1195 (N_1195,N_522,N_825);
or U1196 (N_1196,N_906,N_762);
nand U1197 (N_1197,N_727,N_830);
and U1198 (N_1198,N_964,N_653);
nor U1199 (N_1199,N_733,N_993);
nand U1200 (N_1200,N_669,N_810);
or U1201 (N_1201,N_624,N_842);
and U1202 (N_1202,N_983,N_597);
xor U1203 (N_1203,N_921,N_937);
xnor U1204 (N_1204,N_644,N_822);
nor U1205 (N_1205,N_903,N_801);
nand U1206 (N_1206,N_875,N_594);
nor U1207 (N_1207,N_955,N_611);
nor U1208 (N_1208,N_748,N_900);
xor U1209 (N_1209,N_910,N_749);
nor U1210 (N_1210,N_917,N_738);
or U1211 (N_1211,N_640,N_556);
nand U1212 (N_1212,N_533,N_896);
xnor U1213 (N_1213,N_633,N_722);
xor U1214 (N_1214,N_846,N_737);
nand U1215 (N_1215,N_799,N_934);
and U1216 (N_1216,N_883,N_878);
nand U1217 (N_1217,N_892,N_768);
or U1218 (N_1218,N_734,N_859);
and U1219 (N_1219,N_901,N_572);
or U1220 (N_1220,N_933,N_757);
and U1221 (N_1221,N_945,N_507);
or U1222 (N_1222,N_667,N_960);
and U1223 (N_1223,N_617,N_959);
nor U1224 (N_1224,N_712,N_824);
or U1225 (N_1225,N_931,N_831);
and U1226 (N_1226,N_926,N_596);
and U1227 (N_1227,N_602,N_521);
nor U1228 (N_1228,N_577,N_838);
nand U1229 (N_1229,N_686,N_929);
nor U1230 (N_1230,N_655,N_502);
xnor U1231 (N_1231,N_604,N_545);
or U1232 (N_1232,N_676,N_689);
and U1233 (N_1233,N_804,N_654);
or U1234 (N_1234,N_845,N_726);
or U1235 (N_1235,N_504,N_869);
and U1236 (N_1236,N_639,N_750);
and U1237 (N_1237,N_997,N_938);
or U1238 (N_1238,N_607,N_854);
nand U1239 (N_1239,N_922,N_730);
xor U1240 (N_1240,N_940,N_965);
nor U1241 (N_1241,N_570,N_740);
nand U1242 (N_1242,N_795,N_691);
nor U1243 (N_1243,N_898,N_638);
nand U1244 (N_1244,N_503,N_679);
nor U1245 (N_1245,N_909,N_670);
nor U1246 (N_1246,N_608,N_867);
and U1247 (N_1247,N_879,N_723);
nand U1248 (N_1248,N_948,N_752);
or U1249 (N_1249,N_715,N_781);
nand U1250 (N_1250,N_896,N_664);
and U1251 (N_1251,N_840,N_971);
nand U1252 (N_1252,N_683,N_984);
xor U1253 (N_1253,N_794,N_904);
and U1254 (N_1254,N_579,N_959);
nand U1255 (N_1255,N_575,N_737);
and U1256 (N_1256,N_942,N_553);
and U1257 (N_1257,N_943,N_830);
and U1258 (N_1258,N_560,N_801);
nand U1259 (N_1259,N_863,N_836);
nand U1260 (N_1260,N_798,N_757);
xnor U1261 (N_1261,N_808,N_680);
and U1262 (N_1262,N_945,N_588);
or U1263 (N_1263,N_525,N_664);
nand U1264 (N_1264,N_882,N_948);
or U1265 (N_1265,N_818,N_975);
nor U1266 (N_1266,N_562,N_832);
nor U1267 (N_1267,N_840,N_803);
nand U1268 (N_1268,N_743,N_826);
nand U1269 (N_1269,N_981,N_503);
nor U1270 (N_1270,N_850,N_785);
nand U1271 (N_1271,N_586,N_897);
nand U1272 (N_1272,N_661,N_640);
nor U1273 (N_1273,N_878,N_979);
and U1274 (N_1274,N_631,N_855);
or U1275 (N_1275,N_876,N_659);
nand U1276 (N_1276,N_909,N_897);
nor U1277 (N_1277,N_558,N_794);
or U1278 (N_1278,N_904,N_752);
nand U1279 (N_1279,N_534,N_562);
or U1280 (N_1280,N_892,N_898);
and U1281 (N_1281,N_836,N_780);
and U1282 (N_1282,N_953,N_821);
xnor U1283 (N_1283,N_941,N_583);
and U1284 (N_1284,N_783,N_681);
nand U1285 (N_1285,N_662,N_781);
or U1286 (N_1286,N_938,N_743);
nor U1287 (N_1287,N_936,N_507);
nand U1288 (N_1288,N_803,N_953);
and U1289 (N_1289,N_970,N_759);
and U1290 (N_1290,N_651,N_791);
nand U1291 (N_1291,N_705,N_571);
nor U1292 (N_1292,N_578,N_750);
and U1293 (N_1293,N_691,N_943);
nor U1294 (N_1294,N_634,N_654);
nand U1295 (N_1295,N_775,N_797);
nor U1296 (N_1296,N_677,N_703);
and U1297 (N_1297,N_842,N_746);
xnor U1298 (N_1298,N_921,N_526);
or U1299 (N_1299,N_913,N_530);
nor U1300 (N_1300,N_608,N_718);
and U1301 (N_1301,N_537,N_657);
or U1302 (N_1302,N_734,N_824);
xor U1303 (N_1303,N_743,N_954);
xnor U1304 (N_1304,N_862,N_533);
or U1305 (N_1305,N_648,N_599);
and U1306 (N_1306,N_931,N_756);
or U1307 (N_1307,N_771,N_979);
nand U1308 (N_1308,N_849,N_717);
xnor U1309 (N_1309,N_726,N_583);
and U1310 (N_1310,N_574,N_715);
nor U1311 (N_1311,N_992,N_695);
nor U1312 (N_1312,N_683,N_549);
nand U1313 (N_1313,N_619,N_636);
or U1314 (N_1314,N_829,N_975);
and U1315 (N_1315,N_616,N_841);
nand U1316 (N_1316,N_582,N_927);
nor U1317 (N_1317,N_724,N_876);
or U1318 (N_1318,N_954,N_679);
and U1319 (N_1319,N_719,N_502);
nand U1320 (N_1320,N_840,N_660);
and U1321 (N_1321,N_732,N_813);
nand U1322 (N_1322,N_702,N_798);
nor U1323 (N_1323,N_536,N_939);
nand U1324 (N_1324,N_550,N_979);
nor U1325 (N_1325,N_810,N_950);
and U1326 (N_1326,N_983,N_740);
nand U1327 (N_1327,N_652,N_768);
and U1328 (N_1328,N_612,N_789);
nor U1329 (N_1329,N_553,N_629);
and U1330 (N_1330,N_876,N_819);
nand U1331 (N_1331,N_561,N_889);
xor U1332 (N_1332,N_949,N_851);
or U1333 (N_1333,N_866,N_696);
nand U1334 (N_1334,N_818,N_951);
or U1335 (N_1335,N_844,N_505);
or U1336 (N_1336,N_635,N_916);
nor U1337 (N_1337,N_855,N_951);
nor U1338 (N_1338,N_989,N_699);
nor U1339 (N_1339,N_811,N_949);
and U1340 (N_1340,N_650,N_575);
nor U1341 (N_1341,N_977,N_992);
nand U1342 (N_1342,N_892,N_957);
and U1343 (N_1343,N_996,N_590);
or U1344 (N_1344,N_687,N_564);
or U1345 (N_1345,N_722,N_766);
and U1346 (N_1346,N_875,N_547);
and U1347 (N_1347,N_582,N_762);
nor U1348 (N_1348,N_849,N_781);
and U1349 (N_1349,N_831,N_920);
nand U1350 (N_1350,N_991,N_855);
or U1351 (N_1351,N_879,N_609);
and U1352 (N_1352,N_820,N_863);
nor U1353 (N_1353,N_846,N_629);
nand U1354 (N_1354,N_932,N_739);
nor U1355 (N_1355,N_643,N_518);
or U1356 (N_1356,N_655,N_831);
nand U1357 (N_1357,N_940,N_975);
and U1358 (N_1358,N_848,N_531);
and U1359 (N_1359,N_890,N_516);
nand U1360 (N_1360,N_787,N_702);
or U1361 (N_1361,N_738,N_623);
or U1362 (N_1362,N_968,N_749);
or U1363 (N_1363,N_754,N_728);
or U1364 (N_1364,N_843,N_739);
and U1365 (N_1365,N_526,N_501);
nor U1366 (N_1366,N_972,N_678);
nor U1367 (N_1367,N_539,N_591);
xor U1368 (N_1368,N_537,N_738);
nand U1369 (N_1369,N_569,N_694);
nor U1370 (N_1370,N_757,N_721);
nor U1371 (N_1371,N_932,N_980);
nand U1372 (N_1372,N_549,N_993);
and U1373 (N_1373,N_873,N_832);
nor U1374 (N_1374,N_805,N_896);
and U1375 (N_1375,N_744,N_774);
nand U1376 (N_1376,N_653,N_800);
xor U1377 (N_1377,N_838,N_947);
nor U1378 (N_1378,N_579,N_832);
nor U1379 (N_1379,N_663,N_576);
xnor U1380 (N_1380,N_734,N_706);
and U1381 (N_1381,N_652,N_633);
or U1382 (N_1382,N_533,N_553);
nor U1383 (N_1383,N_722,N_742);
or U1384 (N_1384,N_585,N_900);
or U1385 (N_1385,N_936,N_540);
or U1386 (N_1386,N_690,N_595);
and U1387 (N_1387,N_692,N_969);
xnor U1388 (N_1388,N_622,N_634);
and U1389 (N_1389,N_929,N_606);
or U1390 (N_1390,N_568,N_873);
nor U1391 (N_1391,N_874,N_813);
xor U1392 (N_1392,N_612,N_694);
nand U1393 (N_1393,N_673,N_556);
or U1394 (N_1394,N_950,N_641);
nand U1395 (N_1395,N_512,N_580);
and U1396 (N_1396,N_942,N_854);
or U1397 (N_1397,N_798,N_908);
and U1398 (N_1398,N_842,N_700);
or U1399 (N_1399,N_788,N_577);
xnor U1400 (N_1400,N_689,N_701);
xor U1401 (N_1401,N_719,N_693);
or U1402 (N_1402,N_641,N_535);
nor U1403 (N_1403,N_920,N_847);
or U1404 (N_1404,N_881,N_542);
nand U1405 (N_1405,N_834,N_818);
or U1406 (N_1406,N_528,N_563);
nor U1407 (N_1407,N_909,N_747);
or U1408 (N_1408,N_548,N_784);
xor U1409 (N_1409,N_740,N_836);
or U1410 (N_1410,N_599,N_593);
or U1411 (N_1411,N_667,N_743);
nand U1412 (N_1412,N_672,N_898);
or U1413 (N_1413,N_887,N_738);
nand U1414 (N_1414,N_796,N_690);
or U1415 (N_1415,N_646,N_953);
xnor U1416 (N_1416,N_521,N_802);
or U1417 (N_1417,N_669,N_911);
or U1418 (N_1418,N_754,N_758);
nor U1419 (N_1419,N_808,N_633);
nor U1420 (N_1420,N_724,N_616);
xor U1421 (N_1421,N_755,N_858);
nor U1422 (N_1422,N_906,N_939);
nor U1423 (N_1423,N_980,N_912);
nand U1424 (N_1424,N_889,N_725);
and U1425 (N_1425,N_584,N_618);
xnor U1426 (N_1426,N_984,N_997);
and U1427 (N_1427,N_894,N_753);
or U1428 (N_1428,N_785,N_618);
xnor U1429 (N_1429,N_752,N_575);
nor U1430 (N_1430,N_895,N_891);
nor U1431 (N_1431,N_503,N_639);
and U1432 (N_1432,N_848,N_610);
nor U1433 (N_1433,N_961,N_519);
nand U1434 (N_1434,N_507,N_793);
and U1435 (N_1435,N_950,N_649);
and U1436 (N_1436,N_856,N_556);
nor U1437 (N_1437,N_780,N_541);
or U1438 (N_1438,N_623,N_506);
and U1439 (N_1439,N_605,N_799);
nand U1440 (N_1440,N_901,N_674);
nor U1441 (N_1441,N_857,N_991);
or U1442 (N_1442,N_971,N_919);
nor U1443 (N_1443,N_590,N_865);
xor U1444 (N_1444,N_511,N_605);
or U1445 (N_1445,N_664,N_851);
or U1446 (N_1446,N_643,N_776);
nor U1447 (N_1447,N_740,N_968);
nand U1448 (N_1448,N_902,N_728);
or U1449 (N_1449,N_991,N_979);
nand U1450 (N_1450,N_689,N_672);
and U1451 (N_1451,N_636,N_740);
nand U1452 (N_1452,N_936,N_572);
or U1453 (N_1453,N_973,N_764);
and U1454 (N_1454,N_521,N_985);
nand U1455 (N_1455,N_882,N_885);
nand U1456 (N_1456,N_637,N_860);
nand U1457 (N_1457,N_719,N_659);
or U1458 (N_1458,N_629,N_573);
or U1459 (N_1459,N_845,N_751);
nand U1460 (N_1460,N_910,N_718);
nor U1461 (N_1461,N_502,N_979);
nand U1462 (N_1462,N_920,N_718);
xor U1463 (N_1463,N_899,N_768);
nand U1464 (N_1464,N_597,N_717);
and U1465 (N_1465,N_934,N_591);
nor U1466 (N_1466,N_935,N_686);
and U1467 (N_1467,N_666,N_965);
xor U1468 (N_1468,N_557,N_653);
xor U1469 (N_1469,N_930,N_563);
nor U1470 (N_1470,N_673,N_865);
nor U1471 (N_1471,N_761,N_544);
nand U1472 (N_1472,N_885,N_585);
nor U1473 (N_1473,N_541,N_600);
nor U1474 (N_1474,N_556,N_525);
and U1475 (N_1475,N_575,N_828);
nand U1476 (N_1476,N_515,N_956);
xnor U1477 (N_1477,N_760,N_983);
and U1478 (N_1478,N_653,N_841);
or U1479 (N_1479,N_985,N_810);
and U1480 (N_1480,N_967,N_705);
xnor U1481 (N_1481,N_850,N_722);
xnor U1482 (N_1482,N_801,N_552);
nor U1483 (N_1483,N_682,N_547);
nor U1484 (N_1484,N_731,N_744);
and U1485 (N_1485,N_628,N_950);
nor U1486 (N_1486,N_798,N_647);
or U1487 (N_1487,N_765,N_845);
and U1488 (N_1488,N_699,N_834);
nor U1489 (N_1489,N_794,N_704);
nand U1490 (N_1490,N_756,N_760);
nand U1491 (N_1491,N_937,N_783);
nand U1492 (N_1492,N_606,N_861);
xor U1493 (N_1493,N_610,N_886);
nor U1494 (N_1494,N_539,N_740);
and U1495 (N_1495,N_514,N_958);
and U1496 (N_1496,N_563,N_967);
nor U1497 (N_1497,N_937,N_888);
nand U1498 (N_1498,N_781,N_610);
or U1499 (N_1499,N_565,N_889);
nor U1500 (N_1500,N_1041,N_1371);
or U1501 (N_1501,N_1035,N_1289);
xor U1502 (N_1502,N_1475,N_1384);
or U1503 (N_1503,N_1395,N_1140);
nor U1504 (N_1504,N_1160,N_1147);
nor U1505 (N_1505,N_1150,N_1367);
and U1506 (N_1506,N_1365,N_1252);
nand U1507 (N_1507,N_1232,N_1452);
or U1508 (N_1508,N_1369,N_1443);
or U1509 (N_1509,N_1057,N_1357);
and U1510 (N_1510,N_1014,N_1427);
nand U1511 (N_1511,N_1469,N_1394);
nor U1512 (N_1512,N_1348,N_1319);
nor U1513 (N_1513,N_1176,N_1327);
nor U1514 (N_1514,N_1355,N_1080);
and U1515 (N_1515,N_1163,N_1448);
nand U1516 (N_1516,N_1333,N_1434);
nor U1517 (N_1517,N_1216,N_1105);
or U1518 (N_1518,N_1118,N_1485);
and U1519 (N_1519,N_1456,N_1288);
or U1520 (N_1520,N_1422,N_1330);
or U1521 (N_1521,N_1317,N_1286);
nor U1522 (N_1522,N_1130,N_1197);
nand U1523 (N_1523,N_1438,N_1164);
or U1524 (N_1524,N_1174,N_1334);
or U1525 (N_1525,N_1049,N_1316);
xnor U1526 (N_1526,N_1226,N_1133);
or U1527 (N_1527,N_1496,N_1124);
nor U1528 (N_1528,N_1341,N_1185);
nand U1529 (N_1529,N_1337,N_1213);
and U1530 (N_1530,N_1490,N_1038);
nand U1531 (N_1531,N_1064,N_1137);
nor U1532 (N_1532,N_1378,N_1351);
nand U1533 (N_1533,N_1109,N_1195);
or U1534 (N_1534,N_1476,N_1208);
nor U1535 (N_1535,N_1062,N_1361);
nand U1536 (N_1536,N_1203,N_1396);
or U1537 (N_1537,N_1447,N_1120);
and U1538 (N_1538,N_1444,N_1171);
and U1539 (N_1539,N_1054,N_1007);
xnor U1540 (N_1540,N_1435,N_1240);
and U1541 (N_1541,N_1315,N_1459);
nand U1542 (N_1542,N_1128,N_1220);
nor U1543 (N_1543,N_1373,N_1260);
nand U1544 (N_1544,N_1112,N_1473);
nor U1545 (N_1545,N_1470,N_1324);
and U1546 (N_1546,N_1051,N_1374);
or U1547 (N_1547,N_1217,N_1101);
nand U1548 (N_1548,N_1169,N_1451);
nor U1549 (N_1549,N_1067,N_1186);
nor U1550 (N_1550,N_1097,N_1159);
and U1551 (N_1551,N_1460,N_1403);
and U1552 (N_1552,N_1268,N_1088);
and U1553 (N_1553,N_1425,N_1415);
nor U1554 (N_1554,N_1453,N_1366);
xor U1555 (N_1555,N_1249,N_1360);
nand U1556 (N_1556,N_1295,N_1344);
and U1557 (N_1557,N_1222,N_1497);
nor U1558 (N_1558,N_1023,N_1325);
nand U1559 (N_1559,N_1099,N_1328);
and U1560 (N_1560,N_1000,N_1264);
or U1561 (N_1561,N_1162,N_1257);
xnor U1562 (N_1562,N_1040,N_1441);
or U1563 (N_1563,N_1291,N_1044);
xnor U1564 (N_1564,N_1270,N_1326);
and U1565 (N_1565,N_1281,N_1429);
and U1566 (N_1566,N_1003,N_1407);
nand U1567 (N_1567,N_1294,N_1066);
and U1568 (N_1568,N_1404,N_1179);
nor U1569 (N_1569,N_1034,N_1301);
and U1570 (N_1570,N_1241,N_1078);
nor U1571 (N_1571,N_1290,N_1380);
or U1572 (N_1572,N_1455,N_1103);
or U1573 (N_1573,N_1010,N_1458);
or U1574 (N_1574,N_1206,N_1280);
or U1575 (N_1575,N_1246,N_1187);
nor U1576 (N_1576,N_1022,N_1356);
nand U1577 (N_1577,N_1011,N_1474);
nor U1578 (N_1578,N_1061,N_1091);
nor U1579 (N_1579,N_1461,N_1125);
nor U1580 (N_1580,N_1293,N_1311);
xor U1581 (N_1581,N_1157,N_1214);
nor U1582 (N_1582,N_1183,N_1370);
or U1583 (N_1583,N_1170,N_1030);
and U1584 (N_1584,N_1466,N_1440);
nand U1585 (N_1585,N_1298,N_1234);
or U1586 (N_1586,N_1321,N_1024);
xnor U1587 (N_1587,N_1153,N_1437);
nand U1588 (N_1588,N_1457,N_1012);
nand U1589 (N_1589,N_1494,N_1020);
nand U1590 (N_1590,N_1205,N_1454);
and U1591 (N_1591,N_1306,N_1237);
nand U1592 (N_1592,N_1145,N_1190);
nor U1593 (N_1593,N_1083,N_1383);
or U1594 (N_1594,N_1409,N_1379);
and U1595 (N_1595,N_1184,N_1484);
nor U1596 (N_1596,N_1247,N_1146);
nand U1597 (N_1597,N_1305,N_1221);
nand U1598 (N_1598,N_1292,N_1135);
and U1599 (N_1599,N_1393,N_1063);
nor U1600 (N_1600,N_1148,N_1352);
nand U1601 (N_1601,N_1201,N_1033);
nor U1602 (N_1602,N_1211,N_1047);
nor U1603 (N_1603,N_1055,N_1087);
xnor U1604 (N_1604,N_1028,N_1468);
or U1605 (N_1605,N_1445,N_1006);
and U1606 (N_1606,N_1092,N_1228);
xnor U1607 (N_1607,N_1134,N_1350);
xnor U1608 (N_1608,N_1155,N_1419);
xor U1609 (N_1609,N_1013,N_1483);
nor U1610 (N_1610,N_1359,N_1106);
or U1611 (N_1611,N_1081,N_1102);
nor U1612 (N_1612,N_1271,N_1200);
nor U1613 (N_1613,N_1071,N_1165);
nand U1614 (N_1614,N_1225,N_1412);
nand U1615 (N_1615,N_1230,N_1123);
and U1616 (N_1616,N_1224,N_1115);
or U1617 (N_1617,N_1077,N_1189);
nor U1618 (N_1618,N_1154,N_1262);
nand U1619 (N_1619,N_1245,N_1388);
and U1620 (N_1620,N_1343,N_1110);
and U1621 (N_1621,N_1026,N_1263);
and U1622 (N_1622,N_1486,N_1417);
and U1623 (N_1623,N_1347,N_1482);
nor U1624 (N_1624,N_1242,N_1113);
and U1625 (N_1625,N_1039,N_1089);
or U1626 (N_1626,N_1052,N_1235);
nand U1627 (N_1627,N_1439,N_1219);
nor U1628 (N_1628,N_1210,N_1119);
nand U1629 (N_1629,N_1420,N_1489);
xor U1630 (N_1630,N_1060,N_1336);
or U1631 (N_1631,N_1277,N_1314);
and U1632 (N_1632,N_1107,N_1285);
or U1633 (N_1633,N_1358,N_1131);
xor U1634 (N_1634,N_1032,N_1363);
and U1635 (N_1635,N_1498,N_1266);
nor U1636 (N_1636,N_1025,N_1309);
or U1637 (N_1637,N_1346,N_1495);
nor U1638 (N_1638,N_1430,N_1244);
nand U1639 (N_1639,N_1202,N_1178);
nand U1640 (N_1640,N_1300,N_1181);
nor U1641 (N_1641,N_1094,N_1446);
nand U1642 (N_1642,N_1001,N_1009);
and U1643 (N_1643,N_1215,N_1070);
nor U1644 (N_1644,N_1488,N_1098);
and U1645 (N_1645,N_1273,N_1398);
nor U1646 (N_1646,N_1413,N_1085);
nand U1647 (N_1647,N_1372,N_1046);
nand U1648 (N_1648,N_1076,N_1050);
xor U1649 (N_1649,N_1019,N_1376);
xor U1650 (N_1650,N_1053,N_1467);
or U1651 (N_1651,N_1391,N_1389);
or U1652 (N_1652,N_1307,N_1411);
nand U1653 (N_1653,N_1254,N_1096);
xnor U1654 (N_1654,N_1279,N_1093);
xor U1655 (N_1655,N_1390,N_1037);
nand U1656 (N_1656,N_1255,N_1408);
nor U1657 (N_1657,N_1036,N_1410);
nor U1658 (N_1658,N_1122,N_1045);
nor U1659 (N_1659,N_1068,N_1114);
or U1660 (N_1660,N_1209,N_1168);
or U1661 (N_1661,N_1382,N_1192);
nor U1662 (N_1662,N_1338,N_1079);
xor U1663 (N_1663,N_1303,N_1207);
nand U1664 (N_1664,N_1269,N_1004);
or U1665 (N_1665,N_1199,N_1243);
nor U1666 (N_1666,N_1075,N_1017);
and U1667 (N_1667,N_1354,N_1158);
nor U1668 (N_1668,N_1117,N_1274);
or U1669 (N_1669,N_1177,N_1227);
nand U1670 (N_1670,N_1322,N_1335);
nor U1671 (N_1671,N_1251,N_1223);
nor U1672 (N_1672,N_1231,N_1392);
and U1673 (N_1673,N_1116,N_1016);
or U1674 (N_1674,N_1059,N_1431);
nand U1675 (N_1675,N_1329,N_1141);
and U1676 (N_1676,N_1377,N_1397);
or U1677 (N_1677,N_1250,N_1308);
nor U1678 (N_1678,N_1126,N_1127);
and U1679 (N_1679,N_1381,N_1021);
nand U1680 (N_1680,N_1058,N_1121);
and U1681 (N_1681,N_1471,N_1368);
nor U1682 (N_1682,N_1090,N_1065);
or U1683 (N_1683,N_1188,N_1421);
nand U1684 (N_1684,N_1478,N_1161);
xor U1685 (N_1685,N_1401,N_1212);
and U1686 (N_1686,N_1259,N_1005);
xor U1687 (N_1687,N_1464,N_1275);
nor U1688 (N_1688,N_1072,N_1472);
and U1689 (N_1689,N_1084,N_1043);
nor U1690 (N_1690,N_1320,N_1256);
or U1691 (N_1691,N_1276,N_1287);
and U1692 (N_1692,N_1074,N_1129);
nor U1693 (N_1693,N_1175,N_1082);
nand U1694 (N_1694,N_1349,N_1493);
nor U1695 (N_1695,N_1139,N_1191);
nor U1696 (N_1696,N_1152,N_1104);
nand U1697 (N_1697,N_1239,N_1364);
and U1698 (N_1698,N_1265,N_1339);
and U1699 (N_1699,N_1193,N_1151);
and U1700 (N_1700,N_1302,N_1402);
nand U1701 (N_1701,N_1149,N_1198);
and U1702 (N_1702,N_1172,N_1428);
or U1703 (N_1703,N_1166,N_1436);
nand U1704 (N_1704,N_1282,N_1462);
and U1705 (N_1705,N_1386,N_1353);
xor U1706 (N_1706,N_1424,N_1048);
nand U1707 (N_1707,N_1414,N_1296);
nand U1708 (N_1708,N_1233,N_1261);
nor U1709 (N_1709,N_1313,N_1056);
nand U1710 (N_1710,N_1156,N_1465);
nor U1711 (N_1711,N_1086,N_1433);
and U1712 (N_1712,N_1399,N_1267);
and U1713 (N_1713,N_1229,N_1108);
or U1714 (N_1714,N_1111,N_1018);
and U1715 (N_1715,N_1432,N_1480);
and U1716 (N_1716,N_1304,N_1238);
nor U1717 (N_1717,N_1463,N_1069);
and U1718 (N_1718,N_1132,N_1312);
nand U1719 (N_1719,N_1385,N_1008);
nand U1720 (N_1720,N_1442,N_1318);
nand U1721 (N_1721,N_1073,N_1477);
or U1722 (N_1722,N_1095,N_1499);
xor U1723 (N_1723,N_1491,N_1180);
and U1724 (N_1724,N_1297,N_1387);
or U1725 (N_1725,N_1345,N_1167);
nand U1726 (N_1726,N_1218,N_1029);
nor U1727 (N_1727,N_1342,N_1027);
nor U1728 (N_1728,N_1299,N_1418);
or U1729 (N_1729,N_1492,N_1406);
nand U1730 (N_1730,N_1258,N_1002);
nand U1731 (N_1731,N_1331,N_1015);
nand U1732 (N_1732,N_1487,N_1143);
xor U1733 (N_1733,N_1194,N_1196);
and U1734 (N_1734,N_1362,N_1031);
xnor U1735 (N_1735,N_1278,N_1481);
or U1736 (N_1736,N_1248,N_1173);
nor U1737 (N_1737,N_1253,N_1284);
and U1738 (N_1738,N_1204,N_1405);
or U1739 (N_1739,N_1182,N_1332);
or U1740 (N_1740,N_1136,N_1449);
and U1741 (N_1741,N_1375,N_1272);
xnor U1742 (N_1742,N_1416,N_1144);
or U1743 (N_1743,N_1042,N_1479);
and U1744 (N_1744,N_1236,N_1310);
or U1745 (N_1745,N_1426,N_1283);
nor U1746 (N_1746,N_1340,N_1100);
nand U1747 (N_1747,N_1400,N_1423);
xnor U1748 (N_1748,N_1323,N_1142);
nand U1749 (N_1749,N_1138,N_1450);
or U1750 (N_1750,N_1456,N_1418);
xnor U1751 (N_1751,N_1243,N_1153);
xnor U1752 (N_1752,N_1222,N_1266);
or U1753 (N_1753,N_1433,N_1101);
xnor U1754 (N_1754,N_1295,N_1382);
and U1755 (N_1755,N_1250,N_1356);
xnor U1756 (N_1756,N_1353,N_1411);
or U1757 (N_1757,N_1098,N_1467);
nand U1758 (N_1758,N_1317,N_1229);
nand U1759 (N_1759,N_1302,N_1222);
nor U1760 (N_1760,N_1160,N_1173);
or U1761 (N_1761,N_1042,N_1194);
nand U1762 (N_1762,N_1297,N_1489);
and U1763 (N_1763,N_1246,N_1001);
and U1764 (N_1764,N_1405,N_1238);
nor U1765 (N_1765,N_1013,N_1253);
nor U1766 (N_1766,N_1259,N_1051);
or U1767 (N_1767,N_1217,N_1412);
or U1768 (N_1768,N_1319,N_1133);
and U1769 (N_1769,N_1432,N_1106);
nand U1770 (N_1770,N_1154,N_1316);
nor U1771 (N_1771,N_1010,N_1029);
nand U1772 (N_1772,N_1422,N_1230);
nor U1773 (N_1773,N_1164,N_1283);
nor U1774 (N_1774,N_1262,N_1444);
nand U1775 (N_1775,N_1190,N_1259);
and U1776 (N_1776,N_1376,N_1295);
or U1777 (N_1777,N_1235,N_1063);
and U1778 (N_1778,N_1375,N_1345);
nand U1779 (N_1779,N_1295,N_1279);
and U1780 (N_1780,N_1202,N_1457);
nor U1781 (N_1781,N_1220,N_1211);
nor U1782 (N_1782,N_1412,N_1091);
nor U1783 (N_1783,N_1377,N_1412);
nor U1784 (N_1784,N_1249,N_1083);
and U1785 (N_1785,N_1169,N_1496);
nor U1786 (N_1786,N_1422,N_1406);
or U1787 (N_1787,N_1309,N_1391);
nand U1788 (N_1788,N_1269,N_1027);
xor U1789 (N_1789,N_1351,N_1387);
nor U1790 (N_1790,N_1041,N_1062);
nor U1791 (N_1791,N_1214,N_1357);
xor U1792 (N_1792,N_1459,N_1108);
nor U1793 (N_1793,N_1336,N_1476);
xnor U1794 (N_1794,N_1165,N_1095);
nand U1795 (N_1795,N_1242,N_1481);
and U1796 (N_1796,N_1206,N_1155);
xor U1797 (N_1797,N_1405,N_1240);
nor U1798 (N_1798,N_1361,N_1007);
nand U1799 (N_1799,N_1109,N_1444);
and U1800 (N_1800,N_1476,N_1051);
nand U1801 (N_1801,N_1029,N_1451);
and U1802 (N_1802,N_1346,N_1403);
nand U1803 (N_1803,N_1303,N_1103);
nor U1804 (N_1804,N_1045,N_1080);
nand U1805 (N_1805,N_1354,N_1487);
or U1806 (N_1806,N_1451,N_1020);
or U1807 (N_1807,N_1098,N_1013);
or U1808 (N_1808,N_1161,N_1066);
or U1809 (N_1809,N_1395,N_1124);
and U1810 (N_1810,N_1313,N_1373);
nand U1811 (N_1811,N_1440,N_1010);
nand U1812 (N_1812,N_1499,N_1433);
nor U1813 (N_1813,N_1100,N_1184);
or U1814 (N_1814,N_1284,N_1035);
or U1815 (N_1815,N_1419,N_1104);
and U1816 (N_1816,N_1450,N_1230);
nand U1817 (N_1817,N_1471,N_1297);
or U1818 (N_1818,N_1092,N_1005);
or U1819 (N_1819,N_1386,N_1190);
or U1820 (N_1820,N_1305,N_1493);
and U1821 (N_1821,N_1130,N_1122);
and U1822 (N_1822,N_1212,N_1047);
and U1823 (N_1823,N_1289,N_1103);
nand U1824 (N_1824,N_1435,N_1181);
xor U1825 (N_1825,N_1348,N_1197);
and U1826 (N_1826,N_1343,N_1182);
nand U1827 (N_1827,N_1088,N_1299);
and U1828 (N_1828,N_1309,N_1010);
and U1829 (N_1829,N_1162,N_1087);
and U1830 (N_1830,N_1053,N_1459);
nor U1831 (N_1831,N_1464,N_1251);
and U1832 (N_1832,N_1046,N_1445);
nor U1833 (N_1833,N_1046,N_1462);
nand U1834 (N_1834,N_1108,N_1064);
or U1835 (N_1835,N_1312,N_1298);
nor U1836 (N_1836,N_1494,N_1257);
and U1837 (N_1837,N_1114,N_1338);
nor U1838 (N_1838,N_1374,N_1129);
nand U1839 (N_1839,N_1461,N_1488);
nand U1840 (N_1840,N_1215,N_1048);
nand U1841 (N_1841,N_1445,N_1352);
xnor U1842 (N_1842,N_1137,N_1357);
or U1843 (N_1843,N_1299,N_1001);
and U1844 (N_1844,N_1218,N_1095);
nand U1845 (N_1845,N_1103,N_1165);
nand U1846 (N_1846,N_1045,N_1232);
nand U1847 (N_1847,N_1132,N_1428);
and U1848 (N_1848,N_1313,N_1101);
or U1849 (N_1849,N_1373,N_1024);
and U1850 (N_1850,N_1112,N_1375);
and U1851 (N_1851,N_1187,N_1280);
nor U1852 (N_1852,N_1432,N_1406);
xnor U1853 (N_1853,N_1332,N_1071);
nor U1854 (N_1854,N_1418,N_1167);
or U1855 (N_1855,N_1242,N_1098);
and U1856 (N_1856,N_1410,N_1300);
nand U1857 (N_1857,N_1087,N_1298);
and U1858 (N_1858,N_1294,N_1269);
nor U1859 (N_1859,N_1327,N_1495);
and U1860 (N_1860,N_1063,N_1456);
nor U1861 (N_1861,N_1429,N_1161);
and U1862 (N_1862,N_1154,N_1258);
nor U1863 (N_1863,N_1402,N_1076);
nand U1864 (N_1864,N_1184,N_1182);
nor U1865 (N_1865,N_1173,N_1133);
nand U1866 (N_1866,N_1039,N_1299);
and U1867 (N_1867,N_1302,N_1130);
and U1868 (N_1868,N_1367,N_1336);
nor U1869 (N_1869,N_1455,N_1087);
nand U1870 (N_1870,N_1495,N_1254);
and U1871 (N_1871,N_1020,N_1116);
xor U1872 (N_1872,N_1437,N_1364);
or U1873 (N_1873,N_1078,N_1405);
and U1874 (N_1874,N_1076,N_1406);
and U1875 (N_1875,N_1088,N_1155);
and U1876 (N_1876,N_1352,N_1293);
or U1877 (N_1877,N_1407,N_1088);
or U1878 (N_1878,N_1442,N_1263);
nand U1879 (N_1879,N_1243,N_1023);
and U1880 (N_1880,N_1276,N_1396);
or U1881 (N_1881,N_1475,N_1009);
and U1882 (N_1882,N_1034,N_1368);
xor U1883 (N_1883,N_1011,N_1286);
nand U1884 (N_1884,N_1424,N_1263);
nand U1885 (N_1885,N_1475,N_1218);
or U1886 (N_1886,N_1154,N_1430);
and U1887 (N_1887,N_1018,N_1379);
and U1888 (N_1888,N_1210,N_1322);
nand U1889 (N_1889,N_1361,N_1249);
nand U1890 (N_1890,N_1454,N_1199);
nand U1891 (N_1891,N_1388,N_1267);
nor U1892 (N_1892,N_1453,N_1075);
and U1893 (N_1893,N_1495,N_1208);
or U1894 (N_1894,N_1397,N_1468);
nor U1895 (N_1895,N_1088,N_1325);
and U1896 (N_1896,N_1463,N_1080);
nor U1897 (N_1897,N_1399,N_1152);
xor U1898 (N_1898,N_1297,N_1159);
or U1899 (N_1899,N_1043,N_1382);
and U1900 (N_1900,N_1049,N_1071);
nor U1901 (N_1901,N_1188,N_1326);
nand U1902 (N_1902,N_1467,N_1175);
or U1903 (N_1903,N_1177,N_1076);
xnor U1904 (N_1904,N_1032,N_1277);
nand U1905 (N_1905,N_1063,N_1126);
or U1906 (N_1906,N_1100,N_1290);
and U1907 (N_1907,N_1406,N_1147);
or U1908 (N_1908,N_1047,N_1209);
nand U1909 (N_1909,N_1320,N_1123);
and U1910 (N_1910,N_1058,N_1189);
nand U1911 (N_1911,N_1246,N_1212);
nor U1912 (N_1912,N_1121,N_1302);
or U1913 (N_1913,N_1002,N_1094);
and U1914 (N_1914,N_1022,N_1324);
or U1915 (N_1915,N_1100,N_1094);
or U1916 (N_1916,N_1409,N_1416);
nand U1917 (N_1917,N_1104,N_1125);
and U1918 (N_1918,N_1342,N_1133);
or U1919 (N_1919,N_1374,N_1196);
nor U1920 (N_1920,N_1416,N_1476);
and U1921 (N_1921,N_1474,N_1473);
or U1922 (N_1922,N_1225,N_1256);
and U1923 (N_1923,N_1088,N_1273);
and U1924 (N_1924,N_1307,N_1173);
nor U1925 (N_1925,N_1147,N_1339);
nand U1926 (N_1926,N_1461,N_1272);
or U1927 (N_1927,N_1086,N_1082);
nand U1928 (N_1928,N_1214,N_1388);
nor U1929 (N_1929,N_1288,N_1372);
and U1930 (N_1930,N_1147,N_1411);
nand U1931 (N_1931,N_1416,N_1264);
nand U1932 (N_1932,N_1398,N_1349);
nor U1933 (N_1933,N_1260,N_1086);
and U1934 (N_1934,N_1342,N_1468);
or U1935 (N_1935,N_1263,N_1176);
or U1936 (N_1936,N_1406,N_1457);
and U1937 (N_1937,N_1020,N_1429);
nor U1938 (N_1938,N_1220,N_1124);
nand U1939 (N_1939,N_1434,N_1069);
nand U1940 (N_1940,N_1143,N_1097);
or U1941 (N_1941,N_1165,N_1037);
nand U1942 (N_1942,N_1104,N_1160);
or U1943 (N_1943,N_1180,N_1220);
or U1944 (N_1944,N_1230,N_1393);
and U1945 (N_1945,N_1341,N_1251);
or U1946 (N_1946,N_1326,N_1341);
nand U1947 (N_1947,N_1321,N_1105);
and U1948 (N_1948,N_1225,N_1454);
or U1949 (N_1949,N_1346,N_1190);
or U1950 (N_1950,N_1281,N_1326);
nor U1951 (N_1951,N_1089,N_1213);
nor U1952 (N_1952,N_1297,N_1152);
nand U1953 (N_1953,N_1222,N_1404);
nand U1954 (N_1954,N_1332,N_1133);
or U1955 (N_1955,N_1306,N_1331);
and U1956 (N_1956,N_1202,N_1375);
nor U1957 (N_1957,N_1025,N_1282);
xor U1958 (N_1958,N_1146,N_1214);
nand U1959 (N_1959,N_1230,N_1069);
nand U1960 (N_1960,N_1090,N_1494);
nand U1961 (N_1961,N_1477,N_1458);
and U1962 (N_1962,N_1478,N_1134);
nor U1963 (N_1963,N_1319,N_1067);
and U1964 (N_1964,N_1009,N_1350);
nand U1965 (N_1965,N_1372,N_1016);
nor U1966 (N_1966,N_1462,N_1060);
and U1967 (N_1967,N_1317,N_1182);
and U1968 (N_1968,N_1048,N_1482);
and U1969 (N_1969,N_1373,N_1309);
or U1970 (N_1970,N_1186,N_1188);
or U1971 (N_1971,N_1121,N_1341);
nor U1972 (N_1972,N_1305,N_1263);
and U1973 (N_1973,N_1252,N_1026);
xnor U1974 (N_1974,N_1412,N_1374);
and U1975 (N_1975,N_1207,N_1069);
nand U1976 (N_1976,N_1329,N_1170);
nor U1977 (N_1977,N_1027,N_1215);
or U1978 (N_1978,N_1346,N_1052);
nor U1979 (N_1979,N_1398,N_1298);
or U1980 (N_1980,N_1395,N_1183);
nor U1981 (N_1981,N_1206,N_1040);
nor U1982 (N_1982,N_1394,N_1059);
nor U1983 (N_1983,N_1185,N_1463);
or U1984 (N_1984,N_1333,N_1163);
and U1985 (N_1985,N_1026,N_1283);
and U1986 (N_1986,N_1010,N_1122);
nor U1987 (N_1987,N_1206,N_1435);
or U1988 (N_1988,N_1115,N_1325);
or U1989 (N_1989,N_1366,N_1055);
nor U1990 (N_1990,N_1112,N_1350);
xor U1991 (N_1991,N_1395,N_1297);
nand U1992 (N_1992,N_1023,N_1448);
xnor U1993 (N_1993,N_1020,N_1147);
and U1994 (N_1994,N_1051,N_1483);
or U1995 (N_1995,N_1380,N_1276);
nor U1996 (N_1996,N_1352,N_1372);
nand U1997 (N_1997,N_1419,N_1378);
xnor U1998 (N_1998,N_1040,N_1182);
nand U1999 (N_1999,N_1181,N_1194);
nand U2000 (N_2000,N_1893,N_1990);
xor U2001 (N_2001,N_1996,N_1519);
nor U2002 (N_2002,N_1634,N_1584);
or U2003 (N_2003,N_1505,N_1909);
or U2004 (N_2004,N_1737,N_1745);
and U2005 (N_2005,N_1550,N_1541);
and U2006 (N_2006,N_1768,N_1794);
nor U2007 (N_2007,N_1670,N_1774);
or U2008 (N_2008,N_1583,N_1718);
and U2009 (N_2009,N_1714,N_1753);
nor U2010 (N_2010,N_1624,N_1559);
or U2011 (N_2011,N_1651,N_1594);
nand U2012 (N_2012,N_1972,N_1969);
nor U2013 (N_2013,N_1540,N_1925);
and U2014 (N_2014,N_1542,N_1915);
nand U2015 (N_2015,N_1604,N_1770);
nor U2016 (N_2016,N_1784,N_1952);
nand U2017 (N_2017,N_1937,N_1597);
or U2018 (N_2018,N_1611,N_1798);
xor U2019 (N_2019,N_1892,N_1942);
xor U2020 (N_2020,N_1822,N_1772);
nor U2021 (N_2021,N_1631,N_1521);
or U2022 (N_2022,N_1810,N_1852);
nor U2023 (N_2023,N_1544,N_1755);
and U2024 (N_2024,N_1730,N_1527);
or U2025 (N_2025,N_1586,N_1968);
and U2026 (N_2026,N_1535,N_1713);
nand U2027 (N_2027,N_1816,N_1648);
nand U2028 (N_2028,N_1639,N_1865);
and U2029 (N_2029,N_1828,N_1596);
or U2030 (N_2030,N_1791,N_1543);
nand U2031 (N_2031,N_1805,N_1802);
or U2032 (N_2032,N_1607,N_1979);
or U2033 (N_2033,N_1891,N_1684);
xnor U2034 (N_2034,N_1855,N_1556);
nand U2035 (N_2035,N_1613,N_1854);
nand U2036 (N_2036,N_1553,N_1970);
or U2037 (N_2037,N_1652,N_1796);
xnor U2038 (N_2038,N_1832,N_1529);
or U2039 (N_2039,N_1633,N_1610);
and U2040 (N_2040,N_1706,N_1693);
or U2041 (N_2041,N_1803,N_1766);
nor U2042 (N_2042,N_1973,N_1675);
or U2043 (N_2043,N_1691,N_1662);
nor U2044 (N_2044,N_1821,N_1819);
nor U2045 (N_2045,N_1874,N_1643);
or U2046 (N_2046,N_1524,N_1710);
or U2047 (N_2047,N_1621,N_1561);
or U2048 (N_2048,N_1692,N_1590);
nor U2049 (N_2049,N_1548,N_1762);
nor U2050 (N_2050,N_1956,N_1917);
nor U2051 (N_2051,N_1726,N_1653);
or U2052 (N_2052,N_1789,N_1797);
nor U2053 (N_2053,N_1793,N_1674);
and U2054 (N_2054,N_1767,N_1575);
xor U2055 (N_2055,N_1589,N_1904);
nor U2056 (N_2056,N_1506,N_1591);
nor U2057 (N_2057,N_1955,N_1786);
and U2058 (N_2058,N_1871,N_1655);
and U2059 (N_2059,N_1598,N_1775);
or U2060 (N_2060,N_1567,N_1962);
xor U2061 (N_2061,N_1795,N_1649);
or U2062 (N_2062,N_1830,N_1509);
or U2063 (N_2063,N_1659,N_1685);
nand U2064 (N_2064,N_1546,N_1729);
nor U2065 (N_2065,N_1637,N_1841);
and U2066 (N_2066,N_1552,N_1974);
nand U2067 (N_2067,N_1698,N_1769);
nor U2068 (N_2068,N_1587,N_1715);
nand U2069 (N_2069,N_1950,N_1987);
nand U2070 (N_2070,N_1977,N_1924);
or U2071 (N_2071,N_1686,N_1688);
or U2072 (N_2072,N_1673,N_1627);
or U2073 (N_2073,N_1751,N_1885);
xor U2074 (N_2074,N_1746,N_1672);
or U2075 (N_2075,N_1733,N_1824);
nand U2076 (N_2076,N_1579,N_1890);
and U2077 (N_2077,N_1765,N_1616);
nand U2078 (N_2078,N_1554,N_1776);
xnor U2079 (N_2079,N_1750,N_1603);
xor U2080 (N_2080,N_1878,N_1916);
nor U2081 (N_2081,N_1933,N_1964);
nand U2082 (N_2082,N_1787,N_1722);
and U2083 (N_2083,N_1630,N_1880);
or U2084 (N_2084,N_1581,N_1719);
and U2085 (N_2085,N_1833,N_1615);
and U2086 (N_2086,N_1941,N_1985);
or U2087 (N_2087,N_1981,N_1759);
or U2088 (N_2088,N_1504,N_1600);
nor U2089 (N_2089,N_1647,N_1585);
nand U2090 (N_2090,N_1839,N_1758);
nor U2091 (N_2091,N_1635,N_1701);
nor U2092 (N_2092,N_1592,N_1809);
nand U2093 (N_2093,N_1831,N_1568);
nor U2094 (N_2094,N_1522,N_1626);
or U2095 (N_2095,N_1571,N_1677);
nand U2096 (N_2096,N_1945,N_1650);
and U2097 (N_2097,N_1682,N_1953);
and U2098 (N_2098,N_1525,N_1728);
nor U2099 (N_2099,N_1551,N_1507);
and U2100 (N_2100,N_1708,N_1593);
nand U2101 (N_2101,N_1947,N_1752);
and U2102 (N_2102,N_1864,N_1994);
nand U2103 (N_2103,N_1837,N_1760);
or U2104 (N_2104,N_1508,N_1595);
nor U2105 (N_2105,N_1898,N_1939);
and U2106 (N_2106,N_1560,N_1608);
nand U2107 (N_2107,N_1599,N_1573);
or U2108 (N_2108,N_1811,N_1853);
nand U2109 (N_2109,N_1920,N_1788);
or U2110 (N_2110,N_1748,N_1857);
xor U2111 (N_2111,N_1804,N_1623);
nand U2112 (N_2112,N_1842,N_1515);
and U2113 (N_2113,N_1518,N_1817);
and U2114 (N_2114,N_1702,N_1834);
and U2115 (N_2115,N_1886,N_1761);
nor U2116 (N_2116,N_1922,N_1547);
or U2117 (N_2117,N_1948,N_1875);
nand U2118 (N_2118,N_1844,N_1533);
nand U2119 (N_2119,N_1888,N_1840);
xor U2120 (N_2120,N_1849,N_1555);
and U2121 (N_2121,N_1929,N_1982);
nor U2122 (N_2122,N_1792,N_1778);
nand U2123 (N_2123,N_1731,N_1618);
or U2124 (N_2124,N_1724,N_1565);
nand U2125 (N_2125,N_1779,N_1712);
nand U2126 (N_2126,N_1502,N_1666);
nand U2127 (N_2127,N_1870,N_1873);
nor U2128 (N_2128,N_1738,N_1602);
or U2129 (N_2129,N_1928,N_1539);
xor U2130 (N_2130,N_1869,N_1850);
and U2131 (N_2131,N_1995,N_1801);
and U2132 (N_2132,N_1520,N_1757);
nand U2133 (N_2133,N_1658,N_1512);
nor U2134 (N_2134,N_1534,N_1894);
and U2135 (N_2135,N_1771,N_1903);
nor U2136 (N_2136,N_1663,N_1829);
and U2137 (N_2137,N_1967,N_1808);
nor U2138 (N_2138,N_1989,N_1545);
or U2139 (N_2139,N_1669,N_1566);
nand U2140 (N_2140,N_1697,N_1911);
nand U2141 (N_2141,N_1835,N_1501);
nor U2142 (N_2142,N_1934,N_1511);
and U2143 (N_2143,N_1935,N_1636);
nand U2144 (N_2144,N_1656,N_1763);
nand U2145 (N_2145,N_1695,N_1689);
or U2146 (N_2146,N_1851,N_1734);
and U2147 (N_2147,N_1510,N_1913);
nor U2148 (N_2148,N_1998,N_1879);
or U2149 (N_2149,N_1707,N_1676);
nand U2150 (N_2150,N_1951,N_1971);
nor U2151 (N_2151,N_1667,N_1881);
or U2152 (N_2152,N_1743,N_1699);
and U2153 (N_2153,N_1632,N_1619);
xor U2154 (N_2154,N_1749,N_1780);
or U2155 (N_2155,N_1912,N_1537);
xor U2156 (N_2156,N_1711,N_1826);
nor U2157 (N_2157,N_1988,N_1843);
xnor U2158 (N_2158,N_1949,N_1739);
nor U2159 (N_2159,N_1740,N_1961);
nand U2160 (N_2160,N_1862,N_1549);
nor U2161 (N_2161,N_1813,N_1896);
or U2162 (N_2162,N_1687,N_1580);
and U2163 (N_2163,N_1668,N_1984);
xnor U2164 (N_2164,N_1946,N_1642);
nor U2165 (N_2165,N_1628,N_1754);
and U2166 (N_2166,N_1516,N_1742);
and U2167 (N_2167,N_1756,N_1577);
nor U2168 (N_2168,N_1721,N_1578);
nor U2169 (N_2169,N_1538,N_1572);
xor U2170 (N_2170,N_1965,N_1908);
nor U2171 (N_2171,N_1694,N_1944);
or U2172 (N_2172,N_1536,N_1806);
nor U2173 (N_2173,N_1918,N_1563);
nor U2174 (N_2174,N_1785,N_1588);
nor U2175 (N_2175,N_1861,N_1679);
or U2176 (N_2176,N_1847,N_1836);
nor U2177 (N_2177,N_1732,N_1601);
nor U2178 (N_2178,N_1725,N_1680);
xnor U2179 (N_2179,N_1901,N_1897);
nor U2180 (N_2180,N_1859,N_1614);
nand U2181 (N_2181,N_1564,N_1605);
and U2182 (N_2182,N_1863,N_1856);
or U2183 (N_2183,N_1558,N_1993);
and U2184 (N_2184,N_1902,N_1514);
or U2185 (N_2185,N_1530,N_1629);
or U2186 (N_2186,N_1528,N_1976);
nand U2187 (N_2187,N_1526,N_1884);
and U2188 (N_2188,N_1954,N_1921);
or U2189 (N_2189,N_1574,N_1696);
nand U2190 (N_2190,N_1709,N_1531);
nor U2191 (N_2191,N_1503,N_1704);
and U2192 (N_2192,N_1815,N_1899);
xor U2193 (N_2193,N_1997,N_1930);
xnor U2194 (N_2194,N_1609,N_1812);
and U2195 (N_2195,N_1943,N_1741);
and U2196 (N_2196,N_1678,N_1764);
xor U2197 (N_2197,N_1638,N_1654);
or U2198 (N_2198,N_1848,N_1958);
nor U2199 (N_2199,N_1681,N_1716);
nor U2200 (N_2200,N_1700,N_1523);
nor U2201 (N_2201,N_1980,N_1957);
nand U2202 (N_2202,N_1661,N_1646);
xnor U2203 (N_2203,N_1622,N_1513);
xor U2204 (N_2204,N_1705,N_1999);
or U2205 (N_2205,N_1986,N_1877);
or U2206 (N_2206,N_1966,N_1790);
nand U2207 (N_2207,N_1895,N_1781);
nand U2208 (N_2208,N_1959,N_1889);
xor U2209 (N_2209,N_1906,N_1910);
nor U2210 (N_2210,N_1747,N_1690);
or U2211 (N_2211,N_1671,N_1625);
nand U2212 (N_2212,N_1978,N_1991);
or U2213 (N_2213,N_1975,N_1807);
nand U2214 (N_2214,N_1825,N_1872);
nand U2215 (N_2215,N_1620,N_1683);
and U2216 (N_2216,N_1644,N_1799);
xnor U2217 (N_2217,N_1983,N_1645);
and U2218 (N_2218,N_1818,N_1938);
and U2219 (N_2219,N_1612,N_1919);
nand U2220 (N_2220,N_1783,N_1744);
or U2221 (N_2221,N_1882,N_1569);
nor U2222 (N_2222,N_1582,N_1777);
xor U2223 (N_2223,N_1992,N_1641);
nand U2224 (N_2224,N_1500,N_1867);
nand U2225 (N_2225,N_1838,N_1963);
or U2226 (N_2226,N_1665,N_1823);
nor U2227 (N_2227,N_1723,N_1814);
xnor U2228 (N_2228,N_1782,N_1570);
nand U2229 (N_2229,N_1905,N_1517);
xnor U2230 (N_2230,N_1703,N_1932);
and U2231 (N_2231,N_1926,N_1660);
xnor U2232 (N_2232,N_1914,N_1735);
nor U2233 (N_2233,N_1820,N_1845);
or U2234 (N_2234,N_1562,N_1576);
nor U2235 (N_2235,N_1773,N_1736);
or U2236 (N_2236,N_1720,N_1927);
nor U2237 (N_2237,N_1907,N_1868);
nand U2238 (N_2238,N_1640,N_1923);
nand U2239 (N_2239,N_1960,N_1800);
nand U2240 (N_2240,N_1883,N_1617);
nand U2241 (N_2241,N_1532,N_1940);
xor U2242 (N_2242,N_1664,N_1846);
or U2243 (N_2243,N_1900,N_1866);
nand U2244 (N_2244,N_1860,N_1876);
nand U2245 (N_2245,N_1727,N_1557);
or U2246 (N_2246,N_1858,N_1657);
or U2247 (N_2247,N_1931,N_1936);
nor U2248 (N_2248,N_1887,N_1827);
nand U2249 (N_2249,N_1606,N_1717);
nor U2250 (N_2250,N_1676,N_1512);
xor U2251 (N_2251,N_1717,N_1629);
and U2252 (N_2252,N_1913,N_1940);
or U2253 (N_2253,N_1794,N_1773);
or U2254 (N_2254,N_1983,N_1878);
or U2255 (N_2255,N_1596,N_1722);
or U2256 (N_2256,N_1625,N_1812);
nand U2257 (N_2257,N_1627,N_1612);
and U2258 (N_2258,N_1737,N_1899);
xor U2259 (N_2259,N_1825,N_1866);
and U2260 (N_2260,N_1745,N_1627);
nor U2261 (N_2261,N_1997,N_1826);
nor U2262 (N_2262,N_1885,N_1594);
and U2263 (N_2263,N_1565,N_1607);
nand U2264 (N_2264,N_1972,N_1661);
nand U2265 (N_2265,N_1781,N_1897);
or U2266 (N_2266,N_1632,N_1618);
and U2267 (N_2267,N_1858,N_1891);
nor U2268 (N_2268,N_1744,N_1632);
nand U2269 (N_2269,N_1690,N_1938);
xnor U2270 (N_2270,N_1952,N_1914);
nand U2271 (N_2271,N_1921,N_1812);
or U2272 (N_2272,N_1993,N_1561);
xnor U2273 (N_2273,N_1585,N_1595);
nor U2274 (N_2274,N_1542,N_1875);
nor U2275 (N_2275,N_1719,N_1890);
xor U2276 (N_2276,N_1685,N_1820);
or U2277 (N_2277,N_1567,N_1569);
or U2278 (N_2278,N_1543,N_1680);
or U2279 (N_2279,N_1937,N_1680);
or U2280 (N_2280,N_1781,N_1505);
or U2281 (N_2281,N_1899,N_1703);
nor U2282 (N_2282,N_1505,N_1511);
and U2283 (N_2283,N_1856,N_1814);
nand U2284 (N_2284,N_1603,N_1593);
and U2285 (N_2285,N_1586,N_1832);
and U2286 (N_2286,N_1713,N_1815);
xor U2287 (N_2287,N_1911,N_1527);
and U2288 (N_2288,N_1692,N_1788);
nor U2289 (N_2289,N_1686,N_1559);
or U2290 (N_2290,N_1653,N_1644);
nand U2291 (N_2291,N_1558,N_1829);
nor U2292 (N_2292,N_1954,N_1625);
or U2293 (N_2293,N_1834,N_1749);
or U2294 (N_2294,N_1828,N_1584);
and U2295 (N_2295,N_1737,N_1688);
nand U2296 (N_2296,N_1825,N_1514);
nand U2297 (N_2297,N_1987,N_1630);
or U2298 (N_2298,N_1675,N_1924);
xnor U2299 (N_2299,N_1533,N_1512);
nor U2300 (N_2300,N_1510,N_1617);
and U2301 (N_2301,N_1851,N_1607);
xnor U2302 (N_2302,N_1731,N_1975);
or U2303 (N_2303,N_1510,N_1585);
and U2304 (N_2304,N_1608,N_1987);
nand U2305 (N_2305,N_1510,N_1909);
nand U2306 (N_2306,N_1632,N_1637);
or U2307 (N_2307,N_1933,N_1839);
and U2308 (N_2308,N_1852,N_1668);
or U2309 (N_2309,N_1748,N_1970);
nor U2310 (N_2310,N_1536,N_1880);
nor U2311 (N_2311,N_1916,N_1512);
or U2312 (N_2312,N_1756,N_1751);
or U2313 (N_2313,N_1974,N_1936);
and U2314 (N_2314,N_1779,N_1785);
and U2315 (N_2315,N_1972,N_1925);
nor U2316 (N_2316,N_1513,N_1989);
nor U2317 (N_2317,N_1725,N_1860);
nor U2318 (N_2318,N_1874,N_1861);
or U2319 (N_2319,N_1546,N_1963);
or U2320 (N_2320,N_1847,N_1586);
nor U2321 (N_2321,N_1960,N_1900);
or U2322 (N_2322,N_1715,N_1921);
or U2323 (N_2323,N_1863,N_1604);
or U2324 (N_2324,N_1561,N_1988);
or U2325 (N_2325,N_1623,N_1890);
or U2326 (N_2326,N_1660,N_1861);
nand U2327 (N_2327,N_1689,N_1913);
or U2328 (N_2328,N_1756,N_1878);
nand U2329 (N_2329,N_1768,N_1781);
and U2330 (N_2330,N_1639,N_1789);
nor U2331 (N_2331,N_1994,N_1524);
xnor U2332 (N_2332,N_1542,N_1917);
nor U2333 (N_2333,N_1967,N_1986);
nor U2334 (N_2334,N_1939,N_1714);
or U2335 (N_2335,N_1738,N_1941);
nand U2336 (N_2336,N_1891,N_1647);
and U2337 (N_2337,N_1859,N_1740);
xor U2338 (N_2338,N_1801,N_1775);
and U2339 (N_2339,N_1605,N_1621);
and U2340 (N_2340,N_1567,N_1927);
and U2341 (N_2341,N_1729,N_1932);
and U2342 (N_2342,N_1709,N_1886);
and U2343 (N_2343,N_1590,N_1765);
and U2344 (N_2344,N_1711,N_1888);
or U2345 (N_2345,N_1721,N_1913);
or U2346 (N_2346,N_1855,N_1627);
and U2347 (N_2347,N_1944,N_1678);
or U2348 (N_2348,N_1838,N_1849);
nor U2349 (N_2349,N_1538,N_1820);
or U2350 (N_2350,N_1977,N_1569);
and U2351 (N_2351,N_1919,N_1867);
nor U2352 (N_2352,N_1554,N_1759);
nand U2353 (N_2353,N_1601,N_1933);
and U2354 (N_2354,N_1541,N_1984);
nor U2355 (N_2355,N_1703,N_1675);
nand U2356 (N_2356,N_1998,N_1602);
nor U2357 (N_2357,N_1874,N_1941);
and U2358 (N_2358,N_1899,N_1517);
nor U2359 (N_2359,N_1784,N_1580);
or U2360 (N_2360,N_1994,N_1690);
and U2361 (N_2361,N_1682,N_1887);
and U2362 (N_2362,N_1587,N_1583);
and U2363 (N_2363,N_1701,N_1848);
nand U2364 (N_2364,N_1882,N_1732);
nand U2365 (N_2365,N_1618,N_1955);
and U2366 (N_2366,N_1576,N_1864);
nor U2367 (N_2367,N_1822,N_1892);
and U2368 (N_2368,N_1856,N_1512);
nor U2369 (N_2369,N_1552,N_1913);
and U2370 (N_2370,N_1848,N_1949);
or U2371 (N_2371,N_1887,N_1944);
and U2372 (N_2372,N_1523,N_1655);
nor U2373 (N_2373,N_1987,N_1833);
xnor U2374 (N_2374,N_1517,N_1997);
xnor U2375 (N_2375,N_1824,N_1561);
nand U2376 (N_2376,N_1535,N_1707);
and U2377 (N_2377,N_1554,N_1917);
or U2378 (N_2378,N_1535,N_1874);
or U2379 (N_2379,N_1831,N_1769);
xor U2380 (N_2380,N_1631,N_1801);
xor U2381 (N_2381,N_1530,N_1674);
and U2382 (N_2382,N_1869,N_1689);
or U2383 (N_2383,N_1803,N_1903);
nor U2384 (N_2384,N_1676,N_1620);
nor U2385 (N_2385,N_1639,N_1988);
xnor U2386 (N_2386,N_1531,N_1783);
nand U2387 (N_2387,N_1599,N_1905);
or U2388 (N_2388,N_1626,N_1596);
or U2389 (N_2389,N_1839,N_1958);
nor U2390 (N_2390,N_1632,N_1500);
and U2391 (N_2391,N_1575,N_1708);
nand U2392 (N_2392,N_1766,N_1777);
and U2393 (N_2393,N_1920,N_1535);
xor U2394 (N_2394,N_1914,N_1930);
or U2395 (N_2395,N_1787,N_1883);
nor U2396 (N_2396,N_1912,N_1614);
nand U2397 (N_2397,N_1647,N_1765);
or U2398 (N_2398,N_1553,N_1967);
xor U2399 (N_2399,N_1697,N_1576);
nor U2400 (N_2400,N_1834,N_1658);
and U2401 (N_2401,N_1684,N_1888);
and U2402 (N_2402,N_1778,N_1820);
nand U2403 (N_2403,N_1688,N_1545);
and U2404 (N_2404,N_1846,N_1623);
or U2405 (N_2405,N_1847,N_1597);
or U2406 (N_2406,N_1982,N_1526);
and U2407 (N_2407,N_1606,N_1772);
nor U2408 (N_2408,N_1990,N_1644);
or U2409 (N_2409,N_1770,N_1829);
or U2410 (N_2410,N_1630,N_1912);
and U2411 (N_2411,N_1586,N_1851);
and U2412 (N_2412,N_1910,N_1928);
xor U2413 (N_2413,N_1748,N_1914);
nand U2414 (N_2414,N_1699,N_1831);
and U2415 (N_2415,N_1507,N_1653);
or U2416 (N_2416,N_1574,N_1612);
and U2417 (N_2417,N_1778,N_1991);
or U2418 (N_2418,N_1648,N_1975);
and U2419 (N_2419,N_1804,N_1960);
nor U2420 (N_2420,N_1760,N_1928);
or U2421 (N_2421,N_1973,N_1747);
and U2422 (N_2422,N_1504,N_1869);
nor U2423 (N_2423,N_1649,N_1737);
nand U2424 (N_2424,N_1913,N_1688);
nand U2425 (N_2425,N_1576,N_1995);
or U2426 (N_2426,N_1564,N_1772);
or U2427 (N_2427,N_1563,N_1841);
and U2428 (N_2428,N_1856,N_1765);
nor U2429 (N_2429,N_1810,N_1959);
and U2430 (N_2430,N_1905,N_1611);
and U2431 (N_2431,N_1689,N_1824);
and U2432 (N_2432,N_1717,N_1936);
and U2433 (N_2433,N_1649,N_1970);
nand U2434 (N_2434,N_1942,N_1803);
nand U2435 (N_2435,N_1987,N_1745);
nand U2436 (N_2436,N_1897,N_1564);
and U2437 (N_2437,N_1868,N_1599);
nand U2438 (N_2438,N_1875,N_1531);
nor U2439 (N_2439,N_1509,N_1735);
or U2440 (N_2440,N_1749,N_1750);
xor U2441 (N_2441,N_1771,N_1696);
and U2442 (N_2442,N_1698,N_1915);
or U2443 (N_2443,N_1893,N_1832);
xor U2444 (N_2444,N_1752,N_1737);
or U2445 (N_2445,N_1832,N_1668);
nand U2446 (N_2446,N_1884,N_1547);
nand U2447 (N_2447,N_1867,N_1909);
and U2448 (N_2448,N_1819,N_1547);
or U2449 (N_2449,N_1578,N_1628);
and U2450 (N_2450,N_1621,N_1977);
and U2451 (N_2451,N_1843,N_1756);
nand U2452 (N_2452,N_1642,N_1806);
nand U2453 (N_2453,N_1946,N_1573);
nor U2454 (N_2454,N_1739,N_1818);
and U2455 (N_2455,N_1667,N_1817);
and U2456 (N_2456,N_1860,N_1534);
and U2457 (N_2457,N_1782,N_1674);
nand U2458 (N_2458,N_1946,N_1880);
nand U2459 (N_2459,N_1964,N_1701);
or U2460 (N_2460,N_1518,N_1654);
nor U2461 (N_2461,N_1662,N_1545);
nor U2462 (N_2462,N_1719,N_1534);
nor U2463 (N_2463,N_1602,N_1966);
and U2464 (N_2464,N_1569,N_1970);
or U2465 (N_2465,N_1723,N_1812);
nor U2466 (N_2466,N_1693,N_1836);
and U2467 (N_2467,N_1618,N_1662);
nand U2468 (N_2468,N_1518,N_1626);
or U2469 (N_2469,N_1527,N_1983);
or U2470 (N_2470,N_1947,N_1553);
or U2471 (N_2471,N_1752,N_1993);
and U2472 (N_2472,N_1665,N_1842);
and U2473 (N_2473,N_1929,N_1962);
and U2474 (N_2474,N_1914,N_1650);
xor U2475 (N_2475,N_1858,N_1879);
and U2476 (N_2476,N_1795,N_1568);
or U2477 (N_2477,N_1929,N_1904);
nand U2478 (N_2478,N_1993,N_1963);
xnor U2479 (N_2479,N_1761,N_1606);
nor U2480 (N_2480,N_1718,N_1790);
nor U2481 (N_2481,N_1924,N_1783);
xnor U2482 (N_2482,N_1598,N_1767);
or U2483 (N_2483,N_1620,N_1755);
nand U2484 (N_2484,N_1902,N_1658);
nand U2485 (N_2485,N_1613,N_1721);
nor U2486 (N_2486,N_1901,N_1543);
or U2487 (N_2487,N_1685,N_1635);
and U2488 (N_2488,N_1514,N_1521);
or U2489 (N_2489,N_1828,N_1515);
and U2490 (N_2490,N_1566,N_1833);
nand U2491 (N_2491,N_1964,N_1867);
nand U2492 (N_2492,N_1972,N_1754);
or U2493 (N_2493,N_1837,N_1654);
nand U2494 (N_2494,N_1529,N_1628);
and U2495 (N_2495,N_1851,N_1510);
and U2496 (N_2496,N_1715,N_1954);
and U2497 (N_2497,N_1959,N_1700);
and U2498 (N_2498,N_1693,N_1920);
or U2499 (N_2499,N_1993,N_1565);
xor U2500 (N_2500,N_2000,N_2412);
and U2501 (N_2501,N_2005,N_2159);
or U2502 (N_2502,N_2182,N_2025);
and U2503 (N_2503,N_2057,N_2314);
and U2504 (N_2504,N_2041,N_2114);
and U2505 (N_2505,N_2020,N_2332);
xnor U2506 (N_2506,N_2304,N_2483);
or U2507 (N_2507,N_2298,N_2148);
and U2508 (N_2508,N_2046,N_2054);
or U2509 (N_2509,N_2018,N_2341);
and U2510 (N_2510,N_2176,N_2282);
and U2511 (N_2511,N_2416,N_2215);
and U2512 (N_2512,N_2402,N_2224);
xor U2513 (N_2513,N_2197,N_2070);
nor U2514 (N_2514,N_2239,N_2385);
and U2515 (N_2515,N_2093,N_2082);
or U2516 (N_2516,N_2134,N_2151);
nor U2517 (N_2517,N_2033,N_2276);
nor U2518 (N_2518,N_2245,N_2119);
nor U2519 (N_2519,N_2100,N_2060);
and U2520 (N_2520,N_2226,N_2342);
or U2521 (N_2521,N_2091,N_2129);
nor U2522 (N_2522,N_2450,N_2372);
or U2523 (N_2523,N_2301,N_2002);
nor U2524 (N_2524,N_2455,N_2438);
and U2525 (N_2525,N_2133,N_2166);
and U2526 (N_2526,N_2294,N_2260);
nand U2527 (N_2527,N_2475,N_2424);
and U2528 (N_2528,N_2448,N_2307);
and U2529 (N_2529,N_2272,N_2045);
nand U2530 (N_2530,N_2136,N_2181);
xnor U2531 (N_2531,N_2300,N_2189);
nor U2532 (N_2532,N_2135,N_2081);
nand U2533 (N_2533,N_2343,N_2496);
and U2534 (N_2534,N_2482,N_2132);
xor U2535 (N_2535,N_2037,N_2234);
xor U2536 (N_2536,N_2406,N_2117);
nand U2537 (N_2537,N_2269,N_2139);
nand U2538 (N_2538,N_2280,N_2191);
or U2539 (N_2539,N_2101,N_2375);
nor U2540 (N_2540,N_2327,N_2285);
and U2541 (N_2541,N_2195,N_2398);
nor U2542 (N_2542,N_2437,N_2079);
nand U2543 (N_2543,N_2319,N_2497);
nor U2544 (N_2544,N_2334,N_2076);
nor U2545 (N_2545,N_2083,N_2479);
nand U2546 (N_2546,N_2032,N_2262);
or U2547 (N_2547,N_2316,N_2255);
and U2548 (N_2548,N_2378,N_2487);
or U2549 (N_2549,N_2042,N_2030);
xor U2550 (N_2550,N_2321,N_2222);
nand U2551 (N_2551,N_2328,N_2290);
and U2552 (N_2552,N_2221,N_2146);
or U2553 (N_2553,N_2111,N_2348);
nor U2554 (N_2554,N_2305,N_2165);
xor U2555 (N_2555,N_2205,N_2423);
nor U2556 (N_2556,N_2072,N_2038);
nor U2557 (N_2557,N_2333,N_2175);
xor U2558 (N_2558,N_2329,N_2335);
nor U2559 (N_2559,N_2434,N_2388);
or U2560 (N_2560,N_2264,N_2295);
nor U2561 (N_2561,N_2212,N_2024);
nor U2562 (N_2562,N_2408,N_2391);
nor U2563 (N_2563,N_2379,N_2026);
nor U2564 (N_2564,N_2273,N_2248);
nand U2565 (N_2565,N_2346,N_2097);
nor U2566 (N_2566,N_2049,N_2315);
nand U2567 (N_2567,N_2481,N_2095);
and U2568 (N_2568,N_2432,N_2188);
or U2569 (N_2569,N_2251,N_2204);
and U2570 (N_2570,N_2124,N_2358);
nor U2571 (N_2571,N_2330,N_2246);
nand U2572 (N_2572,N_2089,N_2207);
nor U2573 (N_2573,N_2397,N_2064);
nor U2574 (N_2574,N_2061,N_2278);
xor U2575 (N_2575,N_2445,N_2323);
nand U2576 (N_2576,N_2302,N_2013);
nand U2577 (N_2577,N_2162,N_2011);
and U2578 (N_2578,N_2190,N_2494);
nor U2579 (N_2579,N_2185,N_2271);
or U2580 (N_2580,N_2365,N_2471);
and U2581 (N_2581,N_2073,N_2056);
and U2582 (N_2582,N_2150,N_2228);
xor U2583 (N_2583,N_2259,N_2227);
nor U2584 (N_2584,N_2160,N_2126);
and U2585 (N_2585,N_2058,N_2044);
or U2586 (N_2586,N_2270,N_2377);
nand U2587 (N_2587,N_2443,N_2383);
xor U2588 (N_2588,N_2431,N_2485);
or U2589 (N_2589,N_2409,N_2169);
xor U2590 (N_2590,N_2429,N_2313);
nor U2591 (N_2591,N_2229,N_2367);
or U2592 (N_2592,N_2401,N_2156);
nand U2593 (N_2593,N_2480,N_2094);
or U2594 (N_2594,N_2456,N_2015);
and U2595 (N_2595,N_2363,N_2137);
nand U2596 (N_2596,N_2452,N_2027);
nand U2597 (N_2597,N_2065,N_2220);
nor U2598 (N_2598,N_2312,N_2345);
nand U2599 (N_2599,N_2462,N_2153);
and U2600 (N_2600,N_2236,N_2410);
or U2601 (N_2601,N_2145,N_2127);
or U2602 (N_2602,N_2467,N_2394);
nand U2603 (N_2603,N_2143,N_2357);
or U2604 (N_2604,N_2318,N_2187);
or U2605 (N_2605,N_2068,N_2104);
or U2606 (N_2606,N_2130,N_2173);
nand U2607 (N_2607,N_2303,N_2172);
xnor U2608 (N_2608,N_2336,N_2012);
nand U2609 (N_2609,N_2405,N_2115);
xnor U2610 (N_2610,N_2426,N_2006);
nor U2611 (N_2611,N_2324,N_2347);
nor U2612 (N_2612,N_2419,N_2288);
nor U2613 (N_2613,N_2418,N_2493);
nand U2614 (N_2614,N_2427,N_2351);
and U2615 (N_2615,N_2466,N_2233);
xnor U2616 (N_2616,N_2309,N_2370);
nand U2617 (N_2617,N_2266,N_2225);
nand U2618 (N_2618,N_2053,N_2337);
or U2619 (N_2619,N_2362,N_2086);
and U2620 (N_2620,N_2194,N_2003);
and U2621 (N_2621,N_2157,N_2177);
nor U2622 (N_2622,N_2352,N_2014);
nand U2623 (N_2623,N_2240,N_2308);
nor U2624 (N_2624,N_2199,N_2474);
nor U2625 (N_2625,N_2414,N_2052);
nand U2626 (N_2626,N_2433,N_2339);
and U2627 (N_2627,N_2110,N_2031);
nor U2628 (N_2628,N_2368,N_2219);
nor U2629 (N_2629,N_2010,N_2320);
nand U2630 (N_2630,N_2249,N_2059);
nor U2631 (N_2631,N_2254,N_2184);
and U2632 (N_2632,N_2296,N_2161);
or U2633 (N_2633,N_2265,N_2499);
nand U2634 (N_2634,N_2369,N_2193);
nand U2635 (N_2635,N_2277,N_2460);
or U2636 (N_2636,N_2232,N_2491);
or U2637 (N_2637,N_2353,N_2380);
and U2638 (N_2638,N_2472,N_2490);
nor U2639 (N_2639,N_2090,N_2322);
nor U2640 (N_2640,N_2170,N_2441);
and U2641 (N_2641,N_2361,N_2218);
nand U2642 (N_2642,N_2284,N_2373);
and U2643 (N_2643,N_2164,N_2449);
nor U2644 (N_2644,N_2261,N_2461);
and U2645 (N_2645,N_2454,N_2286);
and U2646 (N_2646,N_2442,N_2067);
nand U2647 (N_2647,N_2469,N_2268);
and U2648 (N_2648,N_2075,N_2393);
nand U2649 (N_2649,N_2144,N_2274);
nand U2650 (N_2650,N_2007,N_2167);
nor U2651 (N_2651,N_2048,N_2242);
and U2652 (N_2652,N_2349,N_2087);
xor U2653 (N_2653,N_2413,N_2022);
or U2654 (N_2654,N_2140,N_2108);
or U2655 (N_2655,N_2258,N_2213);
nor U2656 (N_2656,N_2201,N_2325);
and U2657 (N_2657,N_2297,N_2211);
nand U2658 (N_2658,N_2063,N_2237);
nand U2659 (N_2659,N_2092,N_2340);
xor U2660 (N_2660,N_2241,N_2123);
nand U2661 (N_2661,N_2390,N_2436);
nor U2662 (N_2662,N_2206,N_2484);
and U2663 (N_2663,N_2055,N_2492);
and U2664 (N_2664,N_2384,N_2399);
nor U2665 (N_2665,N_2495,N_2250);
or U2666 (N_2666,N_2389,N_2102);
or U2667 (N_2667,N_2338,N_2120);
nand U2668 (N_2668,N_2196,N_2203);
and U2669 (N_2669,N_2216,N_2252);
xnor U2670 (N_2670,N_2138,N_2407);
nor U2671 (N_2671,N_2096,N_2451);
nor U2672 (N_2672,N_2458,N_2085);
and U2673 (N_2673,N_2478,N_2214);
nand U2674 (N_2674,N_2421,N_2306);
and U2675 (N_2675,N_2198,N_2404);
or U2676 (N_2676,N_2453,N_2381);
nor U2677 (N_2677,N_2403,N_2208);
nand U2678 (N_2678,N_2289,N_2200);
nor U2679 (N_2679,N_2444,N_2174);
nand U2680 (N_2680,N_2062,N_2465);
xor U2681 (N_2681,N_2105,N_2019);
nand U2682 (N_2682,N_2040,N_2178);
and U2683 (N_2683,N_2077,N_2287);
or U2684 (N_2684,N_2217,N_2470);
and U2685 (N_2685,N_2107,N_2446);
nor U2686 (N_2686,N_2179,N_2422);
xor U2687 (N_2687,N_2125,N_2168);
or U2688 (N_2688,N_2017,N_2310);
xor U2689 (N_2689,N_2035,N_2428);
nor U2690 (N_2690,N_2354,N_2311);
and U2691 (N_2691,N_2078,N_2163);
nor U2692 (N_2692,N_2036,N_2489);
or U2693 (N_2693,N_2039,N_2344);
nor U2694 (N_2694,N_2435,N_2326);
xnor U2695 (N_2695,N_2350,N_2074);
or U2696 (N_2696,N_2155,N_2149);
nand U2697 (N_2697,N_2231,N_2147);
nor U2698 (N_2698,N_2299,N_2080);
or U2699 (N_2699,N_2417,N_2034);
nand U2700 (N_2700,N_2008,N_2281);
nor U2701 (N_2701,N_2392,N_2235);
nor U2702 (N_2702,N_2243,N_2047);
nand U2703 (N_2703,N_2459,N_2230);
nand U2704 (N_2704,N_2050,N_2128);
nand U2705 (N_2705,N_2158,N_2376);
and U2706 (N_2706,N_2263,N_2425);
xor U2707 (N_2707,N_2066,N_2430);
nor U2708 (N_2708,N_2486,N_2386);
and U2709 (N_2709,N_2247,N_2366);
or U2710 (N_2710,N_2291,N_2400);
and U2711 (N_2711,N_2118,N_2238);
nand U2712 (N_2712,N_2071,N_2463);
and U2713 (N_2713,N_2279,N_2088);
and U2714 (N_2714,N_2477,N_2192);
or U2715 (N_2715,N_2457,N_2021);
xnor U2716 (N_2716,N_2382,N_2253);
nor U2717 (N_2717,N_2488,N_2069);
or U2718 (N_2718,N_2099,N_2275);
or U2719 (N_2719,N_2396,N_2331);
and U2720 (N_2720,N_2223,N_2356);
nand U2721 (N_2721,N_2473,N_2364);
nand U2722 (N_2722,N_2009,N_2317);
and U2723 (N_2723,N_2043,N_2028);
xnor U2724 (N_2724,N_2103,N_2256);
nor U2725 (N_2725,N_2004,N_2476);
nor U2726 (N_2726,N_2371,N_2374);
or U2727 (N_2727,N_2210,N_2186);
nor U2728 (N_2728,N_2106,N_2447);
nand U2729 (N_2729,N_2109,N_2098);
and U2730 (N_2730,N_2051,N_2420);
nor U2731 (N_2731,N_2141,N_2283);
nor U2732 (N_2732,N_2116,N_2411);
nand U2733 (N_2733,N_2293,N_2112);
or U2734 (N_2734,N_2180,N_2142);
nand U2735 (N_2735,N_2440,N_2121);
or U2736 (N_2736,N_2171,N_2498);
or U2737 (N_2737,N_2244,N_2359);
nor U2738 (N_2738,N_2292,N_2029);
nand U2739 (N_2739,N_2202,N_2084);
nor U2740 (N_2740,N_2468,N_2267);
and U2741 (N_2741,N_2152,N_2209);
nand U2742 (N_2742,N_2016,N_2113);
and U2743 (N_2743,N_2395,N_2415);
or U2744 (N_2744,N_2355,N_2131);
nand U2745 (N_2745,N_2387,N_2464);
nand U2746 (N_2746,N_2360,N_2023);
nor U2747 (N_2747,N_2183,N_2257);
or U2748 (N_2748,N_2001,N_2439);
or U2749 (N_2749,N_2122,N_2154);
nand U2750 (N_2750,N_2258,N_2019);
nor U2751 (N_2751,N_2424,N_2462);
xnor U2752 (N_2752,N_2400,N_2218);
nand U2753 (N_2753,N_2043,N_2100);
or U2754 (N_2754,N_2092,N_2430);
or U2755 (N_2755,N_2492,N_2034);
and U2756 (N_2756,N_2210,N_2198);
or U2757 (N_2757,N_2247,N_2425);
xnor U2758 (N_2758,N_2118,N_2185);
or U2759 (N_2759,N_2492,N_2013);
nor U2760 (N_2760,N_2320,N_2432);
and U2761 (N_2761,N_2295,N_2115);
or U2762 (N_2762,N_2072,N_2394);
xnor U2763 (N_2763,N_2341,N_2181);
nand U2764 (N_2764,N_2190,N_2248);
and U2765 (N_2765,N_2100,N_2106);
or U2766 (N_2766,N_2295,N_2410);
xnor U2767 (N_2767,N_2086,N_2224);
or U2768 (N_2768,N_2011,N_2045);
xor U2769 (N_2769,N_2097,N_2431);
and U2770 (N_2770,N_2241,N_2220);
or U2771 (N_2771,N_2319,N_2087);
nor U2772 (N_2772,N_2180,N_2466);
or U2773 (N_2773,N_2426,N_2162);
and U2774 (N_2774,N_2122,N_2279);
nand U2775 (N_2775,N_2047,N_2175);
xor U2776 (N_2776,N_2277,N_2400);
and U2777 (N_2777,N_2110,N_2177);
and U2778 (N_2778,N_2497,N_2143);
and U2779 (N_2779,N_2151,N_2257);
xor U2780 (N_2780,N_2435,N_2123);
and U2781 (N_2781,N_2118,N_2152);
nor U2782 (N_2782,N_2459,N_2417);
nor U2783 (N_2783,N_2482,N_2222);
and U2784 (N_2784,N_2309,N_2105);
nand U2785 (N_2785,N_2050,N_2167);
nand U2786 (N_2786,N_2475,N_2131);
and U2787 (N_2787,N_2251,N_2401);
nor U2788 (N_2788,N_2211,N_2196);
or U2789 (N_2789,N_2065,N_2192);
nor U2790 (N_2790,N_2040,N_2172);
nor U2791 (N_2791,N_2241,N_2371);
and U2792 (N_2792,N_2276,N_2206);
nor U2793 (N_2793,N_2253,N_2347);
nand U2794 (N_2794,N_2219,N_2210);
or U2795 (N_2795,N_2159,N_2244);
xnor U2796 (N_2796,N_2196,N_2071);
nand U2797 (N_2797,N_2415,N_2457);
nor U2798 (N_2798,N_2497,N_2092);
nand U2799 (N_2799,N_2314,N_2262);
xnor U2800 (N_2800,N_2278,N_2190);
or U2801 (N_2801,N_2370,N_2195);
or U2802 (N_2802,N_2255,N_2207);
nor U2803 (N_2803,N_2481,N_2034);
and U2804 (N_2804,N_2011,N_2003);
or U2805 (N_2805,N_2366,N_2484);
or U2806 (N_2806,N_2051,N_2199);
nor U2807 (N_2807,N_2151,N_2287);
nand U2808 (N_2808,N_2096,N_2238);
xor U2809 (N_2809,N_2160,N_2469);
nand U2810 (N_2810,N_2244,N_2343);
or U2811 (N_2811,N_2369,N_2260);
xor U2812 (N_2812,N_2105,N_2301);
and U2813 (N_2813,N_2352,N_2284);
or U2814 (N_2814,N_2187,N_2358);
or U2815 (N_2815,N_2069,N_2269);
and U2816 (N_2816,N_2039,N_2175);
nand U2817 (N_2817,N_2482,N_2029);
and U2818 (N_2818,N_2123,N_2484);
and U2819 (N_2819,N_2124,N_2388);
xor U2820 (N_2820,N_2181,N_2369);
and U2821 (N_2821,N_2166,N_2211);
and U2822 (N_2822,N_2273,N_2127);
and U2823 (N_2823,N_2408,N_2047);
or U2824 (N_2824,N_2341,N_2409);
nor U2825 (N_2825,N_2029,N_2215);
nand U2826 (N_2826,N_2022,N_2237);
nand U2827 (N_2827,N_2405,N_2181);
nor U2828 (N_2828,N_2099,N_2339);
or U2829 (N_2829,N_2481,N_2156);
and U2830 (N_2830,N_2431,N_2216);
nand U2831 (N_2831,N_2190,N_2249);
nor U2832 (N_2832,N_2388,N_2130);
and U2833 (N_2833,N_2424,N_2327);
and U2834 (N_2834,N_2460,N_2054);
nand U2835 (N_2835,N_2044,N_2411);
nor U2836 (N_2836,N_2491,N_2414);
and U2837 (N_2837,N_2295,N_2322);
xor U2838 (N_2838,N_2278,N_2405);
or U2839 (N_2839,N_2401,N_2112);
nor U2840 (N_2840,N_2488,N_2085);
and U2841 (N_2841,N_2432,N_2441);
or U2842 (N_2842,N_2242,N_2433);
nor U2843 (N_2843,N_2049,N_2491);
xnor U2844 (N_2844,N_2476,N_2332);
or U2845 (N_2845,N_2454,N_2089);
nor U2846 (N_2846,N_2172,N_2226);
nor U2847 (N_2847,N_2135,N_2311);
xor U2848 (N_2848,N_2149,N_2415);
and U2849 (N_2849,N_2052,N_2476);
nor U2850 (N_2850,N_2112,N_2241);
and U2851 (N_2851,N_2489,N_2038);
and U2852 (N_2852,N_2492,N_2198);
nand U2853 (N_2853,N_2057,N_2085);
and U2854 (N_2854,N_2353,N_2408);
and U2855 (N_2855,N_2463,N_2274);
xnor U2856 (N_2856,N_2293,N_2226);
nand U2857 (N_2857,N_2325,N_2285);
nand U2858 (N_2858,N_2174,N_2406);
and U2859 (N_2859,N_2027,N_2147);
xnor U2860 (N_2860,N_2006,N_2170);
nand U2861 (N_2861,N_2369,N_2443);
or U2862 (N_2862,N_2498,N_2045);
or U2863 (N_2863,N_2297,N_2038);
or U2864 (N_2864,N_2448,N_2405);
and U2865 (N_2865,N_2393,N_2284);
and U2866 (N_2866,N_2416,N_2394);
nor U2867 (N_2867,N_2191,N_2486);
nand U2868 (N_2868,N_2444,N_2484);
nand U2869 (N_2869,N_2043,N_2413);
nand U2870 (N_2870,N_2260,N_2202);
nand U2871 (N_2871,N_2204,N_2440);
nand U2872 (N_2872,N_2308,N_2127);
or U2873 (N_2873,N_2084,N_2075);
or U2874 (N_2874,N_2372,N_2083);
nor U2875 (N_2875,N_2261,N_2116);
nand U2876 (N_2876,N_2027,N_2433);
nor U2877 (N_2877,N_2160,N_2009);
nor U2878 (N_2878,N_2216,N_2155);
or U2879 (N_2879,N_2370,N_2412);
or U2880 (N_2880,N_2448,N_2301);
and U2881 (N_2881,N_2091,N_2006);
or U2882 (N_2882,N_2293,N_2289);
and U2883 (N_2883,N_2118,N_2102);
or U2884 (N_2884,N_2490,N_2294);
nand U2885 (N_2885,N_2181,N_2305);
or U2886 (N_2886,N_2408,N_2287);
nor U2887 (N_2887,N_2301,N_2049);
or U2888 (N_2888,N_2450,N_2020);
and U2889 (N_2889,N_2078,N_2139);
and U2890 (N_2890,N_2127,N_2078);
and U2891 (N_2891,N_2249,N_2332);
or U2892 (N_2892,N_2483,N_2154);
nor U2893 (N_2893,N_2197,N_2181);
or U2894 (N_2894,N_2202,N_2362);
and U2895 (N_2895,N_2343,N_2024);
nor U2896 (N_2896,N_2119,N_2094);
nor U2897 (N_2897,N_2482,N_2499);
or U2898 (N_2898,N_2020,N_2102);
nor U2899 (N_2899,N_2023,N_2481);
or U2900 (N_2900,N_2242,N_2489);
nand U2901 (N_2901,N_2168,N_2476);
nand U2902 (N_2902,N_2295,N_2157);
and U2903 (N_2903,N_2216,N_2171);
nor U2904 (N_2904,N_2255,N_2231);
and U2905 (N_2905,N_2109,N_2202);
nor U2906 (N_2906,N_2392,N_2010);
nor U2907 (N_2907,N_2051,N_2189);
nand U2908 (N_2908,N_2280,N_2201);
or U2909 (N_2909,N_2253,N_2008);
and U2910 (N_2910,N_2069,N_2262);
and U2911 (N_2911,N_2093,N_2346);
nand U2912 (N_2912,N_2375,N_2285);
or U2913 (N_2913,N_2271,N_2230);
or U2914 (N_2914,N_2222,N_2121);
or U2915 (N_2915,N_2361,N_2267);
nand U2916 (N_2916,N_2472,N_2487);
xor U2917 (N_2917,N_2180,N_2288);
nor U2918 (N_2918,N_2169,N_2178);
or U2919 (N_2919,N_2294,N_2407);
or U2920 (N_2920,N_2123,N_2233);
nor U2921 (N_2921,N_2019,N_2234);
nand U2922 (N_2922,N_2009,N_2294);
nor U2923 (N_2923,N_2107,N_2289);
or U2924 (N_2924,N_2475,N_2353);
and U2925 (N_2925,N_2169,N_2134);
and U2926 (N_2926,N_2422,N_2128);
nand U2927 (N_2927,N_2498,N_2255);
and U2928 (N_2928,N_2248,N_2403);
nand U2929 (N_2929,N_2200,N_2420);
nand U2930 (N_2930,N_2039,N_2107);
xor U2931 (N_2931,N_2499,N_2401);
nand U2932 (N_2932,N_2219,N_2153);
or U2933 (N_2933,N_2220,N_2377);
nor U2934 (N_2934,N_2011,N_2316);
and U2935 (N_2935,N_2305,N_2469);
and U2936 (N_2936,N_2378,N_2209);
nand U2937 (N_2937,N_2035,N_2234);
nor U2938 (N_2938,N_2262,N_2338);
or U2939 (N_2939,N_2002,N_2274);
nor U2940 (N_2940,N_2428,N_2407);
nor U2941 (N_2941,N_2296,N_2280);
or U2942 (N_2942,N_2362,N_2124);
and U2943 (N_2943,N_2193,N_2174);
nand U2944 (N_2944,N_2452,N_2073);
and U2945 (N_2945,N_2373,N_2291);
nand U2946 (N_2946,N_2368,N_2395);
and U2947 (N_2947,N_2237,N_2438);
xor U2948 (N_2948,N_2391,N_2223);
nand U2949 (N_2949,N_2023,N_2202);
and U2950 (N_2950,N_2495,N_2353);
or U2951 (N_2951,N_2033,N_2334);
or U2952 (N_2952,N_2482,N_2255);
or U2953 (N_2953,N_2071,N_2261);
and U2954 (N_2954,N_2186,N_2333);
or U2955 (N_2955,N_2145,N_2232);
xnor U2956 (N_2956,N_2169,N_2474);
or U2957 (N_2957,N_2244,N_2076);
or U2958 (N_2958,N_2117,N_2187);
nand U2959 (N_2959,N_2117,N_2414);
and U2960 (N_2960,N_2160,N_2398);
nand U2961 (N_2961,N_2488,N_2336);
nand U2962 (N_2962,N_2202,N_2096);
nand U2963 (N_2963,N_2482,N_2124);
nand U2964 (N_2964,N_2189,N_2052);
or U2965 (N_2965,N_2148,N_2158);
and U2966 (N_2966,N_2439,N_2020);
nand U2967 (N_2967,N_2200,N_2394);
nor U2968 (N_2968,N_2461,N_2471);
or U2969 (N_2969,N_2381,N_2292);
and U2970 (N_2970,N_2184,N_2249);
or U2971 (N_2971,N_2419,N_2444);
or U2972 (N_2972,N_2176,N_2223);
xor U2973 (N_2973,N_2326,N_2277);
and U2974 (N_2974,N_2037,N_2163);
nor U2975 (N_2975,N_2397,N_2471);
nor U2976 (N_2976,N_2143,N_2370);
and U2977 (N_2977,N_2019,N_2153);
and U2978 (N_2978,N_2359,N_2066);
xnor U2979 (N_2979,N_2495,N_2262);
or U2980 (N_2980,N_2428,N_2021);
and U2981 (N_2981,N_2188,N_2414);
or U2982 (N_2982,N_2130,N_2180);
nor U2983 (N_2983,N_2141,N_2267);
nand U2984 (N_2984,N_2431,N_2198);
nand U2985 (N_2985,N_2432,N_2269);
or U2986 (N_2986,N_2230,N_2297);
or U2987 (N_2987,N_2206,N_2378);
nand U2988 (N_2988,N_2074,N_2348);
or U2989 (N_2989,N_2090,N_2458);
nand U2990 (N_2990,N_2381,N_2089);
nor U2991 (N_2991,N_2461,N_2347);
xnor U2992 (N_2992,N_2086,N_2201);
nand U2993 (N_2993,N_2043,N_2453);
nor U2994 (N_2994,N_2293,N_2217);
nor U2995 (N_2995,N_2000,N_2099);
and U2996 (N_2996,N_2049,N_2119);
nand U2997 (N_2997,N_2409,N_2056);
or U2998 (N_2998,N_2399,N_2354);
or U2999 (N_2999,N_2446,N_2356);
and U3000 (N_3000,N_2764,N_2859);
or U3001 (N_3001,N_2666,N_2996);
nand U3002 (N_3002,N_2789,N_2541);
nor U3003 (N_3003,N_2627,N_2951);
and U3004 (N_3004,N_2604,N_2932);
or U3005 (N_3005,N_2842,N_2655);
or U3006 (N_3006,N_2620,N_2853);
nand U3007 (N_3007,N_2813,N_2690);
xor U3008 (N_3008,N_2714,N_2664);
and U3009 (N_3009,N_2800,N_2829);
and U3010 (N_3010,N_2687,N_2740);
nor U3011 (N_3011,N_2774,N_2886);
xor U3012 (N_3012,N_2706,N_2625);
and U3013 (N_3013,N_2905,N_2963);
and U3014 (N_3014,N_2956,N_2894);
nand U3015 (N_3015,N_2978,N_2937);
nand U3016 (N_3016,N_2761,N_2626);
nor U3017 (N_3017,N_2839,N_2724);
and U3018 (N_3018,N_2518,N_2936);
and U3019 (N_3019,N_2890,N_2713);
nor U3020 (N_3020,N_2535,N_2867);
and U3021 (N_3021,N_2781,N_2691);
and U3022 (N_3022,N_2969,N_2955);
and U3023 (N_3023,N_2903,N_2716);
nand U3024 (N_3024,N_2505,N_2682);
or U3025 (N_3025,N_2985,N_2995);
and U3026 (N_3026,N_2756,N_2762);
and U3027 (N_3027,N_2838,N_2614);
and U3028 (N_3028,N_2863,N_2929);
nor U3029 (N_3029,N_2844,N_2934);
and U3030 (N_3030,N_2887,N_2515);
or U3031 (N_3031,N_2900,N_2583);
and U3032 (N_3032,N_2982,N_2775);
and U3033 (N_3033,N_2733,N_2790);
or U3034 (N_3034,N_2984,N_2763);
and U3035 (N_3035,N_2631,N_2603);
nor U3036 (N_3036,N_2953,N_2814);
and U3037 (N_3037,N_2538,N_2731);
xor U3038 (N_3038,N_2876,N_2952);
and U3039 (N_3039,N_2926,N_2547);
and U3040 (N_3040,N_2571,N_2941);
or U3041 (N_3041,N_2546,N_2924);
nand U3042 (N_3042,N_2992,N_2909);
nand U3043 (N_3043,N_2578,N_2928);
nor U3044 (N_3044,N_2531,N_2870);
or U3045 (N_3045,N_2826,N_2661);
and U3046 (N_3046,N_2702,N_2968);
and U3047 (N_3047,N_2824,N_2750);
nand U3048 (N_3048,N_2739,N_2720);
nand U3049 (N_3049,N_2574,N_2657);
or U3050 (N_3050,N_2637,N_2757);
nor U3051 (N_3051,N_2721,N_2732);
or U3052 (N_3052,N_2563,N_2516);
xor U3053 (N_3053,N_2660,N_2769);
and U3054 (N_3054,N_2689,N_2704);
nor U3055 (N_3055,N_2792,N_2597);
xor U3056 (N_3056,N_2827,N_2787);
nor U3057 (N_3057,N_2967,N_2680);
xor U3058 (N_3058,N_2526,N_2849);
nor U3059 (N_3059,N_2519,N_2570);
or U3060 (N_3060,N_2972,N_2530);
nor U3061 (N_3061,N_2523,N_2635);
nor U3062 (N_3062,N_2933,N_2577);
and U3063 (N_3063,N_2809,N_2788);
xor U3064 (N_3064,N_2923,N_2866);
and U3065 (N_3065,N_2913,N_2674);
nor U3066 (N_3066,N_2819,N_2513);
and U3067 (N_3067,N_2554,N_2884);
or U3068 (N_3068,N_2940,N_2893);
nand U3069 (N_3069,N_2556,N_2807);
nor U3070 (N_3070,N_2676,N_2634);
and U3071 (N_3071,N_2795,N_2847);
nand U3072 (N_3072,N_2633,N_2507);
xor U3073 (N_3073,N_2889,N_2537);
and U3074 (N_3074,N_2935,N_2745);
nand U3075 (N_3075,N_2586,N_2865);
and U3076 (N_3076,N_2548,N_2916);
nor U3077 (N_3077,N_2860,N_2931);
and U3078 (N_3078,N_2970,N_2669);
nand U3079 (N_3079,N_2754,N_2699);
and U3080 (N_3080,N_2854,N_2649);
nor U3081 (N_3081,N_2881,N_2709);
or U3082 (N_3082,N_2718,N_2652);
nor U3083 (N_3083,N_2551,N_2725);
or U3084 (N_3084,N_2601,N_2918);
and U3085 (N_3085,N_2653,N_2852);
and U3086 (N_3086,N_2991,N_2812);
nand U3087 (N_3087,N_2642,N_2540);
nand U3088 (N_3088,N_2743,N_2607);
xnor U3089 (N_3089,N_2901,N_2677);
nand U3090 (N_3090,N_2834,N_2836);
or U3091 (N_3091,N_2623,N_2736);
or U3092 (N_3092,N_2988,N_2786);
nor U3093 (N_3093,N_2710,N_2802);
and U3094 (N_3094,N_2545,N_2938);
nor U3095 (N_3095,N_2784,N_2755);
nand U3096 (N_3096,N_2590,N_2701);
nand U3097 (N_3097,N_2528,N_2939);
nor U3098 (N_3098,N_2843,N_2947);
nand U3099 (N_3099,N_2667,N_2751);
or U3100 (N_3100,N_2793,N_2919);
and U3101 (N_3101,N_2668,N_2692);
and U3102 (N_3102,N_2695,N_2562);
nor U3103 (N_3103,N_2688,N_2595);
nor U3104 (N_3104,N_2617,N_2640);
nand U3105 (N_3105,N_2521,N_2553);
nor U3106 (N_3106,N_2773,N_2568);
nand U3107 (N_3107,N_2632,N_2708);
or U3108 (N_3108,N_2871,N_2981);
and U3109 (N_3109,N_2550,N_2662);
or U3110 (N_3110,N_2850,N_2845);
and U3111 (N_3111,N_2921,N_2976);
and U3112 (N_3112,N_2711,N_2946);
nand U3113 (N_3113,N_2639,N_2767);
nand U3114 (N_3114,N_2971,N_2615);
and U3115 (N_3115,N_2703,N_2780);
xor U3116 (N_3116,N_2651,N_2804);
nand U3117 (N_3117,N_2821,N_2559);
nor U3118 (N_3118,N_2799,N_2593);
xor U3119 (N_3119,N_2980,N_2927);
or U3120 (N_3120,N_2833,N_2758);
and U3121 (N_3121,N_2672,N_2656);
and U3122 (N_3122,N_2644,N_2645);
or U3123 (N_3123,N_2581,N_2908);
nor U3124 (N_3124,N_2678,N_2864);
nand U3125 (N_3125,N_2748,N_2734);
and U3126 (N_3126,N_2694,N_2797);
and U3127 (N_3127,N_2501,N_2742);
or U3128 (N_3128,N_2879,N_2875);
and U3129 (N_3129,N_2712,N_2608);
or U3130 (N_3130,N_2914,N_2509);
nor U3131 (N_3131,N_2828,N_2636);
and U3132 (N_3132,N_2555,N_2591);
or U3133 (N_3133,N_2848,N_2539);
nor U3134 (N_3134,N_2857,N_2993);
nand U3135 (N_3135,N_2630,N_2594);
or U3136 (N_3136,N_2511,N_2587);
or U3137 (N_3137,N_2723,N_2785);
nor U3138 (N_3138,N_2726,N_2650);
or U3139 (N_3139,N_2965,N_2948);
nand U3140 (N_3140,N_2565,N_2765);
and U3141 (N_3141,N_2575,N_2917);
and U3142 (N_3142,N_2749,N_2517);
xor U3143 (N_3143,N_2883,N_2840);
nor U3144 (N_3144,N_2612,N_2794);
or U3145 (N_3145,N_2782,N_2572);
nor U3146 (N_3146,N_2524,N_2616);
nand U3147 (N_3147,N_2512,N_2869);
or U3148 (N_3148,N_2874,N_2600);
and U3149 (N_3149,N_2618,N_2670);
or U3150 (N_3150,N_2979,N_2675);
and U3151 (N_3151,N_2500,N_2862);
xor U3152 (N_3152,N_2659,N_2610);
or U3153 (N_3153,N_2798,N_2567);
or U3154 (N_3154,N_2728,N_2783);
nor U3155 (N_3155,N_2558,N_2841);
nand U3156 (N_3156,N_2719,N_2779);
or U3157 (N_3157,N_2529,N_2647);
and U3158 (N_3158,N_2638,N_2902);
nor U3159 (N_3159,N_2504,N_2861);
xor U3160 (N_3160,N_2646,N_2506);
xor U3161 (N_3161,N_2958,N_2997);
nand U3162 (N_3162,N_2741,N_2592);
or U3163 (N_3163,N_2705,N_2609);
nand U3164 (N_3164,N_2974,N_2846);
nor U3165 (N_3165,N_2912,N_2697);
and U3166 (N_3166,N_2685,N_2760);
xnor U3167 (N_3167,N_2598,N_2684);
nand U3168 (N_3168,N_2573,N_2817);
and U3169 (N_3169,N_2681,N_2915);
or U3170 (N_3170,N_2977,N_2960);
nand U3171 (N_3171,N_2975,N_2907);
nand U3172 (N_3172,N_2791,N_2801);
nand U3173 (N_3173,N_2772,N_2520);
nand U3174 (N_3174,N_2959,N_2527);
nand U3175 (N_3175,N_2599,N_2855);
nor U3176 (N_3176,N_2543,N_2858);
nand U3177 (N_3177,N_2549,N_2832);
nand U3178 (N_3178,N_2904,N_2696);
nor U3179 (N_3179,N_2942,N_2525);
xnor U3180 (N_3180,N_2544,N_2722);
or U3181 (N_3181,N_2897,N_2679);
nand U3182 (N_3182,N_2698,N_2746);
nor U3183 (N_3183,N_2619,N_2822);
or U3184 (N_3184,N_2514,N_2579);
nor U3185 (N_3185,N_2925,N_2628);
or U3186 (N_3186,N_2777,N_2534);
or U3187 (N_3187,N_2588,N_2665);
or U3188 (N_3188,N_2753,N_2747);
nor U3189 (N_3189,N_2683,N_2727);
nor U3190 (N_3190,N_2737,N_2584);
nand U3191 (N_3191,N_2999,N_2943);
or U3192 (N_3192,N_2818,N_2877);
nor U3193 (N_3193,N_2816,N_2560);
xor U3194 (N_3194,N_2820,N_2983);
and U3195 (N_3195,N_2503,N_2738);
nor U3196 (N_3196,N_2880,N_2717);
and U3197 (N_3197,N_2654,N_2533);
or U3198 (N_3198,N_2966,N_2811);
and U3199 (N_3199,N_2766,N_2557);
nor U3200 (N_3200,N_2837,N_2911);
nand U3201 (N_3201,N_2989,N_2805);
nand U3202 (N_3202,N_2987,N_2532);
or U3203 (N_3203,N_2868,N_2998);
or U3204 (N_3204,N_2658,N_2508);
or U3205 (N_3205,N_2851,N_2806);
nand U3206 (N_3206,N_2873,N_2602);
or U3207 (N_3207,N_2808,N_2891);
nor U3208 (N_3208,N_2830,N_2752);
nor U3209 (N_3209,N_2643,N_2693);
or U3210 (N_3210,N_2606,N_2823);
or U3211 (N_3211,N_2906,N_2552);
nor U3212 (N_3212,N_2957,N_2648);
xor U3213 (N_3213,N_2831,N_2629);
and U3214 (N_3214,N_2536,N_2796);
nand U3215 (N_3215,N_2707,N_2856);
and U3216 (N_3216,N_2569,N_2810);
nand U3217 (N_3217,N_2589,N_2542);
nand U3218 (N_3218,N_2729,N_2895);
nand U3219 (N_3219,N_2744,N_2964);
nand U3220 (N_3220,N_2910,N_2611);
or U3221 (N_3221,N_2768,N_2778);
or U3222 (N_3222,N_2510,N_2585);
or U3223 (N_3223,N_2994,N_2624);
nor U3224 (N_3224,N_2613,N_2759);
xnor U3225 (N_3225,N_2673,N_2825);
or U3226 (N_3226,N_2582,N_2990);
xor U3227 (N_3227,N_2641,N_2899);
nor U3228 (N_3228,N_2835,N_2715);
nand U3229 (N_3229,N_2621,N_2885);
or U3230 (N_3230,N_2502,N_2663);
or U3231 (N_3231,N_2896,N_2962);
and U3232 (N_3232,N_2986,N_2878);
xor U3233 (N_3233,N_2671,N_2882);
and U3234 (N_3234,N_2566,N_2920);
or U3235 (N_3235,N_2522,N_2954);
and U3236 (N_3236,N_2949,N_2580);
and U3237 (N_3237,N_2770,N_2700);
or U3238 (N_3238,N_2950,N_2564);
nor U3239 (N_3239,N_2735,N_2803);
or U3240 (N_3240,N_2944,N_2945);
nand U3241 (N_3241,N_2771,N_2930);
and U3242 (N_3242,N_2922,N_2872);
nor U3243 (N_3243,N_2605,N_2961);
and U3244 (N_3244,N_2622,N_2730);
or U3245 (N_3245,N_2561,N_2576);
nor U3246 (N_3246,N_2776,N_2596);
nand U3247 (N_3247,N_2892,N_2686);
nor U3248 (N_3248,N_2973,N_2898);
nand U3249 (N_3249,N_2888,N_2815);
or U3250 (N_3250,N_2984,N_2902);
and U3251 (N_3251,N_2576,N_2662);
nor U3252 (N_3252,N_2722,N_2508);
nand U3253 (N_3253,N_2973,N_2702);
nand U3254 (N_3254,N_2885,N_2889);
xor U3255 (N_3255,N_2631,N_2574);
xor U3256 (N_3256,N_2795,N_2863);
nor U3257 (N_3257,N_2640,N_2535);
xor U3258 (N_3258,N_2793,N_2799);
or U3259 (N_3259,N_2545,N_2556);
nand U3260 (N_3260,N_2544,N_2933);
nor U3261 (N_3261,N_2926,N_2806);
or U3262 (N_3262,N_2982,N_2587);
or U3263 (N_3263,N_2540,N_2668);
nor U3264 (N_3264,N_2873,N_2836);
and U3265 (N_3265,N_2813,N_2788);
xor U3266 (N_3266,N_2838,N_2875);
nand U3267 (N_3267,N_2993,N_2862);
nor U3268 (N_3268,N_2514,N_2500);
or U3269 (N_3269,N_2748,N_2620);
nor U3270 (N_3270,N_2511,N_2596);
and U3271 (N_3271,N_2644,N_2515);
or U3272 (N_3272,N_2557,N_2611);
and U3273 (N_3273,N_2817,N_2626);
and U3274 (N_3274,N_2668,N_2866);
or U3275 (N_3275,N_2697,N_2878);
or U3276 (N_3276,N_2522,N_2854);
or U3277 (N_3277,N_2675,N_2537);
and U3278 (N_3278,N_2807,N_2957);
xnor U3279 (N_3279,N_2802,N_2674);
nand U3280 (N_3280,N_2589,N_2989);
nor U3281 (N_3281,N_2859,N_2799);
and U3282 (N_3282,N_2844,N_2521);
and U3283 (N_3283,N_2915,N_2939);
and U3284 (N_3284,N_2528,N_2676);
and U3285 (N_3285,N_2576,N_2523);
nand U3286 (N_3286,N_2937,N_2598);
nor U3287 (N_3287,N_2696,N_2860);
or U3288 (N_3288,N_2803,N_2555);
and U3289 (N_3289,N_2984,N_2533);
and U3290 (N_3290,N_2510,N_2808);
or U3291 (N_3291,N_2797,N_2902);
nor U3292 (N_3292,N_2737,N_2849);
or U3293 (N_3293,N_2991,N_2810);
and U3294 (N_3294,N_2592,N_2990);
nand U3295 (N_3295,N_2740,N_2777);
and U3296 (N_3296,N_2712,N_2758);
nor U3297 (N_3297,N_2514,N_2664);
or U3298 (N_3298,N_2570,N_2878);
nand U3299 (N_3299,N_2684,N_2519);
or U3300 (N_3300,N_2645,N_2652);
nor U3301 (N_3301,N_2851,N_2754);
or U3302 (N_3302,N_2591,N_2664);
and U3303 (N_3303,N_2892,N_2613);
nand U3304 (N_3304,N_2990,N_2991);
nor U3305 (N_3305,N_2754,N_2891);
and U3306 (N_3306,N_2987,N_2514);
and U3307 (N_3307,N_2920,N_2620);
nor U3308 (N_3308,N_2544,N_2787);
xnor U3309 (N_3309,N_2961,N_2578);
or U3310 (N_3310,N_2868,N_2847);
and U3311 (N_3311,N_2525,N_2938);
and U3312 (N_3312,N_2788,N_2969);
nand U3313 (N_3313,N_2631,N_2897);
xnor U3314 (N_3314,N_2704,N_2673);
and U3315 (N_3315,N_2959,N_2572);
or U3316 (N_3316,N_2796,N_2931);
xor U3317 (N_3317,N_2520,N_2949);
or U3318 (N_3318,N_2671,N_2526);
nor U3319 (N_3319,N_2644,N_2749);
nor U3320 (N_3320,N_2964,N_2516);
xnor U3321 (N_3321,N_2762,N_2549);
or U3322 (N_3322,N_2622,N_2653);
or U3323 (N_3323,N_2888,N_2614);
nand U3324 (N_3324,N_2831,N_2671);
nor U3325 (N_3325,N_2761,N_2579);
and U3326 (N_3326,N_2515,N_2668);
and U3327 (N_3327,N_2670,N_2710);
and U3328 (N_3328,N_2831,N_2716);
xor U3329 (N_3329,N_2947,N_2601);
or U3330 (N_3330,N_2904,N_2877);
nor U3331 (N_3331,N_2772,N_2709);
nand U3332 (N_3332,N_2669,N_2696);
and U3333 (N_3333,N_2530,N_2871);
nor U3334 (N_3334,N_2877,N_2744);
nor U3335 (N_3335,N_2934,N_2635);
or U3336 (N_3336,N_2574,N_2536);
nand U3337 (N_3337,N_2658,N_2773);
xor U3338 (N_3338,N_2985,N_2984);
nand U3339 (N_3339,N_2719,N_2636);
and U3340 (N_3340,N_2599,N_2757);
or U3341 (N_3341,N_2660,N_2664);
and U3342 (N_3342,N_2766,N_2668);
xor U3343 (N_3343,N_2652,N_2884);
or U3344 (N_3344,N_2605,N_2978);
or U3345 (N_3345,N_2520,N_2703);
nor U3346 (N_3346,N_2629,N_2637);
or U3347 (N_3347,N_2815,N_2929);
nor U3348 (N_3348,N_2929,N_2906);
nand U3349 (N_3349,N_2974,N_2715);
and U3350 (N_3350,N_2952,N_2810);
or U3351 (N_3351,N_2792,N_2679);
nand U3352 (N_3352,N_2640,N_2628);
nand U3353 (N_3353,N_2820,N_2591);
nor U3354 (N_3354,N_2551,N_2627);
nand U3355 (N_3355,N_2629,N_2674);
nor U3356 (N_3356,N_2712,N_2905);
nand U3357 (N_3357,N_2642,N_2575);
nor U3358 (N_3358,N_2885,N_2764);
nor U3359 (N_3359,N_2662,N_2689);
nand U3360 (N_3360,N_2642,N_2928);
nor U3361 (N_3361,N_2721,N_2913);
and U3362 (N_3362,N_2796,N_2656);
nand U3363 (N_3363,N_2991,N_2713);
nand U3364 (N_3364,N_2530,N_2562);
nand U3365 (N_3365,N_2632,N_2942);
or U3366 (N_3366,N_2760,N_2959);
or U3367 (N_3367,N_2887,N_2938);
xnor U3368 (N_3368,N_2684,N_2950);
nor U3369 (N_3369,N_2574,N_2884);
and U3370 (N_3370,N_2797,N_2976);
or U3371 (N_3371,N_2603,N_2782);
nand U3372 (N_3372,N_2996,N_2694);
and U3373 (N_3373,N_2805,N_2797);
and U3374 (N_3374,N_2890,N_2845);
or U3375 (N_3375,N_2835,N_2596);
or U3376 (N_3376,N_2746,N_2541);
or U3377 (N_3377,N_2962,N_2818);
or U3378 (N_3378,N_2763,N_2613);
nor U3379 (N_3379,N_2639,N_2655);
nand U3380 (N_3380,N_2843,N_2881);
nor U3381 (N_3381,N_2500,N_2639);
nand U3382 (N_3382,N_2673,N_2543);
nor U3383 (N_3383,N_2777,N_2732);
nand U3384 (N_3384,N_2990,N_2871);
and U3385 (N_3385,N_2948,N_2848);
or U3386 (N_3386,N_2608,N_2863);
nand U3387 (N_3387,N_2608,N_2640);
nand U3388 (N_3388,N_2882,N_2633);
or U3389 (N_3389,N_2967,N_2983);
xnor U3390 (N_3390,N_2593,N_2661);
and U3391 (N_3391,N_2867,N_2590);
xnor U3392 (N_3392,N_2763,N_2997);
and U3393 (N_3393,N_2897,N_2729);
nor U3394 (N_3394,N_2844,N_2757);
or U3395 (N_3395,N_2880,N_2535);
nor U3396 (N_3396,N_2586,N_2561);
nor U3397 (N_3397,N_2585,N_2934);
xnor U3398 (N_3398,N_2874,N_2900);
and U3399 (N_3399,N_2809,N_2621);
or U3400 (N_3400,N_2748,N_2925);
or U3401 (N_3401,N_2959,N_2794);
xor U3402 (N_3402,N_2659,N_2978);
xnor U3403 (N_3403,N_2714,N_2522);
and U3404 (N_3404,N_2694,N_2989);
and U3405 (N_3405,N_2753,N_2957);
or U3406 (N_3406,N_2842,N_2823);
or U3407 (N_3407,N_2801,N_2907);
and U3408 (N_3408,N_2770,N_2545);
or U3409 (N_3409,N_2717,N_2960);
and U3410 (N_3410,N_2782,N_2996);
nor U3411 (N_3411,N_2756,N_2701);
nor U3412 (N_3412,N_2606,N_2811);
and U3413 (N_3413,N_2943,N_2998);
nor U3414 (N_3414,N_2778,N_2705);
nand U3415 (N_3415,N_2543,N_2565);
and U3416 (N_3416,N_2536,N_2974);
xnor U3417 (N_3417,N_2598,N_2554);
and U3418 (N_3418,N_2881,N_2938);
nand U3419 (N_3419,N_2824,N_2872);
nor U3420 (N_3420,N_2606,N_2952);
and U3421 (N_3421,N_2702,N_2588);
nor U3422 (N_3422,N_2885,N_2671);
or U3423 (N_3423,N_2721,N_2589);
and U3424 (N_3424,N_2761,N_2888);
nand U3425 (N_3425,N_2680,N_2973);
and U3426 (N_3426,N_2534,N_2851);
nor U3427 (N_3427,N_2658,N_2872);
nand U3428 (N_3428,N_2790,N_2565);
xnor U3429 (N_3429,N_2731,N_2862);
xor U3430 (N_3430,N_2712,N_2596);
nor U3431 (N_3431,N_2624,N_2604);
nor U3432 (N_3432,N_2612,N_2653);
xnor U3433 (N_3433,N_2621,N_2586);
nand U3434 (N_3434,N_2956,N_2827);
or U3435 (N_3435,N_2770,N_2869);
and U3436 (N_3436,N_2625,N_2524);
and U3437 (N_3437,N_2911,N_2698);
nor U3438 (N_3438,N_2796,N_2716);
nand U3439 (N_3439,N_2661,N_2811);
or U3440 (N_3440,N_2967,N_2829);
or U3441 (N_3441,N_2978,N_2540);
or U3442 (N_3442,N_2823,N_2921);
or U3443 (N_3443,N_2609,N_2960);
nor U3444 (N_3444,N_2666,N_2630);
and U3445 (N_3445,N_2675,N_2548);
nor U3446 (N_3446,N_2889,N_2988);
nand U3447 (N_3447,N_2932,N_2769);
nor U3448 (N_3448,N_2652,N_2513);
nand U3449 (N_3449,N_2900,N_2509);
nand U3450 (N_3450,N_2705,N_2577);
or U3451 (N_3451,N_2667,N_2539);
and U3452 (N_3452,N_2972,N_2691);
or U3453 (N_3453,N_2913,N_2975);
nor U3454 (N_3454,N_2811,N_2989);
xor U3455 (N_3455,N_2550,N_2695);
and U3456 (N_3456,N_2781,N_2728);
or U3457 (N_3457,N_2520,N_2744);
nor U3458 (N_3458,N_2832,N_2820);
or U3459 (N_3459,N_2701,N_2535);
nor U3460 (N_3460,N_2679,N_2526);
or U3461 (N_3461,N_2661,N_2581);
and U3462 (N_3462,N_2917,N_2515);
or U3463 (N_3463,N_2758,N_2984);
and U3464 (N_3464,N_2816,N_2548);
nand U3465 (N_3465,N_2540,N_2992);
and U3466 (N_3466,N_2510,N_2639);
and U3467 (N_3467,N_2818,N_2831);
nand U3468 (N_3468,N_2505,N_2504);
xnor U3469 (N_3469,N_2528,N_2920);
nand U3470 (N_3470,N_2928,N_2683);
nand U3471 (N_3471,N_2766,N_2591);
nand U3472 (N_3472,N_2744,N_2860);
nand U3473 (N_3473,N_2931,N_2840);
and U3474 (N_3474,N_2678,N_2829);
or U3475 (N_3475,N_2950,N_2553);
nor U3476 (N_3476,N_2593,N_2951);
nor U3477 (N_3477,N_2503,N_2909);
xnor U3478 (N_3478,N_2540,N_2587);
nand U3479 (N_3479,N_2886,N_2891);
nor U3480 (N_3480,N_2969,N_2943);
nand U3481 (N_3481,N_2510,N_2903);
and U3482 (N_3482,N_2814,N_2691);
nand U3483 (N_3483,N_2604,N_2966);
nor U3484 (N_3484,N_2908,N_2875);
and U3485 (N_3485,N_2852,N_2832);
and U3486 (N_3486,N_2526,N_2681);
nand U3487 (N_3487,N_2793,N_2576);
nand U3488 (N_3488,N_2697,N_2927);
or U3489 (N_3489,N_2820,N_2798);
or U3490 (N_3490,N_2610,N_2665);
or U3491 (N_3491,N_2890,N_2545);
xnor U3492 (N_3492,N_2875,N_2888);
nor U3493 (N_3493,N_2559,N_2822);
xor U3494 (N_3494,N_2549,N_2932);
nand U3495 (N_3495,N_2547,N_2932);
xnor U3496 (N_3496,N_2683,N_2589);
nand U3497 (N_3497,N_2519,N_2817);
nor U3498 (N_3498,N_2648,N_2834);
or U3499 (N_3499,N_2859,N_2838);
and U3500 (N_3500,N_3458,N_3059);
xor U3501 (N_3501,N_3072,N_3033);
nand U3502 (N_3502,N_3289,N_3073);
nor U3503 (N_3503,N_3367,N_3281);
or U3504 (N_3504,N_3125,N_3435);
nor U3505 (N_3505,N_3455,N_3209);
xor U3506 (N_3506,N_3296,N_3357);
nor U3507 (N_3507,N_3350,N_3321);
and U3508 (N_3508,N_3362,N_3304);
nand U3509 (N_3509,N_3147,N_3473);
nand U3510 (N_3510,N_3268,N_3356);
xor U3511 (N_3511,N_3271,N_3444);
nor U3512 (N_3512,N_3460,N_3194);
and U3513 (N_3513,N_3273,N_3387);
xnor U3514 (N_3514,N_3115,N_3351);
nand U3515 (N_3515,N_3060,N_3323);
nand U3516 (N_3516,N_3173,N_3320);
nand U3517 (N_3517,N_3461,N_3233);
nor U3518 (N_3518,N_3294,N_3011);
xnor U3519 (N_3519,N_3405,N_3463);
or U3520 (N_3520,N_3089,N_3074);
nand U3521 (N_3521,N_3091,N_3383);
nor U3522 (N_3522,N_3347,N_3199);
xor U3523 (N_3523,N_3198,N_3137);
nand U3524 (N_3524,N_3385,N_3242);
or U3525 (N_3525,N_3348,N_3124);
nand U3526 (N_3526,N_3311,N_3017);
xnor U3527 (N_3527,N_3258,N_3433);
nand U3528 (N_3528,N_3181,N_3338);
and U3529 (N_3529,N_3134,N_3226);
or U3530 (N_3530,N_3277,N_3432);
or U3531 (N_3531,N_3167,N_3427);
or U3532 (N_3532,N_3018,N_3007);
and U3533 (N_3533,N_3131,N_3122);
nor U3534 (N_3534,N_3231,N_3392);
nand U3535 (N_3535,N_3299,N_3412);
and U3536 (N_3536,N_3256,N_3334);
nand U3537 (N_3537,N_3439,N_3168);
nor U3538 (N_3538,N_3141,N_3006);
and U3539 (N_3539,N_3228,N_3327);
or U3540 (N_3540,N_3140,N_3036);
nor U3541 (N_3541,N_3152,N_3224);
nor U3542 (N_3542,N_3210,N_3054);
or U3543 (N_3543,N_3428,N_3062);
nor U3544 (N_3544,N_3494,N_3204);
nand U3545 (N_3545,N_3182,N_3021);
or U3546 (N_3546,N_3312,N_3229);
nor U3547 (N_3547,N_3407,N_3093);
xnor U3548 (N_3548,N_3471,N_3041);
nor U3549 (N_3549,N_3274,N_3485);
and U3550 (N_3550,N_3488,N_3113);
nor U3551 (N_3551,N_3213,N_3430);
and U3552 (N_3552,N_3051,N_3175);
nand U3553 (N_3553,N_3102,N_3222);
and U3554 (N_3554,N_3138,N_3365);
and U3555 (N_3555,N_3389,N_3077);
or U3556 (N_3556,N_3090,N_3078);
or U3557 (N_3557,N_3223,N_3450);
or U3558 (N_3558,N_3331,N_3293);
nand U3559 (N_3559,N_3378,N_3086);
xnor U3560 (N_3560,N_3390,N_3163);
and U3561 (N_3561,N_3453,N_3215);
or U3562 (N_3562,N_3470,N_3448);
or U3563 (N_3563,N_3442,N_3434);
or U3564 (N_3564,N_3094,N_3493);
xor U3565 (N_3565,N_3401,N_3447);
xor U3566 (N_3566,N_3451,N_3066);
or U3567 (N_3567,N_3128,N_3449);
nor U3568 (N_3568,N_3219,N_3034);
nand U3569 (N_3569,N_3001,N_3146);
nand U3570 (N_3570,N_3180,N_3285);
nor U3571 (N_3571,N_3216,N_3440);
and U3572 (N_3572,N_3490,N_3329);
and U3573 (N_3573,N_3156,N_3382);
nor U3574 (N_3574,N_3445,N_3040);
or U3575 (N_3575,N_3038,N_3197);
or U3576 (N_3576,N_3068,N_3272);
and U3577 (N_3577,N_3375,N_3190);
nor U3578 (N_3578,N_3349,N_3438);
and U3579 (N_3579,N_3243,N_3298);
or U3580 (N_3580,N_3003,N_3280);
or U3581 (N_3581,N_3368,N_3415);
nand U3582 (N_3582,N_3087,N_3225);
or U3583 (N_3583,N_3227,N_3107);
nor U3584 (N_3584,N_3393,N_3254);
nor U3585 (N_3585,N_3363,N_3101);
nand U3586 (N_3586,N_3238,N_3100);
xor U3587 (N_3587,N_3208,N_3316);
and U3588 (N_3588,N_3241,N_3381);
and U3589 (N_3589,N_3437,N_3446);
and U3590 (N_3590,N_3030,N_3295);
or U3591 (N_3591,N_3014,N_3234);
or U3592 (N_3592,N_3267,N_3178);
nor U3593 (N_3593,N_3015,N_3340);
or U3594 (N_3594,N_3031,N_3307);
and U3595 (N_3595,N_3203,N_3151);
nor U3596 (N_3596,N_3291,N_3145);
nand U3597 (N_3597,N_3333,N_3244);
or U3598 (N_3598,N_3027,N_3478);
nor U3599 (N_3599,N_3499,N_3235);
or U3600 (N_3600,N_3284,N_3290);
nand U3601 (N_3601,N_3118,N_3196);
or U3602 (N_3602,N_3346,N_3045);
or U3603 (N_3603,N_3263,N_3133);
nand U3604 (N_3604,N_3425,N_3026);
and U3605 (N_3605,N_3024,N_3020);
and U3606 (N_3606,N_3332,N_3337);
nand U3607 (N_3607,N_3217,N_3106);
nand U3608 (N_3608,N_3257,N_3098);
and U3609 (N_3609,N_3088,N_3396);
nand U3610 (N_3610,N_3221,N_3220);
and U3611 (N_3611,N_3000,N_3404);
and U3612 (N_3612,N_3050,N_3160);
nand U3613 (N_3613,N_3028,N_3154);
and U3614 (N_3614,N_3370,N_3341);
or U3615 (N_3615,N_3397,N_3399);
or U3616 (N_3616,N_3092,N_3372);
nor U3617 (N_3617,N_3408,N_3322);
or U3618 (N_3618,N_3057,N_3424);
nor U3619 (N_3619,N_3328,N_3358);
or U3620 (N_3620,N_3245,N_3373);
nor U3621 (N_3621,N_3330,N_3179);
nor U3622 (N_3622,N_3207,N_3201);
and U3623 (N_3623,N_3048,N_3162);
xor U3624 (N_3624,N_3039,N_3476);
nor U3625 (N_3625,N_3465,N_3306);
nor U3626 (N_3626,N_3416,N_3459);
or U3627 (N_3627,N_3300,N_3023);
nor U3628 (N_3628,N_3269,N_3161);
or U3629 (N_3629,N_3126,N_3398);
nor U3630 (N_3630,N_3104,N_3343);
and U3631 (N_3631,N_3353,N_3130);
nand U3632 (N_3632,N_3336,N_3409);
and U3633 (N_3633,N_3029,N_3352);
and U3634 (N_3634,N_3276,N_3344);
or U3635 (N_3635,N_3313,N_3315);
nand U3636 (N_3636,N_3139,N_3103);
or U3637 (N_3637,N_3153,N_3487);
or U3638 (N_3638,N_3489,N_3359);
nand U3639 (N_3639,N_3302,N_3135);
nand U3640 (N_3640,N_3261,N_3319);
nor U3641 (N_3641,N_3108,N_3369);
and U3642 (N_3642,N_3114,N_3441);
xnor U3643 (N_3643,N_3195,N_3251);
or U3644 (N_3644,N_3264,N_3046);
and U3645 (N_3645,N_3047,N_3481);
or U3646 (N_3646,N_3468,N_3127);
or U3647 (N_3647,N_3065,N_3394);
xor U3648 (N_3648,N_3165,N_3248);
and U3649 (N_3649,N_3486,N_3009);
or U3650 (N_3650,N_3212,N_3177);
and U3651 (N_3651,N_3454,N_3043);
nand U3652 (N_3652,N_3121,N_3097);
and U3653 (N_3653,N_3288,N_3308);
nor U3654 (N_3654,N_3474,N_3236);
nor U3655 (N_3655,N_3035,N_3022);
xnor U3656 (N_3656,N_3452,N_3200);
or U3657 (N_3657,N_3232,N_3063);
and U3658 (N_3658,N_3374,N_3172);
xnor U3659 (N_3659,N_3037,N_3067);
and U3660 (N_3660,N_3411,N_3426);
and U3661 (N_3661,N_3164,N_3071);
or U3662 (N_3662,N_3052,N_3469);
and U3663 (N_3663,N_3422,N_3270);
or U3664 (N_3664,N_3237,N_3150);
nor U3665 (N_3665,N_3053,N_3082);
or U3666 (N_3666,N_3266,N_3218);
nor U3667 (N_3667,N_3155,N_3191);
nand U3668 (N_3668,N_3070,N_3120);
xnor U3669 (N_3669,N_3230,N_3081);
nor U3670 (N_3670,N_3205,N_3143);
or U3671 (N_3671,N_3119,N_3410);
or U3672 (N_3672,N_3158,N_3123);
nor U3673 (N_3673,N_3297,N_3326);
and U3674 (N_3674,N_3149,N_3008);
xor U3675 (N_3675,N_3477,N_3085);
nor U3676 (N_3676,N_3391,N_3044);
and U3677 (N_3677,N_3166,N_3279);
nand U3678 (N_3678,N_3250,N_3099);
nor U3679 (N_3679,N_3246,N_3169);
or U3680 (N_3680,N_3206,N_3176);
and U3681 (N_3681,N_3325,N_3283);
or U3682 (N_3682,N_3364,N_3116);
or U3683 (N_3683,N_3402,N_3170);
nor U3684 (N_3684,N_3419,N_3292);
and U3685 (N_3685,N_3183,N_3467);
nand U3686 (N_3686,N_3142,N_3324);
nand U3687 (N_3687,N_3380,N_3386);
or U3688 (N_3688,N_3184,N_3260);
or U3689 (N_3689,N_3211,N_3025);
or U3690 (N_3690,N_3032,N_3105);
or U3691 (N_3691,N_3421,N_3443);
and U3692 (N_3692,N_3069,N_3318);
xnor U3693 (N_3693,N_3005,N_3076);
nor U3694 (N_3694,N_3431,N_3472);
xnor U3695 (N_3695,N_3278,N_3482);
and U3696 (N_3696,N_3317,N_3305);
or U3697 (N_3697,N_3335,N_3144);
nor U3698 (N_3698,N_3174,N_3189);
nor U3699 (N_3699,N_3498,N_3188);
or U3700 (N_3700,N_3491,N_3464);
or U3701 (N_3701,N_3019,N_3436);
nor U3702 (N_3702,N_3202,N_3406);
xor U3703 (N_3703,N_3496,N_3186);
nor U3704 (N_3704,N_3012,N_3360);
and U3705 (N_3705,N_3002,N_3016);
nor U3706 (N_3706,N_3010,N_3148);
and U3707 (N_3707,N_3287,N_3379);
and U3708 (N_3708,N_3413,N_3004);
or U3709 (N_3709,N_3282,N_3253);
nand U3710 (N_3710,N_3129,N_3497);
nand U3711 (N_3711,N_3262,N_3495);
and U3712 (N_3712,N_3423,N_3286);
and U3713 (N_3713,N_3310,N_3388);
or U3714 (N_3714,N_3117,N_3420);
or U3715 (N_3715,N_3275,N_3239);
and U3716 (N_3716,N_3171,N_3084);
or U3717 (N_3717,N_3354,N_3042);
xor U3718 (N_3718,N_3214,N_3303);
or U3719 (N_3719,N_3055,N_3058);
nor U3720 (N_3720,N_3249,N_3345);
nor U3721 (N_3721,N_3265,N_3064);
nand U3722 (N_3722,N_3480,N_3457);
or U3723 (N_3723,N_3376,N_3456);
xor U3724 (N_3724,N_3079,N_3403);
nand U3725 (N_3725,N_3483,N_3247);
nand U3726 (N_3726,N_3095,N_3366);
and U3727 (N_3727,N_3429,N_3110);
or U3728 (N_3728,N_3400,N_3484);
or U3729 (N_3729,N_3309,N_3466);
and U3730 (N_3730,N_3395,N_3414);
and U3731 (N_3731,N_3361,N_3240);
nor U3732 (N_3732,N_3462,N_3049);
and U3733 (N_3733,N_3080,N_3112);
nand U3734 (N_3734,N_3061,N_3187);
nor U3735 (N_3735,N_3159,N_3418);
nand U3736 (N_3736,N_3301,N_3192);
nor U3737 (N_3737,N_3083,N_3111);
and U3738 (N_3738,N_3075,N_3384);
xor U3739 (N_3739,N_3096,N_3377);
xnor U3740 (N_3740,N_3371,N_3185);
nand U3741 (N_3741,N_3132,N_3255);
nand U3742 (N_3742,N_3475,N_3109);
or U3743 (N_3743,N_3417,N_3136);
nor U3744 (N_3744,N_3259,N_3342);
or U3745 (N_3745,N_3013,N_3479);
nand U3746 (N_3746,N_3355,N_3492);
nand U3747 (N_3747,N_3252,N_3056);
or U3748 (N_3748,N_3314,N_3193);
or U3749 (N_3749,N_3157,N_3339);
nor U3750 (N_3750,N_3407,N_3066);
xnor U3751 (N_3751,N_3260,N_3353);
and U3752 (N_3752,N_3221,N_3270);
or U3753 (N_3753,N_3015,N_3416);
nor U3754 (N_3754,N_3332,N_3447);
nand U3755 (N_3755,N_3429,N_3387);
and U3756 (N_3756,N_3221,N_3324);
and U3757 (N_3757,N_3223,N_3059);
nor U3758 (N_3758,N_3211,N_3037);
or U3759 (N_3759,N_3369,N_3065);
nand U3760 (N_3760,N_3275,N_3026);
nor U3761 (N_3761,N_3265,N_3360);
nand U3762 (N_3762,N_3086,N_3401);
xnor U3763 (N_3763,N_3090,N_3011);
or U3764 (N_3764,N_3332,N_3037);
and U3765 (N_3765,N_3311,N_3447);
and U3766 (N_3766,N_3142,N_3495);
or U3767 (N_3767,N_3104,N_3192);
or U3768 (N_3768,N_3389,N_3134);
nand U3769 (N_3769,N_3345,N_3369);
and U3770 (N_3770,N_3018,N_3432);
or U3771 (N_3771,N_3436,N_3499);
or U3772 (N_3772,N_3301,N_3422);
or U3773 (N_3773,N_3308,N_3293);
xor U3774 (N_3774,N_3383,N_3405);
and U3775 (N_3775,N_3025,N_3465);
nand U3776 (N_3776,N_3040,N_3420);
nand U3777 (N_3777,N_3252,N_3426);
nand U3778 (N_3778,N_3136,N_3111);
and U3779 (N_3779,N_3065,N_3023);
nor U3780 (N_3780,N_3260,N_3347);
nand U3781 (N_3781,N_3290,N_3095);
and U3782 (N_3782,N_3453,N_3300);
or U3783 (N_3783,N_3247,N_3053);
nor U3784 (N_3784,N_3006,N_3249);
nor U3785 (N_3785,N_3114,N_3346);
and U3786 (N_3786,N_3162,N_3263);
or U3787 (N_3787,N_3411,N_3310);
nor U3788 (N_3788,N_3088,N_3482);
or U3789 (N_3789,N_3458,N_3003);
nor U3790 (N_3790,N_3458,N_3211);
nor U3791 (N_3791,N_3067,N_3062);
and U3792 (N_3792,N_3316,N_3047);
nand U3793 (N_3793,N_3431,N_3486);
xnor U3794 (N_3794,N_3317,N_3399);
nor U3795 (N_3795,N_3103,N_3156);
nand U3796 (N_3796,N_3013,N_3436);
nand U3797 (N_3797,N_3445,N_3140);
and U3798 (N_3798,N_3146,N_3478);
and U3799 (N_3799,N_3172,N_3153);
or U3800 (N_3800,N_3195,N_3182);
and U3801 (N_3801,N_3409,N_3225);
xor U3802 (N_3802,N_3082,N_3469);
nor U3803 (N_3803,N_3068,N_3017);
xnor U3804 (N_3804,N_3119,N_3469);
and U3805 (N_3805,N_3277,N_3274);
and U3806 (N_3806,N_3463,N_3272);
and U3807 (N_3807,N_3172,N_3282);
and U3808 (N_3808,N_3243,N_3258);
nor U3809 (N_3809,N_3408,N_3349);
and U3810 (N_3810,N_3359,N_3402);
nand U3811 (N_3811,N_3342,N_3468);
nor U3812 (N_3812,N_3308,N_3070);
nor U3813 (N_3813,N_3215,N_3214);
nand U3814 (N_3814,N_3413,N_3175);
nor U3815 (N_3815,N_3132,N_3288);
and U3816 (N_3816,N_3164,N_3153);
nand U3817 (N_3817,N_3111,N_3240);
and U3818 (N_3818,N_3096,N_3376);
nor U3819 (N_3819,N_3302,N_3410);
nor U3820 (N_3820,N_3313,N_3163);
nor U3821 (N_3821,N_3214,N_3420);
and U3822 (N_3822,N_3239,N_3479);
and U3823 (N_3823,N_3237,N_3296);
and U3824 (N_3824,N_3242,N_3187);
nand U3825 (N_3825,N_3402,N_3362);
xor U3826 (N_3826,N_3458,N_3244);
and U3827 (N_3827,N_3410,N_3354);
and U3828 (N_3828,N_3128,N_3197);
nand U3829 (N_3829,N_3336,N_3476);
nor U3830 (N_3830,N_3020,N_3028);
xnor U3831 (N_3831,N_3090,N_3043);
and U3832 (N_3832,N_3266,N_3446);
and U3833 (N_3833,N_3340,N_3454);
or U3834 (N_3834,N_3082,N_3013);
or U3835 (N_3835,N_3450,N_3098);
and U3836 (N_3836,N_3016,N_3426);
nor U3837 (N_3837,N_3104,N_3339);
nand U3838 (N_3838,N_3381,N_3020);
nor U3839 (N_3839,N_3305,N_3226);
nor U3840 (N_3840,N_3355,N_3161);
or U3841 (N_3841,N_3451,N_3059);
nor U3842 (N_3842,N_3416,N_3217);
nand U3843 (N_3843,N_3108,N_3495);
and U3844 (N_3844,N_3374,N_3124);
and U3845 (N_3845,N_3134,N_3420);
or U3846 (N_3846,N_3249,N_3273);
or U3847 (N_3847,N_3261,N_3370);
nand U3848 (N_3848,N_3075,N_3095);
or U3849 (N_3849,N_3167,N_3250);
nand U3850 (N_3850,N_3445,N_3422);
nor U3851 (N_3851,N_3072,N_3048);
or U3852 (N_3852,N_3392,N_3199);
and U3853 (N_3853,N_3469,N_3344);
nor U3854 (N_3854,N_3342,N_3244);
xnor U3855 (N_3855,N_3351,N_3259);
or U3856 (N_3856,N_3031,N_3156);
and U3857 (N_3857,N_3337,N_3456);
or U3858 (N_3858,N_3166,N_3028);
nor U3859 (N_3859,N_3224,N_3049);
xor U3860 (N_3860,N_3065,N_3412);
and U3861 (N_3861,N_3067,N_3469);
nand U3862 (N_3862,N_3426,N_3245);
and U3863 (N_3863,N_3368,N_3364);
and U3864 (N_3864,N_3298,N_3439);
or U3865 (N_3865,N_3080,N_3308);
nand U3866 (N_3866,N_3481,N_3042);
or U3867 (N_3867,N_3199,N_3273);
and U3868 (N_3868,N_3204,N_3270);
nand U3869 (N_3869,N_3214,N_3110);
xnor U3870 (N_3870,N_3370,N_3189);
nor U3871 (N_3871,N_3305,N_3299);
or U3872 (N_3872,N_3115,N_3036);
xnor U3873 (N_3873,N_3486,N_3055);
xnor U3874 (N_3874,N_3136,N_3001);
and U3875 (N_3875,N_3195,N_3119);
nand U3876 (N_3876,N_3408,N_3373);
nor U3877 (N_3877,N_3354,N_3323);
nor U3878 (N_3878,N_3347,N_3499);
or U3879 (N_3879,N_3393,N_3331);
or U3880 (N_3880,N_3474,N_3086);
xor U3881 (N_3881,N_3088,N_3169);
or U3882 (N_3882,N_3450,N_3268);
nand U3883 (N_3883,N_3436,N_3326);
nor U3884 (N_3884,N_3357,N_3463);
xnor U3885 (N_3885,N_3405,N_3114);
and U3886 (N_3886,N_3008,N_3496);
xnor U3887 (N_3887,N_3229,N_3329);
xnor U3888 (N_3888,N_3381,N_3364);
or U3889 (N_3889,N_3060,N_3103);
nor U3890 (N_3890,N_3452,N_3106);
and U3891 (N_3891,N_3286,N_3114);
nor U3892 (N_3892,N_3464,N_3037);
nand U3893 (N_3893,N_3162,N_3120);
and U3894 (N_3894,N_3210,N_3172);
or U3895 (N_3895,N_3340,N_3187);
and U3896 (N_3896,N_3364,N_3433);
and U3897 (N_3897,N_3009,N_3307);
xor U3898 (N_3898,N_3174,N_3017);
nand U3899 (N_3899,N_3349,N_3008);
nand U3900 (N_3900,N_3162,N_3336);
xor U3901 (N_3901,N_3116,N_3024);
nor U3902 (N_3902,N_3450,N_3192);
or U3903 (N_3903,N_3240,N_3300);
nand U3904 (N_3904,N_3289,N_3171);
nor U3905 (N_3905,N_3002,N_3396);
and U3906 (N_3906,N_3269,N_3412);
nand U3907 (N_3907,N_3319,N_3376);
and U3908 (N_3908,N_3496,N_3356);
or U3909 (N_3909,N_3187,N_3018);
nor U3910 (N_3910,N_3487,N_3324);
nor U3911 (N_3911,N_3350,N_3183);
nand U3912 (N_3912,N_3098,N_3083);
and U3913 (N_3913,N_3465,N_3429);
nand U3914 (N_3914,N_3138,N_3245);
and U3915 (N_3915,N_3129,N_3136);
or U3916 (N_3916,N_3183,N_3004);
xnor U3917 (N_3917,N_3185,N_3466);
or U3918 (N_3918,N_3148,N_3192);
xor U3919 (N_3919,N_3178,N_3164);
nor U3920 (N_3920,N_3108,N_3405);
and U3921 (N_3921,N_3086,N_3014);
xnor U3922 (N_3922,N_3394,N_3107);
or U3923 (N_3923,N_3493,N_3056);
or U3924 (N_3924,N_3250,N_3031);
nor U3925 (N_3925,N_3152,N_3489);
and U3926 (N_3926,N_3127,N_3464);
or U3927 (N_3927,N_3223,N_3257);
or U3928 (N_3928,N_3156,N_3153);
nor U3929 (N_3929,N_3327,N_3309);
or U3930 (N_3930,N_3204,N_3433);
nand U3931 (N_3931,N_3367,N_3327);
and U3932 (N_3932,N_3178,N_3453);
nand U3933 (N_3933,N_3162,N_3208);
and U3934 (N_3934,N_3397,N_3239);
or U3935 (N_3935,N_3201,N_3142);
nor U3936 (N_3936,N_3246,N_3272);
nor U3937 (N_3937,N_3358,N_3046);
nor U3938 (N_3938,N_3210,N_3372);
nor U3939 (N_3939,N_3105,N_3095);
or U3940 (N_3940,N_3420,N_3494);
xnor U3941 (N_3941,N_3250,N_3366);
nand U3942 (N_3942,N_3132,N_3212);
nand U3943 (N_3943,N_3282,N_3484);
and U3944 (N_3944,N_3188,N_3499);
or U3945 (N_3945,N_3158,N_3431);
or U3946 (N_3946,N_3143,N_3499);
nand U3947 (N_3947,N_3087,N_3329);
or U3948 (N_3948,N_3193,N_3266);
nand U3949 (N_3949,N_3357,N_3281);
xnor U3950 (N_3950,N_3035,N_3376);
xor U3951 (N_3951,N_3250,N_3185);
or U3952 (N_3952,N_3255,N_3042);
or U3953 (N_3953,N_3254,N_3436);
nand U3954 (N_3954,N_3483,N_3140);
or U3955 (N_3955,N_3166,N_3271);
and U3956 (N_3956,N_3118,N_3243);
nor U3957 (N_3957,N_3305,N_3449);
nand U3958 (N_3958,N_3076,N_3031);
xnor U3959 (N_3959,N_3160,N_3250);
and U3960 (N_3960,N_3118,N_3298);
or U3961 (N_3961,N_3000,N_3206);
and U3962 (N_3962,N_3452,N_3272);
and U3963 (N_3963,N_3457,N_3248);
nand U3964 (N_3964,N_3355,N_3262);
nor U3965 (N_3965,N_3044,N_3323);
nand U3966 (N_3966,N_3074,N_3343);
or U3967 (N_3967,N_3181,N_3066);
xnor U3968 (N_3968,N_3267,N_3118);
and U3969 (N_3969,N_3354,N_3006);
nand U3970 (N_3970,N_3495,N_3010);
nand U3971 (N_3971,N_3187,N_3114);
nand U3972 (N_3972,N_3167,N_3477);
nor U3973 (N_3973,N_3041,N_3006);
nor U3974 (N_3974,N_3125,N_3092);
or U3975 (N_3975,N_3027,N_3289);
or U3976 (N_3976,N_3372,N_3406);
xor U3977 (N_3977,N_3440,N_3480);
and U3978 (N_3978,N_3005,N_3160);
or U3979 (N_3979,N_3405,N_3461);
nor U3980 (N_3980,N_3474,N_3432);
and U3981 (N_3981,N_3397,N_3418);
and U3982 (N_3982,N_3143,N_3358);
nand U3983 (N_3983,N_3322,N_3058);
or U3984 (N_3984,N_3163,N_3191);
and U3985 (N_3985,N_3053,N_3073);
xnor U3986 (N_3986,N_3353,N_3189);
nor U3987 (N_3987,N_3120,N_3128);
and U3988 (N_3988,N_3384,N_3480);
nor U3989 (N_3989,N_3203,N_3258);
or U3990 (N_3990,N_3085,N_3248);
and U3991 (N_3991,N_3481,N_3473);
and U3992 (N_3992,N_3475,N_3120);
or U3993 (N_3993,N_3336,N_3118);
nand U3994 (N_3994,N_3285,N_3231);
and U3995 (N_3995,N_3054,N_3273);
nand U3996 (N_3996,N_3433,N_3354);
or U3997 (N_3997,N_3067,N_3036);
nor U3998 (N_3998,N_3309,N_3390);
or U3999 (N_3999,N_3276,N_3197);
or U4000 (N_4000,N_3642,N_3655);
or U4001 (N_4001,N_3966,N_3889);
nor U4002 (N_4002,N_3530,N_3811);
or U4003 (N_4003,N_3837,N_3677);
nand U4004 (N_4004,N_3576,N_3924);
or U4005 (N_4005,N_3518,N_3728);
or U4006 (N_4006,N_3606,N_3796);
or U4007 (N_4007,N_3885,N_3844);
nor U4008 (N_4008,N_3734,N_3534);
nor U4009 (N_4009,N_3639,N_3542);
nor U4010 (N_4010,N_3672,N_3787);
nand U4011 (N_4011,N_3873,N_3520);
nor U4012 (N_4012,N_3570,N_3609);
and U4013 (N_4013,N_3704,N_3775);
nor U4014 (N_4014,N_3824,N_3954);
or U4015 (N_4015,N_3827,N_3745);
or U4016 (N_4016,N_3867,N_3778);
and U4017 (N_4017,N_3963,N_3846);
nand U4018 (N_4018,N_3925,N_3583);
or U4019 (N_4019,N_3644,N_3860);
and U4020 (N_4020,N_3614,N_3607);
nor U4021 (N_4021,N_3983,N_3508);
nand U4022 (N_4022,N_3957,N_3652);
and U4023 (N_4023,N_3633,N_3551);
or U4024 (N_4024,N_3905,N_3658);
or U4025 (N_4025,N_3931,N_3956);
or U4026 (N_4026,N_3955,N_3635);
and U4027 (N_4027,N_3967,N_3808);
or U4028 (N_4028,N_3501,N_3654);
or U4029 (N_4029,N_3690,N_3555);
and U4030 (N_4030,N_3884,N_3562);
nand U4031 (N_4031,N_3737,N_3777);
nand U4032 (N_4032,N_3507,N_3932);
nand U4033 (N_4033,N_3544,N_3820);
nor U4034 (N_4034,N_3726,N_3693);
or U4035 (N_4035,N_3618,N_3865);
or U4036 (N_4036,N_3667,N_3676);
and U4037 (N_4037,N_3664,N_3879);
nand U4038 (N_4038,N_3743,N_3521);
nor U4039 (N_4039,N_3603,N_3733);
or U4040 (N_4040,N_3647,N_3958);
nor U4041 (N_4041,N_3821,N_3622);
or U4042 (N_4042,N_3640,N_3812);
or U4043 (N_4043,N_3691,N_3862);
or U4044 (N_4044,N_3757,N_3941);
nand U4045 (N_4045,N_3526,N_3571);
or U4046 (N_4046,N_3872,N_3561);
and U4047 (N_4047,N_3505,N_3703);
and U4048 (N_4048,N_3522,N_3510);
nor U4049 (N_4049,N_3921,N_3810);
and U4050 (N_4050,N_3517,N_3709);
or U4051 (N_4051,N_3856,N_3786);
nor U4052 (N_4052,N_3926,N_3539);
and U4053 (N_4053,N_3888,N_3572);
or U4054 (N_4054,N_3779,N_3557);
and U4055 (N_4055,N_3999,N_3683);
nand U4056 (N_4056,N_3506,N_3758);
nor U4057 (N_4057,N_3759,N_3797);
or U4058 (N_4058,N_3536,N_3776);
or U4059 (N_4059,N_3886,N_3706);
nor U4060 (N_4060,N_3568,N_3964);
or U4061 (N_4061,N_3574,N_3825);
nor U4062 (N_4062,N_3817,N_3880);
xor U4063 (N_4063,N_3632,N_3752);
or U4064 (N_4064,N_3564,N_3537);
nor U4065 (N_4065,N_3848,N_3951);
or U4066 (N_4066,N_3813,N_3806);
nor U4067 (N_4067,N_3624,N_3826);
and U4068 (N_4068,N_3604,N_3927);
and U4069 (N_4069,N_3515,N_3906);
nand U4070 (N_4070,N_3877,N_3528);
and U4071 (N_4071,N_3849,N_3790);
and U4072 (N_4072,N_3836,N_3689);
nor U4073 (N_4073,N_3765,N_3898);
or U4074 (N_4074,N_3547,N_3535);
and U4075 (N_4075,N_3916,N_3697);
and U4076 (N_4076,N_3795,N_3649);
nand U4077 (N_4077,N_3513,N_3611);
nand U4078 (N_4078,N_3976,N_3519);
or U4079 (N_4079,N_3866,N_3991);
xor U4080 (N_4080,N_3788,N_3558);
and U4081 (N_4081,N_3656,N_3823);
xor U4082 (N_4082,N_3567,N_3679);
or U4083 (N_4083,N_3863,N_3764);
nor U4084 (N_4084,N_3769,N_3628);
nor U4085 (N_4085,N_3504,N_3887);
and U4086 (N_4086,N_3678,N_3590);
or U4087 (N_4087,N_3828,N_3936);
and U4088 (N_4088,N_3735,N_3566);
xnor U4089 (N_4089,N_3587,N_3597);
or U4090 (N_4090,N_3782,N_3629);
or U4091 (N_4091,N_3962,N_3948);
or U4092 (N_4092,N_3917,N_3914);
and U4093 (N_4093,N_3721,N_3741);
or U4094 (N_4094,N_3659,N_3852);
or U4095 (N_4095,N_3708,N_3700);
nor U4096 (N_4096,N_3780,N_3578);
xnor U4097 (N_4097,N_3593,N_3892);
and U4098 (N_4098,N_3601,N_3746);
and U4099 (N_4099,N_3723,N_3938);
xnor U4100 (N_4100,N_3763,N_3935);
or U4101 (N_4101,N_3871,N_3694);
nor U4102 (N_4102,N_3512,N_3615);
nand U4103 (N_4103,N_3992,N_3680);
or U4104 (N_4104,N_3878,N_3750);
nor U4105 (N_4105,N_3563,N_3623);
nand U4106 (N_4106,N_3641,N_3774);
nor U4107 (N_4107,N_3929,N_3793);
nor U4108 (N_4108,N_3696,N_3854);
nand U4109 (N_4109,N_3538,N_3523);
or U4110 (N_4110,N_3684,N_3949);
and U4111 (N_4111,N_3833,N_3977);
nor U4112 (N_4112,N_3897,N_3663);
nand U4113 (N_4113,N_3533,N_3959);
nor U4114 (N_4114,N_3648,N_3748);
and U4115 (N_4115,N_3972,N_3586);
or U4116 (N_4116,N_3993,N_3937);
nand U4117 (N_4117,N_3985,N_3875);
and U4118 (N_4118,N_3612,N_3975);
or U4119 (N_4119,N_3724,N_3822);
nand U4120 (N_4120,N_3725,N_3876);
xor U4121 (N_4121,N_3631,N_3982);
nor U4122 (N_4122,N_3531,N_3702);
or U4123 (N_4123,N_3989,N_3996);
xnor U4124 (N_4124,N_3695,N_3660);
nand U4125 (N_4125,N_3784,N_3969);
and U4126 (N_4126,N_3920,N_3918);
xor U4127 (N_4127,N_3781,N_3843);
or U4128 (N_4128,N_3653,N_3789);
or U4129 (N_4129,N_3747,N_3911);
nor U4130 (N_4130,N_3699,N_3502);
nor U4131 (N_4131,N_3634,N_3850);
and U4132 (N_4132,N_3608,N_3627);
and U4133 (N_4133,N_3908,N_3807);
or U4134 (N_4134,N_3981,N_3870);
and U4135 (N_4135,N_3881,N_3751);
nand U4136 (N_4136,N_3912,N_3580);
nor U4137 (N_4137,N_3541,N_3625);
or U4138 (N_4138,N_3998,N_3895);
nand U4139 (N_4139,N_3891,N_3990);
xnor U4140 (N_4140,N_3543,N_3589);
and U4141 (N_4141,N_3740,N_3718);
nor U4142 (N_4142,N_3668,N_3804);
and U4143 (N_4143,N_3556,N_3939);
nor U4144 (N_4144,N_3902,N_3588);
nor U4145 (N_4145,N_3933,N_3961);
nor U4146 (N_4146,N_3829,N_3753);
or U4147 (N_4147,N_3548,N_3698);
nor U4148 (N_4148,N_3947,N_3711);
nand U4149 (N_4149,N_3591,N_3670);
xnor U4150 (N_4150,N_3730,N_3638);
or U4151 (N_4151,N_3552,N_3979);
nor U4152 (N_4152,N_3688,N_3845);
xor U4153 (N_4153,N_3953,N_3617);
and U4154 (N_4154,N_3995,N_3835);
or U4155 (N_4155,N_3545,N_3864);
nand U4156 (N_4156,N_3525,N_3754);
nand U4157 (N_4157,N_3665,N_3883);
xor U4158 (N_4158,N_3869,N_3859);
xnor U4159 (N_4159,N_3940,N_3681);
nand U4160 (N_4160,N_3626,N_3973);
and U4161 (N_4161,N_3714,N_3994);
nor U4162 (N_4162,N_3692,N_3853);
xnor U4163 (N_4163,N_3942,N_3974);
and U4164 (N_4164,N_3952,N_3838);
nand U4165 (N_4165,N_3645,N_3762);
nand U4166 (N_4166,N_3894,N_3731);
nor U4167 (N_4167,N_3899,N_3636);
or U4168 (N_4168,N_3610,N_3986);
nor U4169 (N_4169,N_3573,N_3705);
nor U4170 (N_4170,N_3621,N_3599);
nor U4171 (N_4171,N_3791,N_3934);
nor U4172 (N_4172,N_3685,N_3858);
nand U4173 (N_4173,N_3799,N_3815);
or U4174 (N_4174,N_3814,N_3945);
nand U4175 (N_4175,N_3546,N_3713);
and U4176 (N_4176,N_3868,N_3801);
nand U4177 (N_4177,N_3749,N_3717);
and U4178 (N_4178,N_3553,N_3630);
nor U4179 (N_4179,N_3549,N_3805);
nand U4180 (N_4180,N_3919,N_3527);
and U4181 (N_4181,N_3594,N_3909);
nor U4182 (N_4182,N_3569,N_3592);
and U4183 (N_4183,N_3893,N_3915);
and U4184 (N_4184,N_3839,N_3651);
nand U4185 (N_4185,N_3896,N_3831);
or U4186 (N_4186,N_3596,N_3930);
nor U4187 (N_4187,N_3840,N_3581);
or U4188 (N_4188,N_3582,N_3857);
and U4189 (N_4189,N_3944,N_3540);
and U4190 (N_4190,N_3971,N_3803);
or U4191 (N_4191,N_3772,N_3524);
or U4192 (N_4192,N_3907,N_3657);
nand U4193 (N_4193,N_3816,N_3675);
or U4194 (N_4194,N_3739,N_3988);
nor U4195 (N_4195,N_3851,N_3965);
or U4196 (N_4196,N_3855,N_3984);
and U4197 (N_4197,N_3619,N_3575);
or U4198 (N_4198,N_3732,N_3736);
xnor U4199 (N_4199,N_3922,N_3605);
and U4200 (N_4200,N_3842,N_3701);
and U4201 (N_4201,N_3903,N_3616);
and U4202 (N_4202,N_3785,N_3529);
nor U4203 (N_4203,N_3650,N_3809);
and U4204 (N_4204,N_3620,N_3514);
nor U4205 (N_4205,N_3904,N_3559);
xnor U4206 (N_4206,N_3643,N_3770);
and U4207 (N_4207,N_3760,N_3767);
and U4208 (N_4208,N_3585,N_3738);
or U4209 (N_4209,N_3755,N_3960);
or U4210 (N_4210,N_3923,N_3554);
nor U4211 (N_4211,N_3834,N_3928);
nand U4212 (N_4212,N_3602,N_3712);
nor U4213 (N_4213,N_3565,N_3729);
nand U4214 (N_4214,N_3673,N_3661);
nand U4215 (N_4215,N_3509,N_3794);
or U4216 (N_4216,N_3874,N_3560);
and U4217 (N_4217,N_3768,N_3727);
nand U4218 (N_4218,N_3800,N_3595);
nor U4219 (N_4219,N_3783,N_3707);
nand U4220 (N_4220,N_3613,N_3771);
and U4221 (N_4221,N_3598,N_3742);
nor U4222 (N_4222,N_3792,N_3997);
nor U4223 (N_4223,N_3671,N_3646);
or U4224 (N_4224,N_3913,N_3950);
or U4225 (N_4225,N_3682,N_3980);
xor U4226 (N_4226,N_3756,N_3968);
and U4227 (N_4227,N_3503,N_3847);
nand U4228 (N_4228,N_3662,N_3818);
nor U4229 (N_4229,N_3830,N_3722);
xor U4230 (N_4230,N_3686,N_3715);
xnor U4231 (N_4231,N_3666,N_3532);
and U4232 (N_4232,N_3766,N_3577);
nand U4233 (N_4233,N_3579,N_3516);
or U4234 (N_4234,N_3773,N_3832);
or U4235 (N_4235,N_3910,N_3719);
xnor U4236 (N_4236,N_3500,N_3798);
nor U4237 (N_4237,N_3901,N_3600);
or U4238 (N_4238,N_3861,N_3987);
xnor U4239 (N_4239,N_3716,N_3900);
and U4240 (N_4240,N_3890,N_3687);
and U4241 (N_4241,N_3761,N_3550);
nor U4242 (N_4242,N_3970,N_3882);
nor U4243 (N_4243,N_3669,N_3584);
nor U4244 (N_4244,N_3637,N_3943);
and U4245 (N_4245,N_3744,N_3710);
or U4246 (N_4246,N_3819,N_3511);
xor U4247 (N_4247,N_3674,N_3802);
nor U4248 (N_4248,N_3946,N_3841);
nor U4249 (N_4249,N_3720,N_3978);
nor U4250 (N_4250,N_3899,N_3504);
or U4251 (N_4251,N_3897,N_3597);
nor U4252 (N_4252,N_3705,N_3525);
nor U4253 (N_4253,N_3760,N_3722);
and U4254 (N_4254,N_3599,N_3689);
or U4255 (N_4255,N_3856,N_3861);
nor U4256 (N_4256,N_3758,N_3573);
nand U4257 (N_4257,N_3546,N_3673);
or U4258 (N_4258,N_3575,N_3887);
nand U4259 (N_4259,N_3939,N_3945);
nand U4260 (N_4260,N_3746,N_3977);
or U4261 (N_4261,N_3685,N_3941);
and U4262 (N_4262,N_3893,N_3548);
nor U4263 (N_4263,N_3959,N_3778);
nand U4264 (N_4264,N_3841,N_3513);
or U4265 (N_4265,N_3618,N_3892);
or U4266 (N_4266,N_3937,N_3582);
nor U4267 (N_4267,N_3827,N_3623);
nor U4268 (N_4268,N_3920,N_3513);
nor U4269 (N_4269,N_3649,N_3908);
nand U4270 (N_4270,N_3990,N_3903);
nand U4271 (N_4271,N_3710,N_3750);
nand U4272 (N_4272,N_3694,N_3842);
or U4273 (N_4273,N_3936,N_3603);
nand U4274 (N_4274,N_3587,N_3764);
nor U4275 (N_4275,N_3783,N_3929);
or U4276 (N_4276,N_3622,N_3781);
or U4277 (N_4277,N_3522,N_3925);
and U4278 (N_4278,N_3941,N_3680);
or U4279 (N_4279,N_3783,N_3830);
nand U4280 (N_4280,N_3600,N_3991);
and U4281 (N_4281,N_3895,N_3888);
nor U4282 (N_4282,N_3869,N_3858);
or U4283 (N_4283,N_3581,N_3703);
nor U4284 (N_4284,N_3644,N_3973);
xor U4285 (N_4285,N_3953,N_3842);
or U4286 (N_4286,N_3961,N_3542);
or U4287 (N_4287,N_3685,N_3629);
or U4288 (N_4288,N_3725,N_3645);
and U4289 (N_4289,N_3524,N_3508);
nor U4290 (N_4290,N_3521,N_3677);
and U4291 (N_4291,N_3932,N_3722);
or U4292 (N_4292,N_3973,N_3811);
or U4293 (N_4293,N_3900,N_3665);
or U4294 (N_4294,N_3567,N_3858);
or U4295 (N_4295,N_3728,N_3845);
and U4296 (N_4296,N_3830,N_3533);
and U4297 (N_4297,N_3570,N_3627);
nor U4298 (N_4298,N_3678,N_3998);
or U4299 (N_4299,N_3954,N_3993);
nor U4300 (N_4300,N_3768,N_3772);
nor U4301 (N_4301,N_3740,N_3629);
and U4302 (N_4302,N_3513,N_3991);
or U4303 (N_4303,N_3803,N_3718);
nand U4304 (N_4304,N_3520,N_3783);
or U4305 (N_4305,N_3615,N_3505);
and U4306 (N_4306,N_3694,N_3548);
xor U4307 (N_4307,N_3707,N_3763);
and U4308 (N_4308,N_3713,N_3738);
and U4309 (N_4309,N_3631,N_3858);
xnor U4310 (N_4310,N_3952,N_3584);
nor U4311 (N_4311,N_3542,N_3804);
nand U4312 (N_4312,N_3734,N_3938);
nand U4313 (N_4313,N_3925,N_3634);
or U4314 (N_4314,N_3760,N_3662);
nor U4315 (N_4315,N_3786,N_3975);
nand U4316 (N_4316,N_3991,N_3910);
and U4317 (N_4317,N_3670,N_3768);
and U4318 (N_4318,N_3835,N_3565);
nor U4319 (N_4319,N_3918,N_3854);
nand U4320 (N_4320,N_3798,N_3556);
or U4321 (N_4321,N_3684,N_3656);
nand U4322 (N_4322,N_3873,N_3817);
and U4323 (N_4323,N_3725,N_3861);
or U4324 (N_4324,N_3547,N_3649);
or U4325 (N_4325,N_3673,N_3875);
nand U4326 (N_4326,N_3957,N_3798);
or U4327 (N_4327,N_3514,N_3573);
and U4328 (N_4328,N_3524,N_3948);
and U4329 (N_4329,N_3583,N_3800);
or U4330 (N_4330,N_3947,N_3624);
nand U4331 (N_4331,N_3726,N_3624);
nor U4332 (N_4332,N_3850,N_3941);
and U4333 (N_4333,N_3735,N_3678);
or U4334 (N_4334,N_3938,N_3922);
nand U4335 (N_4335,N_3520,N_3508);
nand U4336 (N_4336,N_3677,N_3681);
or U4337 (N_4337,N_3569,N_3500);
nor U4338 (N_4338,N_3547,N_3698);
or U4339 (N_4339,N_3567,N_3561);
or U4340 (N_4340,N_3761,N_3760);
nor U4341 (N_4341,N_3754,N_3905);
nand U4342 (N_4342,N_3895,N_3862);
and U4343 (N_4343,N_3753,N_3594);
or U4344 (N_4344,N_3834,N_3902);
nor U4345 (N_4345,N_3862,N_3693);
or U4346 (N_4346,N_3719,N_3988);
xor U4347 (N_4347,N_3670,N_3901);
or U4348 (N_4348,N_3718,N_3935);
nor U4349 (N_4349,N_3743,N_3906);
nand U4350 (N_4350,N_3552,N_3879);
xnor U4351 (N_4351,N_3868,N_3923);
nand U4352 (N_4352,N_3627,N_3544);
nand U4353 (N_4353,N_3502,N_3903);
nor U4354 (N_4354,N_3609,N_3819);
nor U4355 (N_4355,N_3716,N_3966);
or U4356 (N_4356,N_3842,N_3890);
nand U4357 (N_4357,N_3779,N_3517);
or U4358 (N_4358,N_3769,N_3822);
nor U4359 (N_4359,N_3735,N_3734);
and U4360 (N_4360,N_3936,N_3861);
and U4361 (N_4361,N_3752,N_3674);
nor U4362 (N_4362,N_3637,N_3642);
and U4363 (N_4363,N_3633,N_3500);
or U4364 (N_4364,N_3681,N_3924);
and U4365 (N_4365,N_3748,N_3671);
and U4366 (N_4366,N_3858,N_3627);
nor U4367 (N_4367,N_3939,N_3796);
nor U4368 (N_4368,N_3991,N_3581);
nor U4369 (N_4369,N_3555,N_3769);
and U4370 (N_4370,N_3834,N_3824);
and U4371 (N_4371,N_3886,N_3699);
nor U4372 (N_4372,N_3834,N_3712);
and U4373 (N_4373,N_3670,N_3667);
xor U4374 (N_4374,N_3659,N_3706);
or U4375 (N_4375,N_3642,N_3813);
or U4376 (N_4376,N_3629,N_3671);
and U4377 (N_4377,N_3854,N_3942);
and U4378 (N_4378,N_3819,N_3818);
nand U4379 (N_4379,N_3596,N_3876);
or U4380 (N_4380,N_3615,N_3508);
nor U4381 (N_4381,N_3715,N_3756);
nor U4382 (N_4382,N_3765,N_3556);
nand U4383 (N_4383,N_3823,N_3911);
and U4384 (N_4384,N_3557,N_3941);
nand U4385 (N_4385,N_3617,N_3767);
nor U4386 (N_4386,N_3980,N_3788);
nor U4387 (N_4387,N_3859,N_3670);
nand U4388 (N_4388,N_3846,N_3832);
and U4389 (N_4389,N_3742,N_3596);
and U4390 (N_4390,N_3936,N_3941);
nor U4391 (N_4391,N_3959,N_3814);
or U4392 (N_4392,N_3749,N_3524);
and U4393 (N_4393,N_3715,N_3529);
nand U4394 (N_4394,N_3682,N_3777);
and U4395 (N_4395,N_3615,N_3522);
nand U4396 (N_4396,N_3951,N_3956);
nor U4397 (N_4397,N_3518,N_3589);
nand U4398 (N_4398,N_3567,N_3939);
nor U4399 (N_4399,N_3574,N_3726);
or U4400 (N_4400,N_3734,N_3691);
nor U4401 (N_4401,N_3744,N_3866);
nor U4402 (N_4402,N_3508,N_3791);
nor U4403 (N_4403,N_3582,N_3672);
and U4404 (N_4404,N_3861,N_3827);
nand U4405 (N_4405,N_3698,N_3865);
and U4406 (N_4406,N_3695,N_3854);
and U4407 (N_4407,N_3689,N_3598);
and U4408 (N_4408,N_3546,N_3594);
nand U4409 (N_4409,N_3883,N_3761);
nor U4410 (N_4410,N_3970,N_3511);
or U4411 (N_4411,N_3947,N_3983);
or U4412 (N_4412,N_3895,N_3751);
nand U4413 (N_4413,N_3869,N_3616);
nor U4414 (N_4414,N_3845,N_3757);
nor U4415 (N_4415,N_3916,N_3799);
nand U4416 (N_4416,N_3902,N_3890);
and U4417 (N_4417,N_3742,N_3993);
or U4418 (N_4418,N_3638,N_3922);
xor U4419 (N_4419,N_3680,N_3789);
nand U4420 (N_4420,N_3622,N_3924);
nor U4421 (N_4421,N_3833,N_3973);
or U4422 (N_4422,N_3678,N_3702);
or U4423 (N_4423,N_3641,N_3743);
and U4424 (N_4424,N_3939,N_3769);
xnor U4425 (N_4425,N_3700,N_3868);
nand U4426 (N_4426,N_3592,N_3720);
and U4427 (N_4427,N_3875,N_3548);
and U4428 (N_4428,N_3700,N_3978);
nor U4429 (N_4429,N_3611,N_3966);
or U4430 (N_4430,N_3876,N_3749);
or U4431 (N_4431,N_3551,N_3757);
or U4432 (N_4432,N_3932,N_3924);
and U4433 (N_4433,N_3790,N_3694);
and U4434 (N_4434,N_3913,N_3776);
nor U4435 (N_4435,N_3652,N_3657);
and U4436 (N_4436,N_3760,N_3811);
nand U4437 (N_4437,N_3805,N_3923);
and U4438 (N_4438,N_3965,N_3664);
xor U4439 (N_4439,N_3815,N_3990);
and U4440 (N_4440,N_3513,N_3799);
nor U4441 (N_4441,N_3850,N_3676);
and U4442 (N_4442,N_3592,N_3958);
nand U4443 (N_4443,N_3832,N_3523);
and U4444 (N_4444,N_3986,N_3635);
nand U4445 (N_4445,N_3927,N_3554);
nand U4446 (N_4446,N_3819,N_3781);
and U4447 (N_4447,N_3651,N_3780);
nor U4448 (N_4448,N_3727,N_3951);
nand U4449 (N_4449,N_3932,N_3815);
nor U4450 (N_4450,N_3565,N_3511);
nor U4451 (N_4451,N_3734,N_3627);
and U4452 (N_4452,N_3814,N_3912);
nor U4453 (N_4453,N_3503,N_3926);
or U4454 (N_4454,N_3837,N_3904);
nand U4455 (N_4455,N_3749,N_3935);
or U4456 (N_4456,N_3769,N_3854);
nand U4457 (N_4457,N_3782,N_3788);
nor U4458 (N_4458,N_3553,N_3718);
xor U4459 (N_4459,N_3602,N_3845);
nor U4460 (N_4460,N_3980,N_3802);
nor U4461 (N_4461,N_3806,N_3825);
and U4462 (N_4462,N_3800,N_3810);
nor U4463 (N_4463,N_3564,N_3797);
nor U4464 (N_4464,N_3796,N_3789);
nor U4465 (N_4465,N_3633,N_3814);
nand U4466 (N_4466,N_3812,N_3833);
nand U4467 (N_4467,N_3694,N_3922);
nor U4468 (N_4468,N_3853,N_3504);
nor U4469 (N_4469,N_3572,N_3953);
and U4470 (N_4470,N_3641,N_3911);
or U4471 (N_4471,N_3515,N_3743);
and U4472 (N_4472,N_3729,N_3790);
or U4473 (N_4473,N_3861,N_3687);
nand U4474 (N_4474,N_3517,N_3775);
or U4475 (N_4475,N_3940,N_3710);
or U4476 (N_4476,N_3958,N_3874);
and U4477 (N_4477,N_3701,N_3923);
or U4478 (N_4478,N_3767,N_3932);
nand U4479 (N_4479,N_3884,N_3863);
or U4480 (N_4480,N_3885,N_3995);
nand U4481 (N_4481,N_3729,N_3561);
xor U4482 (N_4482,N_3773,N_3654);
nor U4483 (N_4483,N_3769,N_3568);
nand U4484 (N_4484,N_3794,N_3862);
or U4485 (N_4485,N_3947,N_3672);
xnor U4486 (N_4486,N_3979,N_3840);
nand U4487 (N_4487,N_3634,N_3887);
nand U4488 (N_4488,N_3715,N_3538);
or U4489 (N_4489,N_3793,N_3803);
xor U4490 (N_4490,N_3524,N_3845);
nor U4491 (N_4491,N_3641,N_3725);
nor U4492 (N_4492,N_3847,N_3690);
or U4493 (N_4493,N_3935,N_3926);
nand U4494 (N_4494,N_3830,N_3865);
and U4495 (N_4495,N_3957,N_3607);
and U4496 (N_4496,N_3930,N_3891);
or U4497 (N_4497,N_3839,N_3960);
nor U4498 (N_4498,N_3837,N_3814);
or U4499 (N_4499,N_3528,N_3689);
nand U4500 (N_4500,N_4112,N_4397);
nor U4501 (N_4501,N_4214,N_4352);
and U4502 (N_4502,N_4251,N_4118);
nor U4503 (N_4503,N_4243,N_4186);
nor U4504 (N_4504,N_4474,N_4094);
nand U4505 (N_4505,N_4234,N_4269);
and U4506 (N_4506,N_4233,N_4260);
nor U4507 (N_4507,N_4490,N_4329);
or U4508 (N_4508,N_4056,N_4211);
or U4509 (N_4509,N_4014,N_4267);
nor U4510 (N_4510,N_4389,N_4064);
nand U4511 (N_4511,N_4113,N_4404);
and U4512 (N_4512,N_4188,N_4255);
nor U4513 (N_4513,N_4001,N_4364);
xor U4514 (N_4514,N_4458,N_4008);
nor U4515 (N_4515,N_4197,N_4198);
nand U4516 (N_4516,N_4299,N_4320);
or U4517 (N_4517,N_4482,N_4080);
xor U4518 (N_4518,N_4022,N_4163);
or U4519 (N_4519,N_4092,N_4436);
nor U4520 (N_4520,N_4026,N_4229);
and U4521 (N_4521,N_4132,N_4328);
or U4522 (N_4522,N_4074,N_4219);
or U4523 (N_4523,N_4170,N_4433);
nor U4524 (N_4524,N_4345,N_4461);
nand U4525 (N_4525,N_4342,N_4242);
xor U4526 (N_4526,N_4307,N_4346);
and U4527 (N_4527,N_4387,N_4304);
or U4528 (N_4528,N_4138,N_4354);
and U4529 (N_4529,N_4039,N_4456);
nand U4530 (N_4530,N_4446,N_4077);
and U4531 (N_4531,N_4360,N_4273);
and U4532 (N_4532,N_4046,N_4429);
nand U4533 (N_4533,N_4495,N_4489);
nand U4534 (N_4534,N_4462,N_4470);
or U4535 (N_4535,N_4391,N_4376);
nor U4536 (N_4536,N_4449,N_4065);
nand U4537 (N_4537,N_4373,N_4067);
nand U4538 (N_4538,N_4144,N_4348);
or U4539 (N_4539,N_4448,N_4246);
and U4540 (N_4540,N_4393,N_4398);
nand U4541 (N_4541,N_4016,N_4024);
nor U4542 (N_4542,N_4408,N_4488);
or U4543 (N_4543,N_4159,N_4322);
and U4544 (N_4544,N_4083,N_4230);
and U4545 (N_4545,N_4102,N_4225);
or U4546 (N_4546,N_4106,N_4343);
or U4547 (N_4547,N_4468,N_4479);
and U4548 (N_4548,N_4464,N_4097);
and U4549 (N_4549,N_4084,N_4006);
and U4550 (N_4550,N_4244,N_4275);
or U4551 (N_4551,N_4060,N_4162);
or U4552 (N_4552,N_4160,N_4321);
and U4553 (N_4553,N_4435,N_4002);
and U4554 (N_4554,N_4124,N_4156);
and U4555 (N_4555,N_4086,N_4413);
or U4556 (N_4556,N_4210,N_4369);
or U4557 (N_4557,N_4258,N_4075);
and U4558 (N_4558,N_4099,N_4272);
or U4559 (N_4559,N_4045,N_4055);
nor U4560 (N_4560,N_4428,N_4326);
and U4561 (N_4561,N_4204,N_4426);
or U4562 (N_4562,N_4484,N_4451);
and U4563 (N_4563,N_4418,N_4073);
nand U4564 (N_4564,N_4194,N_4311);
nor U4565 (N_4565,N_4287,N_4151);
and U4566 (N_4566,N_4276,N_4334);
nor U4567 (N_4567,N_4057,N_4146);
and U4568 (N_4568,N_4031,N_4410);
nor U4569 (N_4569,N_4147,N_4333);
or U4570 (N_4570,N_4425,N_4177);
nor U4571 (N_4571,N_4175,N_4079);
nand U4572 (N_4572,N_4472,N_4208);
or U4573 (N_4573,N_4293,N_4407);
nor U4574 (N_4574,N_4424,N_4401);
nor U4575 (N_4575,N_4153,N_4103);
nor U4576 (N_4576,N_4028,N_4315);
or U4577 (N_4577,N_4362,N_4378);
and U4578 (N_4578,N_4200,N_4306);
nand U4579 (N_4579,N_4344,N_4161);
nor U4580 (N_4580,N_4480,N_4098);
and U4581 (N_4581,N_4353,N_4372);
nand U4582 (N_4582,N_4236,N_4125);
nor U4583 (N_4583,N_4325,N_4286);
nor U4584 (N_4584,N_4298,N_4432);
nand U4585 (N_4585,N_4120,N_4017);
nand U4586 (N_4586,N_4394,N_4431);
nor U4587 (N_4587,N_4224,N_4202);
or U4588 (N_4588,N_4252,N_4005);
and U4589 (N_4589,N_4173,N_4009);
and U4590 (N_4590,N_4134,N_4121);
or U4591 (N_4591,N_4004,N_4365);
nor U4592 (N_4592,N_4414,N_4136);
nand U4593 (N_4593,N_4148,N_4453);
and U4594 (N_4594,N_4182,N_4058);
or U4595 (N_4595,N_4294,N_4314);
and U4596 (N_4596,N_4018,N_4303);
nor U4597 (N_4597,N_4347,N_4476);
and U4598 (N_4598,N_4382,N_4473);
nand U4599 (N_4599,N_4048,N_4011);
nor U4600 (N_4600,N_4164,N_4167);
and U4601 (N_4601,N_4296,N_4379);
nor U4602 (N_4602,N_4249,N_4049);
and U4603 (N_4603,N_4361,N_4095);
or U4604 (N_4604,N_4062,N_4265);
nor U4605 (N_4605,N_4399,N_4412);
nand U4606 (N_4606,N_4196,N_4078);
and U4607 (N_4607,N_4235,N_4047);
xor U4608 (N_4608,N_4215,N_4076);
and U4609 (N_4609,N_4459,N_4417);
nor U4610 (N_4610,N_4166,N_4123);
nand U4611 (N_4611,N_4290,N_4192);
and U4612 (N_4612,N_4477,N_4288);
or U4613 (N_4613,N_4411,N_4297);
or U4614 (N_4614,N_4218,N_4025);
or U4615 (N_4615,N_4419,N_4171);
or U4616 (N_4616,N_4030,N_4356);
nor U4617 (N_4617,N_4020,N_4444);
and U4618 (N_4618,N_4469,N_4289);
and U4619 (N_4619,N_4331,N_4040);
nand U4620 (N_4620,N_4115,N_4088);
nor U4621 (N_4621,N_4270,N_4220);
or U4622 (N_4622,N_4285,N_4155);
or U4623 (N_4623,N_4059,N_4437);
or U4624 (N_4624,N_4157,N_4341);
and U4625 (N_4625,N_4250,N_4139);
and U4626 (N_4626,N_4466,N_4172);
nand U4627 (N_4627,N_4281,N_4434);
xor U4628 (N_4628,N_4351,N_4261);
nand U4629 (N_4629,N_4305,N_4090);
nand U4630 (N_4630,N_4183,N_4319);
or U4631 (N_4631,N_4338,N_4487);
and U4632 (N_4632,N_4277,N_4452);
nor U4633 (N_4633,N_4033,N_4491);
nand U4634 (N_4634,N_4247,N_4485);
nor U4635 (N_4635,N_4295,N_4191);
nand U4636 (N_4636,N_4359,N_4205);
and U4637 (N_4637,N_4135,N_4300);
and U4638 (N_4638,N_4145,N_4071);
and U4639 (N_4639,N_4122,N_4119);
or U4640 (N_4640,N_4262,N_4388);
nand U4641 (N_4641,N_4093,N_4370);
or U4642 (N_4642,N_4465,N_4037);
and U4643 (N_4643,N_4108,N_4054);
or U4644 (N_4644,N_4126,N_4237);
nor U4645 (N_4645,N_4209,N_4357);
and U4646 (N_4646,N_4110,N_4238);
nor U4647 (N_4647,N_4072,N_4253);
or U4648 (N_4648,N_4085,N_4044);
or U4649 (N_4649,N_4374,N_4130);
nand U4650 (N_4650,N_4133,N_4422);
nand U4651 (N_4651,N_4069,N_4068);
or U4652 (N_4652,N_4248,N_4317);
nor U4653 (N_4653,N_4061,N_4038);
and U4654 (N_4654,N_4027,N_4180);
nor U4655 (N_4655,N_4212,N_4206);
nor U4656 (N_4656,N_4087,N_4385);
nand U4657 (N_4657,N_4179,N_4492);
nand U4658 (N_4658,N_4423,N_4032);
nor U4659 (N_4659,N_4012,N_4131);
or U4660 (N_4660,N_4070,N_4152);
nor U4661 (N_4661,N_4313,N_4137);
or U4662 (N_4662,N_4416,N_4015);
or U4663 (N_4663,N_4050,N_4336);
or U4664 (N_4664,N_4427,N_4041);
nand U4665 (N_4665,N_4447,N_4463);
and U4666 (N_4666,N_4481,N_4400);
nand U4667 (N_4667,N_4190,N_4471);
or U4668 (N_4668,N_4154,N_4284);
nor U4669 (N_4669,N_4363,N_4189);
nand U4670 (N_4670,N_4327,N_4278);
nor U4671 (N_4671,N_4380,N_4104);
nor U4672 (N_4672,N_4127,N_4128);
nand U4673 (N_4673,N_4034,N_4499);
and U4674 (N_4674,N_4310,N_4221);
nor U4675 (N_4675,N_4239,N_4129);
nor U4676 (N_4676,N_4203,N_4213);
nor U4677 (N_4677,N_4178,N_4283);
or U4678 (N_4678,N_4498,N_4402);
and U4679 (N_4679,N_4358,N_4441);
nand U4680 (N_4680,N_4486,N_4256);
or U4681 (N_4681,N_4332,N_4207);
and U4682 (N_4682,N_4114,N_4096);
or U4683 (N_4683,N_4409,N_4043);
or U4684 (N_4684,N_4386,N_4101);
nor U4685 (N_4685,N_4497,N_4063);
or U4686 (N_4686,N_4440,N_4292);
nand U4687 (N_4687,N_4176,N_4308);
nor U4688 (N_4688,N_4259,N_4116);
or U4689 (N_4689,N_4475,N_4454);
xnor U4690 (N_4690,N_4367,N_4366);
nor U4691 (N_4691,N_4187,N_4291);
and U4692 (N_4692,N_4216,N_4339);
nand U4693 (N_4693,N_4280,N_4268);
and U4694 (N_4694,N_4051,N_4340);
and U4695 (N_4695,N_4271,N_4420);
xor U4696 (N_4696,N_4003,N_4241);
or U4697 (N_4697,N_4141,N_4222);
or U4698 (N_4698,N_4117,N_4478);
xor U4699 (N_4699,N_4066,N_4226);
nor U4700 (N_4700,N_4375,N_4330);
and U4701 (N_4701,N_4042,N_4169);
nand U4702 (N_4702,N_4496,N_4406);
and U4703 (N_4703,N_4029,N_4082);
nor U4704 (N_4704,N_4228,N_4430);
nand U4705 (N_4705,N_4355,N_4323);
nor U4706 (N_4706,N_4377,N_4217);
or U4707 (N_4707,N_4309,N_4199);
nor U4708 (N_4708,N_4396,N_4264);
and U4709 (N_4709,N_4010,N_4109);
nor U4710 (N_4710,N_4282,N_4390);
nand U4711 (N_4711,N_4240,N_4231);
nor U4712 (N_4712,N_4195,N_4450);
nor U4713 (N_4713,N_4007,N_4439);
or U4714 (N_4714,N_4384,N_4421);
nor U4715 (N_4715,N_4140,N_4350);
or U4716 (N_4716,N_4081,N_4107);
nor U4717 (N_4717,N_4232,N_4493);
nand U4718 (N_4718,N_4381,N_4368);
nand U4719 (N_4719,N_4185,N_4279);
or U4720 (N_4720,N_4494,N_4223);
or U4721 (N_4721,N_4349,N_4111);
nand U4722 (N_4722,N_4091,N_4337);
nor U4723 (N_4723,N_4467,N_4302);
and U4724 (N_4724,N_4371,N_4405);
nand U4725 (N_4725,N_4000,N_4403);
nor U4726 (N_4726,N_4021,N_4257);
xnor U4727 (N_4727,N_4165,N_4392);
and U4728 (N_4728,N_4013,N_4395);
xnor U4729 (N_4729,N_4035,N_4274);
nor U4730 (N_4730,N_4442,N_4158);
xor U4731 (N_4731,N_4052,N_4245);
nor U4732 (N_4732,N_4142,N_4445);
or U4733 (N_4733,N_4149,N_4460);
and U4734 (N_4734,N_4483,N_4019);
or U4735 (N_4735,N_4100,N_4105);
and U4736 (N_4736,N_4023,N_4181);
or U4737 (N_4737,N_4318,N_4036);
nand U4738 (N_4738,N_4053,N_4383);
nor U4739 (N_4739,N_4312,N_4415);
nand U4740 (N_4740,N_4457,N_4168);
or U4741 (N_4741,N_4201,N_4438);
and U4742 (N_4742,N_4193,N_4316);
or U4743 (N_4743,N_4263,N_4266);
and U4744 (N_4744,N_4455,N_4143);
or U4745 (N_4745,N_4254,N_4174);
or U4746 (N_4746,N_4184,N_4089);
nor U4747 (N_4747,N_4150,N_4227);
or U4748 (N_4748,N_4335,N_4443);
or U4749 (N_4749,N_4324,N_4301);
or U4750 (N_4750,N_4296,N_4300);
nand U4751 (N_4751,N_4498,N_4031);
and U4752 (N_4752,N_4386,N_4100);
and U4753 (N_4753,N_4295,N_4196);
nand U4754 (N_4754,N_4100,N_4396);
and U4755 (N_4755,N_4068,N_4315);
nand U4756 (N_4756,N_4108,N_4407);
or U4757 (N_4757,N_4408,N_4142);
nor U4758 (N_4758,N_4234,N_4317);
nor U4759 (N_4759,N_4159,N_4333);
nor U4760 (N_4760,N_4123,N_4300);
and U4761 (N_4761,N_4124,N_4489);
and U4762 (N_4762,N_4258,N_4122);
nor U4763 (N_4763,N_4024,N_4419);
and U4764 (N_4764,N_4153,N_4034);
nand U4765 (N_4765,N_4260,N_4372);
nand U4766 (N_4766,N_4011,N_4071);
nor U4767 (N_4767,N_4140,N_4383);
nand U4768 (N_4768,N_4072,N_4213);
nor U4769 (N_4769,N_4271,N_4233);
and U4770 (N_4770,N_4034,N_4027);
nand U4771 (N_4771,N_4486,N_4148);
and U4772 (N_4772,N_4057,N_4314);
and U4773 (N_4773,N_4157,N_4325);
or U4774 (N_4774,N_4179,N_4447);
nand U4775 (N_4775,N_4105,N_4047);
xnor U4776 (N_4776,N_4053,N_4338);
nor U4777 (N_4777,N_4073,N_4337);
or U4778 (N_4778,N_4127,N_4320);
or U4779 (N_4779,N_4332,N_4112);
nor U4780 (N_4780,N_4207,N_4022);
nor U4781 (N_4781,N_4085,N_4167);
and U4782 (N_4782,N_4093,N_4484);
nand U4783 (N_4783,N_4374,N_4274);
nand U4784 (N_4784,N_4130,N_4369);
and U4785 (N_4785,N_4122,N_4225);
or U4786 (N_4786,N_4329,N_4278);
nor U4787 (N_4787,N_4468,N_4097);
and U4788 (N_4788,N_4093,N_4224);
or U4789 (N_4789,N_4291,N_4091);
nand U4790 (N_4790,N_4112,N_4037);
or U4791 (N_4791,N_4395,N_4449);
or U4792 (N_4792,N_4030,N_4032);
and U4793 (N_4793,N_4385,N_4023);
nand U4794 (N_4794,N_4217,N_4313);
or U4795 (N_4795,N_4442,N_4203);
or U4796 (N_4796,N_4266,N_4075);
xnor U4797 (N_4797,N_4330,N_4258);
nor U4798 (N_4798,N_4142,N_4312);
and U4799 (N_4799,N_4334,N_4106);
nor U4800 (N_4800,N_4332,N_4131);
nor U4801 (N_4801,N_4278,N_4077);
nand U4802 (N_4802,N_4451,N_4234);
nand U4803 (N_4803,N_4270,N_4115);
or U4804 (N_4804,N_4225,N_4032);
nand U4805 (N_4805,N_4352,N_4187);
and U4806 (N_4806,N_4457,N_4157);
xor U4807 (N_4807,N_4159,N_4438);
nand U4808 (N_4808,N_4074,N_4411);
xnor U4809 (N_4809,N_4272,N_4055);
nor U4810 (N_4810,N_4438,N_4482);
and U4811 (N_4811,N_4077,N_4083);
nand U4812 (N_4812,N_4307,N_4409);
nand U4813 (N_4813,N_4013,N_4029);
nand U4814 (N_4814,N_4171,N_4013);
xnor U4815 (N_4815,N_4063,N_4438);
nand U4816 (N_4816,N_4327,N_4279);
nand U4817 (N_4817,N_4213,N_4184);
nor U4818 (N_4818,N_4221,N_4116);
and U4819 (N_4819,N_4383,N_4030);
or U4820 (N_4820,N_4055,N_4269);
nor U4821 (N_4821,N_4482,N_4327);
nor U4822 (N_4822,N_4453,N_4282);
and U4823 (N_4823,N_4311,N_4295);
or U4824 (N_4824,N_4261,N_4007);
or U4825 (N_4825,N_4223,N_4187);
nor U4826 (N_4826,N_4211,N_4304);
nand U4827 (N_4827,N_4421,N_4252);
nand U4828 (N_4828,N_4453,N_4227);
nand U4829 (N_4829,N_4357,N_4322);
and U4830 (N_4830,N_4191,N_4366);
xnor U4831 (N_4831,N_4218,N_4265);
and U4832 (N_4832,N_4324,N_4407);
nor U4833 (N_4833,N_4273,N_4153);
or U4834 (N_4834,N_4316,N_4417);
or U4835 (N_4835,N_4093,N_4241);
xnor U4836 (N_4836,N_4409,N_4302);
or U4837 (N_4837,N_4329,N_4311);
and U4838 (N_4838,N_4281,N_4091);
nand U4839 (N_4839,N_4445,N_4032);
nor U4840 (N_4840,N_4343,N_4125);
nand U4841 (N_4841,N_4340,N_4117);
and U4842 (N_4842,N_4039,N_4455);
nand U4843 (N_4843,N_4401,N_4358);
and U4844 (N_4844,N_4215,N_4027);
nand U4845 (N_4845,N_4426,N_4241);
xnor U4846 (N_4846,N_4045,N_4497);
or U4847 (N_4847,N_4062,N_4150);
or U4848 (N_4848,N_4455,N_4033);
or U4849 (N_4849,N_4200,N_4179);
or U4850 (N_4850,N_4218,N_4488);
or U4851 (N_4851,N_4458,N_4211);
and U4852 (N_4852,N_4031,N_4123);
nand U4853 (N_4853,N_4230,N_4354);
nand U4854 (N_4854,N_4146,N_4242);
nand U4855 (N_4855,N_4278,N_4206);
nand U4856 (N_4856,N_4447,N_4481);
or U4857 (N_4857,N_4315,N_4312);
nand U4858 (N_4858,N_4118,N_4400);
and U4859 (N_4859,N_4014,N_4005);
or U4860 (N_4860,N_4383,N_4403);
or U4861 (N_4861,N_4056,N_4054);
and U4862 (N_4862,N_4178,N_4045);
nor U4863 (N_4863,N_4059,N_4094);
or U4864 (N_4864,N_4355,N_4076);
nand U4865 (N_4865,N_4272,N_4370);
nor U4866 (N_4866,N_4059,N_4354);
or U4867 (N_4867,N_4045,N_4138);
nor U4868 (N_4868,N_4074,N_4379);
nand U4869 (N_4869,N_4370,N_4433);
nand U4870 (N_4870,N_4332,N_4359);
nand U4871 (N_4871,N_4149,N_4169);
and U4872 (N_4872,N_4126,N_4415);
nor U4873 (N_4873,N_4012,N_4219);
nor U4874 (N_4874,N_4118,N_4056);
and U4875 (N_4875,N_4331,N_4363);
nor U4876 (N_4876,N_4332,N_4209);
nand U4877 (N_4877,N_4291,N_4081);
xnor U4878 (N_4878,N_4334,N_4310);
or U4879 (N_4879,N_4183,N_4479);
and U4880 (N_4880,N_4407,N_4386);
and U4881 (N_4881,N_4169,N_4232);
or U4882 (N_4882,N_4318,N_4371);
or U4883 (N_4883,N_4002,N_4391);
and U4884 (N_4884,N_4089,N_4432);
and U4885 (N_4885,N_4414,N_4282);
nor U4886 (N_4886,N_4435,N_4341);
and U4887 (N_4887,N_4135,N_4340);
nand U4888 (N_4888,N_4362,N_4297);
and U4889 (N_4889,N_4180,N_4078);
nand U4890 (N_4890,N_4345,N_4265);
or U4891 (N_4891,N_4282,N_4002);
and U4892 (N_4892,N_4401,N_4416);
nor U4893 (N_4893,N_4198,N_4370);
and U4894 (N_4894,N_4307,N_4490);
and U4895 (N_4895,N_4299,N_4126);
xor U4896 (N_4896,N_4337,N_4346);
nor U4897 (N_4897,N_4436,N_4358);
or U4898 (N_4898,N_4343,N_4394);
nand U4899 (N_4899,N_4288,N_4014);
and U4900 (N_4900,N_4472,N_4372);
or U4901 (N_4901,N_4166,N_4017);
or U4902 (N_4902,N_4129,N_4179);
or U4903 (N_4903,N_4353,N_4135);
nand U4904 (N_4904,N_4413,N_4390);
or U4905 (N_4905,N_4407,N_4364);
nand U4906 (N_4906,N_4048,N_4308);
nand U4907 (N_4907,N_4236,N_4323);
nand U4908 (N_4908,N_4452,N_4269);
nand U4909 (N_4909,N_4463,N_4125);
nor U4910 (N_4910,N_4208,N_4464);
and U4911 (N_4911,N_4018,N_4247);
or U4912 (N_4912,N_4365,N_4124);
xnor U4913 (N_4913,N_4264,N_4342);
nor U4914 (N_4914,N_4220,N_4348);
xnor U4915 (N_4915,N_4406,N_4322);
or U4916 (N_4916,N_4072,N_4257);
or U4917 (N_4917,N_4459,N_4317);
or U4918 (N_4918,N_4095,N_4245);
nor U4919 (N_4919,N_4101,N_4322);
nor U4920 (N_4920,N_4463,N_4068);
or U4921 (N_4921,N_4379,N_4217);
xor U4922 (N_4922,N_4242,N_4400);
or U4923 (N_4923,N_4391,N_4040);
or U4924 (N_4924,N_4175,N_4296);
and U4925 (N_4925,N_4473,N_4005);
and U4926 (N_4926,N_4357,N_4025);
xnor U4927 (N_4927,N_4261,N_4124);
or U4928 (N_4928,N_4198,N_4426);
nor U4929 (N_4929,N_4295,N_4044);
or U4930 (N_4930,N_4450,N_4131);
or U4931 (N_4931,N_4177,N_4090);
nand U4932 (N_4932,N_4058,N_4049);
or U4933 (N_4933,N_4473,N_4404);
nor U4934 (N_4934,N_4239,N_4117);
nor U4935 (N_4935,N_4022,N_4210);
nor U4936 (N_4936,N_4051,N_4440);
and U4937 (N_4937,N_4215,N_4015);
nor U4938 (N_4938,N_4409,N_4353);
nor U4939 (N_4939,N_4151,N_4103);
nor U4940 (N_4940,N_4364,N_4285);
nor U4941 (N_4941,N_4063,N_4267);
and U4942 (N_4942,N_4160,N_4415);
nand U4943 (N_4943,N_4493,N_4076);
nor U4944 (N_4944,N_4021,N_4026);
nor U4945 (N_4945,N_4451,N_4471);
xnor U4946 (N_4946,N_4440,N_4306);
or U4947 (N_4947,N_4073,N_4336);
nor U4948 (N_4948,N_4381,N_4075);
or U4949 (N_4949,N_4155,N_4182);
and U4950 (N_4950,N_4048,N_4228);
xor U4951 (N_4951,N_4304,N_4422);
nor U4952 (N_4952,N_4247,N_4238);
nand U4953 (N_4953,N_4163,N_4092);
and U4954 (N_4954,N_4456,N_4484);
nor U4955 (N_4955,N_4289,N_4478);
xnor U4956 (N_4956,N_4293,N_4048);
nand U4957 (N_4957,N_4220,N_4166);
or U4958 (N_4958,N_4443,N_4499);
nor U4959 (N_4959,N_4471,N_4071);
nor U4960 (N_4960,N_4093,N_4138);
nor U4961 (N_4961,N_4047,N_4418);
nor U4962 (N_4962,N_4484,N_4049);
and U4963 (N_4963,N_4273,N_4457);
or U4964 (N_4964,N_4083,N_4480);
or U4965 (N_4965,N_4240,N_4402);
or U4966 (N_4966,N_4058,N_4045);
nand U4967 (N_4967,N_4351,N_4055);
nand U4968 (N_4968,N_4013,N_4027);
or U4969 (N_4969,N_4462,N_4023);
nor U4970 (N_4970,N_4312,N_4214);
and U4971 (N_4971,N_4397,N_4342);
nand U4972 (N_4972,N_4330,N_4435);
or U4973 (N_4973,N_4208,N_4294);
xor U4974 (N_4974,N_4248,N_4071);
or U4975 (N_4975,N_4003,N_4215);
nor U4976 (N_4976,N_4195,N_4306);
or U4977 (N_4977,N_4139,N_4361);
and U4978 (N_4978,N_4150,N_4416);
or U4979 (N_4979,N_4266,N_4397);
nor U4980 (N_4980,N_4120,N_4461);
nand U4981 (N_4981,N_4376,N_4025);
nor U4982 (N_4982,N_4082,N_4304);
nor U4983 (N_4983,N_4187,N_4067);
or U4984 (N_4984,N_4493,N_4444);
nor U4985 (N_4985,N_4392,N_4434);
nand U4986 (N_4986,N_4087,N_4282);
nand U4987 (N_4987,N_4423,N_4044);
nor U4988 (N_4988,N_4193,N_4100);
nand U4989 (N_4989,N_4112,N_4455);
and U4990 (N_4990,N_4499,N_4454);
and U4991 (N_4991,N_4014,N_4232);
or U4992 (N_4992,N_4186,N_4380);
nor U4993 (N_4993,N_4108,N_4470);
nor U4994 (N_4994,N_4240,N_4205);
nand U4995 (N_4995,N_4339,N_4094);
nor U4996 (N_4996,N_4010,N_4188);
and U4997 (N_4997,N_4261,N_4492);
xnor U4998 (N_4998,N_4386,N_4219);
xor U4999 (N_4999,N_4287,N_4159);
or UO_0 (O_0,N_4545,N_4948);
or UO_1 (O_1,N_4638,N_4747);
or UO_2 (O_2,N_4610,N_4565);
nand UO_3 (O_3,N_4943,N_4862);
or UO_4 (O_4,N_4578,N_4762);
nand UO_5 (O_5,N_4768,N_4991);
nand UO_6 (O_6,N_4647,N_4916);
xor UO_7 (O_7,N_4870,N_4789);
nor UO_8 (O_8,N_4844,N_4693);
or UO_9 (O_9,N_4871,N_4531);
nor UO_10 (O_10,N_4960,N_4535);
nor UO_11 (O_11,N_4533,N_4767);
xor UO_12 (O_12,N_4745,N_4669);
and UO_13 (O_13,N_4655,N_4616);
nand UO_14 (O_14,N_4567,N_4918);
nand UO_15 (O_15,N_4922,N_4750);
and UO_16 (O_16,N_4564,N_4725);
nand UO_17 (O_17,N_4778,N_4681);
or UO_18 (O_18,N_4780,N_4597);
nand UO_19 (O_19,N_4521,N_4878);
and UO_20 (O_20,N_4675,N_4574);
nor UO_21 (O_21,N_4884,N_4636);
or UO_22 (O_22,N_4794,N_4596);
nand UO_23 (O_23,N_4555,N_4631);
nand UO_24 (O_24,N_4841,N_4959);
nor UO_25 (O_25,N_4686,N_4880);
or UO_26 (O_26,N_4585,N_4912);
nand UO_27 (O_27,N_4623,N_4713);
or UO_28 (O_28,N_4997,N_4718);
nand UO_29 (O_29,N_4553,N_4698);
nand UO_30 (O_30,N_4532,N_4798);
nand UO_31 (O_31,N_4809,N_4732);
nand UO_32 (O_32,N_4832,N_4771);
nand UO_33 (O_33,N_4924,N_4885);
and UO_34 (O_34,N_4607,N_4865);
nand UO_35 (O_35,N_4996,N_4920);
and UO_36 (O_36,N_4867,N_4528);
nand UO_37 (O_37,N_4509,N_4682);
xor UO_38 (O_38,N_4606,N_4559);
and UO_39 (O_39,N_4632,N_4807);
nand UO_40 (O_40,N_4861,N_4538);
nand UO_41 (O_41,N_4856,N_4801);
nand UO_42 (O_42,N_4548,N_4744);
or UO_43 (O_43,N_4571,N_4942);
nor UO_44 (O_44,N_4608,N_4985);
or UO_45 (O_45,N_4770,N_4982);
nand UO_46 (O_46,N_4705,N_4691);
or UO_47 (O_47,N_4530,N_4733);
nand UO_48 (O_48,N_4579,N_4969);
nand UO_49 (O_49,N_4726,N_4722);
and UO_50 (O_50,N_4864,N_4989);
and UO_51 (O_51,N_4629,N_4816);
or UO_52 (O_52,N_4536,N_4843);
nand UO_53 (O_53,N_4605,N_4749);
or UO_54 (O_54,N_4627,N_4519);
nor UO_55 (O_55,N_4620,N_4526);
and UO_56 (O_56,N_4769,N_4668);
or UO_57 (O_57,N_4847,N_4926);
nand UO_58 (O_58,N_4562,N_4908);
nand UO_59 (O_59,N_4783,N_4764);
and UO_60 (O_60,N_4554,N_4803);
or UO_61 (O_61,N_4566,N_4848);
nor UO_62 (O_62,N_4966,N_4950);
nand UO_63 (O_63,N_4857,N_4793);
and UO_64 (O_64,N_4734,N_4973);
xnor UO_65 (O_65,N_4677,N_4586);
nand UO_66 (O_66,N_4729,N_4992);
nor UO_67 (O_67,N_4712,N_4952);
and UO_68 (O_68,N_4874,N_4637);
or UO_69 (O_69,N_4674,N_4859);
and UO_70 (O_70,N_4701,N_4609);
or UO_71 (O_71,N_4853,N_4970);
and UO_72 (O_72,N_4648,N_4613);
and UO_73 (O_73,N_4928,N_4588);
nor UO_74 (O_74,N_4662,N_4800);
or UO_75 (O_75,N_4557,N_4806);
or UO_76 (O_76,N_4510,N_4965);
and UO_77 (O_77,N_4976,N_4808);
xor UO_78 (O_78,N_4706,N_4537);
nor UO_79 (O_79,N_4502,N_4819);
or UO_80 (O_80,N_4940,N_4879);
xor UO_81 (O_81,N_4898,N_4963);
nand UO_82 (O_82,N_4738,N_4736);
nor UO_83 (O_83,N_4855,N_4890);
and UO_84 (O_84,N_4813,N_4891);
nor UO_85 (O_85,N_4915,N_4820);
nor UO_86 (O_86,N_4672,N_4782);
nand UO_87 (O_87,N_4641,N_4508);
or UO_88 (O_88,N_4727,N_4645);
or UO_89 (O_89,N_4600,N_4709);
nor UO_90 (O_90,N_4739,N_4561);
nor UO_91 (O_91,N_4748,N_4756);
nor UO_92 (O_92,N_4773,N_4866);
nand UO_93 (O_93,N_4906,N_4741);
nor UO_94 (O_94,N_4883,N_4877);
xnor UO_95 (O_95,N_4573,N_4830);
and UO_96 (O_96,N_4518,N_4889);
nor UO_97 (O_97,N_4743,N_4904);
xnor UO_98 (O_98,N_4619,N_4507);
nand UO_99 (O_99,N_4897,N_4882);
and UO_100 (O_100,N_4849,N_4525);
or UO_101 (O_101,N_4978,N_4503);
nand UO_102 (O_102,N_4961,N_4643);
or UO_103 (O_103,N_4946,N_4994);
nor UO_104 (O_104,N_4580,N_4583);
xor UO_105 (O_105,N_4760,N_4863);
nand UO_106 (O_106,N_4551,N_4735);
xnor UO_107 (O_107,N_4504,N_4506);
nand UO_108 (O_108,N_4602,N_4524);
nor UO_109 (O_109,N_4569,N_4979);
nor UO_110 (O_110,N_4575,N_4595);
nand UO_111 (O_111,N_4810,N_4667);
or UO_112 (O_112,N_4663,N_4740);
or UO_113 (O_113,N_4714,N_4746);
nand UO_114 (O_114,N_4707,N_4850);
and UO_115 (O_115,N_4917,N_4825);
or UO_116 (O_116,N_4921,N_4781);
xnor UO_117 (O_117,N_4945,N_4792);
or UO_118 (O_118,N_4671,N_4517);
nand UO_119 (O_119,N_4990,N_4776);
nand UO_120 (O_120,N_4910,N_4710);
or UO_121 (O_121,N_4765,N_4761);
or UO_122 (O_122,N_4639,N_4986);
nand UO_123 (O_123,N_4618,N_4685);
nor UO_124 (O_124,N_4872,N_4817);
and UO_125 (O_125,N_4887,N_4520);
xnor UO_126 (O_126,N_4993,N_4589);
nor UO_127 (O_127,N_4811,N_4822);
nand UO_128 (O_128,N_4649,N_4755);
or UO_129 (O_129,N_4752,N_4543);
and UO_130 (O_130,N_4913,N_4983);
nor UO_131 (O_131,N_4611,N_4688);
nand UO_132 (O_132,N_4689,N_4988);
and UO_133 (O_133,N_4951,N_4975);
or UO_134 (O_134,N_4544,N_4967);
or UO_135 (O_135,N_4786,N_4716);
nor UO_136 (O_136,N_4679,N_4823);
or UO_137 (O_137,N_4790,N_4614);
and UO_138 (O_138,N_4888,N_4552);
nor UO_139 (O_139,N_4927,N_4893);
nand UO_140 (O_140,N_4980,N_4836);
or UO_141 (O_141,N_4604,N_4628);
nand UO_142 (O_142,N_4923,N_4795);
or UO_143 (O_143,N_4742,N_4840);
nor UO_144 (O_144,N_4542,N_4995);
nand UO_145 (O_145,N_4895,N_4899);
or UO_146 (O_146,N_4834,N_4695);
or UO_147 (O_147,N_4657,N_4894);
xnor UO_148 (O_148,N_4515,N_4772);
or UO_149 (O_149,N_4653,N_4652);
nand UO_150 (O_150,N_4935,N_4534);
or UO_151 (O_151,N_4720,N_4560);
nor UO_152 (O_152,N_4594,N_4852);
and UO_153 (O_153,N_4584,N_4612);
nand UO_154 (O_154,N_4625,N_4939);
and UO_155 (O_155,N_4958,N_4858);
nand UO_156 (O_156,N_4696,N_4824);
nand UO_157 (O_157,N_4998,N_4955);
or UO_158 (O_158,N_4576,N_4914);
or UO_159 (O_159,N_4724,N_4837);
xor UO_160 (O_160,N_4666,N_4796);
or UO_161 (O_161,N_4896,N_4708);
and UO_162 (O_162,N_4876,N_4757);
nand UO_163 (O_163,N_4972,N_4717);
nand UO_164 (O_164,N_4953,N_4590);
or UO_165 (O_165,N_4687,N_4875);
and UO_166 (O_166,N_4670,N_4947);
and UO_167 (O_167,N_4974,N_4881);
and UO_168 (O_168,N_4673,N_4805);
nand UO_169 (O_169,N_4591,N_4501);
or UO_170 (O_170,N_4635,N_4617);
and UO_171 (O_171,N_4941,N_4868);
nand UO_172 (O_172,N_4886,N_4572);
nand UO_173 (O_173,N_4582,N_4541);
nor UO_174 (O_174,N_4802,N_4621);
nor UO_175 (O_175,N_4640,N_4799);
nand UO_176 (O_176,N_4911,N_4821);
or UO_177 (O_177,N_4642,N_4683);
and UO_178 (O_178,N_4690,N_4547);
nand UO_179 (O_179,N_4784,N_4930);
nand UO_180 (O_180,N_4815,N_4633);
xnor UO_181 (O_181,N_4842,N_4660);
and UO_182 (O_182,N_4615,N_4558);
and UO_183 (O_183,N_4925,N_4936);
and UO_184 (O_184,N_4758,N_4829);
nand UO_185 (O_185,N_4984,N_4546);
or UO_186 (O_186,N_4909,N_4719);
or UO_187 (O_187,N_4754,N_4753);
nand UO_188 (O_188,N_4661,N_4599);
nand UO_189 (O_189,N_4905,N_4540);
nor UO_190 (O_190,N_4937,N_4563);
xnor UO_191 (O_191,N_4634,N_4791);
or UO_192 (O_192,N_4839,N_4646);
or UO_193 (O_193,N_4964,N_4723);
and UO_194 (O_194,N_4827,N_4826);
nand UO_195 (O_195,N_4812,N_4680);
xnor UO_196 (O_196,N_4804,N_4968);
or UO_197 (O_197,N_4644,N_4846);
or UO_198 (O_198,N_4651,N_4833);
or UO_199 (O_199,N_4938,N_4570);
nand UO_200 (O_200,N_4539,N_4919);
nand UO_201 (O_201,N_4932,N_4656);
and UO_202 (O_202,N_4626,N_4700);
nand UO_203 (O_203,N_4511,N_4901);
and UO_204 (O_204,N_4715,N_4957);
nand UO_205 (O_205,N_4512,N_4987);
nand UO_206 (O_206,N_4624,N_4676);
or UO_207 (O_207,N_4731,N_4721);
nand UO_208 (O_208,N_4654,N_4500);
or UO_209 (O_209,N_4854,N_4702);
xnor UO_210 (O_210,N_4873,N_4902);
nand UO_211 (O_211,N_4737,N_4598);
nor UO_212 (O_212,N_4704,N_4766);
xor UO_213 (O_213,N_4814,N_4699);
nor UO_214 (O_214,N_4581,N_4835);
nor UO_215 (O_215,N_4697,N_4659);
nand UO_216 (O_216,N_4514,N_4777);
or UO_217 (O_217,N_4949,N_4977);
nor UO_218 (O_218,N_4650,N_4587);
or UO_219 (O_219,N_4944,N_4785);
and UO_220 (O_220,N_4892,N_4971);
nor UO_221 (O_221,N_4999,N_4711);
nand UO_222 (O_222,N_4929,N_4845);
nor UO_223 (O_223,N_4549,N_4664);
and UO_224 (O_224,N_4522,N_4556);
and UO_225 (O_225,N_4730,N_4931);
xnor UO_226 (O_226,N_4592,N_4818);
and UO_227 (O_227,N_4831,N_4779);
or UO_228 (O_228,N_4907,N_4665);
nand UO_229 (O_229,N_4934,N_4981);
or UO_230 (O_230,N_4513,N_4568);
and UO_231 (O_231,N_4759,N_4787);
xor UO_232 (O_232,N_4603,N_4678);
xnor UO_233 (O_233,N_4903,N_4851);
nand UO_234 (O_234,N_4775,N_4860);
or UO_235 (O_235,N_4529,N_4954);
and UO_236 (O_236,N_4658,N_4763);
nor UO_237 (O_237,N_4703,N_4728);
or UO_238 (O_238,N_4933,N_4962);
nor UO_239 (O_239,N_4838,N_4516);
and UO_240 (O_240,N_4774,N_4692);
nand UO_241 (O_241,N_4828,N_4684);
or UO_242 (O_242,N_4694,N_4751);
and UO_243 (O_243,N_4630,N_4622);
nand UO_244 (O_244,N_4869,N_4601);
nor UO_245 (O_245,N_4527,N_4900);
xnor UO_246 (O_246,N_4956,N_4788);
nor UO_247 (O_247,N_4550,N_4577);
nand UO_248 (O_248,N_4523,N_4797);
nor UO_249 (O_249,N_4593,N_4505);
and UO_250 (O_250,N_4864,N_4501);
or UO_251 (O_251,N_4844,N_4644);
nand UO_252 (O_252,N_4933,N_4596);
or UO_253 (O_253,N_4647,N_4989);
nand UO_254 (O_254,N_4678,N_4773);
nor UO_255 (O_255,N_4544,N_4633);
xnor UO_256 (O_256,N_4989,N_4760);
and UO_257 (O_257,N_4609,N_4680);
or UO_258 (O_258,N_4517,N_4535);
or UO_259 (O_259,N_4539,N_4534);
nand UO_260 (O_260,N_4872,N_4745);
and UO_261 (O_261,N_4604,N_4508);
and UO_262 (O_262,N_4809,N_4581);
and UO_263 (O_263,N_4724,N_4733);
xor UO_264 (O_264,N_4702,N_4907);
and UO_265 (O_265,N_4888,N_4555);
and UO_266 (O_266,N_4865,N_4614);
nor UO_267 (O_267,N_4691,N_4656);
nor UO_268 (O_268,N_4625,N_4992);
xnor UO_269 (O_269,N_4758,N_4666);
or UO_270 (O_270,N_4776,N_4702);
nor UO_271 (O_271,N_4900,N_4834);
and UO_272 (O_272,N_4534,N_4971);
or UO_273 (O_273,N_4647,N_4898);
nand UO_274 (O_274,N_4558,N_4860);
nand UO_275 (O_275,N_4969,N_4544);
xor UO_276 (O_276,N_4773,N_4988);
nand UO_277 (O_277,N_4674,N_4724);
nor UO_278 (O_278,N_4963,N_4628);
nand UO_279 (O_279,N_4554,N_4666);
xor UO_280 (O_280,N_4658,N_4895);
xor UO_281 (O_281,N_4767,N_4845);
and UO_282 (O_282,N_4959,N_4696);
or UO_283 (O_283,N_4649,N_4753);
xnor UO_284 (O_284,N_4995,N_4893);
or UO_285 (O_285,N_4900,N_4581);
or UO_286 (O_286,N_4684,N_4765);
nor UO_287 (O_287,N_4897,N_4764);
or UO_288 (O_288,N_4596,N_4808);
or UO_289 (O_289,N_4709,N_4663);
and UO_290 (O_290,N_4673,N_4545);
and UO_291 (O_291,N_4818,N_4893);
nor UO_292 (O_292,N_4762,N_4985);
nand UO_293 (O_293,N_4695,N_4749);
nor UO_294 (O_294,N_4970,N_4923);
xnor UO_295 (O_295,N_4549,N_4827);
or UO_296 (O_296,N_4775,N_4725);
or UO_297 (O_297,N_4548,N_4814);
and UO_298 (O_298,N_4672,N_4868);
nor UO_299 (O_299,N_4651,N_4515);
nor UO_300 (O_300,N_4723,N_4886);
or UO_301 (O_301,N_4914,N_4700);
xor UO_302 (O_302,N_4928,N_4769);
and UO_303 (O_303,N_4901,N_4742);
or UO_304 (O_304,N_4757,N_4506);
nand UO_305 (O_305,N_4996,N_4679);
and UO_306 (O_306,N_4595,N_4915);
and UO_307 (O_307,N_4807,N_4692);
or UO_308 (O_308,N_4738,N_4829);
and UO_309 (O_309,N_4597,N_4637);
and UO_310 (O_310,N_4847,N_4713);
nor UO_311 (O_311,N_4532,N_4866);
xnor UO_312 (O_312,N_4819,N_4658);
nor UO_313 (O_313,N_4650,N_4959);
nand UO_314 (O_314,N_4599,N_4788);
nand UO_315 (O_315,N_4840,N_4854);
xnor UO_316 (O_316,N_4814,N_4684);
nand UO_317 (O_317,N_4591,N_4531);
or UO_318 (O_318,N_4692,N_4697);
nor UO_319 (O_319,N_4558,N_4786);
or UO_320 (O_320,N_4904,N_4568);
nor UO_321 (O_321,N_4911,N_4792);
and UO_322 (O_322,N_4979,N_4531);
nor UO_323 (O_323,N_4704,N_4978);
nor UO_324 (O_324,N_4715,N_4649);
or UO_325 (O_325,N_4500,N_4956);
and UO_326 (O_326,N_4924,N_4673);
xor UO_327 (O_327,N_4812,N_4611);
nand UO_328 (O_328,N_4501,N_4969);
or UO_329 (O_329,N_4573,N_4713);
nor UO_330 (O_330,N_4618,N_4828);
nor UO_331 (O_331,N_4907,N_4636);
nor UO_332 (O_332,N_4527,N_4833);
nand UO_333 (O_333,N_4685,N_4954);
nor UO_334 (O_334,N_4566,N_4931);
or UO_335 (O_335,N_4560,N_4697);
nor UO_336 (O_336,N_4804,N_4524);
and UO_337 (O_337,N_4539,N_4596);
nor UO_338 (O_338,N_4925,N_4995);
nor UO_339 (O_339,N_4622,N_4706);
xnor UO_340 (O_340,N_4516,N_4638);
nor UO_341 (O_341,N_4554,N_4678);
or UO_342 (O_342,N_4556,N_4869);
or UO_343 (O_343,N_4765,N_4976);
and UO_344 (O_344,N_4558,N_4546);
and UO_345 (O_345,N_4681,N_4504);
nand UO_346 (O_346,N_4706,N_4923);
and UO_347 (O_347,N_4844,N_4819);
or UO_348 (O_348,N_4608,N_4982);
nand UO_349 (O_349,N_4796,N_4779);
nor UO_350 (O_350,N_4726,N_4847);
nand UO_351 (O_351,N_4810,N_4760);
and UO_352 (O_352,N_4630,N_4814);
nand UO_353 (O_353,N_4730,N_4821);
xor UO_354 (O_354,N_4774,N_4653);
or UO_355 (O_355,N_4845,N_4977);
and UO_356 (O_356,N_4677,N_4703);
nand UO_357 (O_357,N_4940,N_4788);
nand UO_358 (O_358,N_4573,N_4947);
and UO_359 (O_359,N_4645,N_4668);
or UO_360 (O_360,N_4853,N_4576);
nand UO_361 (O_361,N_4752,N_4890);
nand UO_362 (O_362,N_4553,N_4600);
nor UO_363 (O_363,N_4607,N_4668);
nor UO_364 (O_364,N_4815,N_4681);
and UO_365 (O_365,N_4881,N_4623);
nand UO_366 (O_366,N_4903,N_4597);
or UO_367 (O_367,N_4960,N_4942);
nor UO_368 (O_368,N_4933,N_4857);
nand UO_369 (O_369,N_4555,N_4745);
nand UO_370 (O_370,N_4649,N_4783);
or UO_371 (O_371,N_4690,N_4865);
nor UO_372 (O_372,N_4723,N_4596);
and UO_373 (O_373,N_4554,N_4936);
and UO_374 (O_374,N_4905,N_4693);
or UO_375 (O_375,N_4730,N_4645);
and UO_376 (O_376,N_4546,N_4624);
nor UO_377 (O_377,N_4998,N_4664);
nand UO_378 (O_378,N_4534,N_4631);
or UO_379 (O_379,N_4750,N_4506);
nand UO_380 (O_380,N_4688,N_4717);
nor UO_381 (O_381,N_4765,N_4873);
nor UO_382 (O_382,N_4829,N_4936);
and UO_383 (O_383,N_4595,N_4597);
nand UO_384 (O_384,N_4625,N_4904);
nor UO_385 (O_385,N_4972,N_4575);
and UO_386 (O_386,N_4682,N_4957);
xnor UO_387 (O_387,N_4576,N_4511);
and UO_388 (O_388,N_4978,N_4553);
and UO_389 (O_389,N_4960,N_4929);
or UO_390 (O_390,N_4820,N_4640);
and UO_391 (O_391,N_4547,N_4966);
nor UO_392 (O_392,N_4748,N_4720);
xor UO_393 (O_393,N_4781,N_4528);
xor UO_394 (O_394,N_4972,N_4823);
xor UO_395 (O_395,N_4533,N_4625);
nor UO_396 (O_396,N_4652,N_4924);
nand UO_397 (O_397,N_4602,N_4919);
nand UO_398 (O_398,N_4994,N_4516);
and UO_399 (O_399,N_4761,N_4588);
or UO_400 (O_400,N_4538,N_4582);
nand UO_401 (O_401,N_4849,N_4632);
nand UO_402 (O_402,N_4645,N_4619);
and UO_403 (O_403,N_4756,N_4995);
nor UO_404 (O_404,N_4786,N_4881);
and UO_405 (O_405,N_4991,N_4536);
nand UO_406 (O_406,N_4804,N_4831);
nor UO_407 (O_407,N_4646,N_4816);
nand UO_408 (O_408,N_4531,N_4752);
nand UO_409 (O_409,N_4903,N_4869);
xnor UO_410 (O_410,N_4720,N_4638);
nor UO_411 (O_411,N_4555,N_4573);
or UO_412 (O_412,N_4521,N_4544);
and UO_413 (O_413,N_4892,N_4870);
or UO_414 (O_414,N_4856,N_4639);
nand UO_415 (O_415,N_4777,N_4678);
nor UO_416 (O_416,N_4997,N_4802);
nor UO_417 (O_417,N_4931,N_4783);
xor UO_418 (O_418,N_4565,N_4912);
or UO_419 (O_419,N_4827,N_4673);
and UO_420 (O_420,N_4632,N_4664);
xnor UO_421 (O_421,N_4640,N_4952);
and UO_422 (O_422,N_4676,N_4831);
or UO_423 (O_423,N_4776,N_4550);
xor UO_424 (O_424,N_4531,N_4634);
or UO_425 (O_425,N_4598,N_4879);
xnor UO_426 (O_426,N_4671,N_4549);
or UO_427 (O_427,N_4765,N_4746);
nor UO_428 (O_428,N_4654,N_4679);
or UO_429 (O_429,N_4589,N_4610);
nor UO_430 (O_430,N_4560,N_4686);
nor UO_431 (O_431,N_4662,N_4959);
and UO_432 (O_432,N_4897,N_4738);
or UO_433 (O_433,N_4790,N_4749);
nor UO_434 (O_434,N_4976,N_4789);
or UO_435 (O_435,N_4510,N_4624);
and UO_436 (O_436,N_4782,N_4780);
nor UO_437 (O_437,N_4913,N_4698);
or UO_438 (O_438,N_4993,N_4810);
nand UO_439 (O_439,N_4839,N_4708);
and UO_440 (O_440,N_4548,N_4712);
nand UO_441 (O_441,N_4516,N_4955);
or UO_442 (O_442,N_4770,N_4913);
nand UO_443 (O_443,N_4906,N_4900);
nor UO_444 (O_444,N_4987,N_4607);
and UO_445 (O_445,N_4537,N_4755);
nand UO_446 (O_446,N_4696,N_4958);
nor UO_447 (O_447,N_4827,N_4907);
nand UO_448 (O_448,N_4628,N_4681);
nand UO_449 (O_449,N_4612,N_4951);
nor UO_450 (O_450,N_4772,N_4511);
or UO_451 (O_451,N_4704,N_4767);
nor UO_452 (O_452,N_4759,N_4766);
and UO_453 (O_453,N_4661,N_4999);
and UO_454 (O_454,N_4506,N_4744);
and UO_455 (O_455,N_4969,N_4897);
nor UO_456 (O_456,N_4936,N_4758);
xor UO_457 (O_457,N_4915,N_4664);
nor UO_458 (O_458,N_4795,N_4856);
nand UO_459 (O_459,N_4528,N_4593);
nand UO_460 (O_460,N_4741,N_4937);
and UO_461 (O_461,N_4791,N_4940);
nor UO_462 (O_462,N_4901,N_4782);
nand UO_463 (O_463,N_4668,N_4987);
or UO_464 (O_464,N_4546,N_4968);
nand UO_465 (O_465,N_4899,N_4699);
nand UO_466 (O_466,N_4854,N_4692);
xor UO_467 (O_467,N_4957,N_4714);
xor UO_468 (O_468,N_4972,N_4977);
nor UO_469 (O_469,N_4772,N_4623);
and UO_470 (O_470,N_4642,N_4860);
or UO_471 (O_471,N_4661,N_4772);
or UO_472 (O_472,N_4542,N_4908);
xor UO_473 (O_473,N_4554,N_4559);
xnor UO_474 (O_474,N_4981,N_4539);
nand UO_475 (O_475,N_4822,N_4581);
nor UO_476 (O_476,N_4760,N_4595);
and UO_477 (O_477,N_4908,N_4705);
xor UO_478 (O_478,N_4974,N_4777);
or UO_479 (O_479,N_4597,N_4998);
nand UO_480 (O_480,N_4557,N_4693);
nand UO_481 (O_481,N_4556,N_4518);
or UO_482 (O_482,N_4627,N_4762);
xnor UO_483 (O_483,N_4653,N_4709);
nand UO_484 (O_484,N_4833,N_4918);
nand UO_485 (O_485,N_4505,N_4592);
nand UO_486 (O_486,N_4691,N_4732);
or UO_487 (O_487,N_4746,N_4776);
xor UO_488 (O_488,N_4808,N_4776);
and UO_489 (O_489,N_4969,N_4752);
nor UO_490 (O_490,N_4504,N_4622);
and UO_491 (O_491,N_4947,N_4504);
and UO_492 (O_492,N_4500,N_4998);
and UO_493 (O_493,N_4576,N_4789);
nand UO_494 (O_494,N_4751,N_4834);
xor UO_495 (O_495,N_4961,N_4681);
nand UO_496 (O_496,N_4721,N_4681);
and UO_497 (O_497,N_4611,N_4974);
and UO_498 (O_498,N_4870,N_4901);
xnor UO_499 (O_499,N_4559,N_4634);
xor UO_500 (O_500,N_4747,N_4855);
nor UO_501 (O_501,N_4532,N_4959);
nor UO_502 (O_502,N_4924,N_4730);
nand UO_503 (O_503,N_4848,N_4800);
and UO_504 (O_504,N_4800,N_4964);
nand UO_505 (O_505,N_4955,N_4848);
nor UO_506 (O_506,N_4551,N_4672);
and UO_507 (O_507,N_4943,N_4515);
and UO_508 (O_508,N_4834,N_4671);
or UO_509 (O_509,N_4632,N_4801);
nand UO_510 (O_510,N_4888,N_4751);
nor UO_511 (O_511,N_4851,N_4595);
nor UO_512 (O_512,N_4536,N_4655);
xnor UO_513 (O_513,N_4969,N_4576);
nand UO_514 (O_514,N_4835,N_4607);
and UO_515 (O_515,N_4672,N_4539);
or UO_516 (O_516,N_4569,N_4517);
and UO_517 (O_517,N_4841,N_4948);
or UO_518 (O_518,N_4698,N_4703);
xnor UO_519 (O_519,N_4627,N_4909);
nand UO_520 (O_520,N_4664,N_4851);
nor UO_521 (O_521,N_4540,N_4819);
nand UO_522 (O_522,N_4893,N_4796);
xnor UO_523 (O_523,N_4641,N_4739);
nand UO_524 (O_524,N_4638,N_4713);
nor UO_525 (O_525,N_4780,N_4624);
and UO_526 (O_526,N_4619,N_4791);
and UO_527 (O_527,N_4528,N_4628);
nor UO_528 (O_528,N_4570,N_4820);
xor UO_529 (O_529,N_4900,N_4996);
nand UO_530 (O_530,N_4589,N_4804);
xor UO_531 (O_531,N_4773,N_4774);
and UO_532 (O_532,N_4788,N_4946);
nor UO_533 (O_533,N_4758,N_4996);
nand UO_534 (O_534,N_4948,N_4983);
nor UO_535 (O_535,N_4527,N_4666);
xnor UO_536 (O_536,N_4926,N_4610);
nand UO_537 (O_537,N_4992,N_4668);
and UO_538 (O_538,N_4643,N_4571);
or UO_539 (O_539,N_4755,N_4869);
nand UO_540 (O_540,N_4865,N_4764);
nand UO_541 (O_541,N_4926,N_4973);
nor UO_542 (O_542,N_4847,N_4685);
nor UO_543 (O_543,N_4990,N_4522);
and UO_544 (O_544,N_4799,N_4808);
or UO_545 (O_545,N_4994,N_4913);
nor UO_546 (O_546,N_4770,N_4501);
or UO_547 (O_547,N_4621,N_4920);
and UO_548 (O_548,N_4897,N_4599);
xnor UO_549 (O_549,N_4930,N_4838);
nor UO_550 (O_550,N_4506,N_4786);
nor UO_551 (O_551,N_4536,N_4930);
nor UO_552 (O_552,N_4933,N_4951);
nor UO_553 (O_553,N_4993,N_4687);
nand UO_554 (O_554,N_4752,N_4931);
nand UO_555 (O_555,N_4501,N_4776);
xor UO_556 (O_556,N_4938,N_4535);
and UO_557 (O_557,N_4872,N_4542);
xor UO_558 (O_558,N_4988,N_4588);
nand UO_559 (O_559,N_4564,N_4720);
nor UO_560 (O_560,N_4671,N_4991);
nand UO_561 (O_561,N_4987,N_4775);
xnor UO_562 (O_562,N_4977,N_4937);
or UO_563 (O_563,N_4565,N_4555);
nor UO_564 (O_564,N_4742,N_4533);
or UO_565 (O_565,N_4618,N_4514);
and UO_566 (O_566,N_4901,N_4555);
and UO_567 (O_567,N_4776,N_4738);
nand UO_568 (O_568,N_4530,N_4678);
nor UO_569 (O_569,N_4981,N_4704);
nor UO_570 (O_570,N_4932,N_4509);
and UO_571 (O_571,N_4747,N_4509);
nor UO_572 (O_572,N_4599,N_4813);
nor UO_573 (O_573,N_4680,N_4840);
xnor UO_574 (O_574,N_4974,N_4737);
nor UO_575 (O_575,N_4723,N_4830);
and UO_576 (O_576,N_4651,N_4790);
and UO_577 (O_577,N_4925,N_4798);
nor UO_578 (O_578,N_4871,N_4932);
nand UO_579 (O_579,N_4796,N_4979);
and UO_580 (O_580,N_4981,N_4558);
and UO_581 (O_581,N_4505,N_4678);
nand UO_582 (O_582,N_4806,N_4702);
nand UO_583 (O_583,N_4927,N_4669);
and UO_584 (O_584,N_4670,N_4807);
nand UO_585 (O_585,N_4664,N_4968);
nand UO_586 (O_586,N_4674,N_4808);
and UO_587 (O_587,N_4883,N_4516);
xnor UO_588 (O_588,N_4711,N_4841);
or UO_589 (O_589,N_4971,N_4895);
nand UO_590 (O_590,N_4938,N_4658);
or UO_591 (O_591,N_4744,N_4878);
nand UO_592 (O_592,N_4658,N_4887);
or UO_593 (O_593,N_4650,N_4535);
nor UO_594 (O_594,N_4765,N_4554);
nor UO_595 (O_595,N_4838,N_4604);
nand UO_596 (O_596,N_4616,N_4597);
nand UO_597 (O_597,N_4590,N_4653);
or UO_598 (O_598,N_4658,N_4703);
and UO_599 (O_599,N_4827,N_4574);
xnor UO_600 (O_600,N_4705,N_4791);
and UO_601 (O_601,N_4809,N_4687);
xor UO_602 (O_602,N_4771,N_4567);
xor UO_603 (O_603,N_4651,N_4996);
nor UO_604 (O_604,N_4753,N_4679);
nand UO_605 (O_605,N_4687,N_4754);
nand UO_606 (O_606,N_4904,N_4883);
nand UO_607 (O_607,N_4696,N_4825);
nand UO_608 (O_608,N_4934,N_4841);
nand UO_609 (O_609,N_4682,N_4508);
or UO_610 (O_610,N_4810,N_4756);
and UO_611 (O_611,N_4810,N_4715);
xor UO_612 (O_612,N_4949,N_4779);
nand UO_613 (O_613,N_4886,N_4524);
or UO_614 (O_614,N_4586,N_4927);
or UO_615 (O_615,N_4525,N_4829);
and UO_616 (O_616,N_4996,N_4946);
nor UO_617 (O_617,N_4586,N_4617);
nor UO_618 (O_618,N_4654,N_4540);
or UO_619 (O_619,N_4785,N_4723);
xor UO_620 (O_620,N_4970,N_4771);
and UO_621 (O_621,N_4944,N_4744);
xnor UO_622 (O_622,N_4841,N_4675);
xnor UO_623 (O_623,N_4792,N_4601);
nor UO_624 (O_624,N_4578,N_4740);
nand UO_625 (O_625,N_4691,N_4896);
or UO_626 (O_626,N_4769,N_4999);
nand UO_627 (O_627,N_4798,N_4703);
and UO_628 (O_628,N_4882,N_4833);
nor UO_629 (O_629,N_4612,N_4991);
nand UO_630 (O_630,N_4812,N_4551);
nor UO_631 (O_631,N_4831,N_4719);
or UO_632 (O_632,N_4973,N_4612);
and UO_633 (O_633,N_4644,N_4920);
or UO_634 (O_634,N_4519,N_4591);
nand UO_635 (O_635,N_4652,N_4768);
nand UO_636 (O_636,N_4781,N_4569);
or UO_637 (O_637,N_4769,N_4701);
or UO_638 (O_638,N_4697,N_4698);
and UO_639 (O_639,N_4871,N_4764);
xnor UO_640 (O_640,N_4635,N_4653);
xor UO_641 (O_641,N_4664,N_4653);
nor UO_642 (O_642,N_4842,N_4929);
nor UO_643 (O_643,N_4592,N_4642);
and UO_644 (O_644,N_4950,N_4904);
nand UO_645 (O_645,N_4957,N_4502);
nor UO_646 (O_646,N_4557,N_4592);
nand UO_647 (O_647,N_4600,N_4652);
and UO_648 (O_648,N_4793,N_4671);
nand UO_649 (O_649,N_4900,N_4839);
and UO_650 (O_650,N_4599,N_4982);
nand UO_651 (O_651,N_4963,N_4660);
nand UO_652 (O_652,N_4687,N_4677);
xor UO_653 (O_653,N_4999,N_4782);
nor UO_654 (O_654,N_4872,N_4786);
and UO_655 (O_655,N_4511,N_4913);
nor UO_656 (O_656,N_4717,N_4602);
nor UO_657 (O_657,N_4666,N_4801);
nand UO_658 (O_658,N_4933,N_4869);
xor UO_659 (O_659,N_4979,N_4593);
xor UO_660 (O_660,N_4786,N_4531);
nor UO_661 (O_661,N_4968,N_4985);
nor UO_662 (O_662,N_4768,N_4803);
nor UO_663 (O_663,N_4742,N_4525);
and UO_664 (O_664,N_4933,N_4631);
or UO_665 (O_665,N_4856,N_4971);
or UO_666 (O_666,N_4581,N_4709);
and UO_667 (O_667,N_4609,N_4541);
and UO_668 (O_668,N_4791,N_4742);
and UO_669 (O_669,N_4596,N_4935);
and UO_670 (O_670,N_4849,N_4556);
or UO_671 (O_671,N_4684,N_4594);
or UO_672 (O_672,N_4802,N_4518);
and UO_673 (O_673,N_4515,N_4951);
nand UO_674 (O_674,N_4506,N_4930);
and UO_675 (O_675,N_4826,N_4994);
nand UO_676 (O_676,N_4677,N_4662);
or UO_677 (O_677,N_4879,N_4919);
nor UO_678 (O_678,N_4765,N_4849);
nor UO_679 (O_679,N_4908,N_4579);
or UO_680 (O_680,N_4528,N_4673);
nand UO_681 (O_681,N_4923,N_4723);
nor UO_682 (O_682,N_4957,N_4813);
nand UO_683 (O_683,N_4612,N_4893);
nand UO_684 (O_684,N_4868,N_4910);
or UO_685 (O_685,N_4657,N_4634);
and UO_686 (O_686,N_4708,N_4856);
nand UO_687 (O_687,N_4994,N_4857);
nand UO_688 (O_688,N_4611,N_4737);
nand UO_689 (O_689,N_4737,N_4560);
and UO_690 (O_690,N_4733,N_4532);
xor UO_691 (O_691,N_4598,N_4990);
nand UO_692 (O_692,N_4861,N_4985);
nand UO_693 (O_693,N_4972,N_4502);
xnor UO_694 (O_694,N_4902,N_4846);
or UO_695 (O_695,N_4589,N_4793);
nor UO_696 (O_696,N_4800,N_4547);
nand UO_697 (O_697,N_4548,N_4886);
and UO_698 (O_698,N_4606,N_4687);
nand UO_699 (O_699,N_4626,N_4797);
nor UO_700 (O_700,N_4957,N_4601);
or UO_701 (O_701,N_4599,N_4943);
and UO_702 (O_702,N_4932,N_4898);
nand UO_703 (O_703,N_4762,N_4503);
nand UO_704 (O_704,N_4637,N_4817);
or UO_705 (O_705,N_4721,N_4801);
or UO_706 (O_706,N_4741,N_4966);
and UO_707 (O_707,N_4691,N_4923);
and UO_708 (O_708,N_4587,N_4681);
xnor UO_709 (O_709,N_4673,N_4503);
nand UO_710 (O_710,N_4720,N_4770);
nand UO_711 (O_711,N_4547,N_4840);
nand UO_712 (O_712,N_4945,N_4714);
nor UO_713 (O_713,N_4908,N_4624);
nand UO_714 (O_714,N_4987,N_4507);
or UO_715 (O_715,N_4717,N_4701);
nor UO_716 (O_716,N_4513,N_4760);
nand UO_717 (O_717,N_4522,N_4666);
nand UO_718 (O_718,N_4778,N_4586);
xor UO_719 (O_719,N_4906,N_4670);
and UO_720 (O_720,N_4629,N_4812);
nand UO_721 (O_721,N_4996,N_4674);
and UO_722 (O_722,N_4722,N_4715);
and UO_723 (O_723,N_4707,N_4784);
nor UO_724 (O_724,N_4542,N_4554);
or UO_725 (O_725,N_4598,N_4502);
nand UO_726 (O_726,N_4541,N_4894);
or UO_727 (O_727,N_4608,N_4922);
nand UO_728 (O_728,N_4746,N_4860);
or UO_729 (O_729,N_4716,N_4876);
xnor UO_730 (O_730,N_4682,N_4598);
nand UO_731 (O_731,N_4988,N_4547);
or UO_732 (O_732,N_4930,N_4552);
nor UO_733 (O_733,N_4976,N_4703);
nand UO_734 (O_734,N_4715,N_4778);
nand UO_735 (O_735,N_4759,N_4935);
nor UO_736 (O_736,N_4984,N_4783);
xnor UO_737 (O_737,N_4909,N_4532);
or UO_738 (O_738,N_4866,N_4637);
nand UO_739 (O_739,N_4585,N_4532);
nand UO_740 (O_740,N_4830,N_4683);
or UO_741 (O_741,N_4775,N_4515);
nand UO_742 (O_742,N_4806,N_4826);
and UO_743 (O_743,N_4770,N_4553);
and UO_744 (O_744,N_4514,N_4703);
nor UO_745 (O_745,N_4577,N_4551);
and UO_746 (O_746,N_4511,N_4537);
nor UO_747 (O_747,N_4981,N_4914);
or UO_748 (O_748,N_4679,N_4928);
and UO_749 (O_749,N_4603,N_4578);
xnor UO_750 (O_750,N_4599,N_4954);
xor UO_751 (O_751,N_4861,N_4940);
and UO_752 (O_752,N_4842,N_4758);
nand UO_753 (O_753,N_4874,N_4557);
nand UO_754 (O_754,N_4963,N_4912);
nand UO_755 (O_755,N_4658,N_4932);
xor UO_756 (O_756,N_4817,N_4967);
and UO_757 (O_757,N_4851,N_4905);
nand UO_758 (O_758,N_4753,N_4995);
nand UO_759 (O_759,N_4976,N_4532);
and UO_760 (O_760,N_4926,N_4711);
and UO_761 (O_761,N_4646,N_4998);
or UO_762 (O_762,N_4708,N_4754);
nand UO_763 (O_763,N_4662,N_4690);
xor UO_764 (O_764,N_4759,N_4971);
nand UO_765 (O_765,N_4673,N_4890);
and UO_766 (O_766,N_4840,N_4767);
and UO_767 (O_767,N_4775,N_4762);
and UO_768 (O_768,N_4619,N_4983);
nor UO_769 (O_769,N_4958,N_4619);
or UO_770 (O_770,N_4790,N_4637);
nand UO_771 (O_771,N_4649,N_4996);
and UO_772 (O_772,N_4542,N_4729);
and UO_773 (O_773,N_4893,N_4691);
nand UO_774 (O_774,N_4529,N_4676);
or UO_775 (O_775,N_4770,N_4594);
or UO_776 (O_776,N_4510,N_4867);
nor UO_777 (O_777,N_4849,N_4736);
nand UO_778 (O_778,N_4513,N_4848);
and UO_779 (O_779,N_4623,N_4917);
xnor UO_780 (O_780,N_4934,N_4689);
nand UO_781 (O_781,N_4835,N_4509);
xor UO_782 (O_782,N_4893,N_4751);
nand UO_783 (O_783,N_4683,N_4597);
and UO_784 (O_784,N_4778,N_4741);
nor UO_785 (O_785,N_4666,N_4635);
nand UO_786 (O_786,N_4704,N_4847);
or UO_787 (O_787,N_4765,N_4704);
or UO_788 (O_788,N_4717,N_4642);
and UO_789 (O_789,N_4614,N_4580);
nor UO_790 (O_790,N_4716,N_4880);
nor UO_791 (O_791,N_4605,N_4992);
nand UO_792 (O_792,N_4635,N_4665);
nor UO_793 (O_793,N_4611,N_4868);
and UO_794 (O_794,N_4938,N_4944);
nand UO_795 (O_795,N_4973,N_4568);
and UO_796 (O_796,N_4973,N_4505);
or UO_797 (O_797,N_4587,N_4856);
and UO_798 (O_798,N_4549,N_4825);
or UO_799 (O_799,N_4974,N_4948);
nand UO_800 (O_800,N_4500,N_4706);
and UO_801 (O_801,N_4798,N_4502);
xor UO_802 (O_802,N_4920,N_4767);
and UO_803 (O_803,N_4933,N_4735);
nand UO_804 (O_804,N_4714,N_4673);
and UO_805 (O_805,N_4601,N_4916);
or UO_806 (O_806,N_4940,N_4955);
nand UO_807 (O_807,N_4975,N_4881);
or UO_808 (O_808,N_4997,N_4703);
nor UO_809 (O_809,N_4819,N_4558);
xnor UO_810 (O_810,N_4728,N_4642);
nand UO_811 (O_811,N_4543,N_4844);
nand UO_812 (O_812,N_4597,N_4972);
or UO_813 (O_813,N_4645,N_4969);
nand UO_814 (O_814,N_4886,N_4820);
and UO_815 (O_815,N_4737,N_4699);
xor UO_816 (O_816,N_4688,N_4589);
nand UO_817 (O_817,N_4886,N_4962);
nand UO_818 (O_818,N_4954,N_4856);
nor UO_819 (O_819,N_4917,N_4513);
nand UO_820 (O_820,N_4867,N_4625);
or UO_821 (O_821,N_4727,N_4870);
nand UO_822 (O_822,N_4997,N_4644);
and UO_823 (O_823,N_4601,N_4556);
or UO_824 (O_824,N_4818,N_4621);
and UO_825 (O_825,N_4810,N_4723);
xnor UO_826 (O_826,N_4874,N_4697);
or UO_827 (O_827,N_4690,N_4890);
nand UO_828 (O_828,N_4956,N_4508);
and UO_829 (O_829,N_4659,N_4574);
and UO_830 (O_830,N_4753,N_4747);
nand UO_831 (O_831,N_4739,N_4801);
and UO_832 (O_832,N_4940,N_4679);
or UO_833 (O_833,N_4626,N_4705);
and UO_834 (O_834,N_4659,N_4736);
xnor UO_835 (O_835,N_4789,N_4921);
or UO_836 (O_836,N_4639,N_4623);
nor UO_837 (O_837,N_4572,N_4930);
or UO_838 (O_838,N_4761,N_4980);
and UO_839 (O_839,N_4827,N_4678);
or UO_840 (O_840,N_4776,N_4646);
nand UO_841 (O_841,N_4703,N_4550);
xnor UO_842 (O_842,N_4873,N_4954);
nor UO_843 (O_843,N_4686,N_4705);
or UO_844 (O_844,N_4804,N_4502);
xor UO_845 (O_845,N_4807,N_4822);
nand UO_846 (O_846,N_4709,N_4975);
and UO_847 (O_847,N_4584,N_4932);
nor UO_848 (O_848,N_4897,N_4772);
nand UO_849 (O_849,N_4723,N_4674);
and UO_850 (O_850,N_4993,N_4633);
xor UO_851 (O_851,N_4809,N_4924);
nand UO_852 (O_852,N_4643,N_4895);
or UO_853 (O_853,N_4793,N_4983);
or UO_854 (O_854,N_4758,N_4667);
nor UO_855 (O_855,N_4744,N_4719);
and UO_856 (O_856,N_4582,N_4946);
or UO_857 (O_857,N_4851,N_4538);
or UO_858 (O_858,N_4990,N_4671);
nor UO_859 (O_859,N_4676,N_4619);
and UO_860 (O_860,N_4650,N_4606);
and UO_861 (O_861,N_4667,N_4843);
xor UO_862 (O_862,N_4669,N_4935);
and UO_863 (O_863,N_4962,N_4714);
nand UO_864 (O_864,N_4964,N_4999);
nand UO_865 (O_865,N_4545,N_4748);
or UO_866 (O_866,N_4988,N_4896);
and UO_867 (O_867,N_4647,N_4777);
or UO_868 (O_868,N_4953,N_4600);
nor UO_869 (O_869,N_4914,N_4612);
nor UO_870 (O_870,N_4750,N_4700);
or UO_871 (O_871,N_4562,N_4527);
nand UO_872 (O_872,N_4951,N_4725);
or UO_873 (O_873,N_4562,N_4531);
nand UO_874 (O_874,N_4520,N_4996);
and UO_875 (O_875,N_4832,N_4756);
nor UO_876 (O_876,N_4914,N_4861);
nor UO_877 (O_877,N_4624,N_4558);
nor UO_878 (O_878,N_4814,N_4615);
or UO_879 (O_879,N_4842,N_4587);
nor UO_880 (O_880,N_4971,N_4772);
and UO_881 (O_881,N_4839,N_4957);
or UO_882 (O_882,N_4688,N_4641);
nor UO_883 (O_883,N_4964,N_4562);
xnor UO_884 (O_884,N_4695,N_4923);
xor UO_885 (O_885,N_4938,N_4884);
nor UO_886 (O_886,N_4901,N_4842);
nand UO_887 (O_887,N_4628,N_4838);
nor UO_888 (O_888,N_4512,N_4647);
nand UO_889 (O_889,N_4648,N_4527);
nor UO_890 (O_890,N_4832,N_4992);
or UO_891 (O_891,N_4503,N_4512);
nand UO_892 (O_892,N_4820,N_4774);
nor UO_893 (O_893,N_4506,N_4527);
or UO_894 (O_894,N_4981,N_4811);
and UO_895 (O_895,N_4940,N_4715);
nor UO_896 (O_896,N_4989,N_4805);
and UO_897 (O_897,N_4693,N_4854);
and UO_898 (O_898,N_4784,N_4619);
and UO_899 (O_899,N_4588,N_4890);
or UO_900 (O_900,N_4871,N_4891);
nand UO_901 (O_901,N_4648,N_4669);
or UO_902 (O_902,N_4682,N_4773);
nor UO_903 (O_903,N_4911,N_4777);
or UO_904 (O_904,N_4594,N_4571);
nor UO_905 (O_905,N_4523,N_4999);
nor UO_906 (O_906,N_4846,N_4934);
and UO_907 (O_907,N_4719,N_4687);
nand UO_908 (O_908,N_4826,N_4608);
and UO_909 (O_909,N_4826,N_4991);
or UO_910 (O_910,N_4780,N_4833);
nor UO_911 (O_911,N_4730,N_4690);
nand UO_912 (O_912,N_4654,N_4993);
xnor UO_913 (O_913,N_4760,N_4963);
or UO_914 (O_914,N_4812,N_4817);
xor UO_915 (O_915,N_4787,N_4612);
and UO_916 (O_916,N_4666,N_4633);
and UO_917 (O_917,N_4615,N_4971);
and UO_918 (O_918,N_4959,N_4647);
and UO_919 (O_919,N_4743,N_4948);
nand UO_920 (O_920,N_4556,N_4964);
nand UO_921 (O_921,N_4699,N_4689);
nand UO_922 (O_922,N_4625,N_4813);
and UO_923 (O_923,N_4663,N_4988);
or UO_924 (O_924,N_4620,N_4720);
nand UO_925 (O_925,N_4544,N_4637);
or UO_926 (O_926,N_4570,N_4845);
nand UO_927 (O_927,N_4531,N_4530);
nand UO_928 (O_928,N_4632,N_4613);
and UO_929 (O_929,N_4891,N_4549);
nor UO_930 (O_930,N_4890,N_4995);
or UO_931 (O_931,N_4929,N_4672);
or UO_932 (O_932,N_4710,N_4600);
or UO_933 (O_933,N_4583,N_4783);
nand UO_934 (O_934,N_4606,N_4875);
nor UO_935 (O_935,N_4880,N_4675);
and UO_936 (O_936,N_4521,N_4907);
and UO_937 (O_937,N_4533,N_4600);
and UO_938 (O_938,N_4543,N_4504);
nand UO_939 (O_939,N_4638,N_4666);
nor UO_940 (O_940,N_4809,N_4985);
nand UO_941 (O_941,N_4567,N_4967);
nor UO_942 (O_942,N_4997,N_4832);
nor UO_943 (O_943,N_4593,N_4503);
nor UO_944 (O_944,N_4897,N_4884);
and UO_945 (O_945,N_4988,N_4501);
and UO_946 (O_946,N_4543,N_4583);
and UO_947 (O_947,N_4514,N_4773);
and UO_948 (O_948,N_4740,N_4521);
and UO_949 (O_949,N_4940,N_4783);
and UO_950 (O_950,N_4703,N_4814);
and UO_951 (O_951,N_4801,N_4764);
nand UO_952 (O_952,N_4776,N_4958);
nand UO_953 (O_953,N_4845,N_4565);
and UO_954 (O_954,N_4576,N_4769);
or UO_955 (O_955,N_4742,N_4703);
or UO_956 (O_956,N_4953,N_4843);
or UO_957 (O_957,N_4813,N_4543);
nand UO_958 (O_958,N_4811,N_4781);
and UO_959 (O_959,N_4539,N_4689);
nand UO_960 (O_960,N_4861,N_4728);
nand UO_961 (O_961,N_4703,N_4835);
or UO_962 (O_962,N_4987,N_4852);
or UO_963 (O_963,N_4809,N_4683);
xor UO_964 (O_964,N_4515,N_4659);
and UO_965 (O_965,N_4921,N_4829);
and UO_966 (O_966,N_4798,N_4546);
nor UO_967 (O_967,N_4964,N_4935);
nor UO_968 (O_968,N_4751,N_4716);
nand UO_969 (O_969,N_4964,N_4766);
nor UO_970 (O_970,N_4586,N_4668);
and UO_971 (O_971,N_4587,N_4640);
and UO_972 (O_972,N_4859,N_4913);
nand UO_973 (O_973,N_4946,N_4674);
nand UO_974 (O_974,N_4901,N_4835);
or UO_975 (O_975,N_4546,N_4752);
nor UO_976 (O_976,N_4807,N_4741);
and UO_977 (O_977,N_4522,N_4678);
xnor UO_978 (O_978,N_4738,N_4755);
and UO_979 (O_979,N_4833,N_4554);
and UO_980 (O_980,N_4664,N_4786);
or UO_981 (O_981,N_4792,N_4955);
nor UO_982 (O_982,N_4959,N_4969);
nor UO_983 (O_983,N_4532,N_4560);
nand UO_984 (O_984,N_4856,N_4852);
xnor UO_985 (O_985,N_4872,N_4951);
xor UO_986 (O_986,N_4522,N_4939);
xor UO_987 (O_987,N_4850,N_4959);
xor UO_988 (O_988,N_4707,N_4772);
nand UO_989 (O_989,N_4768,N_4685);
or UO_990 (O_990,N_4560,N_4791);
nand UO_991 (O_991,N_4662,N_4657);
and UO_992 (O_992,N_4705,N_4816);
or UO_993 (O_993,N_4758,N_4873);
nand UO_994 (O_994,N_4903,N_4760);
nand UO_995 (O_995,N_4949,N_4594);
and UO_996 (O_996,N_4899,N_4797);
nand UO_997 (O_997,N_4619,N_4599);
nor UO_998 (O_998,N_4659,N_4786);
nor UO_999 (O_999,N_4535,N_4525);
endmodule