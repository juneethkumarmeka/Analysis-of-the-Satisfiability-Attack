module basic_2500_25000_3000_100_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_2434,In_1526);
xor U1 (N_1,In_1837,In_1174);
and U2 (N_2,In_1424,In_914);
nor U3 (N_3,In_1401,In_1196);
xnor U4 (N_4,In_2047,In_2346);
and U5 (N_5,In_1370,In_1659);
xnor U6 (N_6,In_1362,In_2254);
nand U7 (N_7,In_635,In_1682);
nand U8 (N_8,In_76,In_644);
nor U9 (N_9,In_579,In_1316);
xor U10 (N_10,In_529,In_1958);
and U11 (N_11,In_1122,In_1304);
or U12 (N_12,In_2228,In_303);
or U13 (N_13,In_818,In_246);
nand U14 (N_14,In_1431,In_1386);
and U15 (N_15,In_1675,In_2327);
nor U16 (N_16,In_881,In_2258);
and U17 (N_17,In_2481,In_1282);
xor U18 (N_18,In_2038,In_402);
or U19 (N_19,In_1758,In_1228);
nand U20 (N_20,In_1392,In_1467);
nor U21 (N_21,In_779,In_549);
or U22 (N_22,In_742,In_532);
nand U23 (N_23,In_634,In_2362);
or U24 (N_24,In_774,In_1644);
nor U25 (N_25,In_1986,In_1398);
and U26 (N_26,In_2242,In_1396);
or U27 (N_27,In_253,In_1119);
and U28 (N_28,In_2154,In_684);
or U29 (N_29,In_1046,In_839);
or U30 (N_30,In_2227,In_5);
or U31 (N_31,In_985,In_1676);
or U32 (N_32,In_796,In_1246);
and U33 (N_33,In_636,In_1110);
or U34 (N_34,In_2009,In_135);
or U35 (N_35,In_1505,In_1479);
nand U36 (N_36,In_641,In_1480);
nor U37 (N_37,In_1691,In_1579);
xor U38 (N_38,In_2283,In_1887);
xor U39 (N_39,In_2135,In_2066);
and U40 (N_40,In_1694,In_2005);
and U41 (N_41,In_625,In_187);
and U42 (N_42,In_1210,In_2472);
nand U43 (N_43,In_723,In_2131);
nand U44 (N_44,In_995,In_314);
or U45 (N_45,In_631,In_627);
nor U46 (N_46,In_281,In_1634);
xnor U47 (N_47,In_2160,In_991);
nand U48 (N_48,In_2319,In_316);
nor U49 (N_49,In_1017,In_1495);
or U50 (N_50,In_486,In_1413);
nor U51 (N_51,In_1762,In_570);
nor U52 (N_52,In_275,In_1609);
and U53 (N_53,In_950,In_1870);
or U54 (N_54,In_1306,In_1523);
and U55 (N_55,In_1716,In_1351);
or U56 (N_56,In_507,In_1819);
or U57 (N_57,In_1143,In_971);
or U58 (N_58,In_415,In_2074);
or U59 (N_59,In_2496,In_675);
xnor U60 (N_60,In_1845,In_1563);
and U61 (N_61,In_201,In_2337);
or U62 (N_62,In_876,In_2050);
nor U63 (N_63,In_537,In_55);
nor U64 (N_64,In_864,In_988);
nand U65 (N_65,In_280,In_390);
or U66 (N_66,In_1452,In_2100);
nor U67 (N_67,In_2121,In_1948);
nor U68 (N_68,In_2381,In_1060);
xnor U69 (N_69,In_2352,In_1188);
or U70 (N_70,In_1273,In_1920);
nand U71 (N_71,In_1408,In_364);
or U72 (N_72,In_2322,In_761);
xor U73 (N_73,In_1337,In_2029);
nor U74 (N_74,In_138,In_77);
nor U75 (N_75,In_2139,In_480);
nand U76 (N_76,In_722,In_899);
xor U77 (N_77,In_856,In_1965);
nor U78 (N_78,In_660,In_1685);
nor U79 (N_79,In_1750,In_2358);
nand U80 (N_80,In_1836,In_756);
or U81 (N_81,In_1735,In_1902);
xor U82 (N_82,In_1772,In_2188);
and U83 (N_83,In_1132,In_928);
nand U84 (N_84,In_1292,In_847);
and U85 (N_85,In_2378,In_1739);
xor U86 (N_86,In_749,In_1451);
or U87 (N_87,In_2264,In_1142);
xor U88 (N_88,In_438,In_1420);
xor U89 (N_89,In_313,In_1256);
nor U90 (N_90,In_2442,In_2141);
nand U91 (N_91,In_2349,In_230);
or U92 (N_92,In_808,In_1215);
nand U93 (N_93,In_49,In_1339);
or U94 (N_94,In_1532,In_1194);
and U95 (N_95,In_447,In_1347);
nand U96 (N_96,In_229,In_2189);
or U97 (N_97,In_397,In_937);
or U98 (N_98,In_1521,In_545);
and U99 (N_99,In_8,In_1624);
and U100 (N_100,In_330,In_1348);
and U101 (N_101,In_1258,In_1906);
or U102 (N_102,In_1001,In_952);
or U103 (N_103,In_1697,In_2048);
nand U104 (N_104,In_2069,In_2382);
or U105 (N_105,In_1049,In_1155);
or U106 (N_106,In_1140,In_895);
and U107 (N_107,In_1741,In_86);
xor U108 (N_108,In_2394,In_643);
or U109 (N_109,In_2476,In_44);
nor U110 (N_110,In_287,In_1120);
and U111 (N_111,In_2208,In_813);
nor U112 (N_112,In_737,In_2302);
nor U113 (N_113,In_1326,In_2392);
nand U114 (N_114,In_48,In_2178);
nand U115 (N_115,In_2343,In_594);
xnor U116 (N_116,In_1918,In_944);
nand U117 (N_117,In_852,In_263);
nor U118 (N_118,In_1933,In_1874);
and U119 (N_119,In_786,In_1176);
nor U120 (N_120,In_787,In_1193);
nand U121 (N_121,In_2391,In_894);
nand U122 (N_122,In_1813,In_1529);
or U123 (N_123,In_243,In_2180);
xor U124 (N_124,In_1240,In_2300);
or U125 (N_125,In_1296,In_1898);
nand U126 (N_126,In_1821,In_1357);
nand U127 (N_127,In_2197,In_1630);
or U128 (N_128,In_341,In_593);
nand U129 (N_129,In_2195,In_1071);
nor U130 (N_130,In_543,In_1222);
and U131 (N_131,In_1514,In_2078);
or U132 (N_132,In_2176,In_1656);
nor U133 (N_133,In_785,In_491);
xor U134 (N_134,In_106,In_191);
or U135 (N_135,In_652,In_166);
xor U136 (N_136,In_994,In_1148);
nand U137 (N_137,In_1710,In_412);
or U138 (N_138,In_202,In_1007);
xor U139 (N_139,In_753,In_423);
nand U140 (N_140,In_884,In_38);
or U141 (N_141,In_696,In_2444);
or U142 (N_142,In_354,In_1573);
or U143 (N_143,In_861,In_2292);
xnor U144 (N_144,In_2452,In_613);
or U145 (N_145,In_1065,In_765);
or U146 (N_146,In_850,In_1009);
nand U147 (N_147,In_139,In_160);
or U148 (N_148,In_87,In_1253);
nand U149 (N_149,In_81,In_2310);
xor U150 (N_150,In_1700,In_2179);
or U151 (N_151,In_1914,In_1012);
nor U152 (N_152,In_1552,In_2018);
nand U153 (N_153,In_2276,In_1338);
or U154 (N_154,In_359,In_1225);
nor U155 (N_155,In_1779,In_755);
or U156 (N_156,In_1738,In_1928);
nand U157 (N_157,In_1878,In_1982);
nand U158 (N_158,In_2341,In_783);
xnor U159 (N_159,In_121,In_1719);
xnor U160 (N_160,In_169,In_274);
nand U161 (N_161,In_2022,In_554);
nor U162 (N_162,In_1542,In_1803);
xnor U163 (N_163,In_347,In_496);
and U164 (N_164,In_499,In_1355);
nand U165 (N_165,In_1156,In_1592);
nand U166 (N_166,In_1454,In_2446);
nand U167 (N_167,In_1620,In_816);
nand U168 (N_168,In_1736,In_1519);
nor U169 (N_169,In_705,In_2130);
nand U170 (N_170,In_297,In_1608);
and U171 (N_171,In_493,In_1987);
xor U172 (N_172,In_2093,In_2136);
and U173 (N_173,In_1418,In_1033);
or U174 (N_174,In_2203,In_107);
and U175 (N_175,In_2303,In_124);
xor U176 (N_176,In_2207,In_1770);
nor U177 (N_177,In_1254,In_1707);
or U178 (N_178,In_964,In_1834);
nand U179 (N_179,In_1056,In_2320);
xor U180 (N_180,In_271,In_807);
nand U181 (N_181,In_2413,In_987);
nor U182 (N_182,In_739,In_1767);
or U183 (N_183,In_222,In_383);
nor U184 (N_184,In_1020,In_1476);
and U185 (N_185,In_1379,In_918);
nand U186 (N_186,In_1714,In_597);
nand U187 (N_187,In_1513,In_2417);
and U188 (N_188,In_830,In_2110);
nand U189 (N_189,In_814,In_79);
xor U190 (N_190,In_110,In_1782);
nand U191 (N_191,In_1016,In_2196);
or U192 (N_192,In_2487,In_118);
or U193 (N_193,In_2479,In_1212);
nand U194 (N_194,In_420,In_310);
or U195 (N_195,In_978,In_245);
nor U196 (N_196,In_621,In_395);
nand U197 (N_197,In_1249,In_2247);
nand U198 (N_198,In_2367,In_1875);
xor U199 (N_199,In_936,In_2223);
nand U200 (N_200,In_1080,In_798);
and U201 (N_201,In_2012,In_1124);
nor U202 (N_202,In_630,In_773);
and U203 (N_203,In_172,In_687);
nand U204 (N_204,In_780,In_815);
xnor U205 (N_205,In_508,In_424);
nand U206 (N_206,In_2166,In_302);
xnor U207 (N_207,In_535,In_1187);
xor U208 (N_208,In_1548,In_2281);
nor U209 (N_209,In_827,In_150);
and U210 (N_210,In_91,In_1239);
nor U211 (N_211,In_1761,In_1209);
nand U212 (N_212,In_2017,In_1462);
and U213 (N_213,In_1810,In_285);
xnor U214 (N_214,In_1863,In_1531);
and U215 (N_215,In_2266,In_812);
xor U216 (N_216,In_1121,In_2256);
and U217 (N_217,In_2084,In_154);
nand U218 (N_218,In_1891,In_1516);
nand U219 (N_219,In_1236,In_880);
nand U220 (N_220,In_1035,In_902);
xnor U221 (N_221,In_299,In_1076);
and U222 (N_222,In_209,In_1565);
nand U223 (N_223,In_130,In_214);
nor U224 (N_224,In_718,In_671);
xnor U225 (N_225,In_2328,In_41);
nand U226 (N_226,In_1733,In_1997);
nand U227 (N_227,In_2422,In_972);
nor U228 (N_228,In_1399,In_2355);
nor U229 (N_229,In_674,In_1151);
or U230 (N_230,In_1655,In_1089);
nor U231 (N_231,In_1108,In_1594);
xnor U232 (N_232,In_1090,In_269);
and U233 (N_233,In_1667,In_1876);
nand U234 (N_234,In_410,In_519);
xnor U235 (N_235,In_1045,In_362);
nand U236 (N_236,In_1536,In_2014);
or U237 (N_237,In_1680,In_1031);
and U238 (N_238,In_392,In_2370);
and U239 (N_239,In_1104,In_1547);
and U240 (N_240,In_2152,In_1072);
and U241 (N_241,In_1162,In_261);
or U242 (N_242,In_834,In_497);
xor U243 (N_243,In_350,In_1590);
or U244 (N_244,In_1449,In_2268);
and U245 (N_245,In_1577,In_1947);
nor U246 (N_246,In_1260,In_1062);
and U247 (N_247,In_1383,In_58);
xor U248 (N_248,In_1722,In_2272);
or U249 (N_249,In_1358,In_2306);
nor U250 (N_250,In_896,In_2026);
nand U251 (N_251,In_1091,In_1843);
or U252 (N_252,In_1402,In_1558);
and U253 (N_253,In_2257,In_2395);
xor U254 (N_254,In_709,In_963);
and U255 (N_255,In_958,N_75);
xor U256 (N_256,In_679,In_1423);
xnor U257 (N_257,In_975,In_26);
or U258 (N_258,In_1028,In_1956);
nand U259 (N_259,In_458,In_940);
nor U260 (N_260,N_156,In_851);
xor U261 (N_261,In_1393,In_1695);
and U262 (N_262,In_1665,In_2144);
and U263 (N_263,N_91,In_2153);
nor U264 (N_264,In_733,In_1864);
or U265 (N_265,In_1293,In_247);
xor U266 (N_266,In_1786,N_201);
xnor U267 (N_267,In_1734,In_1061);
nor U268 (N_268,In_970,In_1311);
nor U269 (N_269,In_1973,In_2353);
and U270 (N_270,In_1745,In_73);
nor U271 (N_271,In_581,N_207);
nand U272 (N_272,In_1456,In_826);
or U273 (N_273,In_859,In_2478);
nor U274 (N_274,In_112,In_1468);
xnor U275 (N_275,In_1923,In_113);
and U276 (N_276,In_295,In_1527);
xnor U277 (N_277,In_1400,In_463);
nand U278 (N_278,In_2471,In_211);
xor U279 (N_279,In_2222,In_1972);
nand U280 (N_280,In_158,In_1959);
nand U281 (N_281,In_1998,In_2046);
nor U282 (N_282,In_587,In_1627);
nand U283 (N_283,In_1520,In_1429);
nor U284 (N_284,In_1650,In_1838);
nand U285 (N_285,In_734,In_1753);
xnor U286 (N_286,In_920,In_1158);
xnor U287 (N_287,In_373,In_1578);
nor U288 (N_288,In_1818,In_1751);
or U289 (N_289,In_2194,In_1599);
nor U290 (N_290,In_1335,In_1300);
xnor U291 (N_291,In_2102,In_221);
nor U292 (N_292,In_1244,In_555);
nor U293 (N_293,In_1967,In_82);
nand U294 (N_294,N_180,In_2275);
or U295 (N_295,In_1006,In_664);
nand U296 (N_296,In_715,In_1833);
xor U297 (N_297,In_1191,In_2072);
or U298 (N_298,In_288,In_673);
and U299 (N_299,N_160,In_1534);
xnor U300 (N_300,In_939,In_695);
nand U301 (N_301,In_418,In_968);
xnor U302 (N_302,In_665,In_1471);
nor U303 (N_303,In_682,In_1201);
nor U304 (N_304,In_1078,In_102);
nor U305 (N_305,In_71,N_30);
and U306 (N_306,In_1961,In_2056);
xnor U307 (N_307,In_2165,In_1098);
and U308 (N_308,In_2229,In_572);
nor U309 (N_309,In_452,In_1999);
and U310 (N_310,In_1276,In_1904);
nand U311 (N_311,In_534,In_513);
or U312 (N_312,In_1605,In_2067);
or U313 (N_313,In_1952,In_1795);
and U314 (N_314,In_460,In_132);
nand U315 (N_315,In_721,In_1231);
nand U316 (N_316,In_345,In_2339);
xor U317 (N_317,In_2334,In_1086);
xnor U318 (N_318,In_1678,In_2285);
nand U319 (N_319,In_1224,In_2435);
or U320 (N_320,In_672,In_1628);
xor U321 (N_321,N_136,In_942);
nor U322 (N_322,In_1882,In_547);
xnor U323 (N_323,In_2250,In_1286);
or U324 (N_324,In_490,In_925);
nand U325 (N_325,In_738,In_1549);
nor U326 (N_326,N_104,In_1032);
xnor U327 (N_327,In_1217,In_459);
or U328 (N_328,In_680,In_1905);
or U329 (N_329,In_1406,In_1903);
nand U330 (N_330,In_2145,In_2364);
or U331 (N_331,In_436,In_259);
or U332 (N_332,In_1629,N_190);
xnor U333 (N_333,N_196,N_177);
and U334 (N_334,In_2255,In_2430);
nor U335 (N_335,N_24,In_1820);
or U336 (N_336,In_2298,In_1546);
nor U337 (N_337,In_967,In_368);
or U338 (N_338,In_277,In_916);
and U339 (N_339,N_152,In_2488);
nor U340 (N_340,In_254,In_1152);
nor U341 (N_341,In_2201,In_366);
or U342 (N_342,N_114,In_1617);
nand U343 (N_343,In_292,In_111);
nor U344 (N_344,In_203,In_589);
and U345 (N_345,In_1178,In_772);
nand U346 (N_346,In_1434,In_1912);
xnor U347 (N_347,In_2260,In_1291);
and U348 (N_348,In_1030,N_170);
xnor U349 (N_349,In_1499,In_2015);
nor U350 (N_350,In_348,In_1689);
xor U351 (N_351,In_1352,In_1789);
xor U352 (N_352,In_1374,In_1910);
nor U353 (N_353,N_172,In_1704);
and U354 (N_354,N_225,In_2384);
xnor U355 (N_355,In_1248,In_1283);
or U356 (N_356,In_809,In_741);
xor U357 (N_357,In_2027,In_784);
nor U358 (N_358,In_1669,In_699);
nand U359 (N_359,In_2467,In_1146);
nand U360 (N_360,In_114,In_335);
or U361 (N_361,In_1332,In_462);
nor U362 (N_362,In_552,In_2405);
and U363 (N_363,In_320,N_4);
nand U364 (N_364,N_203,In_540);
xnor U365 (N_365,In_2385,In_1058);
nor U366 (N_366,In_912,In_1356);
nand U367 (N_367,In_2315,In_367);
xnor U368 (N_368,In_1488,In_36);
nand U369 (N_369,In_1709,In_1614);
xor U370 (N_370,In_290,In_878);
or U371 (N_371,In_1389,N_44);
and U372 (N_372,In_1189,In_2082);
and U373 (N_373,In_913,In_601);
xnor U374 (N_374,In_1341,In_1953);
nand U375 (N_375,In_1443,In_1315);
nand U376 (N_376,In_1437,N_1);
and U377 (N_377,In_2108,In_42);
or U378 (N_378,In_1302,In_223);
or U379 (N_379,In_21,In_2170);
xor U380 (N_380,In_2297,In_276);
xnor U381 (N_381,In_1472,In_1498);
nand U382 (N_382,In_833,In_871);
nor U383 (N_383,In_560,In_678);
nor U384 (N_384,In_1583,In_2473);
or U385 (N_385,In_1872,In_874);
nand U386 (N_386,In_1721,In_2374);
xor U387 (N_387,N_189,In_1359);
nand U388 (N_388,In_161,In_1190);
or U389 (N_389,In_88,In_1633);
nor U390 (N_390,In_760,In_1464);
and U391 (N_391,In_1482,In_1053);
nor U392 (N_392,In_2482,In_1003);
nor U393 (N_393,In_580,In_385);
or U394 (N_394,In_1993,In_1981);
nor U395 (N_395,N_18,In_1388);
nor U396 (N_396,In_2323,In_2184);
or U397 (N_397,In_1699,In_1074);
nor U398 (N_398,In_576,In_54);
nand U399 (N_399,In_2049,In_1539);
nor U400 (N_400,N_58,In_1705);
and U401 (N_401,In_401,In_2494);
nor U402 (N_402,In_1417,In_2010);
nor U403 (N_403,N_223,In_2149);
or U404 (N_404,N_92,In_322);
nand U405 (N_405,In_1175,In_657);
nor U406 (N_406,In_866,In_2286);
xor U407 (N_407,In_1307,N_41);
nand U408 (N_408,In_1600,In_1641);
nand U409 (N_409,In_1963,In_2044);
or U410 (N_410,In_1112,In_1823);
nor U411 (N_411,In_1892,N_240);
xor U412 (N_412,N_173,In_109);
nand U413 (N_413,In_2090,In_1483);
nand U414 (N_414,In_2282,In_2345);
nor U415 (N_415,N_31,N_205);
and U416 (N_416,N_0,In_710);
or U417 (N_417,N_118,In_2025);
or U418 (N_418,In_1899,In_591);
nand U419 (N_419,In_1501,In_1005);
nor U420 (N_420,In_575,In_1346);
xnor U421 (N_421,In_855,In_2486);
nor U422 (N_422,In_1202,N_80);
nor U423 (N_423,In_437,In_2340);
nand U424 (N_424,In_23,In_2347);
and U425 (N_425,In_1343,N_234);
nor U426 (N_426,In_1491,In_2344);
or U427 (N_427,In_1131,In_1754);
or U428 (N_428,In_2037,In_2342);
nand U429 (N_429,In_1092,N_134);
or U430 (N_430,N_56,In_2371);
xor U431 (N_431,In_2036,In_638);
xor U432 (N_432,In_19,In_1512);
and U433 (N_433,In_2380,In_1869);
xnor U434 (N_434,In_569,In_308);
or U435 (N_435,In_1668,In_1208);
nand U436 (N_436,In_2104,In_1756);
nor U437 (N_437,In_1432,In_1002);
nor U438 (N_438,In_2398,In_104);
xnor U439 (N_439,In_1852,In_2277);
nor U440 (N_440,In_1730,In_1136);
nand U441 (N_441,N_88,In_1584);
nand U442 (N_442,In_441,In_2267);
xnor U443 (N_443,In_2311,In_860);
xnor U444 (N_444,In_488,In_2457);
nand U445 (N_445,In_1141,In_2428);
xor U446 (N_446,In_1824,In_1220);
or U447 (N_447,In_1281,N_16);
xnor U448 (N_448,N_9,In_1846);
nor U449 (N_449,In_1455,In_477);
or U450 (N_450,In_1197,In_697);
nand U451 (N_451,In_1144,In_1944);
nor U452 (N_452,In_2312,In_771);
and U453 (N_453,In_242,In_841);
and U454 (N_454,N_148,In_1069);
nand U455 (N_455,In_2226,In_623);
xnor U456 (N_456,In_1647,In_1114);
nor U457 (N_457,In_1368,In_740);
xnor U458 (N_458,N_49,In_283);
nor U459 (N_459,In_328,In_533);
xnor U460 (N_460,In_2237,In_2138);
nor U461 (N_461,In_100,In_1740);
nand U462 (N_462,In_571,In_1744);
xor U463 (N_463,In_1257,In_1507);
or U464 (N_464,In_228,In_1635);
nor U465 (N_465,In_2220,In_241);
nand U466 (N_466,In_754,In_1849);
or U467 (N_467,In_2273,In_2363);
nor U468 (N_468,In_311,In_911);
xor U469 (N_469,In_1595,In_175);
xnor U470 (N_470,In_1545,In_382);
xor U471 (N_471,In_1211,In_521);
xor U472 (N_472,In_1572,In_1977);
nor U473 (N_473,N_208,In_193);
or U474 (N_474,In_618,In_344);
and U475 (N_475,In_1497,In_1232);
nand U476 (N_476,N_121,In_1980);
and U477 (N_477,In_207,In_2333);
and U478 (N_478,In_2451,In_51);
or U479 (N_479,In_658,In_237);
and U480 (N_480,In_1662,In_1781);
and U481 (N_481,In_1792,In_470);
nor U482 (N_482,N_210,In_2495);
and U483 (N_483,In_1990,In_2239);
nand U484 (N_484,In_1796,In_1067);
xnor U485 (N_485,In_946,In_1791);
and U486 (N_486,In_1113,In_649);
or U487 (N_487,In_2271,In_1459);
and U488 (N_488,N_10,In_986);
nor U489 (N_489,In_1177,In_596);
nor U490 (N_490,In_2115,In_1469);
xnor U491 (N_491,In_1702,In_732);
nand U492 (N_492,In_1123,In_333);
or U493 (N_493,In_1252,In_2175);
xor U494 (N_494,In_2313,In_1496);
nand U495 (N_495,In_2023,In_1262);
xor U496 (N_496,In_1672,N_98);
xnor U497 (N_497,In_380,In_1706);
nor U498 (N_498,In_1757,In_1227);
nor U499 (N_499,In_1289,In_2142);
xnor U500 (N_500,N_157,In_2419);
nand U501 (N_501,In_1732,In_563);
nand U502 (N_502,In_1317,In_1510);
and U503 (N_503,In_762,N_119);
xor U504 (N_504,In_1385,In_2489);
xnor U505 (N_505,In_1242,In_1461);
or U506 (N_506,In_2007,In_352);
xnor U507 (N_507,N_374,In_182);
xnor U508 (N_508,N_200,In_1556);
nor U509 (N_509,In_2096,N_341);
or U510 (N_510,In_406,In_2172);
xnor U511 (N_511,In_1942,In_2061);
nor U512 (N_512,N_237,In_1099);
nor U513 (N_513,N_452,In_1908);
nand U514 (N_514,In_67,In_1107);
or U515 (N_515,In_28,In_962);
xnor U516 (N_516,N_451,In_1036);
xor U517 (N_517,N_378,In_2021);
and U518 (N_518,In_1743,In_1640);
or U519 (N_519,In_666,In_727);
xor U520 (N_520,In_472,In_751);
nor U521 (N_521,N_425,In_1083);
or U522 (N_522,In_1128,In_1660);
nor U523 (N_523,In_481,In_2377);
nand U524 (N_524,In_1159,In_2134);
or U525 (N_525,In_1487,N_391);
xnor U526 (N_526,In_2006,N_11);
nor U527 (N_527,N_274,N_140);
nand U528 (N_528,In_1237,N_97);
and U529 (N_529,In_719,N_473);
nor U530 (N_530,N_79,In_1873);
or U531 (N_531,In_1611,In_1686);
nor U532 (N_532,In_1830,In_566);
xnor U533 (N_533,In_2307,In_231);
nor U534 (N_534,In_1364,In_249);
xor U535 (N_535,In_2293,In_2402);
nor U536 (N_536,In_1580,In_2461);
and U537 (N_537,In_1251,In_1204);
nor U538 (N_538,In_1426,In_872);
xnor U539 (N_539,In_1777,N_213);
nor U540 (N_540,In_178,In_965);
and U541 (N_541,In_1439,In_1427);
or U542 (N_542,In_1460,In_1788);
nor U543 (N_543,In_1897,In_1784);
or U544 (N_544,In_1925,In_1199);
or U545 (N_545,N_112,In_1992);
or U546 (N_546,In_1149,In_1206);
and U547 (N_547,In_922,N_310);
or U548 (N_548,N_366,In_1715);
and U549 (N_549,N_212,In_1862);
and U550 (N_550,In_1305,In_2284);
nand U551 (N_551,In_1935,N_246);
nand U552 (N_552,N_306,In_2098);
or U553 (N_553,In_1771,In_484);
xor U554 (N_554,N_47,N_247);
xnor U555 (N_555,N_166,N_286);
nand U556 (N_556,N_17,In_2243);
and U557 (N_557,In_2232,N_52);
xnor U558 (N_558,In_89,In_1118);
or U559 (N_559,In_479,In_1941);
nand U560 (N_560,In_1749,N_192);
or U561 (N_561,N_403,In_900);
nand U562 (N_562,In_234,N_411);
xnor U563 (N_563,In_1991,N_328);
xnor U564 (N_564,In_2087,In_2173);
and U565 (N_565,In_1748,In_59);
xor U566 (N_566,In_2214,In_993);
nor U567 (N_567,In_2458,In_1737);
and U568 (N_568,In_1787,In_9);
nand U569 (N_569,In_40,N_362);
nand U570 (N_570,In_69,In_1453);
or U571 (N_571,In_128,In_2064);
nand U572 (N_572,In_747,In_1485);
or U573 (N_573,In_1154,In_2350);
and U574 (N_574,In_2369,In_731);
or U575 (N_575,In_1111,In_386);
or U576 (N_576,In_548,In_953);
and U577 (N_577,In_1226,N_340);
nand U578 (N_578,In_1566,N_355);
or U579 (N_579,N_493,In_251);
and U580 (N_580,In_63,In_2089);
nor U581 (N_581,In_842,In_2071);
nand U582 (N_582,In_421,N_399);
and U583 (N_583,In_2008,In_917);
or U584 (N_584,In_485,In_1570);
and U585 (N_585,In_1890,N_272);
xor U586 (N_586,In_1533,In_1809);
and U587 (N_587,In_849,In_1047);
xnor U588 (N_588,In_2301,In_1975);
nor U589 (N_589,In_1394,In_2101);
and U590 (N_590,In_1994,In_883);
or U591 (N_591,In_1681,In_1085);
xnor U592 (N_592,In_1860,N_113);
xnor U593 (N_593,In_353,In_162);
nor U594 (N_594,N_143,N_326);
nor U595 (N_595,In_2356,In_518);
and U596 (N_596,In_2414,In_30);
xor U597 (N_597,In_233,In_232);
nand U598 (N_598,In_4,In_157);
or U599 (N_599,N_316,N_431);
nor U600 (N_600,In_1538,N_158);
xor U601 (N_601,In_973,In_85);
nor U602 (N_602,In_2424,In_615);
nor U603 (N_603,In_177,N_266);
and U604 (N_604,In_901,In_1448);
or U605 (N_605,N_164,In_1932);
xor U606 (N_606,N_490,In_1901);
xor U607 (N_607,In_1806,In_1511);
xnor U608 (N_608,N_12,N_99);
nor U609 (N_609,In_1692,N_314);
and U610 (N_610,In_204,In_2183);
xnor U611 (N_611,In_585,N_171);
xnor U612 (N_612,In_351,In_256);
nor U613 (N_613,In_1591,In_1278);
or U614 (N_614,In_1802,In_167);
and U615 (N_615,N_381,In_1841);
xor U616 (N_616,N_255,N_321);
or U617 (N_617,In_417,In_538);
or U618 (N_618,N_393,N_462);
and U619 (N_619,N_131,In_1517);
or U620 (N_620,N_179,In_1391);
nand U621 (N_621,In_1308,In_123);
nand U622 (N_622,In_1164,In_938);
xnor U623 (N_623,In_45,In_1909);
nand U624 (N_624,In_2146,In_494);
or U625 (N_625,N_108,In_2287);
or U626 (N_626,N_69,In_305);
xnor U627 (N_627,In_1015,N_3);
or U628 (N_628,In_255,In_1569);
xor U629 (N_629,In_2338,In_736);
or U630 (N_630,In_464,N_468);
or U631 (N_631,In_337,N_147);
or U632 (N_632,In_2147,In_1314);
nor U633 (N_633,In_474,In_1275);
or U634 (N_634,In_2278,N_402);
or U635 (N_635,In_1250,In_2456);
or U636 (N_636,In_189,In_2474);
nand U637 (N_637,In_966,In_2198);
nor U638 (N_638,In_1318,In_1951);
nand U639 (N_639,N_139,In_434);
nand U640 (N_640,In_1334,N_351);
or U641 (N_641,In_924,In_1798);
nand U642 (N_642,In_206,In_1342);
nand U643 (N_643,In_2477,In_642);
or U644 (N_644,In_2070,In_1983);
nand U645 (N_645,N_342,N_299);
and U646 (N_646,In_1814,In_164);
and U647 (N_647,In_1822,In_1857);
nand U648 (N_648,In_306,In_655);
or U649 (N_649,In_1481,In_802);
or U650 (N_650,In_1117,In_843);
xor U651 (N_651,In_2455,In_2217);
xor U652 (N_652,In_606,N_35);
nand U653 (N_653,In_2033,In_194);
xor U654 (N_654,In_365,In_600);
nor U655 (N_655,N_400,In_1631);
or U656 (N_656,In_465,In_1267);
xnor U657 (N_657,In_550,In_473);
and U658 (N_658,In_592,N_27);
and U659 (N_659,In_1200,In_2321);
nand U660 (N_660,In_869,In_831);
nor U661 (N_661,In_1747,N_232);
nand U662 (N_662,In_527,In_1027);
or U663 (N_663,In_151,In_183);
xor U664 (N_664,In_1422,N_423);
xnor U665 (N_665,In_1502,N_392);
or U666 (N_666,In_1052,In_147);
or U667 (N_667,In_1717,In_1970);
and U668 (N_668,N_494,N_243);
nor U669 (N_669,N_467,In_1405);
nor U670 (N_670,In_610,In_1038);
or U671 (N_671,In_744,In_2234);
nor U672 (N_672,N_453,In_1153);
or U673 (N_673,In_768,In_577);
or U674 (N_674,N_22,In_1598);
and U675 (N_675,In_1198,N_256);
nand U676 (N_676,In_2081,In_957);
xnor U677 (N_677,N_318,In_886);
xor U678 (N_678,In_2410,N_464);
nand U679 (N_679,N_487,In_2236);
and U680 (N_680,In_405,In_717);
nand U681 (N_681,In_1589,In_1518);
nor U682 (N_682,N_382,In_2140);
nand U683 (N_683,In_1412,In_94);
nand U684 (N_684,In_141,N_73);
nand U685 (N_685,In_294,N_449);
and U686 (N_686,In_304,In_120);
nor U687 (N_687,N_277,N_436);
nand U688 (N_688,In_1082,In_64);
and U689 (N_689,In_1588,In_2028);
and U690 (N_690,In_2427,In_530);
and U691 (N_691,In_948,In_805);
and U692 (N_692,N_168,In_2043);
nor U693 (N_693,In_1720,In_2167);
xor U694 (N_694,In_215,In_1900);
nand U695 (N_695,In_456,In_1515);
and U696 (N_696,In_1575,In_2244);
or U697 (N_697,N_394,In_7);
xor U698 (N_698,In_1698,In_159);
and U699 (N_699,In_1494,In_2432);
nand U700 (N_700,In_1026,N_454);
xnor U701 (N_701,N_260,In_453);
or U702 (N_702,In_1444,In_536);
and U703 (N_703,In_2274,N_275);
nand U704 (N_704,In_1827,In_1323);
or U705 (N_705,In_2304,N_458);
or U706 (N_706,N_161,In_2483);
and U707 (N_707,N_132,N_130);
nor U708 (N_708,N_339,N_373);
and U709 (N_709,In_148,In_2426);
nand U710 (N_710,In_301,N_40);
and U711 (N_711,N_276,N_202);
and U712 (N_712,In_979,N_477);
or U713 (N_713,In_52,In_2128);
nand U714 (N_714,In_265,N_224);
or U715 (N_715,In_716,In_804);
or U716 (N_716,In_1157,In_956);
and U717 (N_717,N_43,In_1486);
nand U718 (N_718,N_417,In_6);
nand U719 (N_719,N_67,In_2042);
nand U720 (N_720,In_504,N_174);
nand U721 (N_721,In_210,In_1182);
nand U722 (N_722,N_144,In_1025);
nand U723 (N_723,In_1509,In_2155);
nand U724 (N_724,In_790,In_1245);
and U725 (N_725,In_2498,In_1350);
or U726 (N_726,N_48,In_1430);
and U727 (N_727,In_1057,In_309);
nor U728 (N_728,In_2120,N_499);
nand U729 (N_729,In_33,In_2094);
xor U730 (N_730,In_662,N_450);
nor U731 (N_731,In_1713,In_857);
nand U732 (N_732,In_31,In_2492);
nor U733 (N_733,In_1327,N_288);
or U734 (N_734,In_1995,N_74);
nor U735 (N_735,In_2468,In_801);
and U736 (N_736,In_404,In_983);
or U737 (N_737,In_1138,In_757);
and U738 (N_738,In_1329,In_1435);
or U739 (N_739,In_1653,In_2045);
nor U740 (N_740,In_2168,In_2365);
or U741 (N_741,In_639,In_1557);
nor U742 (N_742,In_286,N_145);
xor U743 (N_743,In_604,In_2433);
or U744 (N_744,In_1223,N_386);
and U745 (N_745,N_109,In_1186);
nand U746 (N_746,In_116,In_1850);
or U747 (N_747,In_605,In_1560);
and U748 (N_748,In_1978,N_182);
nand U749 (N_749,In_764,In_2289);
and U750 (N_750,In_890,In_1938);
and U751 (N_751,In_326,In_445);
and U752 (N_752,N_267,N_688);
nand U753 (N_753,N_418,In_562);
or U754 (N_754,In_1247,N_740);
or U755 (N_755,N_501,N_239);
or U756 (N_756,In_476,In_1492);
or U757 (N_757,In_945,In_1382);
and U758 (N_758,N_691,In_2469);
and U759 (N_759,N_549,In_1103);
and U760 (N_760,In_457,N_509);
or U761 (N_761,In_1416,N_258);
and U762 (N_762,N_422,In_1812);
or U763 (N_763,N_154,In_239);
xor U764 (N_764,In_2125,In_2251);
xor U765 (N_765,In_1029,N_347);
nand U766 (N_766,In_1645,In_848);
nand U767 (N_767,N_345,N_405);
xnor U768 (N_768,In_2454,N_714);
nor U769 (N_769,In_1506,In_769);
nor U770 (N_770,In_670,In_1116);
and U771 (N_771,N_481,N_187);
nor U772 (N_772,In_1039,N_741);
xnor U773 (N_773,N_331,In_1303);
nand U774 (N_774,In_1213,In_1299);
or U775 (N_775,In_837,In_2035);
xnor U776 (N_776,In_1203,In_218);
xnor U777 (N_777,N_638,In_517);
nand U778 (N_778,N_33,In_74);
and U779 (N_779,In_609,In_117);
nor U780 (N_780,In_1181,In_2412);
nor U781 (N_781,In_2218,N_59);
nor U782 (N_782,In_1133,N_653);
or U783 (N_783,In_403,N_435);
nor U784 (N_784,In_146,N_229);
xor U785 (N_785,N_544,In_1800);
nor U786 (N_786,In_399,In_278);
and U787 (N_787,N_732,In_1279);
and U788 (N_788,In_980,N_36);
nor U789 (N_789,In_266,In_692);
nand U790 (N_790,N_427,In_57);
and U791 (N_791,In_730,In_1625);
nor U792 (N_792,N_311,N_528);
and U793 (N_793,In_541,In_1018);
xor U794 (N_794,In_2124,In_2114);
xnor U795 (N_795,N_543,In_1969);
nand U796 (N_796,In_407,In_419);
nand U797 (N_797,In_378,In_746);
and U798 (N_798,In_645,N_547);
and U799 (N_799,In_525,In_2441);
nand U800 (N_800,N_244,In_2443);
xor U801 (N_801,In_1989,In_1054);
xnor U802 (N_802,In_1433,N_517);
and U803 (N_803,In_1671,In_1503);
nand U804 (N_804,N_619,In_334);
or U805 (N_805,In_1331,N_372);
xor U806 (N_806,In_2485,In_2253);
and U807 (N_807,N_410,N_39);
or U808 (N_808,In_2493,In_1478);
xor U809 (N_809,N_536,N_669);
xnor U810 (N_810,N_293,N_644);
xnor U811 (N_811,N_261,In_2409);
and U812 (N_812,In_1541,N_78);
or U813 (N_813,In_1214,N_568);
and U814 (N_814,In_954,N_424);
and U815 (N_815,In_1372,N_383);
nand U816 (N_816,N_730,In_2418);
nor U817 (N_817,In_1233,In_2366);
nand U818 (N_818,In_1855,In_1270);
nand U819 (N_819,In_1917,In_388);
nor U820 (N_820,N_61,In_1934);
nor U821 (N_821,N_279,In_1839);
and U822 (N_822,In_941,In_1263);
and U823 (N_823,In_1390,In_1369);
and U824 (N_824,In_224,In_2294);
or U825 (N_825,In_1438,In_1937);
xnor U826 (N_826,In_1664,In_2156);
xor U827 (N_827,In_2215,In_2295);
or U828 (N_828,In_1137,N_265);
nand U829 (N_829,N_287,In_2460);
and U830 (N_830,In_2054,N_106);
and U831 (N_831,In_929,In_500);
nor U832 (N_832,N_656,N_657);
xnor U833 (N_833,In_510,In_1550);
or U834 (N_834,In_1893,In_844);
or U835 (N_835,In_1219,N_515);
or U836 (N_836,N_336,In_574);
or U837 (N_837,N_483,In_694);
nand U838 (N_838,In_2265,In_904);
nor U839 (N_839,In_923,In_142);
nor U840 (N_840,N_505,In_384);
nor U841 (N_841,N_550,N_330);
and U842 (N_842,In_2032,In_626);
and U843 (N_843,In_2235,In_1436);
and U844 (N_844,In_1924,In_526);
or U845 (N_845,In_2126,In_1616);
nor U846 (N_846,In_2396,In_1553);
and U847 (N_847,In_188,N_551);
nor U848 (N_848,N_15,In_1752);
nand U849 (N_849,In_1593,N_661);
and U850 (N_850,N_54,In_685);
xor U851 (N_851,N_169,In_272);
and U852 (N_852,In_1055,N_683);
and U853 (N_853,In_56,N_724);
and U854 (N_854,N_510,N_221);
or U855 (N_855,In_586,N_233);
or U856 (N_856,N_564,In_422);
nand U857 (N_857,In_1790,In_1854);
or U858 (N_858,N_262,In_1606);
xor U859 (N_859,In_882,N_28);
nor U860 (N_860,N_296,N_334);
nand U861 (N_861,In_1075,In_1105);
and U862 (N_862,In_134,In_2439);
or U863 (N_863,In_551,In_1024);
and U864 (N_864,In_959,In_1765);
nand U865 (N_865,In_845,In_92);
xnor U866 (N_866,In_825,N_472);
nor U867 (N_867,N_709,N_13);
or U868 (N_868,In_2375,In_72);
xor U869 (N_869,N_401,In_369);
nand U870 (N_870,In_777,In_1421);
xnor U871 (N_871,N_120,N_349);
nand U872 (N_872,N_292,In_346);
or U873 (N_873,N_512,N_502);
nand U874 (N_874,In_323,In_2075);
nand U875 (N_875,In_544,In_588);
or U876 (N_876,N_682,In_62);
and U877 (N_877,N_406,In_163);
nor U878 (N_878,In_284,N_664);
and U879 (N_879,N_557,N_364);
xnor U880 (N_880,N_667,In_1294);
nor U881 (N_881,In_2261,In_1868);
nor U882 (N_882,In_1703,In_240);
nand U883 (N_883,In_217,N_188);
or U884 (N_884,In_1930,N_281);
nand U885 (N_885,N_433,In_2361);
xor U886 (N_886,N_250,In_2209);
and U887 (N_887,In_1807,N_748);
xnor U888 (N_888,In_2397,In_778);
xor U889 (N_889,In_1095,In_2448);
nor U890 (N_890,N_511,In_1106);
or U891 (N_891,N_304,In_506);
nand U892 (N_892,In_2262,In_1646);
or U893 (N_893,N_589,N_398);
nand U894 (N_894,In_1829,In_1794);
or U895 (N_895,N_489,In_1102);
or U896 (N_896,In_1950,In_1309);
nand U897 (N_897,N_630,In_2205);
or U898 (N_898,In_1377,In_176);
nor U899 (N_899,In_2324,N_238);
xnor U900 (N_900,In_961,In_1643);
nand U901 (N_901,N_601,In_509);
and U902 (N_902,N_526,In_1450);
xor U903 (N_903,N_746,N_242);
nand U904 (N_904,N_722,N_445);
nor U905 (N_905,In_799,In_1371);
nand U906 (N_906,N_519,In_1879);
or U907 (N_907,N_465,In_955);
xnor U908 (N_908,N_46,In_95);
nand U909 (N_909,In_1168,In_152);
nand U910 (N_910,In_27,N_555);
and U911 (N_911,N_747,In_1817);
and U912 (N_912,In_1163,In_2270);
or U913 (N_913,In_838,N_68);
nor U914 (N_914,In_2252,In_2200);
or U915 (N_915,In_1321,In_400);
xor U916 (N_916,In_446,In_416);
xor U917 (N_917,In_1298,In_512);
or U918 (N_918,N_111,In_2230);
xnor U919 (N_919,N_325,N_598);
xnor U920 (N_920,In_1384,In_628);
or U921 (N_921,N_461,In_877);
or U922 (N_922,In_616,In_1865);
or U923 (N_923,In_1648,In_1508);
or U924 (N_924,In_885,In_1828);
xor U925 (N_925,In_794,N_470);
and U926 (N_926,N_86,N_395);
xnor U927 (N_927,In_766,In_467);
or U928 (N_928,In_515,In_854);
nor U929 (N_929,In_1216,In_726);
xnor U930 (N_930,In_676,In_264);
xnor U931 (N_931,In_84,In_1363);
xnor U932 (N_932,In_501,N_605);
or U933 (N_933,In_559,N_514);
nor U934 (N_934,In_1185,In_2053);
nor U935 (N_935,In_1125,In_216);
nand U936 (N_936,In_2088,In_568);
nor U937 (N_937,N_60,N_123);
and U938 (N_938,N_214,In_1657);
xor U939 (N_939,In_1353,N_579);
or U940 (N_940,N_358,In_2425);
nor U941 (N_941,In_2336,In_1880);
and U942 (N_942,In_2299,In_1976);
or U943 (N_943,N_642,In_2357);
nand U944 (N_944,In_2158,In_475);
or U945 (N_945,In_2030,In_1411);
or U946 (N_946,N_610,N_251);
nand U947 (N_947,N_53,In_1729);
and U948 (N_948,In_1943,In_298);
nor U949 (N_949,In_1621,N_673);
nor U950 (N_950,N_29,N_117);
nand U951 (N_951,N_652,In_868);
or U952 (N_952,In_2105,N_122);
nor U953 (N_953,In_179,In_450);
xnor U954 (N_954,In_565,In_1447);
xor U955 (N_955,In_1776,N_649);
nor U956 (N_956,In_573,N_540);
xnor U957 (N_957,In_1457,In_2400);
xor U958 (N_958,In_200,N_315);
nor U959 (N_959,In_1601,In_1964);
nor U960 (N_960,In_1130,In_1780);
nand U961 (N_961,In_2288,In_663);
nor U962 (N_962,In_131,N_631);
or U963 (N_963,N_2,In_1084);
nand U964 (N_964,N_26,N_678);
nor U965 (N_965,In_846,In_192);
xor U966 (N_966,N_126,In_1238);
nand U967 (N_967,In_2440,In_381);
and U968 (N_968,In_1725,In_524);
nor U969 (N_969,N_666,N_107);
or U970 (N_970,In_797,N_298);
nor U971 (N_971,In_1192,In_196);
xor U972 (N_972,N_63,In_1070);
or U973 (N_973,N_377,In_1856);
xnor U974 (N_974,N_85,In_1683);
xor U975 (N_975,In_461,In_478);
xnor U976 (N_976,In_46,N_459);
or U977 (N_977,N_566,N_222);
nor U978 (N_978,In_832,In_80);
xnor U979 (N_979,In_149,In_1173);
and U980 (N_980,In_440,N_181);
nand U981 (N_981,In_219,N_660);
and U982 (N_982,In_1778,In_1066);
xor U983 (N_983,N_72,N_151);
nor U984 (N_984,In_336,In_103);
or U985 (N_985,N_138,N_681);
nor U986 (N_986,In_2407,In_653);
nor U987 (N_987,In_1921,N_686);
or U988 (N_988,In_840,In_542);
nand U989 (N_989,In_1775,In_1773);
nand U990 (N_990,In_324,N_127);
xnor U991 (N_991,In_1597,In_279);
nand U992 (N_992,N_90,In_1261);
and U993 (N_993,In_1871,In_776);
xnor U994 (N_994,In_1927,In_1759);
nand U995 (N_995,In_879,In_35);
nor U996 (N_996,N_273,N_554);
nor U997 (N_997,In_823,In_1050);
or U998 (N_998,N_737,In_25);
nand U999 (N_999,N_45,In_1376);
xnor U1000 (N_1000,In_992,N_840);
nand U1001 (N_1001,In_1008,In_1473);
and U1002 (N_1002,N_482,In_1916);
nand U1003 (N_1003,In_293,In_1718);
and U1004 (N_1004,N_64,N_404);
xnor U1005 (N_1005,N_744,N_795);
nor U1006 (N_1006,In_1183,N_415);
xor U1007 (N_1007,In_2150,N_845);
and U1008 (N_1008,N_996,N_283);
nor U1009 (N_1009,N_892,In_633);
and U1010 (N_1010,In_1607,In_651);
or U1011 (N_1011,In_1755,N_198);
and U1012 (N_1012,In_98,In_108);
and U1013 (N_1013,In_1442,N_794);
or U1014 (N_1014,N_824,N_542);
xnor U1015 (N_1015,In_1769,N_115);
or U1016 (N_1016,N_284,N_186);
or U1017 (N_1017,In_2192,N_66);
and U1018 (N_1018,In_1403,In_2453);
and U1019 (N_1019,N_989,In_898);
and U1020 (N_1020,In_1381,In_607);
xor U1021 (N_1021,In_2040,In_1832);
and U1022 (N_1022,N_497,In_1723);
xor U1023 (N_1023,In_153,N_909);
xnor U1024 (N_1024,In_947,In_707);
or U1025 (N_1025,In_1974,In_1724);
and U1026 (N_1026,In_2159,In_1325);
xnor U1027 (N_1027,In_1064,In_656);
or U1028 (N_1028,In_329,In_2129);
and U1029 (N_1029,N_777,In_1465);
or U1030 (N_1030,N_885,In_1096);
xor U1031 (N_1031,N_215,N_670);
or U1032 (N_1032,N_167,In_981);
and U1033 (N_1033,In_1243,N_70);
and U1034 (N_1034,In_1285,In_595);
and U1035 (N_1035,N_324,In_523);
or U1036 (N_1036,In_1167,In_414);
nor U1037 (N_1037,N_76,In_1684);
or U1038 (N_1038,N_818,N_191);
xor U1039 (N_1039,In_2073,In_2041);
xor U1040 (N_1040,In_1345,In_2316);
xor U1041 (N_1041,In_910,In_2466);
or U1042 (N_1042,N_842,N_165);
nand U1043 (N_1043,In_140,N_954);
or U1044 (N_1044,N_853,In_659);
xnor U1045 (N_1045,In_612,In_1484);
xnor U1046 (N_1046,In_1654,In_2177);
xor U1047 (N_1047,In_448,N_721);
xor U1048 (N_1048,N_767,In_1626);
nand U1049 (N_1049,In_213,N_823);
nand U1050 (N_1050,In_1059,N_887);
or U1051 (N_1051,In_16,N_816);
or U1052 (N_1052,N_443,In_1555);
and U1053 (N_1053,N_434,N_368);
nor U1054 (N_1054,In_743,N_591);
nor U1055 (N_1055,In_2436,N_783);
or U1056 (N_1056,In_1979,In_1234);
nand U1057 (N_1057,In_1147,In_260);
and U1058 (N_1058,In_1763,In_708);
nor U1059 (N_1059,In_720,In_792);
or U1060 (N_1060,N_980,N_614);
xnor U1061 (N_1061,N_677,In_2182);
or U1062 (N_1062,In_1241,In_1021);
nand U1063 (N_1063,N_14,In_119);
and U1064 (N_1064,In_1493,In_2003);
and U1065 (N_1065,N_931,In_1885);
xor U1066 (N_1066,N_300,N_129);
and U1067 (N_1067,In_439,N_291);
nand U1068 (N_1068,N_62,N_371);
xnor U1069 (N_1069,In_1540,N_492);
xor U1070 (N_1070,In_1410,In_2132);
xnor U1071 (N_1071,In_2112,In_70);
xnor U1072 (N_1072,In_1742,In_1161);
nor U1073 (N_1073,In_1568,N_698);
and U1074 (N_1074,N_674,N_854);
and U1075 (N_1075,In_2020,N_197);
nand U1076 (N_1076,In_1373,In_469);
and U1077 (N_1077,In_2404,N_175);
nand U1078 (N_1078,In_1847,N_574);
or U1079 (N_1079,In_1883,In_489);
or U1080 (N_1080,In_1446,In_2137);
nand U1081 (N_1081,In_321,N_697);
and U1082 (N_1082,In_1543,N_982);
or U1083 (N_1083,In_2065,In_725);
or U1084 (N_1084,N_82,In_998);
nor U1085 (N_1085,N_159,In_1929);
or U1086 (N_1086,N_184,N_530);
or U1087 (N_1087,N_253,N_533);
nand U1088 (N_1088,N_877,N_622);
nand U1089 (N_1089,In_889,N_432);
and U1090 (N_1090,N_969,In_1661);
or U1091 (N_1091,N_739,In_282);
and U1092 (N_1092,N_507,N_301);
or U1093 (N_1093,N_137,In_431);
and U1094 (N_1094,N_597,In_1835);
or U1095 (N_1095,In_1889,N_966);
nor U1096 (N_1096,N_5,N_414);
xor U1097 (N_1097,In_220,In_396);
and U1098 (N_1098,N_720,N_848);
and U1099 (N_1099,In_1344,N_791);
nand U1100 (N_1100,In_2212,N_801);
nand U1101 (N_1101,In_1115,In_691);
or U1102 (N_1102,In_1160,N_624);
nand U1103 (N_1103,In_788,In_1019);
nor U1104 (N_1104,N_590,In_2111);
or U1105 (N_1105,N_940,N_934);
nor U1106 (N_1106,In_1586,N_227);
or U1107 (N_1107,In_90,In_319);
nor U1108 (N_1108,In_20,In_1658);
or U1109 (N_1109,N_430,N_476);
nand U1110 (N_1110,In_650,In_498);
nor U1111 (N_1111,N_319,In_2024);
xor U1112 (N_1112,In_1619,In_2360);
and U1113 (N_1113,In_0,N_919);
and U1114 (N_1114,N_937,N_805);
nor U1115 (N_1115,In_2429,In_977);
or U1116 (N_1116,N_596,In_1272);
nand U1117 (N_1117,In_226,In_300);
and U1118 (N_1118,N_782,In_2193);
and U1119 (N_1119,In_858,N_367);
nor U1120 (N_1120,In_408,N_929);
nand U1121 (N_1121,N_539,In_2376);
and U1122 (N_1122,In_974,In_190);
nor U1123 (N_1123,In_2401,N_305);
and U1124 (N_1124,In_1310,In_2186);
xnor U1125 (N_1125,N_663,In_262);
xnor U1126 (N_1126,N_992,N_799);
and U1127 (N_1127,In_1048,N_689);
xnor U1128 (N_1128,In_1295,In_1623);
or U1129 (N_1129,In_2415,In_398);
or U1130 (N_1130,In_315,In_2462);
nor U1131 (N_1131,N_77,N_914);
and U1132 (N_1132,In_1322,N_986);
nand U1133 (N_1133,N_380,N_755);
or U1134 (N_1134,In_1962,N_811);
nand U1135 (N_1135,In_2431,N_906);
xor U1136 (N_1136,In_137,In_2406);
and U1137 (N_1137,In_342,In_905);
nor U1138 (N_1138,In_1971,N_21);
xnor U1139 (N_1139,In_647,N_268);
xnor U1140 (N_1140,In_829,N_524);
nor U1141 (N_1141,In_133,In_53);
or U1142 (N_1142,N_859,In_1011);
and U1143 (N_1143,In_2000,In_1287);
xnor U1144 (N_1144,N_495,In_1268);
nor U1145 (N_1145,N_295,In_690);
or U1146 (N_1146,In_2122,N_508);
xnor U1147 (N_1147,In_2,N_344);
and U1148 (N_1148,N_817,N_646);
nand U1149 (N_1149,N_738,N_270);
nor U1150 (N_1150,In_1040,N_778);
xor U1151 (N_1151,In_2190,N_776);
nor U1152 (N_1152,In_582,In_101);
nand U1153 (N_1153,In_686,N_908);
xnor U1154 (N_1154,N_486,In_2238);
xnor U1155 (N_1155,N_910,N_680);
and U1156 (N_1156,In_1333,N_765);
xnor U1157 (N_1157,In_1097,In_1696);
nand U1158 (N_1158,In_83,N_559);
or U1159 (N_1159,N_608,In_1931);
nand U1160 (N_1160,In_1858,N_89);
nand U1161 (N_1161,In_97,In_425);
and U1162 (N_1162,In_943,N_650);
or U1163 (N_1163,N_729,N_572);
nand U1164 (N_1164,N_488,In_409);
nor U1165 (N_1165,N_149,In_2309);
and U1166 (N_1166,In_668,N_998);
xnor U1167 (N_1167,In_2470,In_2459);
xor U1168 (N_1168,In_1799,In_2117);
xor U1169 (N_1169,N_754,In_2143);
nor U1170 (N_1170,N_379,In_1853);
nand U1171 (N_1171,In_2151,In_893);
xnor U1172 (N_1172,N_8,In_339);
and U1173 (N_1173,N_807,In_969);
and U1174 (N_1174,In_1666,In_471);
nor U1175 (N_1175,N_926,N_142);
nor U1176 (N_1176,N_850,N_705);
xnor U1177 (N_1177,In_1419,N_333);
nand U1178 (N_1178,In_598,N_659);
nor U1179 (N_1179,N_684,In_759);
or U1180 (N_1180,In_2291,In_1109);
and U1181 (N_1181,In_371,N_907);
and U1182 (N_1182,In_1544,N_643);
nand U1183 (N_1183,N_413,In_1288);
nand U1184 (N_1184,N_951,In_1826);
xor U1185 (N_1185,In_443,In_1602);
or U1186 (N_1186,N_613,N_868);
nor U1187 (N_1187,In_1041,N_651);
and U1188 (N_1188,In_689,In_556);
and U1189 (N_1189,N_949,N_878);
xor U1190 (N_1190,In_1632,N_847);
and U1191 (N_1191,N_771,N_409);
and U1192 (N_1192,N_975,In_171);
nor U1193 (N_1193,In_2379,N_491);
nand U1194 (N_1194,N_821,In_583);
nor U1195 (N_1195,N_902,N_731);
nand U1196 (N_1196,N_569,In_1677);
and U1197 (N_1197,N_662,In_567);
xnor U1198 (N_1198,In_122,N_357);
nor U1199 (N_1199,In_1407,In_1063);
nor U1200 (N_1200,N_150,N_625);
nor U1201 (N_1201,In_669,In_539);
xor U1202 (N_1202,In_2308,N_356);
nor U1203 (N_1203,In_199,N_20);
and U1204 (N_1204,In_1825,N_105);
nand U1205 (N_1205,In_389,In_1205);
nor U1206 (N_1206,In_332,In_376);
xor U1207 (N_1207,N_585,N_984);
xor U1208 (N_1208,In_466,N_580);
nand U1209 (N_1209,In_1349,In_758);
or U1210 (N_1210,In_2317,N_50);
and U1211 (N_1211,In_1673,N_780);
and U1212 (N_1212,N_51,In_1077);
or U1213 (N_1213,In_363,In_13);
or U1214 (N_1214,In_2231,N_827);
nand U1215 (N_1215,N_690,In_2450);
xnor U1216 (N_1216,N_719,In_1139);
or U1217 (N_1217,N_133,N_781);
and U1218 (N_1218,In_817,In_361);
or U1219 (N_1219,In_1269,In_2202);
or U1220 (N_1220,In_1087,N_498);
or U1221 (N_1221,N_895,In_767);
nor U1222 (N_1222,N_429,In_356);
nor U1223 (N_1223,N_883,In_1808);
nand U1224 (N_1224,N_475,N_930);
nor U1225 (N_1225,In_2447,In_1895);
nand U1226 (N_1226,In_909,In_1966);
or U1227 (N_1227,N_545,In_267);
or U1228 (N_1228,In_37,N_571);
or U1229 (N_1229,In_906,In_1336);
xnor U1230 (N_1230,In_1375,In_430);
nor U1231 (N_1231,In_2497,N_441);
xnor U1232 (N_1232,In_770,N_360);
xor U1233 (N_1233,In_1867,N_894);
xnor U1234 (N_1234,N_363,In_1831);
nor U1235 (N_1235,In_2051,N_658);
xnor U1236 (N_1236,In_867,In_1652);
nor U1237 (N_1237,In_2325,In_248);
nand U1238 (N_1238,N_898,N_570);
xor U1239 (N_1239,In_1081,N_871);
and U1240 (N_1240,N_806,In_887);
nor U1241 (N_1241,N_773,In_921);
or U1242 (N_1242,In_2210,N_594);
and U1243 (N_1243,In_863,In_693);
xnor U1244 (N_1244,In_667,N_668);
or U1245 (N_1245,N_125,In_155);
or U1246 (N_1246,In_273,N_970);
or U1247 (N_1247,N_578,N_768);
xnor U1248 (N_1248,In_173,N_506);
xnor U1249 (N_1249,N_618,In_821);
nor U1250 (N_1250,In_317,In_1184);
and U1251 (N_1251,N_1124,N_974);
nor U1252 (N_1252,N_1040,N_1085);
or U1253 (N_1253,In_327,N_1123);
and U1254 (N_1254,N_626,N_1011);
xor U1255 (N_1255,In_1955,In_2211);
nor U1256 (N_1256,N_407,In_1440);
or U1257 (N_1257,N_442,In_2181);
or U1258 (N_1258,In_291,In_1378);
and U1259 (N_1259,In_143,In_875);
xor U1260 (N_1260,N_757,In_2245);
or U1261 (N_1261,In_1280,N_1177);
nand U1262 (N_1262,In_2057,N_558);
and U1263 (N_1263,In_236,N_1207);
or U1264 (N_1264,N_957,In_1380);
and U1265 (N_1265,N_706,In_2221);
nor U1266 (N_1266,In_1907,N_1147);
or U1267 (N_1267,In_411,In_873);
xor U1268 (N_1268,N_522,N_110);
nor U1269 (N_1269,In_2002,N_387);
xnor U1270 (N_1270,In_996,In_244);
xor U1271 (N_1271,In_862,In_1324);
nor U1272 (N_1272,N_1070,N_1016);
or U1273 (N_1273,N_303,N_733);
xnor U1274 (N_1274,In_32,N_1115);
or U1275 (N_1275,N_282,N_1121);
xor U1276 (N_1276,N_390,In_1731);
and U1277 (N_1277,In_2092,N_193);
and U1278 (N_1278,N_567,In_2116);
xor U1279 (N_1279,In_1764,In_2076);
nand U1280 (N_1280,In_1604,In_129);
or U1281 (N_1281,In_1297,In_1649);
nor U1282 (N_1282,In_1271,N_1151);
nor U1283 (N_1283,N_855,N_874);
nand U1284 (N_1284,In_2335,N_725);
nand U1285 (N_1285,N_361,N_924);
nor U1286 (N_1286,In_495,N_1222);
nand U1287 (N_1287,In_2118,N_1138);
and U1288 (N_1288,N_775,N_987);
xnor U1289 (N_1289,N_831,In_646);
xor U1290 (N_1290,In_1466,In_1688);
nor U1291 (N_1291,In_1044,In_1985);
xor U1292 (N_1292,In_681,N_876);
xor U1293 (N_1293,N_124,In_2199);
nor U1294 (N_1294,In_180,In_2204);
nand U1295 (N_1295,N_1174,N_128);
nor U1296 (N_1296,N_972,N_1243);
nand U1297 (N_1297,N_421,In_558);
or U1298 (N_1298,N_789,N_1128);
nand U1299 (N_1299,In_1093,In_1458);
nor U1300 (N_1300,N_1066,N_736);
nand U1301 (N_1301,N_577,In_1221);
and U1302 (N_1302,In_1265,In_1365);
nor U1303 (N_1303,In_528,N_849);
nand U1304 (N_1304,In_1968,N_1045);
nand U1305 (N_1305,N_1002,N_890);
xor U1306 (N_1306,In_1535,N_183);
or U1307 (N_1307,In_1101,In_1042);
xor U1308 (N_1308,N_712,In_1946);
or U1309 (N_1309,N_309,N_57);
or U1310 (N_1310,N_1193,N_307);
nor U1311 (N_1311,In_1727,N_1005);
or U1312 (N_1312,In_96,N_703);
and U1313 (N_1313,N_815,N_766);
nand U1314 (N_1314,In_1859,N_1248);
nor U1315 (N_1315,N_636,N_338);
or U1316 (N_1316,N_1061,In_1815);
nor U1317 (N_1317,N_1188,In_1218);
or U1318 (N_1318,N_1140,N_1249);
or U1319 (N_1319,N_479,N_1169);
nor U1320 (N_1320,N_252,N_1136);
nor U1321 (N_1321,In_502,N_582);
or U1322 (N_1322,N_685,N_921);
and U1323 (N_1323,In_61,In_935);
nand U1324 (N_1324,N_707,N_478);
nor U1325 (N_1325,N_162,In_729);
or U1326 (N_1326,N_1246,In_78);
xnor U1327 (N_1327,In_2001,N_838);
nor U1328 (N_1328,In_1612,In_270);
and U1329 (N_1329,N_375,N_796);
xor U1330 (N_1330,In_2499,In_892);
xnor U1331 (N_1331,N_312,N_1015);
or U1332 (N_1332,In_2034,N_416);
nor U1333 (N_1333,In_22,N_1095);
nand U1334 (N_1334,In_252,In_449);
and U1335 (N_1335,N_1187,N_764);
nor U1336 (N_1336,In_1135,N_918);
nand U1337 (N_1337,In_29,N_38);
or U1338 (N_1338,N_1113,In_608);
xnor U1339 (N_1339,In_1134,N_1240);
nor U1340 (N_1340,In_413,In_1768);
and U1341 (N_1341,In_546,N_1146);
and U1342 (N_1342,N_178,N_259);
or U1343 (N_1343,N_750,N_155);
and U1344 (N_1344,N_1159,N_1046);
and U1345 (N_1345,In_835,N_950);
nor U1346 (N_1346,In_227,In_1034);
xor U1347 (N_1347,N_235,In_791);
nor U1348 (N_1348,In_1945,N_216);
nand U1349 (N_1349,N_611,In_564);
xor U1350 (N_1350,In_355,N_369);
or U1351 (N_1351,In_1954,In_2329);
xor U1352 (N_1352,In_2248,In_1094);
xnor U1353 (N_1353,N_1106,N_1160);
xor U1354 (N_1354,In_1129,In_1610);
nand U1355 (N_1355,N_218,In_1940);
xor U1356 (N_1356,In_1881,N_1111);
nor U1357 (N_1357,N_332,In_1919);
and U1358 (N_1358,N_873,N_863);
or U1359 (N_1359,In_603,N_1232);
xor U1360 (N_1360,N_786,N_1148);
nor U1361 (N_1361,In_1079,N_886);
nor U1362 (N_1362,N_808,N_1129);
nand U1363 (N_1363,N_802,In_2097);
xor U1364 (N_1364,N_1189,N_1211);
or U1365 (N_1365,N_856,N_388);
xnor U1366 (N_1366,In_1474,N_944);
xor U1367 (N_1367,N_676,N_1026);
nand U1368 (N_1368,N_1035,N_647);
or U1369 (N_1369,N_1057,In_503);
xor U1370 (N_1370,N_617,N_1197);
or U1371 (N_1371,N_1074,N_1133);
nand U1372 (N_1372,N_1024,In_1712);
nor U1373 (N_1373,In_105,In_1804);
and U1374 (N_1374,N_941,In_688);
or U1375 (N_1375,In_432,In_296);
or U1376 (N_1376,N_1053,N_348);
or U1377 (N_1377,N_621,In_1255);
xor U1378 (N_1378,In_557,In_372);
or U1379 (N_1379,In_819,In_1425);
and U1380 (N_1380,N_916,In_2224);
or U1381 (N_1381,In_763,In_435);
or U1382 (N_1382,N_1201,In_1319);
xnor U1383 (N_1383,In_926,In_181);
or U1384 (N_1384,N_726,N_553);
nand U1385 (N_1385,N_32,In_1284);
and U1386 (N_1386,N_297,In_997);
xor U1387 (N_1387,N_1150,In_1230);
and U1388 (N_1388,In_888,N_599);
and U1389 (N_1389,N_102,In_1679);
or U1390 (N_1390,In_1866,In_511);
nor U1391 (N_1391,In_1051,N_444);
or U1392 (N_1392,N_1067,N_420);
or U1393 (N_1393,In_2157,In_2463);
nor U1394 (N_1394,N_23,In_1);
or U1395 (N_1395,In_1361,In_2216);
nand U1396 (N_1396,N_763,N_1076);
nand U1397 (N_1397,N_1110,N_904);
nor U1398 (N_1398,N_1226,N_1097);
and U1399 (N_1399,N_879,N_912);
nand U1400 (N_1400,N_19,N_1091);
and U1401 (N_1401,N_959,N_1209);
xor U1402 (N_1402,N_335,N_903);
nor U1403 (N_1403,N_525,In_505);
nor U1404 (N_1404,N_627,In_184);
or U1405 (N_1405,N_83,In_1525);
xnor U1406 (N_1406,N_843,In_15);
and U1407 (N_1407,N_1099,N_1120);
xor U1408 (N_1408,N_199,In_1596);
or U1409 (N_1409,In_1340,N_993);
or U1410 (N_1410,N_751,In_1229);
nor U1411 (N_1411,N_728,N_933);
and U1412 (N_1412,N_503,N_752);
and U1413 (N_1413,In_1766,N_389);
nor U1414 (N_1414,In_360,N_922);
nor U1415 (N_1415,In_2416,N_1227);
xor U1416 (N_1416,N_897,N_308);
and U1417 (N_1417,N_1204,In_2420);
nand U1418 (N_1418,N_290,N_632);
nor U1419 (N_1419,N_758,In_531);
or U1420 (N_1420,N_520,N_977);
nand U1421 (N_1421,N_1114,In_208);
and U1422 (N_1422,In_2213,N_742);
xnor U1423 (N_1423,In_1259,N_93);
nor U1424 (N_1424,In_865,N_865);
nor U1425 (N_1425,In_1957,N_826);
xor U1426 (N_1426,N_1050,In_127);
nor U1427 (N_1427,N_397,In_2330);
or U1428 (N_1428,In_1554,N_1142);
or U1429 (N_1429,N_1027,N_245);
or U1430 (N_1430,N_586,N_1105);
xnor U1431 (N_1431,In_2389,N_439);
nand U1432 (N_1432,N_981,N_759);
nor U1433 (N_1433,In_584,N_1213);
and U1434 (N_1434,In_1576,N_206);
nor U1435 (N_1435,In_2077,N_1182);
nand U1436 (N_1436,N_484,In_2169);
or U1437 (N_1437,In_1489,N_264);
xnor U1438 (N_1438,In_250,In_2059);
nand U1439 (N_1439,N_1172,In_2246);
nor U1440 (N_1440,In_1561,In_1585);
nor U1441 (N_1441,In_442,In_1797);
nand U1442 (N_1442,In_1264,In_2062);
or U1443 (N_1443,In_1562,N_254);
xnor U1444 (N_1444,In_828,N_803);
nand U1445 (N_1445,N_1198,In_951);
xor U1446 (N_1446,N_226,N_1089);
nor U1447 (N_1447,In_989,In_2171);
xnor U1448 (N_1448,N_323,In_1022);
and U1449 (N_1449,N_1244,N_994);
nor U1450 (N_1450,In_156,N_1088);
nand U1451 (N_1451,N_991,N_1191);
and U1452 (N_1452,N_1205,In_1530);
xor U1453 (N_1453,N_1039,N_915);
nand U1454 (N_1454,In_2438,N_997);
and U1455 (N_1455,N_1208,N_936);
and U1456 (N_1456,N_851,N_715);
nor U1457 (N_1457,In_1179,N_1131);
and U1458 (N_1458,N_370,N_1071);
nor U1459 (N_1459,N_65,N_1109);
xor U1460 (N_1460,In_1984,N_1055);
xnor U1461 (N_1461,N_1059,N_900);
and U1462 (N_1462,In_590,In_2148);
xor U1463 (N_1463,In_1811,In_1785);
or U1464 (N_1464,In_126,In_728);
or U1465 (N_1465,N_101,In_2019);
nand U1466 (N_1466,In_39,N_576);
nor U1467 (N_1467,N_988,N_327);
xor U1468 (N_1468,N_964,N_735);
and U1469 (N_1469,In_632,N_1168);
xor U1470 (N_1470,In_1088,In_12);
nand U1471 (N_1471,In_599,N_645);
nand U1472 (N_1472,In_2269,N_426);
nor U1473 (N_1473,In_933,N_953);
nor U1474 (N_1474,N_100,N_447);
nand U1475 (N_1475,N_1180,N_911);
nand U1476 (N_1476,N_230,In_387);
nor U1477 (N_1477,N_761,N_146);
or U1478 (N_1478,In_325,In_115);
and U1479 (N_1479,N_455,N_1044);
and U1480 (N_1480,In_2411,N_790);
nor U1481 (N_1481,In_990,N_1043);
nand U1482 (N_1482,N_620,In_1500);
nand U1483 (N_1483,N_1103,N_1192);
xor U1484 (N_1484,In_2060,In_700);
or U1485 (N_1485,N_628,In_1690);
xor U1486 (N_1486,In_136,N_204);
nand U1487 (N_1487,N_973,In_2354);
or U1488 (N_1488,N_535,N_852);
and U1489 (N_1489,N_1185,N_1073);
nor U1490 (N_1490,In_2331,In_2174);
nor U1491 (N_1491,In_2185,N_438);
nand U1492 (N_1492,N_337,N_702);
nor U1493 (N_1493,N_1152,N_1122);
nor U1494 (N_1494,N_846,N_1052);
and U1495 (N_1495,In_1409,In_1266);
and U1496 (N_1496,N_965,N_376);
or U1497 (N_1497,N_562,N_548);
and U1498 (N_1498,In_1470,In_1884);
and U1499 (N_1499,N_1100,In_487);
and U1500 (N_1500,N_280,N_836);
or U1501 (N_1501,N_471,N_412);
nand U1502 (N_1502,N_1282,N_194);
xor U1503 (N_1503,In_2475,N_983);
or U1504 (N_1504,N_990,N_1096);
and U1505 (N_1505,In_810,In_1397);
nand U1506 (N_1506,N_1276,N_385);
and U1507 (N_1507,N_1153,N_592);
xor U1508 (N_1508,N_1499,N_195);
and U1509 (N_1509,In_1023,In_1638);
xnor U1510 (N_1510,N_1342,N_1229);
or U1511 (N_1511,N_1346,N_858);
nor U1512 (N_1512,N_437,N_1063);
and U1513 (N_1513,N_749,In_34);
xnor U1514 (N_1514,In_793,N_448);
nand U1515 (N_1515,N_1242,In_1603);
xnor U1516 (N_1516,N_1056,N_1477);
nor U1517 (N_1517,N_1331,N_1462);
nor U1518 (N_1518,N_1281,In_750);
or U1519 (N_1519,N_639,N_1286);
nand U1520 (N_1520,N_655,N_606);
nand U1521 (N_1521,N_257,N_285);
xnor U1522 (N_1522,In_1524,N_971);
or U1523 (N_1523,N_1183,In_318);
and U1524 (N_1524,N_7,N_716);
nor U1525 (N_1525,N_460,In_11);
or U1526 (N_1526,N_1217,N_1403);
and U1527 (N_1527,N_1196,N_1234);
nor U1528 (N_1528,In_703,N_870);
or U1529 (N_1529,N_1326,In_903);
nand U1530 (N_1530,In_698,In_68);
nand U1531 (N_1531,N_1223,N_1141);
or U1532 (N_1532,N_948,N_1195);
nand U1533 (N_1533,N_1333,In_1013);
nand U1534 (N_1534,N_692,In_1441);
nor U1535 (N_1535,In_553,N_1479);
nand U1536 (N_1536,N_711,In_1537);
or U1537 (N_1537,N_968,N_935);
or U1538 (N_1538,In_482,N_1054);
or U1539 (N_1539,N_634,N_813);
xnor U1540 (N_1540,In_1615,N_609);
nor U1541 (N_1541,N_1397,N_1225);
or U1542 (N_1542,N_958,In_1793);
nand U1543 (N_1543,N_932,In_1037);
nand U1544 (N_1544,N_563,In_683);
or U1545 (N_1545,N_648,N_1393);
nor U1546 (N_1546,In_1844,N_529);
xor U1547 (N_1547,In_1235,N_1391);
nand U1548 (N_1548,N_1093,In_198);
nand U1549 (N_1549,In_2280,In_2388);
nand U1550 (N_1550,N_1455,N_881);
nand U1551 (N_1551,In_752,N_1300);
xor U1552 (N_1552,N_546,In_1170);
and U1553 (N_1553,In_617,In_451);
xor U1554 (N_1554,N_1202,In_1195);
xnor U1555 (N_1555,N_584,In_2206);
nor U1556 (N_1556,N_1006,N_788);
and U1557 (N_1557,N_263,In_393);
nand U1558 (N_1558,N_1432,N_1360);
nor U1559 (N_1559,N_560,In_2187);
nand U1560 (N_1560,N_860,In_984);
xnor U1561 (N_1561,N_84,N_1154);
and U1562 (N_1562,N_1376,N_1399);
and U1563 (N_1563,N_1363,N_469);
or U1564 (N_1564,In_2305,N_945);
nor U1565 (N_1565,N_1490,N_1303);
nor U1566 (N_1566,N_629,N_346);
or U1567 (N_1567,N_1402,N_1020);
xnor U1568 (N_1568,In_803,In_1587);
nor U1569 (N_1569,N_1190,N_1439);
nand U1570 (N_1570,N_1442,N_521);
nor U1571 (N_1571,In_2393,N_1480);
nand U1572 (N_1572,In_637,N_1075);
or U1573 (N_1573,In_50,In_197);
or U1574 (N_1574,N_1254,N_1162);
xor U1575 (N_1575,In_578,N_1456);
xor U1576 (N_1576,N_1029,N_1062);
nor U1577 (N_1577,N_923,N_701);
or U1578 (N_1578,N_1378,In_185);
and U1579 (N_1579,N_55,In_811);
nand U1580 (N_1580,In_1000,N_1022);
xor U1581 (N_1581,N_1336,N_1436);
nand U1582 (N_1582,N_1384,N_602);
xor U1583 (N_1583,In_444,N_1320);
nor U1584 (N_1584,In_1354,N_1485);
nor U1585 (N_1585,In_1622,N_500);
nand U1586 (N_1586,N_1431,N_1049);
and U1587 (N_1587,N_1112,N_995);
xnor U1588 (N_1588,N_1484,In_982);
nor U1589 (N_1589,N_1012,N_1330);
xnor U1590 (N_1590,N_278,N_1447);
or U1591 (N_1591,N_1175,N_1325);
nor U1592 (N_1592,N_792,N_1350);
nor U1593 (N_1593,N_1472,N_1418);
or U1594 (N_1594,N_623,In_225);
and U1595 (N_1595,In_1567,N_710);
or U1596 (N_1596,N_575,N_665);
xor U1597 (N_1597,N_1135,In_2372);
nand U1598 (N_1598,N_1373,N_1459);
or U1599 (N_1599,N_1394,N_835);
nand U1600 (N_1600,N_888,In_2013);
xnor U1601 (N_1601,In_1913,In_2123);
xor U1602 (N_1602,N_1210,In_782);
nor U1603 (N_1603,In_428,N_1019);
nor U1604 (N_1604,N_1264,In_2219);
xnor U1605 (N_1605,N_837,N_798);
or U1606 (N_1606,N_1440,N_176);
and U1607 (N_1607,N_396,N_516);
and U1608 (N_1608,In_561,In_713);
or U1609 (N_1609,N_875,N_713);
nor U1610 (N_1610,N_893,N_774);
and U1611 (N_1611,In_2490,In_2408);
nor U1612 (N_1612,N_1017,In_1274);
xnor U1613 (N_1613,In_18,In_186);
nor U1614 (N_1614,N_1377,In_2290);
and U1615 (N_1615,N_463,In_426);
nor U1616 (N_1616,N_864,In_377);
xnor U1617 (N_1617,N_1400,N_961);
nand U1618 (N_1618,N_1285,N_95);
nor U1619 (N_1619,N_1163,In_2079);
nand U1620 (N_1620,N_1092,N_869);
xor U1621 (N_1621,N_1473,In_357);
and U1622 (N_1622,N_1353,N_1291);
and U1623 (N_1623,In_2004,N_1139);
or U1624 (N_1624,In_468,In_433);
nand U1625 (N_1625,N_1467,N_1009);
xor U1626 (N_1626,N_1388,In_919);
and U1627 (N_1627,In_1746,N_901);
or U1628 (N_1628,N_734,N_1042);
nand U1629 (N_1629,In_2164,N_1302);
or U1630 (N_1630,N_866,N_384);
xnor U1631 (N_1631,N_1461,N_1345);
nor U1632 (N_1632,N_787,N_236);
nand U1633 (N_1633,N_1423,In_949);
and U1634 (N_1634,In_2279,In_2031);
nor U1635 (N_1635,In_394,N_446);
xor U1636 (N_1636,In_374,In_1330);
xnor U1637 (N_1637,N_1030,N_727);
nor U1638 (N_1638,N_985,In_1551);
or U1639 (N_1639,N_939,N_523);
or U1640 (N_1640,N_474,In_1851);
nor U1641 (N_1641,N_607,In_1366);
and U1642 (N_1642,N_834,In_1915);
nand U1643 (N_1643,In_2083,N_1441);
nor U1644 (N_1644,In_1145,N_1458);
or U1645 (N_1645,In_268,In_1636);
nand U1646 (N_1646,N_704,N_1116);
xor U1647 (N_1647,N_1392,N_1315);
or U1648 (N_1648,N_1215,N_962);
nor U1649 (N_1649,In_2039,N_1424);
and U1650 (N_1650,N_1161,In_1395);
or U1651 (N_1651,N_675,In_2241);
xnor U1652 (N_1652,In_1127,N_1448);
nand U1653 (N_1653,In_1760,N_228);
and U1654 (N_1654,N_717,N_612);
nor U1655 (N_1655,N_1272,N_820);
xor U1656 (N_1656,N_699,N_1433);
xnor U1657 (N_1657,In_1642,N_756);
or U1658 (N_1658,N_1289,N_153);
and U1659 (N_1659,In_238,N_1260);
nand U1660 (N_1660,In_2263,N_693);
nand U1661 (N_1661,N_1381,In_258);
xor U1662 (N_1662,N_1498,N_952);
and U1663 (N_1663,N_211,In_897);
or U1664 (N_1664,N_1176,N_1481);
or U1665 (N_1665,In_2437,In_1877);
xnor U1666 (N_1666,N_1343,In_343);
nand U1667 (N_1667,N_947,N_1310);
nand U1668 (N_1668,N_365,N_71);
xor U1669 (N_1669,In_1687,N_249);
and U1670 (N_1670,N_1033,In_257);
xnor U1671 (N_1671,N_1416,In_60);
or U1672 (N_1672,N_1396,N_1003);
or U1673 (N_1673,N_518,In_2011);
nor U1674 (N_1674,In_960,N_679);
and U1675 (N_1675,N_1446,In_2491);
or U1676 (N_1676,N_1233,N_687);
nand U1677 (N_1677,N_1395,N_1094);
xor U1678 (N_1678,In_1445,In_2103);
nand U1679 (N_1679,N_534,In_2161);
xor U1680 (N_1680,N_1426,N_804);
and U1681 (N_1681,In_1693,In_1171);
nand U1682 (N_1682,In_1528,N_1134);
and U1683 (N_1683,In_1711,In_934);
and U1684 (N_1684,In_1166,N_770);
or U1685 (N_1685,N_1256,N_1230);
or U1686 (N_1686,N_561,N_1224);
or U1687 (N_1687,N_1058,In_1848);
nor U1688 (N_1688,N_1438,In_2465);
or U1689 (N_1689,In_822,In_358);
nand U1690 (N_1690,N_1468,In_125);
and U1691 (N_1691,N_1463,N_1380);
nor U1692 (N_1692,In_2445,N_1238);
nand U1693 (N_1693,N_1284,N_1312);
nand U1694 (N_1694,In_711,In_331);
and U1695 (N_1695,N_1453,N_819);
xnor U1696 (N_1696,N_1130,N_640);
xnor U1697 (N_1697,In_2016,N_1322);
and U1698 (N_1698,N_1298,N_1087);
xnor U1699 (N_1699,N_1069,N_1299);
nor U1700 (N_1700,N_1068,N_1104);
xor U1701 (N_1701,In_379,In_1180);
or U1702 (N_1702,N_1495,N_1445);
and U1703 (N_1703,In_853,N_880);
and U1704 (N_1704,N_1265,N_779);
or U1705 (N_1705,N_1082,N_891);
and U1706 (N_1706,N_822,N_1367);
or U1707 (N_1707,N_1412,N_1164);
nor U1708 (N_1708,In_1774,N_905);
and U1709 (N_1709,N_1270,N_920);
nand U1710 (N_1710,In_2386,N_350);
nand U1711 (N_1711,N_1166,N_1170);
nand U1712 (N_1712,N_313,N_1356);
and U1713 (N_1713,In_1581,N_784);
nand U1714 (N_1714,In_338,N_466);
xnor U1715 (N_1715,In_706,N_1023);
nand U1716 (N_1716,N_1351,N_1494);
nor U1717 (N_1717,N_353,In_514);
nor U1718 (N_1718,N_1370,N_1171);
or U1719 (N_1719,N_1341,In_1475);
and U1720 (N_1720,In_1165,In_1277);
or U1721 (N_1721,N_1268,N_889);
xor U1722 (N_1722,In_24,N_1469);
or U1723 (N_1723,In_195,N_1263);
xor U1724 (N_1724,In_429,N_1080);
or U1725 (N_1725,N_1247,N_1278);
or U1726 (N_1726,In_2368,N_913);
xnor U1727 (N_1727,In_602,N_1297);
xor U1728 (N_1728,N_1258,In_836);
and U1729 (N_1729,N_800,N_1157);
and U1730 (N_1730,In_520,N_1149);
nor U1731 (N_1731,In_10,N_343);
nor U1732 (N_1732,N_654,N_1337);
nor U1733 (N_1733,In_1169,N_1316);
nor U1734 (N_1734,N_1167,N_1072);
nor U1735 (N_1735,In_1428,N_899);
or U1736 (N_1736,In_1922,N_1206);
or U1737 (N_1737,N_1261,In_1313);
or U1738 (N_1738,In_1949,In_907);
or U1739 (N_1739,N_1334,In_1926);
nor U1740 (N_1740,In_1618,N_1451);
and U1741 (N_1741,N_1245,In_1100);
or U1742 (N_1742,N_1324,N_1010);
nand U1743 (N_1743,N_269,N_1410);
xnor U1744 (N_1744,N_485,N_1079);
or U1745 (N_1745,In_2318,N_1025);
and U1746 (N_1746,N_1060,N_513);
and U1747 (N_1747,N_1000,N_671);
xnor U1748 (N_1748,N_587,N_1077);
xor U1749 (N_1749,In_1571,In_999);
nand U1750 (N_1750,N_1422,N_1522);
or U1751 (N_1751,N_1083,N_616);
nand U1752 (N_1752,N_1102,N_1715);
nor U1753 (N_1753,N_1450,In_654);
nor U1754 (N_1754,N_1406,N_1667);
nand U1755 (N_1755,N_1581,N_1501);
and U1756 (N_1756,In_2085,In_340);
xnor U1757 (N_1757,N_1007,N_1475);
nand U1758 (N_1758,N_1701,N_1567);
xor U1759 (N_1759,N_1532,N_219);
and U1760 (N_1760,N_1572,N_1239);
xnor U1761 (N_1761,N_1713,In_1207);
xnor U1762 (N_1762,N_841,In_43);
and U1763 (N_1763,In_1490,N_1747);
or U1764 (N_1764,In_1988,N_1200);
xnor U1765 (N_1765,N_1724,In_2423);
and U1766 (N_1766,N_1425,N_1119);
nor U1767 (N_1767,N_1327,N_867);
xnor U1768 (N_1768,N_1741,In_205);
xnor U1769 (N_1769,N_1536,In_1522);
nor U1770 (N_1770,N_1428,In_3);
and U1771 (N_1771,N_1497,N_1421);
nor U1772 (N_1772,In_714,N_1681);
or U1773 (N_1773,In_931,N_1735);
nor U1774 (N_1774,In_65,N_1746);
nor U1775 (N_1775,N_1155,N_1408);
or U1776 (N_1776,N_1236,N_217);
or U1777 (N_1777,N_1430,In_1842);
xnor U1778 (N_1778,In_806,N_1538);
xnor U1779 (N_1779,In_2109,N_1587);
nand U1780 (N_1780,N_603,N_637);
nor U1781 (N_1781,N_96,N_718);
or U1782 (N_1782,In_2259,N_967);
and U1783 (N_1783,N_1721,N_1672);
nor U1784 (N_1784,N_1563,In_1414);
or U1785 (N_1785,N_25,N_1317);
xor U1786 (N_1786,N_1637,N_1560);
nand U1787 (N_1787,N_1557,N_588);
and U1788 (N_1788,N_1364,In_93);
and U1789 (N_1789,N_1382,N_1483);
or U1790 (N_1790,N_1551,N_1429);
xor U1791 (N_1791,N_1296,In_1312);
and U1792 (N_1792,In_915,N_1544);
and U1793 (N_1793,N_928,N_1117);
xnor U1794 (N_1794,N_1634,In_1861);
or U1795 (N_1795,N_1535,N_1728);
or U1796 (N_1796,N_1269,N_1098);
and U1797 (N_1797,N_1705,N_231);
nand U1798 (N_1798,N_1253,N_1619);
xnor U1799 (N_1799,N_1658,In_1126);
xnor U1800 (N_1800,N_1528,In_2099);
nor U1801 (N_1801,In_2464,N_1311);
nand U1802 (N_1802,N_1437,N_1048);
and U1803 (N_1803,N_504,N_695);
nand U1804 (N_1804,N_94,N_1645);
nand U1805 (N_1805,In_212,N_769);
xnor U1806 (N_1806,N_593,N_1365);
and U1807 (N_1807,N_1537,In_800);
xnor U1808 (N_1808,N_1457,N_1318);
nor U1809 (N_1809,N_1465,N_1657);
nand U1810 (N_1810,In_1663,N_1613);
xor U1811 (N_1811,N_1585,N_1576);
xnor U1812 (N_1812,In_391,N_1712);
xor U1813 (N_1813,N_1515,N_1569);
or U1814 (N_1814,N_1018,N_1308);
nand U1815 (N_1815,N_1267,N_1127);
nor U1816 (N_1816,N_830,N_1013);
nand U1817 (N_1817,N_1454,N_1578);
and U1818 (N_1818,N_1691,N_1065);
and U1819 (N_1819,N_1434,In_1613);
and U1820 (N_1820,N_1561,N_1216);
and U1821 (N_1821,N_810,N_1693);
xnor U1822 (N_1822,N_809,N_1583);
and U1823 (N_1823,N_1369,In_1801);
nor U1824 (N_1824,In_1415,N_1165);
or U1825 (N_1825,In_1637,N_1487);
xor U1826 (N_1826,N_359,N_1503);
and U1827 (N_1827,In_1559,N_1452);
xor U1828 (N_1828,N_1550,N_1612);
or U1829 (N_1829,N_1476,N_1255);
xor U1830 (N_1830,N_1723,In_516);
and U1831 (N_1831,N_1661,N_1502);
xor U1832 (N_1832,In_170,In_2348);
and U1833 (N_1833,In_1073,In_75);
and U1834 (N_1834,N_1500,N_1571);
and U1835 (N_1835,N_1590,N_1158);
or U1836 (N_1836,In_1805,In_702);
nand U1837 (N_1837,N_428,N_1496);
nand U1838 (N_1838,N_456,In_2058);
or U1839 (N_1839,N_1602,N_1519);
and U1840 (N_1840,N_1386,N_1335);
nor U1841 (N_1841,N_1385,In_1936);
nand U1842 (N_1842,N_87,N_1682);
xnor U1843 (N_1843,N_1004,N_541);
and U1844 (N_1844,In_789,N_1700);
nor U1845 (N_1845,N_583,N_1379);
nor U1846 (N_1846,N_1292,N_1295);
nor U1847 (N_1847,N_1357,In_1816);
nor U1848 (N_1848,In_375,In_1172);
nor U1849 (N_1849,N_1478,N_1314);
or U1850 (N_1850,N_1648,In_427);
xor U1851 (N_1851,In_2107,N_1443);
and U1852 (N_1852,In_775,N_1221);
xor U1853 (N_1853,N_1738,N_581);
or U1854 (N_1854,N_956,N_884);
or U1855 (N_1855,N_289,N_857);
and U1856 (N_1856,In_820,N_1145);
nor U1857 (N_1857,N_1530,In_2113);
nor U1858 (N_1858,N_1358,N_1199);
xnor U1859 (N_1859,N_1540,N_1417);
nand U1860 (N_1860,N_1321,N_812);
nand U1861 (N_1861,N_1608,In_824);
nor U1862 (N_1862,In_2383,N_1579);
nor U1863 (N_1863,N_1703,N_352);
nor U1864 (N_1864,N_1362,N_1504);
nor U1865 (N_1865,N_1374,N_1699);
xor U1866 (N_1866,N_1644,In_2191);
nor U1867 (N_1867,In_1574,In_795);
or U1868 (N_1868,In_1320,In_1387);
nor U1869 (N_1869,In_1896,N_896);
xor U1870 (N_1870,N_1328,N_1525);
nand U1871 (N_1871,N_1307,N_1309);
nor U1872 (N_1872,N_1184,N_1078);
or U1873 (N_1873,N_1553,N_1214);
or U1874 (N_1874,N_1340,N_1737);
xnor U1875 (N_1875,N_1101,N_1616);
nand U1876 (N_1876,In_2390,N_1624);
nor U1877 (N_1877,N_942,In_522);
nand U1878 (N_1878,In_2106,N_1660);
and U1879 (N_1879,N_1632,N_641);
nand U1880 (N_1880,N_1574,In_2359);
nor U1881 (N_1881,N_1694,N_1580);
nand U1882 (N_1882,N_135,N_1420);
xor U1883 (N_1883,N_1520,In_1726);
nor U1884 (N_1884,In_2387,N_317);
nand U1885 (N_1885,N_1556,N_595);
nand U1886 (N_1886,N_1510,N_1552);
xnor U1887 (N_1887,N_1186,In_1939);
and U1888 (N_1888,N_1032,N_1598);
nor U1889 (N_1889,N_1601,N_1031);
xor U1890 (N_1890,In_2091,N_1620);
nand U1891 (N_1891,N_1277,N_1368);
or U1892 (N_1892,N_1257,N_34);
nor U1893 (N_1893,N_1649,N_556);
nand U1894 (N_1894,N_1352,In_1504);
nor U1895 (N_1895,N_1614,N_882);
nand U1896 (N_1896,In_748,N_1558);
nor U1897 (N_1897,In_661,N_1629);
xor U1898 (N_1898,N_938,N_141);
xor U1899 (N_1899,In_870,N_1279);
xnor U1900 (N_1900,In_2119,In_1728);
or U1901 (N_1901,N_1554,N_999);
nand U1902 (N_1902,N_1546,In_2399);
or U1903 (N_1903,N_1283,N_329);
nor U1904 (N_1904,In_927,N_1687);
xnor U1905 (N_1905,N_1132,N_1401);
nor U1906 (N_1906,N_354,In_614);
nand U1907 (N_1907,N_1118,N_1541);
or U1908 (N_1908,N_1599,N_1573);
nor U1909 (N_1909,N_1250,N_1716);
and U1910 (N_1910,N_1647,N_1559);
or U1911 (N_1911,N_1562,N_1241);
nand U1912 (N_1912,N_1375,N_1665);
xor U1913 (N_1913,N_1435,N_1329);
and U1914 (N_1914,N_1274,In_2163);
or U1915 (N_1915,N_839,N_1584);
and U1916 (N_1916,N_527,N_1651);
xor U1917 (N_1917,N_1635,In_1004);
xnor U1918 (N_1918,N_1523,N_979);
and U1919 (N_1919,In_1894,N_6);
or U1920 (N_1920,N_708,N_1742);
xor U1921 (N_1921,In_1043,N_322);
nand U1922 (N_1922,N_1288,N_1680);
nor U1923 (N_1923,N_1470,N_1663);
xor U1924 (N_1924,N_1505,N_1577);
or U1925 (N_1925,N_1692,N_1028);
and U1926 (N_1926,N_1491,N_1178);
xor U1927 (N_1927,In_2240,In_14);
or U1928 (N_1928,In_1960,N_1610);
xor U1929 (N_1929,N_1695,N_946);
nor U1930 (N_1930,N_1512,N_1290);
nor U1931 (N_1931,N_1398,N_1636);
or U1932 (N_1932,N_163,N_1444);
xnor U1933 (N_1933,In_677,N_1575);
or U1934 (N_1934,N_1037,In_1783);
nand U1935 (N_1935,N_496,N_1419);
nand U1936 (N_1936,N_1513,In_1360);
xor U1937 (N_1937,N_1383,N_1228);
xor U1938 (N_1938,In_611,N_861);
or U1939 (N_1939,N_960,N_1547);
and U1940 (N_1940,N_1460,N_37);
and U1941 (N_1941,N_1466,N_1690);
xor U1942 (N_1942,N_1526,N_1626);
nor U1943 (N_1943,In_1639,N_1597);
or U1944 (N_1944,N_1280,In_2055);
and U1945 (N_1945,In_624,In_2403);
and U1946 (N_1946,In_2314,In_1651);
or U1947 (N_1947,N_1339,N_1709);
nand U1948 (N_1948,N_1301,N_1527);
or U1949 (N_1949,N_1294,In_2052);
nor U1950 (N_1950,N_302,N_1488);
or U1951 (N_1951,In_2086,N_1231);
and U1952 (N_1952,N_1137,In_622);
and U1953 (N_1953,N_1733,N_1051);
and U1954 (N_1954,N_1492,N_1749);
nor U1955 (N_1955,N_1021,N_1212);
and U1956 (N_1956,N_1427,N_1354);
xnor U1957 (N_1957,N_1555,N_1565);
or U1958 (N_1958,N_978,N_1084);
xnor U1959 (N_1959,N_1630,N_1305);
xnor U1960 (N_1960,N_1361,In_145);
nand U1961 (N_1961,N_1729,N_1633);
nand U1962 (N_1962,In_2421,N_1507);
xnor U1963 (N_1963,N_1407,In_2233);
or U1964 (N_1964,N_480,N_1349);
or U1965 (N_1965,N_1041,N_829);
and U1966 (N_1966,In_1463,N_1344);
nand U1967 (N_1967,N_635,N_1516);
xor U1968 (N_1968,N_1539,N_832);
xor U1969 (N_1969,N_271,N_1697);
nor U1970 (N_1970,N_1748,N_1194);
nor U1971 (N_1971,N_1219,N_1389);
and U1972 (N_1972,N_1545,In_1888);
nand U1973 (N_1973,In_1010,N_1596);
or U1974 (N_1974,N_1319,In_1150);
nor U1975 (N_1975,N_760,In_1014);
xnor U1976 (N_1976,N_1743,N_1666);
or U1977 (N_1977,N_1144,N_1641);
xnor U1978 (N_1978,N_1621,N_1730);
and U1979 (N_1979,N_1220,N_1404);
or U1980 (N_1980,N_1586,N_1652);
or U1981 (N_1981,In_2095,In_619);
or U1982 (N_1982,N_1603,N_209);
xor U1983 (N_1983,N_1235,N_917);
or U1984 (N_1984,In_976,N_1591);
or U1985 (N_1985,N_925,N_1549);
or U1986 (N_1986,N_797,N_116);
nand U1987 (N_1987,In_1068,In_2225);
xor U1988 (N_1988,N_1531,N_1595);
nor U1989 (N_1989,In_307,N_927);
and U1990 (N_1990,N_1372,In_2484);
nand U1991 (N_1991,N_1543,N_1745);
and U1992 (N_1992,N_1676,In_454);
or U1993 (N_1993,N_1740,N_1355);
nor U1994 (N_1994,N_440,In_781);
nor U1995 (N_1995,In_492,N_1622);
or U1996 (N_1996,In_1886,N_1708);
nand U1997 (N_1997,N_1411,N_408);
nor U1998 (N_1998,N_1486,In_455);
nor U1999 (N_1999,N_963,N_1387);
or U2000 (N_2000,N_1731,N_1972);
nand U2001 (N_2001,N_1850,N_1975);
nor U2002 (N_2002,N_1757,In_2326);
nand U2003 (N_2003,N_1996,N_1933);
nand U2004 (N_2004,N_1237,N_828);
nand U2005 (N_2005,N_1885,N_1871);
and U2006 (N_2006,N_1371,N_1853);
nor U2007 (N_2007,N_1845,N_457);
nor U2008 (N_2008,N_1566,N_1533);
xor U2009 (N_2009,N_1865,N_1706);
and U2010 (N_2010,N_1600,N_1179);
nor U2011 (N_2011,N_772,N_1409);
or U2012 (N_2012,N_1720,In_2373);
xnor U2013 (N_2013,N_1304,N_1756);
and U2014 (N_2014,In_349,In_235);
nand U2015 (N_2015,N_1951,N_1686);
nor U2016 (N_2016,N_1855,N_42);
or U2017 (N_2017,N_1332,N_1888);
nand U2018 (N_2018,N_1777,N_1768);
xor U2019 (N_2019,N_1313,N_1589);
and U2020 (N_2020,N_1086,N_1252);
nor U2021 (N_2021,N_1935,N_1973);
and U2022 (N_2022,N_1932,N_1760);
xnor U2023 (N_2023,N_1919,N_1669);
nor U2024 (N_2024,N_1793,N_1718);
nor U2025 (N_2025,N_538,N_1921);
xnor U2026 (N_2026,N_862,N_1482);
xnor U2027 (N_2027,N_1926,In_1582);
and U2028 (N_2028,N_1826,N_1405);
and U2029 (N_2029,N_1880,N_1848);
and U2030 (N_2030,N_1934,N_552);
or U2031 (N_2031,N_1805,N_1873);
nor U2032 (N_2032,N_1984,In_1301);
and U2033 (N_2033,In_2080,N_1811);
xnor U2034 (N_2034,N_1772,N_1977);
and U2035 (N_2035,N_1664,N_1908);
xnor U2036 (N_2036,N_1754,N_1798);
nor U2037 (N_2037,N_1889,N_1963);
and U2038 (N_2038,In_483,N_1776);
nor U2039 (N_2039,N_955,N_1415);
and U2040 (N_2040,N_1988,N_1625);
xnor U2041 (N_2041,N_1971,N_1967);
nand U2042 (N_2042,N_1588,N_1816);
nor U2043 (N_2043,N_1928,N_1752);
nand U2044 (N_2044,N_1958,N_1414);
and U2045 (N_2045,In_2068,In_1840);
nor U2046 (N_2046,N_1509,N_1994);
nor U2047 (N_2047,N_1471,N_1833);
xnor U2048 (N_2048,N_1789,N_700);
nor U2049 (N_2049,N_1825,N_1771);
and U2050 (N_2050,N_1995,N_1802);
nor U2051 (N_2051,N_1474,N_1837);
nand U2052 (N_2052,N_1689,N_615);
nor U2053 (N_2053,N_220,N_1819);
nor U2054 (N_2054,N_1348,In_1328);
nand U2055 (N_2055,N_1872,N_1203);
and U2056 (N_2056,In_2162,N_1064);
and U2057 (N_2057,N_1834,N_1683);
xor U2058 (N_2058,N_1960,N_1857);
xnor U2059 (N_2059,N_1878,In_2296);
or U2060 (N_2060,N_1987,N_1875);
and U2061 (N_2061,N_1899,In_891);
nand U2062 (N_2062,In_1911,N_1623);
nand U2063 (N_2063,N_1879,N_833);
or U2064 (N_2064,N_1656,N_419);
nand U2065 (N_2065,N_1751,N_1803);
nand U2066 (N_2066,N_1774,N_1911);
nand U2067 (N_2067,N_1755,N_1143);
or U2068 (N_2068,N_1864,N_1108);
or U2069 (N_2069,In_1564,N_1841);
nor U2070 (N_2070,N_1981,N_1654);
nor U2071 (N_2071,N_1787,N_1856);
nor U2072 (N_2072,N_1640,N_1534);
xnor U2073 (N_2073,N_1867,N_531);
xor U2074 (N_2074,N_1790,N_1287);
and U2075 (N_2075,N_1947,N_1852);
and U2076 (N_2076,N_1831,N_1998);
nor U2077 (N_2077,N_1815,N_241);
xor U2078 (N_2078,N_1293,N_81);
nor U2079 (N_2079,N_1677,N_1990);
nor U2080 (N_2080,N_1950,N_1961);
xnor U2081 (N_2081,N_1897,N_1970);
nand U2082 (N_2082,N_1915,N_1814);
and U2083 (N_2083,In_66,N_1854);
nand U2084 (N_2084,N_1125,In_99);
and U2085 (N_2085,N_1924,In_1404);
nand U2086 (N_2086,N_1671,N_1949);
and U2087 (N_2087,N_1993,N_604);
xnor U2088 (N_2088,N_1974,N_1702);
nand U2089 (N_2089,N_1874,In_1674);
nor U2090 (N_2090,In_2249,N_1780);
nor U2091 (N_2091,N_1882,N_1800);
nand U2092 (N_2092,N_1901,In_2351);
and U2093 (N_2093,N_1968,In_620);
or U2094 (N_2094,N_1844,N_1604);
and U2095 (N_2095,N_1955,N_1107);
nand U2096 (N_2096,N_1775,N_1861);
nand U2097 (N_2097,N_1639,N_1034);
xnor U2098 (N_2098,N_1920,N_1863);
nor U2099 (N_2099,N_1824,N_1918);
nor U2100 (N_2100,N_743,In_735);
xnor U2101 (N_2101,N_1714,N_1945);
xor U2102 (N_2102,N_1668,In_701);
nand U2103 (N_2103,N_825,N_1906);
or U2104 (N_2104,N_1883,N_1909);
nand U2105 (N_2105,N_1764,N_1835);
nor U2106 (N_2106,N_1684,N_1937);
or U2107 (N_2107,N_1643,N_1927);
nand U2108 (N_2108,N_1966,N_1758);
nor U2109 (N_2109,N_1860,N_1081);
and U2110 (N_2110,N_844,N_1761);
or U2111 (N_2111,In_1290,N_1753);
nand U2112 (N_2112,In_2449,N_1518);
nor U2113 (N_2113,In_629,N_1047);
xor U2114 (N_2114,N_1778,N_1936);
and U2115 (N_2115,N_1910,N_1851);
xor U2116 (N_2116,N_1895,N_1568);
nor U2117 (N_2117,N_1893,N_103);
nand U2118 (N_2118,N_1799,N_1744);
xor U2119 (N_2119,N_1913,N_1902);
xor U2120 (N_2120,N_1978,N_696);
xor U2121 (N_2121,N_1986,N_1923);
nand U2122 (N_2122,N_1818,N_1765);
nand U2123 (N_2123,N_1840,In_2480);
and U2124 (N_2124,N_1631,N_1763);
xor U2125 (N_2125,N_1907,N_1914);
nand U2126 (N_2126,N_1008,N_943);
nand U2127 (N_2127,N_1628,N_1954);
or U2128 (N_2128,N_694,N_793);
and U2129 (N_2129,N_1791,N_1717);
nor U2130 (N_2130,N_1829,N_1783);
and U2131 (N_2131,In_47,N_1821);
xor U2132 (N_2132,N_1609,N_1592);
and U2133 (N_2133,In_2332,N_573);
nor U2134 (N_2134,N_1982,N_1259);
and U2135 (N_2135,N_1271,N_1605);
xor U2136 (N_2136,N_1090,N_1413);
and U2137 (N_2137,N_1969,N_1734);
or U2138 (N_2138,N_1846,N_1508);
or U2139 (N_2139,N_1941,N_1781);
and U2140 (N_2140,N_1810,N_1014);
nor U2141 (N_2141,N_1795,N_1218);
and U2142 (N_2142,N_1627,N_1957);
and U2143 (N_2143,N_1983,N_1823);
nor U2144 (N_2144,N_1916,N_1646);
nand U2145 (N_2145,N_1891,N_565);
nand U2146 (N_2146,N_1650,N_1570);
and U2147 (N_2147,N_1773,In_165);
nor U2148 (N_2148,N_1670,N_1785);
or U2149 (N_2149,In_745,N_1338);
nor U2150 (N_2150,N_1828,N_1273);
and U2151 (N_2151,N_1842,N_1992);
and U2152 (N_2152,N_248,In_704);
nand U2153 (N_2153,N_1359,N_1940);
xor U2154 (N_2154,N_1894,N_723);
or U2155 (N_2155,N_1807,N_1642);
nor U2156 (N_2156,In_932,N_1722);
or U2157 (N_2157,N_1001,N_1905);
and U2158 (N_2158,In_144,In_2133);
and U2159 (N_2159,N_672,N_1890);
xnor U2160 (N_2160,N_1827,N_1898);
and U2161 (N_2161,N_1948,N_745);
xnor U2162 (N_2162,N_1868,N_1942);
xor U2163 (N_2163,N_1801,N_1696);
nor U2164 (N_2164,N_600,N_1838);
nor U2165 (N_2165,N_1779,N_1710);
nor U2166 (N_2166,In_1701,N_1529);
xnor U2167 (N_2167,N_1959,N_814);
and U2168 (N_2168,N_1653,N_1323);
nand U2169 (N_2169,N_1962,In_312);
nand U2170 (N_2170,N_1675,N_320);
or U2171 (N_2171,N_1877,N_1869);
and U2172 (N_2172,N_1390,N_1514);
or U2173 (N_2173,N_1870,N_1156);
or U2174 (N_2174,N_1506,N_1929);
xnor U2175 (N_2175,N_1953,N_1886);
and U2176 (N_2176,N_1939,N_1678);
xor U2177 (N_2177,N_1900,N_1036);
and U2178 (N_2178,N_1704,N_1449);
nor U2179 (N_2179,N_1711,N_1956);
and U2180 (N_2180,N_1732,N_1615);
nand U2181 (N_2181,N_1564,N_1817);
or U2182 (N_2182,In_1996,N_1809);
and U2183 (N_2183,N_1989,In_1708);
or U2184 (N_2184,N_872,N_1904);
nor U2185 (N_2185,N_1839,N_1750);
or U2186 (N_2186,In_174,N_1979);
or U2187 (N_2187,N_1181,N_1784);
nor U2188 (N_2188,N_1944,N_1674);
nand U2189 (N_2189,N_1769,N_1938);
and U2190 (N_2190,N_1782,In_724);
and U2191 (N_2191,N_1038,N_1849);
or U2192 (N_2192,N_1593,In_2127);
nor U2193 (N_2193,N_1607,N_1611);
nor U2194 (N_2194,N_1822,N_1739);
nand U2195 (N_2195,In_930,N_1943);
and U2196 (N_2196,N_1804,N_1930);
xor U2197 (N_2197,N_1679,N_1859);
and U2198 (N_2198,N_1582,N_1876);
or U2199 (N_2199,N_762,In_640);
xor U2200 (N_2200,N_294,In_1367);
and U2201 (N_2201,N_1638,N_1832);
nor U2202 (N_2202,N_532,N_1511);
xnor U2203 (N_2203,N_1925,N_1727);
or U2204 (N_2204,N_1655,N_1797);
xor U2205 (N_2205,N_1464,N_1976);
xnor U2206 (N_2206,N_1896,N_1251);
or U2207 (N_2207,N_1881,N_1493);
nor U2208 (N_2208,N_633,N_1788);
nor U2209 (N_2209,N_1813,In_370);
nand U2210 (N_2210,In_1670,N_1887);
nor U2211 (N_2211,N_1999,N_1808);
and U2212 (N_2212,N_1725,N_1912);
xnor U2213 (N_2213,N_1698,N_1736);
nor U2214 (N_2214,N_1903,N_1786);
nand U2215 (N_2215,N_1917,N_1892);
xor U2216 (N_2216,N_1673,N_1952);
nand U2217 (N_2217,N_1812,N_1707);
xor U2218 (N_2218,N_1542,N_1946);
nor U2219 (N_2219,N_1173,N_1517);
nand U2220 (N_2220,N_1489,N_1858);
nand U2221 (N_2221,N_1794,N_1266);
nor U2222 (N_2222,N_1662,N_1126);
or U2223 (N_2223,N_1991,In_2063);
xnor U2224 (N_2224,N_1866,N_1766);
and U2225 (N_2225,N_1347,In_1477);
and U2226 (N_2226,N_1719,N_1830);
xnor U2227 (N_2227,N_1997,In_908);
and U2228 (N_2228,N_1965,In_17);
xnor U2229 (N_2229,In_289,N_1618);
xor U2230 (N_2230,N_1964,N_1606);
and U2231 (N_2231,N_1820,N_1884);
or U2232 (N_2232,In_168,N_1980);
nor U2233 (N_2233,N_1521,N_1306);
or U2234 (N_2234,N_1792,N_1931);
nand U2235 (N_2235,N_1796,N_1767);
nand U2236 (N_2236,N_1594,In_648);
or U2237 (N_2237,N_1688,N_1617);
xor U2238 (N_2238,N_1985,N_1726);
or U2239 (N_2239,N_537,N_1836);
nor U2240 (N_2240,N_1548,N_785);
nand U2241 (N_2241,N_1366,N_753);
nor U2242 (N_2242,N_1922,N_1862);
or U2243 (N_2243,N_185,N_1262);
and U2244 (N_2244,In_712,N_1770);
nand U2245 (N_2245,N_1759,N_1275);
and U2246 (N_2246,N_1524,N_1847);
and U2247 (N_2247,N_1685,N_1806);
and U2248 (N_2248,N_976,N_1659);
or U2249 (N_2249,N_1762,N_1843);
xnor U2250 (N_2250,N_2076,N_2187);
nand U2251 (N_2251,N_2167,N_2056);
and U2252 (N_2252,N_2182,N_2104);
nand U2253 (N_2253,N_2203,N_2213);
and U2254 (N_2254,N_2032,N_2127);
nand U2255 (N_2255,N_2095,N_2027);
and U2256 (N_2256,N_2026,N_2066);
or U2257 (N_2257,N_2198,N_2249);
nor U2258 (N_2258,N_2029,N_2061);
and U2259 (N_2259,N_2153,N_2195);
nor U2260 (N_2260,N_2118,N_2156);
or U2261 (N_2261,N_2111,N_2239);
xor U2262 (N_2262,N_2017,N_2045);
or U2263 (N_2263,N_2054,N_2067);
nor U2264 (N_2264,N_2243,N_2129);
xor U2265 (N_2265,N_2171,N_2021);
xnor U2266 (N_2266,N_2141,N_2064);
nor U2267 (N_2267,N_2110,N_2139);
xnor U2268 (N_2268,N_2003,N_2233);
nor U2269 (N_2269,N_2138,N_2150);
and U2270 (N_2270,N_2071,N_2151);
or U2271 (N_2271,N_2157,N_2037);
xnor U2272 (N_2272,N_2245,N_2248);
nand U2273 (N_2273,N_2079,N_2215);
nand U2274 (N_2274,N_2214,N_2193);
and U2275 (N_2275,N_2098,N_2048);
nand U2276 (N_2276,N_2080,N_2180);
and U2277 (N_2277,N_2166,N_2160);
nor U2278 (N_2278,N_2220,N_2238);
nand U2279 (N_2279,N_2042,N_2173);
nand U2280 (N_2280,N_2022,N_2216);
and U2281 (N_2281,N_2190,N_2073);
nor U2282 (N_2282,N_2096,N_2165);
nand U2283 (N_2283,N_2192,N_2212);
xor U2284 (N_2284,N_2132,N_2197);
xnor U2285 (N_2285,N_2047,N_2038);
nand U2286 (N_2286,N_2230,N_2117);
or U2287 (N_2287,N_2170,N_2225);
nor U2288 (N_2288,N_2075,N_2130);
and U2289 (N_2289,N_2217,N_2135);
xnor U2290 (N_2290,N_2128,N_2020);
xor U2291 (N_2291,N_2218,N_2155);
nor U2292 (N_2292,N_2046,N_2202);
xnor U2293 (N_2293,N_2234,N_2224);
or U2294 (N_2294,N_2205,N_2176);
or U2295 (N_2295,N_2068,N_2229);
nor U2296 (N_2296,N_2179,N_2070);
and U2297 (N_2297,N_2201,N_2018);
nand U2298 (N_2298,N_2090,N_2158);
and U2299 (N_2299,N_2199,N_2107);
and U2300 (N_2300,N_2161,N_2102);
and U2301 (N_2301,N_2148,N_2186);
nand U2302 (N_2302,N_2143,N_2231);
nand U2303 (N_2303,N_2236,N_2085);
nor U2304 (N_2304,N_2050,N_2164);
nor U2305 (N_2305,N_2174,N_2108);
or U2306 (N_2306,N_2188,N_2087);
nor U2307 (N_2307,N_2089,N_2007);
or U2308 (N_2308,N_2065,N_2097);
nand U2309 (N_2309,N_2140,N_2126);
and U2310 (N_2310,N_2226,N_2082);
and U2311 (N_2311,N_2222,N_2010);
nand U2312 (N_2312,N_2028,N_2228);
and U2313 (N_2313,N_2105,N_2168);
and U2314 (N_2314,N_2103,N_2206);
and U2315 (N_2315,N_2059,N_2112);
or U2316 (N_2316,N_2039,N_2088);
or U2317 (N_2317,N_2178,N_2169);
xor U2318 (N_2318,N_2172,N_2241);
or U2319 (N_2319,N_2145,N_2083);
or U2320 (N_2320,N_2040,N_2014);
or U2321 (N_2321,N_2019,N_2009);
nand U2322 (N_2322,N_2211,N_2077);
nor U2323 (N_2323,N_2031,N_2005);
nand U2324 (N_2324,N_2024,N_2122);
and U2325 (N_2325,N_2060,N_2147);
and U2326 (N_2326,N_2227,N_2136);
nand U2327 (N_2327,N_2041,N_2081);
and U2328 (N_2328,N_2146,N_2049);
xnor U2329 (N_2329,N_2115,N_2191);
nor U2330 (N_2330,N_2091,N_2247);
or U2331 (N_2331,N_2175,N_2006);
xnor U2332 (N_2332,N_2034,N_2099);
nand U2333 (N_2333,N_2194,N_2052);
and U2334 (N_2334,N_2149,N_2240);
nor U2335 (N_2335,N_2008,N_2134);
and U2336 (N_2336,N_2044,N_2154);
or U2337 (N_2337,N_2053,N_2210);
and U2338 (N_2338,N_2219,N_2235);
nor U2339 (N_2339,N_2237,N_2051);
nand U2340 (N_2340,N_2012,N_2004);
or U2341 (N_2341,N_2058,N_2062);
and U2342 (N_2342,N_2159,N_2133);
or U2343 (N_2343,N_2033,N_2162);
nor U2344 (N_2344,N_2011,N_2124);
or U2345 (N_2345,N_2092,N_2209);
nand U2346 (N_2346,N_2036,N_2183);
nand U2347 (N_2347,N_2184,N_2055);
and U2348 (N_2348,N_2242,N_2137);
and U2349 (N_2349,N_2144,N_2063);
xnor U2350 (N_2350,N_2016,N_2114);
nand U2351 (N_2351,N_2113,N_2000);
and U2352 (N_2352,N_2223,N_2181);
nor U2353 (N_2353,N_2101,N_2119);
and U2354 (N_2354,N_2074,N_2185);
and U2355 (N_2355,N_2025,N_2106);
or U2356 (N_2356,N_2246,N_2116);
and U2357 (N_2357,N_2207,N_2208);
and U2358 (N_2358,N_2232,N_2086);
nand U2359 (N_2359,N_2030,N_2120);
nand U2360 (N_2360,N_2069,N_2013);
nor U2361 (N_2361,N_2189,N_2204);
nor U2362 (N_2362,N_2163,N_2123);
xor U2363 (N_2363,N_2152,N_2131);
nand U2364 (N_2364,N_2125,N_2057);
xor U2365 (N_2365,N_2094,N_2078);
nor U2366 (N_2366,N_2002,N_2244);
nand U2367 (N_2367,N_2043,N_2196);
nor U2368 (N_2368,N_2177,N_2023);
or U2369 (N_2369,N_2001,N_2084);
or U2370 (N_2370,N_2015,N_2221);
or U2371 (N_2371,N_2142,N_2109);
nor U2372 (N_2372,N_2093,N_2035);
xor U2373 (N_2373,N_2200,N_2072);
xnor U2374 (N_2374,N_2121,N_2100);
nand U2375 (N_2375,N_2040,N_2168);
nor U2376 (N_2376,N_2156,N_2102);
or U2377 (N_2377,N_2063,N_2109);
and U2378 (N_2378,N_2224,N_2185);
xnor U2379 (N_2379,N_2026,N_2196);
xnor U2380 (N_2380,N_2222,N_2116);
or U2381 (N_2381,N_2065,N_2163);
or U2382 (N_2382,N_2103,N_2186);
xor U2383 (N_2383,N_2032,N_2149);
and U2384 (N_2384,N_2161,N_2181);
xor U2385 (N_2385,N_2061,N_2098);
xnor U2386 (N_2386,N_2060,N_2107);
and U2387 (N_2387,N_2007,N_2181);
nor U2388 (N_2388,N_2183,N_2151);
or U2389 (N_2389,N_2115,N_2165);
nand U2390 (N_2390,N_2072,N_2217);
xnor U2391 (N_2391,N_2142,N_2111);
and U2392 (N_2392,N_2144,N_2013);
nor U2393 (N_2393,N_2171,N_2137);
xnor U2394 (N_2394,N_2167,N_2120);
nand U2395 (N_2395,N_2217,N_2079);
nand U2396 (N_2396,N_2089,N_2092);
and U2397 (N_2397,N_2122,N_2220);
or U2398 (N_2398,N_2201,N_2112);
or U2399 (N_2399,N_2018,N_2239);
or U2400 (N_2400,N_2109,N_2059);
xor U2401 (N_2401,N_2113,N_2039);
nor U2402 (N_2402,N_2006,N_2126);
nand U2403 (N_2403,N_2245,N_2008);
xnor U2404 (N_2404,N_2160,N_2105);
or U2405 (N_2405,N_2124,N_2238);
or U2406 (N_2406,N_2234,N_2073);
xnor U2407 (N_2407,N_2008,N_2152);
xnor U2408 (N_2408,N_2150,N_2231);
nor U2409 (N_2409,N_2247,N_2050);
or U2410 (N_2410,N_2241,N_2243);
or U2411 (N_2411,N_2113,N_2187);
xnor U2412 (N_2412,N_2038,N_2085);
xor U2413 (N_2413,N_2043,N_2044);
and U2414 (N_2414,N_2113,N_2008);
xnor U2415 (N_2415,N_2246,N_2012);
nor U2416 (N_2416,N_2129,N_2015);
nand U2417 (N_2417,N_2057,N_2005);
and U2418 (N_2418,N_2228,N_2186);
and U2419 (N_2419,N_2244,N_2171);
nor U2420 (N_2420,N_2129,N_2192);
xnor U2421 (N_2421,N_2047,N_2235);
nor U2422 (N_2422,N_2238,N_2142);
or U2423 (N_2423,N_2199,N_2095);
or U2424 (N_2424,N_2046,N_2173);
xor U2425 (N_2425,N_2228,N_2046);
xor U2426 (N_2426,N_2239,N_2159);
xnor U2427 (N_2427,N_2068,N_2116);
xnor U2428 (N_2428,N_2139,N_2119);
nor U2429 (N_2429,N_2031,N_2049);
xnor U2430 (N_2430,N_2090,N_2213);
or U2431 (N_2431,N_2023,N_2142);
nand U2432 (N_2432,N_2053,N_2044);
xor U2433 (N_2433,N_2027,N_2057);
xor U2434 (N_2434,N_2113,N_2074);
xnor U2435 (N_2435,N_2113,N_2018);
and U2436 (N_2436,N_2092,N_2123);
and U2437 (N_2437,N_2194,N_2004);
or U2438 (N_2438,N_2107,N_2157);
and U2439 (N_2439,N_2241,N_2031);
nor U2440 (N_2440,N_2002,N_2115);
or U2441 (N_2441,N_2021,N_2206);
nand U2442 (N_2442,N_2219,N_2171);
nor U2443 (N_2443,N_2040,N_2046);
nand U2444 (N_2444,N_2164,N_2103);
and U2445 (N_2445,N_2176,N_2112);
or U2446 (N_2446,N_2055,N_2052);
or U2447 (N_2447,N_2045,N_2018);
and U2448 (N_2448,N_2014,N_2161);
and U2449 (N_2449,N_2146,N_2170);
xnor U2450 (N_2450,N_2215,N_2248);
and U2451 (N_2451,N_2024,N_2135);
or U2452 (N_2452,N_2016,N_2029);
and U2453 (N_2453,N_2182,N_2232);
or U2454 (N_2454,N_2214,N_2146);
or U2455 (N_2455,N_2048,N_2185);
nor U2456 (N_2456,N_2004,N_2023);
xor U2457 (N_2457,N_2136,N_2014);
nor U2458 (N_2458,N_2158,N_2036);
nor U2459 (N_2459,N_2226,N_2154);
xnor U2460 (N_2460,N_2121,N_2098);
xor U2461 (N_2461,N_2015,N_2234);
xor U2462 (N_2462,N_2041,N_2118);
and U2463 (N_2463,N_2057,N_2213);
nor U2464 (N_2464,N_2243,N_2150);
xnor U2465 (N_2465,N_2200,N_2047);
and U2466 (N_2466,N_2051,N_2180);
or U2467 (N_2467,N_2112,N_2190);
and U2468 (N_2468,N_2213,N_2155);
or U2469 (N_2469,N_2231,N_2065);
or U2470 (N_2470,N_2186,N_2003);
and U2471 (N_2471,N_2157,N_2244);
and U2472 (N_2472,N_2096,N_2027);
and U2473 (N_2473,N_2083,N_2089);
and U2474 (N_2474,N_2085,N_2242);
xnor U2475 (N_2475,N_2084,N_2121);
or U2476 (N_2476,N_2061,N_2123);
nor U2477 (N_2477,N_2049,N_2201);
and U2478 (N_2478,N_2032,N_2028);
and U2479 (N_2479,N_2220,N_2098);
or U2480 (N_2480,N_2024,N_2109);
nand U2481 (N_2481,N_2054,N_2177);
xnor U2482 (N_2482,N_2144,N_2016);
and U2483 (N_2483,N_2180,N_2134);
xnor U2484 (N_2484,N_2237,N_2155);
and U2485 (N_2485,N_2080,N_2104);
nor U2486 (N_2486,N_2154,N_2014);
nand U2487 (N_2487,N_2163,N_2176);
nor U2488 (N_2488,N_2077,N_2178);
nor U2489 (N_2489,N_2081,N_2178);
and U2490 (N_2490,N_2136,N_2184);
and U2491 (N_2491,N_2009,N_2113);
and U2492 (N_2492,N_2169,N_2224);
xor U2493 (N_2493,N_2077,N_2146);
xor U2494 (N_2494,N_2117,N_2237);
xnor U2495 (N_2495,N_2231,N_2014);
nor U2496 (N_2496,N_2195,N_2071);
nor U2497 (N_2497,N_2039,N_2067);
nor U2498 (N_2498,N_2104,N_2020);
xnor U2499 (N_2499,N_2132,N_2242);
nor U2500 (N_2500,N_2270,N_2259);
and U2501 (N_2501,N_2261,N_2316);
nor U2502 (N_2502,N_2306,N_2310);
xnor U2503 (N_2503,N_2326,N_2444);
nor U2504 (N_2504,N_2313,N_2395);
or U2505 (N_2505,N_2285,N_2278);
or U2506 (N_2506,N_2373,N_2391);
xor U2507 (N_2507,N_2354,N_2355);
nor U2508 (N_2508,N_2488,N_2277);
nand U2509 (N_2509,N_2400,N_2311);
nor U2510 (N_2510,N_2439,N_2365);
nand U2511 (N_2511,N_2468,N_2429);
nor U2512 (N_2512,N_2297,N_2383);
nand U2513 (N_2513,N_2472,N_2476);
xor U2514 (N_2514,N_2369,N_2340);
xnor U2515 (N_2515,N_2454,N_2352);
xor U2516 (N_2516,N_2392,N_2314);
nand U2517 (N_2517,N_2327,N_2304);
and U2518 (N_2518,N_2403,N_2273);
nor U2519 (N_2519,N_2371,N_2457);
or U2520 (N_2520,N_2492,N_2417);
or U2521 (N_2521,N_2484,N_2428);
or U2522 (N_2522,N_2296,N_2330);
and U2523 (N_2523,N_2412,N_2291);
or U2524 (N_2524,N_2455,N_2471);
nor U2525 (N_2525,N_2345,N_2299);
nor U2526 (N_2526,N_2387,N_2290);
nand U2527 (N_2527,N_2328,N_2287);
or U2528 (N_2528,N_2267,N_2325);
or U2529 (N_2529,N_2293,N_2350);
xnor U2530 (N_2530,N_2493,N_2446);
or U2531 (N_2531,N_2498,N_2425);
and U2532 (N_2532,N_2307,N_2463);
or U2533 (N_2533,N_2443,N_2283);
xor U2534 (N_2534,N_2281,N_2478);
xnor U2535 (N_2535,N_2384,N_2434);
xnor U2536 (N_2536,N_2436,N_2253);
xnor U2537 (N_2537,N_2295,N_2449);
nor U2538 (N_2538,N_2333,N_2265);
xor U2539 (N_2539,N_2335,N_2289);
nand U2540 (N_2540,N_2469,N_2301);
nand U2541 (N_2541,N_2324,N_2349);
nand U2542 (N_2542,N_2258,N_2421);
nand U2543 (N_2543,N_2275,N_2423);
nor U2544 (N_2544,N_2474,N_2441);
and U2545 (N_2545,N_2485,N_2359);
and U2546 (N_2546,N_2389,N_2491);
nor U2547 (N_2547,N_2495,N_2440);
or U2548 (N_2548,N_2336,N_2338);
or U2549 (N_2549,N_2347,N_2450);
xor U2550 (N_2550,N_2442,N_2264);
nand U2551 (N_2551,N_2317,N_2433);
and U2552 (N_2552,N_2368,N_2353);
xor U2553 (N_2553,N_2394,N_2416);
and U2554 (N_2554,N_2451,N_2453);
nand U2555 (N_2555,N_2305,N_2276);
nand U2556 (N_2556,N_2378,N_2381);
and U2557 (N_2557,N_2464,N_2319);
and U2558 (N_2558,N_2424,N_2407);
and U2559 (N_2559,N_2271,N_2462);
xnor U2560 (N_2560,N_2377,N_2385);
or U2561 (N_2561,N_2337,N_2320);
or U2562 (N_2562,N_2380,N_2358);
xnor U2563 (N_2563,N_2375,N_2419);
xnor U2564 (N_2564,N_2410,N_2279);
or U2565 (N_2565,N_2481,N_2360);
and U2566 (N_2566,N_2362,N_2448);
and U2567 (N_2567,N_2399,N_2386);
or U2568 (N_2568,N_2272,N_2432);
or U2569 (N_2569,N_2366,N_2318);
or U2570 (N_2570,N_2351,N_2341);
nor U2571 (N_2571,N_2300,N_2339);
and U2572 (N_2572,N_2342,N_2269);
nand U2573 (N_2573,N_2274,N_2466);
nand U2574 (N_2574,N_2256,N_2370);
nand U2575 (N_2575,N_2308,N_2262);
nand U2576 (N_2576,N_2334,N_2458);
and U2577 (N_2577,N_2251,N_2465);
nor U2578 (N_2578,N_2376,N_2483);
nor U2579 (N_2579,N_2332,N_2361);
nor U2580 (N_2580,N_2418,N_2288);
nand U2581 (N_2581,N_2401,N_2393);
or U2582 (N_2582,N_2479,N_2286);
nand U2583 (N_2583,N_2315,N_2367);
xnor U2584 (N_2584,N_2473,N_2427);
xor U2585 (N_2585,N_2266,N_2348);
nor U2586 (N_2586,N_2430,N_2363);
or U2587 (N_2587,N_2250,N_2344);
nor U2588 (N_2588,N_2294,N_2343);
or U2589 (N_2589,N_2411,N_2437);
or U2590 (N_2590,N_2438,N_2292);
or U2591 (N_2591,N_2382,N_2257);
nor U2592 (N_2592,N_2467,N_2379);
nand U2593 (N_2593,N_2452,N_2475);
or U2594 (N_2594,N_2331,N_2426);
or U2595 (N_2595,N_2388,N_2357);
nand U2596 (N_2596,N_2477,N_2435);
nand U2597 (N_2597,N_2482,N_2499);
nor U2598 (N_2598,N_2490,N_2497);
xnor U2599 (N_2599,N_2398,N_2397);
nand U2600 (N_2600,N_2461,N_2284);
nand U2601 (N_2601,N_2260,N_2406);
nor U2602 (N_2602,N_2323,N_2364);
nand U2603 (N_2603,N_2329,N_2303);
nand U2604 (N_2604,N_2494,N_2254);
nand U2605 (N_2605,N_2470,N_2486);
nor U2606 (N_2606,N_2346,N_2496);
nor U2607 (N_2607,N_2302,N_2396);
and U2608 (N_2608,N_2489,N_2356);
and U2609 (N_2609,N_2280,N_2447);
and U2610 (N_2610,N_2420,N_2414);
and U2611 (N_2611,N_2322,N_2445);
nor U2612 (N_2612,N_2268,N_2390);
and U2613 (N_2613,N_2298,N_2422);
xor U2614 (N_2614,N_2456,N_2409);
or U2615 (N_2615,N_2413,N_2408);
or U2616 (N_2616,N_2321,N_2460);
and U2617 (N_2617,N_2405,N_2263);
nand U2618 (N_2618,N_2309,N_2404);
xnor U2619 (N_2619,N_2415,N_2402);
nor U2620 (N_2620,N_2374,N_2282);
xor U2621 (N_2621,N_2431,N_2459);
nand U2622 (N_2622,N_2480,N_2252);
or U2623 (N_2623,N_2255,N_2372);
or U2624 (N_2624,N_2487,N_2312);
xor U2625 (N_2625,N_2386,N_2480);
and U2626 (N_2626,N_2368,N_2269);
or U2627 (N_2627,N_2288,N_2305);
and U2628 (N_2628,N_2452,N_2430);
xnor U2629 (N_2629,N_2411,N_2266);
or U2630 (N_2630,N_2324,N_2252);
nor U2631 (N_2631,N_2349,N_2439);
xor U2632 (N_2632,N_2459,N_2303);
xor U2633 (N_2633,N_2488,N_2289);
xor U2634 (N_2634,N_2399,N_2495);
nor U2635 (N_2635,N_2494,N_2289);
nand U2636 (N_2636,N_2481,N_2433);
and U2637 (N_2637,N_2404,N_2301);
and U2638 (N_2638,N_2272,N_2455);
and U2639 (N_2639,N_2418,N_2341);
xnor U2640 (N_2640,N_2443,N_2280);
nand U2641 (N_2641,N_2473,N_2482);
nor U2642 (N_2642,N_2308,N_2309);
or U2643 (N_2643,N_2276,N_2362);
nor U2644 (N_2644,N_2332,N_2381);
nor U2645 (N_2645,N_2437,N_2442);
nor U2646 (N_2646,N_2356,N_2292);
or U2647 (N_2647,N_2283,N_2323);
and U2648 (N_2648,N_2403,N_2385);
and U2649 (N_2649,N_2497,N_2483);
and U2650 (N_2650,N_2339,N_2452);
xor U2651 (N_2651,N_2325,N_2316);
nand U2652 (N_2652,N_2471,N_2380);
and U2653 (N_2653,N_2481,N_2380);
nand U2654 (N_2654,N_2288,N_2372);
and U2655 (N_2655,N_2499,N_2429);
or U2656 (N_2656,N_2296,N_2324);
and U2657 (N_2657,N_2370,N_2265);
nor U2658 (N_2658,N_2372,N_2461);
nor U2659 (N_2659,N_2351,N_2432);
nand U2660 (N_2660,N_2330,N_2301);
and U2661 (N_2661,N_2406,N_2453);
or U2662 (N_2662,N_2383,N_2470);
and U2663 (N_2663,N_2498,N_2268);
nand U2664 (N_2664,N_2421,N_2351);
and U2665 (N_2665,N_2285,N_2462);
xnor U2666 (N_2666,N_2466,N_2474);
nor U2667 (N_2667,N_2413,N_2345);
nand U2668 (N_2668,N_2300,N_2277);
nor U2669 (N_2669,N_2418,N_2431);
and U2670 (N_2670,N_2352,N_2253);
and U2671 (N_2671,N_2489,N_2325);
xnor U2672 (N_2672,N_2265,N_2473);
nand U2673 (N_2673,N_2291,N_2476);
or U2674 (N_2674,N_2257,N_2338);
nor U2675 (N_2675,N_2457,N_2362);
or U2676 (N_2676,N_2471,N_2322);
and U2677 (N_2677,N_2462,N_2289);
nand U2678 (N_2678,N_2428,N_2452);
nand U2679 (N_2679,N_2303,N_2498);
nand U2680 (N_2680,N_2494,N_2472);
nor U2681 (N_2681,N_2446,N_2261);
and U2682 (N_2682,N_2424,N_2342);
and U2683 (N_2683,N_2434,N_2268);
and U2684 (N_2684,N_2452,N_2410);
xor U2685 (N_2685,N_2274,N_2485);
and U2686 (N_2686,N_2401,N_2457);
and U2687 (N_2687,N_2312,N_2481);
nand U2688 (N_2688,N_2378,N_2459);
nor U2689 (N_2689,N_2304,N_2388);
or U2690 (N_2690,N_2305,N_2253);
nand U2691 (N_2691,N_2428,N_2397);
or U2692 (N_2692,N_2293,N_2433);
nor U2693 (N_2693,N_2495,N_2386);
xor U2694 (N_2694,N_2487,N_2275);
or U2695 (N_2695,N_2490,N_2264);
xor U2696 (N_2696,N_2453,N_2314);
nand U2697 (N_2697,N_2277,N_2431);
nand U2698 (N_2698,N_2433,N_2355);
xnor U2699 (N_2699,N_2321,N_2287);
xnor U2700 (N_2700,N_2481,N_2276);
or U2701 (N_2701,N_2498,N_2437);
nor U2702 (N_2702,N_2286,N_2342);
nand U2703 (N_2703,N_2289,N_2452);
nor U2704 (N_2704,N_2339,N_2384);
and U2705 (N_2705,N_2341,N_2465);
and U2706 (N_2706,N_2353,N_2485);
nor U2707 (N_2707,N_2266,N_2359);
nand U2708 (N_2708,N_2342,N_2431);
nor U2709 (N_2709,N_2384,N_2331);
nand U2710 (N_2710,N_2347,N_2448);
nor U2711 (N_2711,N_2495,N_2336);
or U2712 (N_2712,N_2420,N_2369);
and U2713 (N_2713,N_2474,N_2418);
nor U2714 (N_2714,N_2294,N_2338);
xnor U2715 (N_2715,N_2308,N_2340);
nor U2716 (N_2716,N_2329,N_2301);
nand U2717 (N_2717,N_2259,N_2385);
and U2718 (N_2718,N_2299,N_2464);
or U2719 (N_2719,N_2272,N_2453);
and U2720 (N_2720,N_2264,N_2479);
nand U2721 (N_2721,N_2492,N_2433);
nand U2722 (N_2722,N_2487,N_2315);
xor U2723 (N_2723,N_2407,N_2281);
xor U2724 (N_2724,N_2283,N_2499);
nand U2725 (N_2725,N_2426,N_2261);
nor U2726 (N_2726,N_2256,N_2267);
nor U2727 (N_2727,N_2494,N_2403);
nand U2728 (N_2728,N_2389,N_2467);
and U2729 (N_2729,N_2369,N_2260);
or U2730 (N_2730,N_2363,N_2324);
nor U2731 (N_2731,N_2449,N_2354);
and U2732 (N_2732,N_2489,N_2309);
or U2733 (N_2733,N_2330,N_2408);
nor U2734 (N_2734,N_2264,N_2390);
or U2735 (N_2735,N_2468,N_2304);
nand U2736 (N_2736,N_2280,N_2413);
or U2737 (N_2737,N_2375,N_2328);
nor U2738 (N_2738,N_2404,N_2275);
nand U2739 (N_2739,N_2411,N_2498);
or U2740 (N_2740,N_2336,N_2324);
nand U2741 (N_2741,N_2341,N_2261);
or U2742 (N_2742,N_2270,N_2388);
nor U2743 (N_2743,N_2316,N_2466);
and U2744 (N_2744,N_2490,N_2393);
and U2745 (N_2745,N_2323,N_2419);
nand U2746 (N_2746,N_2374,N_2312);
and U2747 (N_2747,N_2380,N_2493);
nand U2748 (N_2748,N_2370,N_2446);
or U2749 (N_2749,N_2434,N_2386);
nand U2750 (N_2750,N_2724,N_2596);
and U2751 (N_2751,N_2642,N_2500);
or U2752 (N_2752,N_2575,N_2705);
xor U2753 (N_2753,N_2628,N_2540);
and U2754 (N_2754,N_2546,N_2733);
and U2755 (N_2755,N_2521,N_2542);
and U2756 (N_2756,N_2600,N_2523);
and U2757 (N_2757,N_2676,N_2688);
and U2758 (N_2758,N_2608,N_2515);
nand U2759 (N_2759,N_2585,N_2650);
and U2760 (N_2760,N_2667,N_2633);
and U2761 (N_2761,N_2597,N_2537);
nor U2762 (N_2762,N_2513,N_2729);
or U2763 (N_2763,N_2570,N_2594);
or U2764 (N_2764,N_2602,N_2538);
nor U2765 (N_2765,N_2530,N_2639);
nor U2766 (N_2766,N_2566,N_2719);
and U2767 (N_2767,N_2534,N_2535);
nand U2768 (N_2768,N_2731,N_2624);
or U2769 (N_2769,N_2657,N_2691);
nor U2770 (N_2770,N_2647,N_2630);
and U2771 (N_2771,N_2622,N_2710);
xor U2772 (N_2772,N_2584,N_2548);
nand U2773 (N_2773,N_2727,N_2663);
nand U2774 (N_2774,N_2562,N_2581);
nor U2775 (N_2775,N_2576,N_2745);
or U2776 (N_2776,N_2699,N_2524);
nand U2777 (N_2777,N_2675,N_2531);
xnor U2778 (N_2778,N_2735,N_2553);
nand U2779 (N_2779,N_2591,N_2682);
xor U2780 (N_2780,N_2641,N_2545);
nor U2781 (N_2781,N_2681,N_2595);
nor U2782 (N_2782,N_2666,N_2572);
and U2783 (N_2783,N_2627,N_2607);
nand U2784 (N_2784,N_2592,N_2706);
or U2785 (N_2785,N_2571,N_2656);
and U2786 (N_2786,N_2632,N_2559);
nor U2787 (N_2787,N_2687,N_2744);
or U2788 (N_2788,N_2659,N_2560);
nor U2789 (N_2789,N_2520,N_2668);
and U2790 (N_2790,N_2723,N_2673);
or U2791 (N_2791,N_2509,N_2743);
and U2792 (N_2792,N_2708,N_2617);
or U2793 (N_2793,N_2590,N_2611);
xnor U2794 (N_2794,N_2737,N_2718);
nor U2795 (N_2795,N_2544,N_2685);
or U2796 (N_2796,N_2589,N_2533);
or U2797 (N_2797,N_2670,N_2742);
nor U2798 (N_2798,N_2623,N_2721);
xor U2799 (N_2799,N_2720,N_2736);
and U2800 (N_2800,N_2514,N_2651);
nor U2801 (N_2801,N_2504,N_2644);
nor U2802 (N_2802,N_2717,N_2588);
or U2803 (N_2803,N_2665,N_2722);
xnor U2804 (N_2804,N_2715,N_2629);
nor U2805 (N_2805,N_2646,N_2679);
nand U2806 (N_2806,N_2558,N_2728);
xor U2807 (N_2807,N_2716,N_2634);
and U2808 (N_2808,N_2677,N_2539);
or U2809 (N_2809,N_2714,N_2583);
xnor U2810 (N_2810,N_2525,N_2577);
and U2811 (N_2811,N_2740,N_2606);
and U2812 (N_2812,N_2593,N_2614);
nand U2813 (N_2813,N_2598,N_2662);
and U2814 (N_2814,N_2746,N_2635);
or U2815 (N_2815,N_2703,N_2574);
xor U2816 (N_2816,N_2686,N_2637);
and U2817 (N_2817,N_2519,N_2573);
nor U2818 (N_2818,N_2610,N_2726);
and U2819 (N_2819,N_2700,N_2587);
or U2820 (N_2820,N_2604,N_2749);
nand U2821 (N_2821,N_2653,N_2618);
nand U2822 (N_2822,N_2620,N_2701);
nor U2823 (N_2823,N_2506,N_2582);
or U2824 (N_2824,N_2580,N_2510);
xor U2825 (N_2825,N_2536,N_2517);
xor U2826 (N_2826,N_2696,N_2730);
nor U2827 (N_2827,N_2645,N_2569);
nand U2828 (N_2828,N_2664,N_2543);
or U2829 (N_2829,N_2621,N_2601);
nor U2830 (N_2830,N_2612,N_2599);
nand U2831 (N_2831,N_2615,N_2638);
or U2832 (N_2832,N_2625,N_2552);
xnor U2833 (N_2833,N_2528,N_2511);
nand U2834 (N_2834,N_2516,N_2563);
or U2835 (N_2835,N_2551,N_2660);
and U2836 (N_2836,N_2671,N_2564);
nand U2837 (N_2837,N_2565,N_2672);
nand U2838 (N_2838,N_2549,N_2655);
or U2839 (N_2839,N_2502,N_2561);
and U2840 (N_2840,N_2661,N_2636);
and U2841 (N_2841,N_2711,N_2674);
nand U2842 (N_2842,N_2709,N_2693);
xnor U2843 (N_2843,N_2609,N_2669);
nand U2844 (N_2844,N_2555,N_2678);
nand U2845 (N_2845,N_2527,N_2748);
or U2846 (N_2846,N_2725,N_2526);
or U2847 (N_2847,N_2713,N_2532);
nand U2848 (N_2848,N_2626,N_2586);
nor U2849 (N_2849,N_2554,N_2738);
nor U2850 (N_2850,N_2658,N_2613);
xor U2851 (N_2851,N_2652,N_2603);
xor U2852 (N_2852,N_2567,N_2689);
nor U2853 (N_2853,N_2707,N_2648);
and U2854 (N_2854,N_2690,N_2508);
or U2855 (N_2855,N_2694,N_2654);
xor U2856 (N_2856,N_2579,N_2732);
and U2857 (N_2857,N_2692,N_2578);
and U2858 (N_2858,N_2512,N_2683);
or U2859 (N_2859,N_2643,N_2529);
or U2860 (N_2860,N_2684,N_2503);
or U2861 (N_2861,N_2507,N_2739);
xnor U2862 (N_2862,N_2702,N_2501);
nand U2863 (N_2863,N_2695,N_2547);
or U2864 (N_2864,N_2616,N_2568);
and U2865 (N_2865,N_2680,N_2631);
and U2866 (N_2866,N_2550,N_2741);
nor U2867 (N_2867,N_2518,N_2522);
or U2868 (N_2868,N_2605,N_2704);
nand U2869 (N_2869,N_2712,N_2640);
nor U2870 (N_2870,N_2734,N_2698);
or U2871 (N_2871,N_2541,N_2619);
nor U2872 (N_2872,N_2556,N_2649);
and U2873 (N_2873,N_2747,N_2505);
and U2874 (N_2874,N_2557,N_2697);
nand U2875 (N_2875,N_2588,N_2531);
or U2876 (N_2876,N_2590,N_2638);
nand U2877 (N_2877,N_2573,N_2593);
nand U2878 (N_2878,N_2620,N_2729);
or U2879 (N_2879,N_2689,N_2589);
and U2880 (N_2880,N_2631,N_2679);
or U2881 (N_2881,N_2731,N_2522);
and U2882 (N_2882,N_2547,N_2724);
xor U2883 (N_2883,N_2585,N_2596);
nor U2884 (N_2884,N_2639,N_2583);
or U2885 (N_2885,N_2706,N_2601);
nor U2886 (N_2886,N_2648,N_2552);
or U2887 (N_2887,N_2540,N_2600);
nand U2888 (N_2888,N_2529,N_2609);
xor U2889 (N_2889,N_2532,N_2638);
xnor U2890 (N_2890,N_2508,N_2595);
nand U2891 (N_2891,N_2517,N_2526);
and U2892 (N_2892,N_2524,N_2655);
nand U2893 (N_2893,N_2685,N_2717);
or U2894 (N_2894,N_2624,N_2550);
nand U2895 (N_2895,N_2531,N_2639);
and U2896 (N_2896,N_2710,N_2736);
xor U2897 (N_2897,N_2695,N_2571);
or U2898 (N_2898,N_2546,N_2621);
nand U2899 (N_2899,N_2748,N_2534);
nor U2900 (N_2900,N_2525,N_2745);
nor U2901 (N_2901,N_2708,N_2620);
nand U2902 (N_2902,N_2717,N_2653);
xnor U2903 (N_2903,N_2613,N_2557);
or U2904 (N_2904,N_2517,N_2621);
nand U2905 (N_2905,N_2549,N_2711);
or U2906 (N_2906,N_2702,N_2597);
nor U2907 (N_2907,N_2741,N_2690);
or U2908 (N_2908,N_2630,N_2625);
and U2909 (N_2909,N_2603,N_2551);
or U2910 (N_2910,N_2647,N_2611);
nor U2911 (N_2911,N_2594,N_2737);
or U2912 (N_2912,N_2574,N_2647);
xor U2913 (N_2913,N_2610,N_2510);
xor U2914 (N_2914,N_2570,N_2520);
nor U2915 (N_2915,N_2650,N_2676);
nand U2916 (N_2916,N_2652,N_2530);
nor U2917 (N_2917,N_2523,N_2700);
and U2918 (N_2918,N_2673,N_2613);
or U2919 (N_2919,N_2532,N_2673);
nand U2920 (N_2920,N_2746,N_2656);
and U2921 (N_2921,N_2608,N_2703);
or U2922 (N_2922,N_2730,N_2601);
nand U2923 (N_2923,N_2652,N_2537);
nand U2924 (N_2924,N_2710,N_2707);
nor U2925 (N_2925,N_2511,N_2715);
nand U2926 (N_2926,N_2647,N_2534);
nand U2927 (N_2927,N_2597,N_2727);
nor U2928 (N_2928,N_2672,N_2688);
nand U2929 (N_2929,N_2652,N_2687);
xnor U2930 (N_2930,N_2700,N_2534);
or U2931 (N_2931,N_2569,N_2626);
xnor U2932 (N_2932,N_2698,N_2696);
nand U2933 (N_2933,N_2552,N_2509);
or U2934 (N_2934,N_2722,N_2682);
nor U2935 (N_2935,N_2510,N_2743);
or U2936 (N_2936,N_2606,N_2641);
and U2937 (N_2937,N_2538,N_2559);
nor U2938 (N_2938,N_2673,N_2684);
nor U2939 (N_2939,N_2732,N_2567);
nand U2940 (N_2940,N_2545,N_2500);
nor U2941 (N_2941,N_2558,N_2732);
nor U2942 (N_2942,N_2626,N_2614);
or U2943 (N_2943,N_2664,N_2642);
nand U2944 (N_2944,N_2648,N_2614);
nor U2945 (N_2945,N_2566,N_2574);
nor U2946 (N_2946,N_2653,N_2616);
xnor U2947 (N_2947,N_2513,N_2518);
nand U2948 (N_2948,N_2631,N_2616);
and U2949 (N_2949,N_2661,N_2689);
xor U2950 (N_2950,N_2670,N_2521);
and U2951 (N_2951,N_2630,N_2686);
and U2952 (N_2952,N_2661,N_2560);
xor U2953 (N_2953,N_2672,N_2694);
xnor U2954 (N_2954,N_2732,N_2629);
nor U2955 (N_2955,N_2595,N_2711);
nor U2956 (N_2956,N_2525,N_2607);
or U2957 (N_2957,N_2710,N_2550);
xnor U2958 (N_2958,N_2688,N_2578);
and U2959 (N_2959,N_2731,N_2516);
or U2960 (N_2960,N_2631,N_2582);
nor U2961 (N_2961,N_2730,N_2514);
nand U2962 (N_2962,N_2692,N_2548);
nor U2963 (N_2963,N_2634,N_2696);
and U2964 (N_2964,N_2606,N_2508);
and U2965 (N_2965,N_2718,N_2629);
or U2966 (N_2966,N_2544,N_2695);
and U2967 (N_2967,N_2597,N_2566);
and U2968 (N_2968,N_2728,N_2617);
xor U2969 (N_2969,N_2596,N_2645);
or U2970 (N_2970,N_2609,N_2682);
and U2971 (N_2971,N_2710,N_2705);
xnor U2972 (N_2972,N_2737,N_2659);
nand U2973 (N_2973,N_2606,N_2743);
and U2974 (N_2974,N_2622,N_2635);
or U2975 (N_2975,N_2559,N_2687);
and U2976 (N_2976,N_2737,N_2612);
or U2977 (N_2977,N_2546,N_2613);
nor U2978 (N_2978,N_2549,N_2709);
xnor U2979 (N_2979,N_2531,N_2554);
xor U2980 (N_2980,N_2577,N_2734);
and U2981 (N_2981,N_2591,N_2504);
or U2982 (N_2982,N_2589,N_2556);
xor U2983 (N_2983,N_2586,N_2501);
nor U2984 (N_2984,N_2629,N_2702);
or U2985 (N_2985,N_2615,N_2639);
and U2986 (N_2986,N_2636,N_2560);
xor U2987 (N_2987,N_2544,N_2637);
and U2988 (N_2988,N_2614,N_2636);
or U2989 (N_2989,N_2724,N_2673);
or U2990 (N_2990,N_2706,N_2665);
xor U2991 (N_2991,N_2519,N_2557);
xor U2992 (N_2992,N_2546,N_2648);
or U2993 (N_2993,N_2539,N_2721);
or U2994 (N_2994,N_2700,N_2515);
and U2995 (N_2995,N_2671,N_2548);
xnor U2996 (N_2996,N_2571,N_2509);
and U2997 (N_2997,N_2693,N_2705);
and U2998 (N_2998,N_2514,N_2512);
nor U2999 (N_2999,N_2620,N_2549);
nand U3000 (N_3000,N_2961,N_2817);
or U3001 (N_3001,N_2956,N_2971);
or U3002 (N_3002,N_2768,N_2894);
xor U3003 (N_3003,N_2902,N_2857);
and U3004 (N_3004,N_2859,N_2887);
xnor U3005 (N_3005,N_2866,N_2919);
nand U3006 (N_3006,N_2910,N_2984);
xor U3007 (N_3007,N_2875,N_2928);
xor U3008 (N_3008,N_2770,N_2751);
and U3009 (N_3009,N_2931,N_2920);
nor U3010 (N_3010,N_2825,N_2991);
nor U3011 (N_3011,N_2900,N_2889);
nor U3012 (N_3012,N_2898,N_2842);
nand U3013 (N_3013,N_2836,N_2790);
xnor U3014 (N_3014,N_2933,N_2802);
or U3015 (N_3015,N_2819,N_2774);
nand U3016 (N_3016,N_2883,N_2880);
and U3017 (N_3017,N_2840,N_2918);
nand U3018 (N_3018,N_2878,N_2899);
and U3019 (N_3019,N_2917,N_2858);
or U3020 (N_3020,N_2789,N_2929);
xor U3021 (N_3021,N_2766,N_2925);
or U3022 (N_3022,N_2980,N_2785);
and U3023 (N_3023,N_2848,N_2800);
and U3024 (N_3024,N_2916,N_2821);
nor U3025 (N_3025,N_2983,N_2813);
xor U3026 (N_3026,N_2937,N_2822);
and U3027 (N_3027,N_2997,N_2752);
nand U3028 (N_3028,N_2993,N_2870);
and U3029 (N_3029,N_2787,N_2760);
and U3030 (N_3030,N_2950,N_2958);
and U3031 (N_3031,N_2845,N_2903);
and U3032 (N_3032,N_2758,N_2976);
or U3033 (N_3033,N_2773,N_2945);
nand U3034 (N_3034,N_2754,N_2904);
and U3035 (N_3035,N_2776,N_2863);
and U3036 (N_3036,N_2926,N_2882);
or U3037 (N_3037,N_2949,N_2994);
or U3038 (N_3038,N_2869,N_2812);
xnor U3039 (N_3039,N_2818,N_2977);
nor U3040 (N_3040,N_2974,N_2885);
or U3041 (N_3041,N_2884,N_2988);
xnor U3042 (N_3042,N_2943,N_2851);
and U3043 (N_3043,N_2948,N_2951);
xor U3044 (N_3044,N_2820,N_2927);
and U3045 (N_3045,N_2897,N_2811);
nor U3046 (N_3046,N_2890,N_2996);
nor U3047 (N_3047,N_2992,N_2841);
nor U3048 (N_3048,N_2839,N_2987);
and U3049 (N_3049,N_2924,N_2968);
nand U3050 (N_3050,N_2886,N_2816);
and U3051 (N_3051,N_2775,N_2864);
nor U3052 (N_3052,N_2901,N_2786);
nand U3053 (N_3053,N_2922,N_2982);
nand U3054 (N_3054,N_2809,N_2966);
nor U3055 (N_3055,N_2761,N_2962);
xnor U3056 (N_3056,N_2810,N_2844);
xnor U3057 (N_3057,N_2801,N_2762);
and U3058 (N_3058,N_2905,N_2792);
and U3059 (N_3059,N_2893,N_2915);
and U3060 (N_3060,N_2756,N_2941);
or U3061 (N_3061,N_2873,N_2938);
xor U3062 (N_3062,N_2876,N_2759);
nor U3063 (N_3063,N_2995,N_2838);
nand U3064 (N_3064,N_2777,N_2803);
xor U3065 (N_3065,N_2881,N_2835);
xor U3066 (N_3066,N_2856,N_2827);
or U3067 (N_3067,N_2771,N_2763);
and U3068 (N_3068,N_2868,N_2963);
xor U3069 (N_3069,N_2837,N_2755);
and U3070 (N_3070,N_2972,N_2834);
nor U3071 (N_3071,N_2874,N_2940);
nand U3072 (N_3072,N_2824,N_2911);
and U3073 (N_3073,N_2990,N_2794);
nand U3074 (N_3074,N_2796,N_2973);
and U3075 (N_3075,N_2960,N_2872);
and U3076 (N_3076,N_2846,N_2954);
xnor U3077 (N_3077,N_2871,N_2828);
or U3078 (N_3078,N_2781,N_2895);
and U3079 (N_3079,N_2860,N_2877);
and U3080 (N_3080,N_2867,N_2765);
and U3081 (N_3081,N_2935,N_2978);
and U3082 (N_3082,N_2879,N_2831);
xnor U3083 (N_3083,N_2896,N_2823);
nor U3084 (N_3084,N_2830,N_2791);
xnor U3085 (N_3085,N_2942,N_2953);
or U3086 (N_3086,N_2815,N_2964);
nor U3087 (N_3087,N_2850,N_2855);
and U3088 (N_3088,N_2969,N_2783);
xnor U3089 (N_3089,N_2861,N_2797);
nor U3090 (N_3090,N_2772,N_2959);
and U3091 (N_3091,N_2975,N_2967);
nor U3092 (N_3092,N_2930,N_2907);
or U3093 (N_3093,N_2852,N_2753);
nor U3094 (N_3094,N_2798,N_2854);
and U3095 (N_3095,N_2932,N_2936);
nor U3096 (N_3096,N_2769,N_2939);
nor U3097 (N_3097,N_2843,N_2957);
nor U3098 (N_3098,N_2757,N_2833);
xor U3099 (N_3099,N_2805,N_2849);
nand U3100 (N_3100,N_2952,N_2806);
and U3101 (N_3101,N_2970,N_2909);
or U3102 (N_3102,N_2981,N_2853);
xor U3103 (N_3103,N_2788,N_2784);
nor U3104 (N_3104,N_2965,N_2847);
nand U3105 (N_3105,N_2778,N_2906);
and U3106 (N_3106,N_2814,N_2921);
and U3107 (N_3107,N_2764,N_2934);
or U3108 (N_3108,N_2892,N_2807);
nor U3109 (N_3109,N_2914,N_2999);
or U3110 (N_3110,N_2912,N_2750);
nor U3111 (N_3111,N_2829,N_2779);
xor U3112 (N_3112,N_2808,N_2862);
nand U3113 (N_3113,N_2780,N_2986);
xor U3114 (N_3114,N_2782,N_2804);
nor U3115 (N_3115,N_2767,N_2955);
and U3116 (N_3116,N_2913,N_2979);
and U3117 (N_3117,N_2908,N_2923);
nor U3118 (N_3118,N_2998,N_2795);
nand U3119 (N_3119,N_2865,N_2891);
xor U3120 (N_3120,N_2946,N_2793);
or U3121 (N_3121,N_2985,N_2944);
nand U3122 (N_3122,N_2888,N_2826);
xnor U3123 (N_3123,N_2989,N_2832);
nand U3124 (N_3124,N_2799,N_2947);
nor U3125 (N_3125,N_2949,N_2959);
or U3126 (N_3126,N_2761,N_2923);
nand U3127 (N_3127,N_2786,N_2915);
nor U3128 (N_3128,N_2927,N_2857);
nand U3129 (N_3129,N_2905,N_2975);
nor U3130 (N_3130,N_2793,N_2752);
nand U3131 (N_3131,N_2815,N_2906);
or U3132 (N_3132,N_2812,N_2913);
and U3133 (N_3133,N_2752,N_2769);
nor U3134 (N_3134,N_2980,N_2827);
xor U3135 (N_3135,N_2952,N_2858);
nor U3136 (N_3136,N_2859,N_2752);
nor U3137 (N_3137,N_2852,N_2975);
and U3138 (N_3138,N_2945,N_2803);
nand U3139 (N_3139,N_2955,N_2881);
nor U3140 (N_3140,N_2952,N_2889);
nor U3141 (N_3141,N_2803,N_2800);
nand U3142 (N_3142,N_2942,N_2962);
or U3143 (N_3143,N_2823,N_2849);
nand U3144 (N_3144,N_2852,N_2939);
nor U3145 (N_3145,N_2899,N_2841);
xnor U3146 (N_3146,N_2984,N_2955);
or U3147 (N_3147,N_2877,N_2876);
and U3148 (N_3148,N_2789,N_2841);
nor U3149 (N_3149,N_2943,N_2799);
nor U3150 (N_3150,N_2879,N_2885);
and U3151 (N_3151,N_2980,N_2789);
and U3152 (N_3152,N_2761,N_2792);
or U3153 (N_3153,N_2898,N_2783);
nand U3154 (N_3154,N_2995,N_2793);
and U3155 (N_3155,N_2881,N_2799);
and U3156 (N_3156,N_2812,N_2970);
nand U3157 (N_3157,N_2997,N_2888);
nor U3158 (N_3158,N_2765,N_2929);
nor U3159 (N_3159,N_2906,N_2807);
nor U3160 (N_3160,N_2792,N_2811);
and U3161 (N_3161,N_2886,N_2983);
nand U3162 (N_3162,N_2787,N_2942);
xor U3163 (N_3163,N_2848,N_2923);
nand U3164 (N_3164,N_2784,N_2969);
xor U3165 (N_3165,N_2999,N_2870);
nand U3166 (N_3166,N_2963,N_2947);
or U3167 (N_3167,N_2797,N_2958);
or U3168 (N_3168,N_2962,N_2988);
and U3169 (N_3169,N_2855,N_2808);
and U3170 (N_3170,N_2874,N_2934);
xnor U3171 (N_3171,N_2952,N_2894);
or U3172 (N_3172,N_2838,N_2928);
nand U3173 (N_3173,N_2769,N_2796);
and U3174 (N_3174,N_2773,N_2860);
nand U3175 (N_3175,N_2897,N_2914);
nor U3176 (N_3176,N_2944,N_2823);
nand U3177 (N_3177,N_2931,N_2769);
nor U3178 (N_3178,N_2835,N_2808);
or U3179 (N_3179,N_2784,N_2822);
xor U3180 (N_3180,N_2980,N_2891);
nand U3181 (N_3181,N_2862,N_2954);
nand U3182 (N_3182,N_2883,N_2869);
and U3183 (N_3183,N_2789,N_2900);
nor U3184 (N_3184,N_2790,N_2972);
and U3185 (N_3185,N_2995,N_2792);
nand U3186 (N_3186,N_2757,N_2951);
nand U3187 (N_3187,N_2857,N_2787);
and U3188 (N_3188,N_2780,N_2769);
nand U3189 (N_3189,N_2778,N_2788);
nor U3190 (N_3190,N_2812,N_2919);
nor U3191 (N_3191,N_2949,N_2850);
or U3192 (N_3192,N_2945,N_2878);
or U3193 (N_3193,N_2979,N_2751);
xor U3194 (N_3194,N_2869,N_2923);
or U3195 (N_3195,N_2913,N_2900);
nor U3196 (N_3196,N_2814,N_2897);
or U3197 (N_3197,N_2896,N_2970);
or U3198 (N_3198,N_2781,N_2872);
xnor U3199 (N_3199,N_2767,N_2832);
and U3200 (N_3200,N_2978,N_2876);
xnor U3201 (N_3201,N_2854,N_2969);
or U3202 (N_3202,N_2823,N_2804);
and U3203 (N_3203,N_2781,N_2946);
or U3204 (N_3204,N_2997,N_2992);
nand U3205 (N_3205,N_2774,N_2834);
xor U3206 (N_3206,N_2855,N_2893);
nand U3207 (N_3207,N_2796,N_2794);
xor U3208 (N_3208,N_2833,N_2957);
and U3209 (N_3209,N_2993,N_2804);
nor U3210 (N_3210,N_2894,N_2803);
and U3211 (N_3211,N_2868,N_2975);
nand U3212 (N_3212,N_2900,N_2765);
or U3213 (N_3213,N_2834,N_2954);
xnor U3214 (N_3214,N_2963,N_2822);
xor U3215 (N_3215,N_2876,N_2769);
or U3216 (N_3216,N_2856,N_2779);
nand U3217 (N_3217,N_2841,N_2924);
or U3218 (N_3218,N_2983,N_2903);
xor U3219 (N_3219,N_2809,N_2808);
or U3220 (N_3220,N_2984,N_2937);
nand U3221 (N_3221,N_2951,N_2908);
or U3222 (N_3222,N_2842,N_2946);
nand U3223 (N_3223,N_2870,N_2796);
or U3224 (N_3224,N_2977,N_2924);
nand U3225 (N_3225,N_2790,N_2838);
nand U3226 (N_3226,N_2834,N_2979);
and U3227 (N_3227,N_2903,N_2785);
nand U3228 (N_3228,N_2791,N_2950);
nor U3229 (N_3229,N_2899,N_2985);
nor U3230 (N_3230,N_2907,N_2873);
and U3231 (N_3231,N_2840,N_2757);
and U3232 (N_3232,N_2986,N_2844);
xor U3233 (N_3233,N_2929,N_2822);
nand U3234 (N_3234,N_2986,N_2935);
or U3235 (N_3235,N_2833,N_2894);
xnor U3236 (N_3236,N_2914,N_2875);
and U3237 (N_3237,N_2841,N_2838);
nor U3238 (N_3238,N_2766,N_2983);
nand U3239 (N_3239,N_2930,N_2954);
nor U3240 (N_3240,N_2930,N_2939);
or U3241 (N_3241,N_2959,N_2858);
or U3242 (N_3242,N_2932,N_2893);
or U3243 (N_3243,N_2832,N_2869);
or U3244 (N_3244,N_2818,N_2996);
and U3245 (N_3245,N_2773,N_2996);
or U3246 (N_3246,N_2917,N_2759);
or U3247 (N_3247,N_2989,N_2943);
xnor U3248 (N_3248,N_2859,N_2964);
or U3249 (N_3249,N_2887,N_2817);
and U3250 (N_3250,N_3118,N_3164);
and U3251 (N_3251,N_3056,N_3064);
or U3252 (N_3252,N_3035,N_3134);
nor U3253 (N_3253,N_3103,N_3194);
xnor U3254 (N_3254,N_3132,N_3068);
xnor U3255 (N_3255,N_3096,N_3129);
nand U3256 (N_3256,N_3143,N_3127);
and U3257 (N_3257,N_3079,N_3063);
and U3258 (N_3258,N_3201,N_3151);
nor U3259 (N_3259,N_3214,N_3159);
xor U3260 (N_3260,N_3228,N_3128);
nor U3261 (N_3261,N_3115,N_3144);
and U3262 (N_3262,N_3003,N_3177);
nand U3263 (N_3263,N_3012,N_3047);
or U3264 (N_3264,N_3204,N_3091);
nor U3265 (N_3265,N_3211,N_3145);
or U3266 (N_3266,N_3190,N_3046);
xnor U3267 (N_3267,N_3111,N_3087);
or U3268 (N_3268,N_3066,N_3155);
or U3269 (N_3269,N_3113,N_3104);
or U3270 (N_3270,N_3075,N_3095);
or U3271 (N_3271,N_3098,N_3033);
or U3272 (N_3272,N_3017,N_3153);
nor U3273 (N_3273,N_3168,N_3061);
nor U3274 (N_3274,N_3001,N_3059);
nand U3275 (N_3275,N_3016,N_3238);
or U3276 (N_3276,N_3032,N_3048);
nor U3277 (N_3277,N_3199,N_3231);
nor U3278 (N_3278,N_3074,N_3185);
nand U3279 (N_3279,N_3026,N_3148);
nor U3280 (N_3280,N_3036,N_3213);
xor U3281 (N_3281,N_3239,N_3212);
xor U3282 (N_3282,N_3116,N_3126);
or U3283 (N_3283,N_3163,N_3099);
and U3284 (N_3284,N_3223,N_3147);
nand U3285 (N_3285,N_3100,N_3043);
xnor U3286 (N_3286,N_3137,N_3092);
xor U3287 (N_3287,N_3067,N_3184);
and U3288 (N_3288,N_3200,N_3023);
xor U3289 (N_3289,N_3205,N_3004);
xor U3290 (N_3290,N_3247,N_3162);
xor U3291 (N_3291,N_3249,N_3021);
xor U3292 (N_3292,N_3229,N_3042);
or U3293 (N_3293,N_3034,N_3101);
or U3294 (N_3294,N_3089,N_3243);
nand U3295 (N_3295,N_3130,N_3172);
or U3296 (N_3296,N_3244,N_3183);
or U3297 (N_3297,N_3090,N_3202);
nor U3298 (N_3298,N_3141,N_3045);
xnor U3299 (N_3299,N_3240,N_3235);
xnor U3300 (N_3300,N_3197,N_3041);
nand U3301 (N_3301,N_3241,N_3076);
xnor U3302 (N_3302,N_3019,N_3071);
nand U3303 (N_3303,N_3233,N_3158);
nor U3304 (N_3304,N_3000,N_3156);
xor U3305 (N_3305,N_3221,N_3139);
nand U3306 (N_3306,N_3133,N_3077);
and U3307 (N_3307,N_3082,N_3246);
or U3308 (N_3308,N_3025,N_3072);
xnor U3309 (N_3309,N_3069,N_3149);
and U3310 (N_3310,N_3031,N_3013);
nor U3311 (N_3311,N_3088,N_3105);
nand U3312 (N_3312,N_3157,N_3039);
and U3313 (N_3313,N_3186,N_3140);
nand U3314 (N_3314,N_3174,N_3054);
and U3315 (N_3315,N_3227,N_3191);
xor U3316 (N_3316,N_3171,N_3119);
xnor U3317 (N_3317,N_3108,N_3085);
and U3318 (N_3318,N_3248,N_3220);
nand U3319 (N_3319,N_3160,N_3022);
nand U3320 (N_3320,N_3169,N_3131);
xnor U3321 (N_3321,N_3230,N_3180);
nand U3322 (N_3322,N_3136,N_3015);
or U3323 (N_3323,N_3135,N_3222);
nor U3324 (N_3324,N_3225,N_3138);
or U3325 (N_3325,N_3107,N_3002);
and U3326 (N_3326,N_3165,N_3217);
xnor U3327 (N_3327,N_3175,N_3049);
or U3328 (N_3328,N_3027,N_3224);
nor U3329 (N_3329,N_3125,N_3030);
or U3330 (N_3330,N_3008,N_3226);
and U3331 (N_3331,N_3106,N_3237);
xor U3332 (N_3332,N_3083,N_3080);
xnor U3333 (N_3333,N_3245,N_3150);
nor U3334 (N_3334,N_3232,N_3114);
xor U3335 (N_3335,N_3121,N_3040);
or U3336 (N_3336,N_3070,N_3206);
nor U3337 (N_3337,N_3018,N_3179);
nor U3338 (N_3338,N_3093,N_3094);
nor U3339 (N_3339,N_3110,N_3193);
nor U3340 (N_3340,N_3053,N_3122);
or U3341 (N_3341,N_3120,N_3242);
xor U3342 (N_3342,N_3189,N_3117);
and U3343 (N_3343,N_3024,N_3006);
nor U3344 (N_3344,N_3218,N_3052);
xor U3345 (N_3345,N_3007,N_3073);
nor U3346 (N_3346,N_3038,N_3055);
or U3347 (N_3347,N_3142,N_3044);
nor U3348 (N_3348,N_3209,N_3167);
nand U3349 (N_3349,N_3161,N_3112);
or U3350 (N_3350,N_3196,N_3078);
and U3351 (N_3351,N_3170,N_3215);
xnor U3352 (N_3352,N_3102,N_3216);
nor U3353 (N_3353,N_3109,N_3203);
nand U3354 (N_3354,N_3198,N_3123);
nand U3355 (N_3355,N_3173,N_3051);
nand U3356 (N_3356,N_3188,N_3028);
nor U3357 (N_3357,N_3219,N_3187);
and U3358 (N_3358,N_3065,N_3084);
and U3359 (N_3359,N_3234,N_3029);
xor U3360 (N_3360,N_3146,N_3005);
or U3361 (N_3361,N_3182,N_3086);
and U3362 (N_3362,N_3210,N_3192);
and U3363 (N_3363,N_3097,N_3176);
and U3364 (N_3364,N_3166,N_3009);
nor U3365 (N_3365,N_3208,N_3058);
nor U3366 (N_3366,N_3154,N_3062);
or U3367 (N_3367,N_3020,N_3011);
nor U3368 (N_3368,N_3014,N_3010);
and U3369 (N_3369,N_3207,N_3195);
xnor U3370 (N_3370,N_3060,N_3236);
nor U3371 (N_3371,N_3124,N_3152);
xnor U3372 (N_3372,N_3057,N_3178);
or U3373 (N_3373,N_3037,N_3181);
nor U3374 (N_3374,N_3050,N_3081);
nand U3375 (N_3375,N_3216,N_3052);
nor U3376 (N_3376,N_3094,N_3153);
and U3377 (N_3377,N_3154,N_3134);
xor U3378 (N_3378,N_3013,N_3161);
and U3379 (N_3379,N_3035,N_3106);
or U3380 (N_3380,N_3225,N_3073);
nor U3381 (N_3381,N_3206,N_3216);
xor U3382 (N_3382,N_3066,N_3233);
nand U3383 (N_3383,N_3044,N_3083);
and U3384 (N_3384,N_3060,N_3203);
nor U3385 (N_3385,N_3003,N_3110);
nand U3386 (N_3386,N_3040,N_3055);
and U3387 (N_3387,N_3117,N_3106);
nor U3388 (N_3388,N_3142,N_3200);
xnor U3389 (N_3389,N_3115,N_3223);
and U3390 (N_3390,N_3104,N_3053);
nor U3391 (N_3391,N_3037,N_3111);
nor U3392 (N_3392,N_3003,N_3099);
nor U3393 (N_3393,N_3100,N_3197);
xor U3394 (N_3394,N_3170,N_3131);
and U3395 (N_3395,N_3163,N_3028);
xor U3396 (N_3396,N_3154,N_3013);
and U3397 (N_3397,N_3112,N_3067);
nor U3398 (N_3398,N_3108,N_3166);
or U3399 (N_3399,N_3127,N_3045);
xor U3400 (N_3400,N_3001,N_3097);
and U3401 (N_3401,N_3088,N_3007);
nor U3402 (N_3402,N_3132,N_3159);
nor U3403 (N_3403,N_3123,N_3189);
nand U3404 (N_3404,N_3246,N_3165);
and U3405 (N_3405,N_3002,N_3136);
xor U3406 (N_3406,N_3091,N_3203);
xor U3407 (N_3407,N_3053,N_3072);
nor U3408 (N_3408,N_3221,N_3207);
nand U3409 (N_3409,N_3031,N_3143);
nand U3410 (N_3410,N_3236,N_3191);
and U3411 (N_3411,N_3075,N_3088);
or U3412 (N_3412,N_3119,N_3170);
xnor U3413 (N_3413,N_3122,N_3198);
or U3414 (N_3414,N_3039,N_3237);
xor U3415 (N_3415,N_3102,N_3209);
xnor U3416 (N_3416,N_3214,N_3218);
xor U3417 (N_3417,N_3218,N_3037);
nand U3418 (N_3418,N_3191,N_3215);
xnor U3419 (N_3419,N_3024,N_3048);
nand U3420 (N_3420,N_3212,N_3245);
nor U3421 (N_3421,N_3052,N_3040);
nand U3422 (N_3422,N_3042,N_3127);
or U3423 (N_3423,N_3071,N_3075);
and U3424 (N_3424,N_3037,N_3157);
nand U3425 (N_3425,N_3010,N_3169);
xor U3426 (N_3426,N_3007,N_3165);
nand U3427 (N_3427,N_3044,N_3212);
and U3428 (N_3428,N_3104,N_3235);
or U3429 (N_3429,N_3110,N_3175);
and U3430 (N_3430,N_3079,N_3107);
xnor U3431 (N_3431,N_3080,N_3248);
and U3432 (N_3432,N_3157,N_3031);
nand U3433 (N_3433,N_3136,N_3030);
xor U3434 (N_3434,N_3147,N_3148);
nand U3435 (N_3435,N_3137,N_3016);
nand U3436 (N_3436,N_3030,N_3021);
nand U3437 (N_3437,N_3228,N_3106);
nor U3438 (N_3438,N_3020,N_3217);
nand U3439 (N_3439,N_3144,N_3008);
nor U3440 (N_3440,N_3018,N_3085);
nand U3441 (N_3441,N_3212,N_3016);
nand U3442 (N_3442,N_3187,N_3078);
or U3443 (N_3443,N_3082,N_3232);
nor U3444 (N_3444,N_3084,N_3240);
nand U3445 (N_3445,N_3233,N_3157);
xor U3446 (N_3446,N_3080,N_3243);
xnor U3447 (N_3447,N_3108,N_3090);
or U3448 (N_3448,N_3240,N_3092);
nor U3449 (N_3449,N_3184,N_3177);
or U3450 (N_3450,N_3052,N_3238);
nand U3451 (N_3451,N_3223,N_3241);
nand U3452 (N_3452,N_3155,N_3164);
nand U3453 (N_3453,N_3131,N_3067);
and U3454 (N_3454,N_3099,N_3013);
nor U3455 (N_3455,N_3126,N_3025);
or U3456 (N_3456,N_3102,N_3147);
nand U3457 (N_3457,N_3233,N_3040);
or U3458 (N_3458,N_3049,N_3176);
or U3459 (N_3459,N_3018,N_3099);
and U3460 (N_3460,N_3096,N_3070);
nand U3461 (N_3461,N_3135,N_3095);
or U3462 (N_3462,N_3217,N_3103);
xor U3463 (N_3463,N_3021,N_3024);
or U3464 (N_3464,N_3187,N_3042);
xor U3465 (N_3465,N_3034,N_3021);
xnor U3466 (N_3466,N_3173,N_3067);
or U3467 (N_3467,N_3116,N_3144);
and U3468 (N_3468,N_3041,N_3209);
xor U3469 (N_3469,N_3040,N_3222);
and U3470 (N_3470,N_3138,N_3102);
xnor U3471 (N_3471,N_3115,N_3067);
nor U3472 (N_3472,N_3034,N_3040);
nand U3473 (N_3473,N_3042,N_3216);
nor U3474 (N_3474,N_3106,N_3083);
nand U3475 (N_3475,N_3181,N_3196);
xnor U3476 (N_3476,N_3037,N_3222);
nand U3477 (N_3477,N_3038,N_3172);
and U3478 (N_3478,N_3134,N_3108);
or U3479 (N_3479,N_3184,N_3047);
nor U3480 (N_3480,N_3179,N_3107);
and U3481 (N_3481,N_3157,N_3129);
nor U3482 (N_3482,N_3231,N_3116);
nand U3483 (N_3483,N_3090,N_3020);
nand U3484 (N_3484,N_3228,N_3118);
nand U3485 (N_3485,N_3231,N_3143);
and U3486 (N_3486,N_3120,N_3127);
xnor U3487 (N_3487,N_3021,N_3144);
nand U3488 (N_3488,N_3066,N_3197);
nand U3489 (N_3489,N_3060,N_3061);
or U3490 (N_3490,N_3176,N_3128);
xor U3491 (N_3491,N_3178,N_3096);
nand U3492 (N_3492,N_3034,N_3043);
and U3493 (N_3493,N_3145,N_3129);
or U3494 (N_3494,N_3165,N_3019);
and U3495 (N_3495,N_3178,N_3106);
and U3496 (N_3496,N_3042,N_3052);
and U3497 (N_3497,N_3023,N_3028);
nor U3498 (N_3498,N_3094,N_3218);
and U3499 (N_3499,N_3079,N_3140);
xor U3500 (N_3500,N_3277,N_3411);
and U3501 (N_3501,N_3357,N_3463);
nor U3502 (N_3502,N_3366,N_3423);
nand U3503 (N_3503,N_3426,N_3368);
or U3504 (N_3504,N_3388,N_3283);
nand U3505 (N_3505,N_3360,N_3498);
or U3506 (N_3506,N_3252,N_3419);
nand U3507 (N_3507,N_3344,N_3375);
or U3508 (N_3508,N_3295,N_3307);
nor U3509 (N_3509,N_3301,N_3269);
nand U3510 (N_3510,N_3403,N_3270);
nand U3511 (N_3511,N_3255,N_3484);
nand U3512 (N_3512,N_3409,N_3313);
and U3513 (N_3513,N_3481,N_3470);
nand U3514 (N_3514,N_3362,N_3381);
nor U3515 (N_3515,N_3385,N_3454);
and U3516 (N_3516,N_3446,N_3397);
nor U3517 (N_3517,N_3414,N_3336);
nor U3518 (N_3518,N_3330,N_3435);
xnor U3519 (N_3519,N_3347,N_3325);
nor U3520 (N_3520,N_3272,N_3392);
and U3521 (N_3521,N_3405,N_3343);
xnor U3522 (N_3522,N_3308,N_3292);
or U3523 (N_3523,N_3445,N_3378);
or U3524 (N_3524,N_3395,N_3437);
nor U3525 (N_3525,N_3492,N_3441);
or U3526 (N_3526,N_3425,N_3333);
nand U3527 (N_3527,N_3465,N_3479);
nand U3528 (N_3528,N_3415,N_3466);
nand U3529 (N_3529,N_3304,N_3447);
nand U3530 (N_3530,N_3494,N_3444);
and U3531 (N_3531,N_3259,N_3471);
nor U3532 (N_3532,N_3299,N_3449);
or U3533 (N_3533,N_3334,N_3458);
nand U3534 (N_3534,N_3251,N_3493);
nand U3535 (N_3535,N_3383,N_3400);
and U3536 (N_3536,N_3398,N_3349);
nand U3537 (N_3537,N_3358,N_3438);
xnor U3538 (N_3538,N_3422,N_3456);
and U3539 (N_3539,N_3496,N_3420);
nor U3540 (N_3540,N_3490,N_3332);
and U3541 (N_3541,N_3469,N_3315);
or U3542 (N_3542,N_3382,N_3285);
or U3543 (N_3543,N_3337,N_3291);
nand U3544 (N_3544,N_3391,N_3340);
xor U3545 (N_3545,N_3394,N_3455);
xnor U3546 (N_3546,N_3254,N_3281);
or U3547 (N_3547,N_3436,N_3316);
or U3548 (N_3548,N_3472,N_3369);
nand U3549 (N_3549,N_3380,N_3341);
nand U3550 (N_3550,N_3312,N_3275);
xnor U3551 (N_3551,N_3488,N_3480);
nor U3552 (N_3552,N_3287,N_3311);
or U3553 (N_3553,N_3250,N_3289);
nor U3554 (N_3554,N_3384,N_3373);
nor U3555 (N_3555,N_3439,N_3489);
xor U3556 (N_3556,N_3278,N_3314);
and U3557 (N_3557,N_3370,N_3342);
nand U3558 (N_3558,N_3457,N_3361);
nor U3559 (N_3559,N_3324,N_3410);
or U3560 (N_3560,N_3267,N_3475);
or U3561 (N_3561,N_3320,N_3377);
and U3562 (N_3562,N_3280,N_3363);
nor U3563 (N_3563,N_3356,N_3430);
nor U3564 (N_3564,N_3263,N_3318);
xor U3565 (N_3565,N_3351,N_3328);
nand U3566 (N_3566,N_3284,N_3339);
nand U3567 (N_3567,N_3294,N_3485);
and U3568 (N_3568,N_3310,N_3468);
or U3569 (N_3569,N_3486,N_3413);
nor U3570 (N_3570,N_3317,N_3302);
or U3571 (N_3571,N_3348,N_3274);
nor U3572 (N_3572,N_3322,N_3404);
or U3573 (N_3573,N_3387,N_3402);
xnor U3574 (N_3574,N_3390,N_3353);
and U3575 (N_3575,N_3467,N_3389);
nor U3576 (N_3576,N_3393,N_3461);
nand U3577 (N_3577,N_3376,N_3323);
xor U3578 (N_3578,N_3386,N_3260);
nor U3579 (N_3579,N_3429,N_3427);
nand U3580 (N_3580,N_3428,N_3477);
or U3581 (N_3581,N_3290,N_3408);
xnor U3582 (N_3582,N_3452,N_3367);
nand U3583 (N_3583,N_3364,N_3483);
nor U3584 (N_3584,N_3288,N_3433);
or U3585 (N_3585,N_3379,N_3431);
or U3586 (N_3586,N_3350,N_3418);
nand U3587 (N_3587,N_3276,N_3497);
and U3588 (N_3588,N_3271,N_3495);
xor U3589 (N_3589,N_3491,N_3293);
xnor U3590 (N_3590,N_3261,N_3268);
nor U3591 (N_3591,N_3406,N_3326);
xnor U3592 (N_3592,N_3371,N_3416);
xnor U3593 (N_3593,N_3499,N_3258);
nor U3594 (N_3594,N_3374,N_3407);
and U3595 (N_3595,N_3412,N_3396);
and U3596 (N_3596,N_3443,N_3346);
nor U3597 (N_3597,N_3296,N_3448);
or U3598 (N_3598,N_3464,N_3352);
nand U3599 (N_3599,N_3321,N_3345);
nor U3600 (N_3600,N_3303,N_3442);
or U3601 (N_3601,N_3262,N_3421);
nand U3602 (N_3602,N_3297,N_3473);
nor U3603 (N_3603,N_3365,N_3253);
and U3604 (N_3604,N_3300,N_3319);
or U3605 (N_3605,N_3453,N_3279);
nand U3606 (N_3606,N_3264,N_3335);
nor U3607 (N_3607,N_3256,N_3399);
nand U3608 (N_3608,N_3432,N_3487);
and U3609 (N_3609,N_3338,N_3298);
nand U3610 (N_3610,N_3355,N_3327);
nor U3611 (N_3611,N_3440,N_3309);
or U3612 (N_3612,N_3482,N_3286);
xnor U3613 (N_3613,N_3354,N_3359);
and U3614 (N_3614,N_3273,N_3305);
nor U3615 (N_3615,N_3401,N_3459);
or U3616 (N_3616,N_3451,N_3265);
nand U3617 (N_3617,N_3434,N_3424);
nor U3618 (N_3618,N_3450,N_3462);
or U3619 (N_3619,N_3306,N_3257);
xnor U3620 (N_3620,N_3266,N_3476);
and U3621 (N_3621,N_3474,N_3282);
or U3622 (N_3622,N_3478,N_3372);
or U3623 (N_3623,N_3331,N_3417);
and U3624 (N_3624,N_3329,N_3460);
xor U3625 (N_3625,N_3460,N_3496);
nand U3626 (N_3626,N_3375,N_3464);
nor U3627 (N_3627,N_3372,N_3425);
nand U3628 (N_3628,N_3314,N_3364);
and U3629 (N_3629,N_3251,N_3355);
and U3630 (N_3630,N_3449,N_3432);
xor U3631 (N_3631,N_3260,N_3404);
xor U3632 (N_3632,N_3316,N_3394);
nand U3633 (N_3633,N_3431,N_3364);
nand U3634 (N_3634,N_3475,N_3407);
nor U3635 (N_3635,N_3326,N_3318);
nor U3636 (N_3636,N_3333,N_3478);
nor U3637 (N_3637,N_3267,N_3323);
or U3638 (N_3638,N_3292,N_3439);
nor U3639 (N_3639,N_3437,N_3385);
or U3640 (N_3640,N_3287,N_3400);
xor U3641 (N_3641,N_3417,N_3307);
nand U3642 (N_3642,N_3416,N_3400);
and U3643 (N_3643,N_3401,N_3295);
nand U3644 (N_3644,N_3253,N_3447);
nor U3645 (N_3645,N_3284,N_3264);
xnor U3646 (N_3646,N_3386,N_3345);
nor U3647 (N_3647,N_3354,N_3380);
nand U3648 (N_3648,N_3448,N_3463);
and U3649 (N_3649,N_3389,N_3365);
nand U3650 (N_3650,N_3478,N_3319);
or U3651 (N_3651,N_3380,N_3404);
and U3652 (N_3652,N_3450,N_3436);
nor U3653 (N_3653,N_3318,N_3441);
and U3654 (N_3654,N_3254,N_3307);
nand U3655 (N_3655,N_3283,N_3374);
nand U3656 (N_3656,N_3371,N_3431);
and U3657 (N_3657,N_3347,N_3486);
nand U3658 (N_3658,N_3365,N_3401);
nand U3659 (N_3659,N_3468,N_3297);
nor U3660 (N_3660,N_3326,N_3290);
nand U3661 (N_3661,N_3267,N_3306);
and U3662 (N_3662,N_3391,N_3385);
and U3663 (N_3663,N_3493,N_3451);
or U3664 (N_3664,N_3265,N_3388);
xnor U3665 (N_3665,N_3478,N_3410);
nor U3666 (N_3666,N_3382,N_3371);
nand U3667 (N_3667,N_3461,N_3418);
and U3668 (N_3668,N_3451,N_3373);
or U3669 (N_3669,N_3257,N_3442);
or U3670 (N_3670,N_3413,N_3334);
xor U3671 (N_3671,N_3294,N_3258);
or U3672 (N_3672,N_3271,N_3460);
nor U3673 (N_3673,N_3322,N_3342);
and U3674 (N_3674,N_3354,N_3490);
nor U3675 (N_3675,N_3442,N_3490);
and U3676 (N_3676,N_3333,N_3251);
or U3677 (N_3677,N_3462,N_3369);
xor U3678 (N_3678,N_3272,N_3312);
and U3679 (N_3679,N_3253,N_3267);
and U3680 (N_3680,N_3381,N_3417);
xnor U3681 (N_3681,N_3405,N_3445);
and U3682 (N_3682,N_3264,N_3281);
nor U3683 (N_3683,N_3288,N_3381);
and U3684 (N_3684,N_3355,N_3401);
and U3685 (N_3685,N_3352,N_3273);
nor U3686 (N_3686,N_3307,N_3357);
nand U3687 (N_3687,N_3296,N_3452);
nor U3688 (N_3688,N_3447,N_3302);
or U3689 (N_3689,N_3477,N_3412);
xor U3690 (N_3690,N_3252,N_3476);
and U3691 (N_3691,N_3309,N_3422);
nor U3692 (N_3692,N_3493,N_3342);
nor U3693 (N_3693,N_3306,N_3488);
or U3694 (N_3694,N_3360,N_3301);
nand U3695 (N_3695,N_3403,N_3463);
or U3696 (N_3696,N_3409,N_3373);
nand U3697 (N_3697,N_3333,N_3483);
or U3698 (N_3698,N_3386,N_3499);
nor U3699 (N_3699,N_3459,N_3323);
xnor U3700 (N_3700,N_3396,N_3381);
nor U3701 (N_3701,N_3407,N_3328);
xnor U3702 (N_3702,N_3458,N_3476);
nand U3703 (N_3703,N_3403,N_3296);
xnor U3704 (N_3704,N_3408,N_3353);
xor U3705 (N_3705,N_3484,N_3300);
nor U3706 (N_3706,N_3430,N_3250);
or U3707 (N_3707,N_3343,N_3366);
xor U3708 (N_3708,N_3259,N_3466);
or U3709 (N_3709,N_3312,N_3256);
nand U3710 (N_3710,N_3455,N_3339);
xor U3711 (N_3711,N_3376,N_3291);
nand U3712 (N_3712,N_3390,N_3269);
xnor U3713 (N_3713,N_3351,N_3292);
and U3714 (N_3714,N_3361,N_3278);
nand U3715 (N_3715,N_3429,N_3374);
xnor U3716 (N_3716,N_3332,N_3457);
or U3717 (N_3717,N_3333,N_3472);
and U3718 (N_3718,N_3272,N_3484);
and U3719 (N_3719,N_3477,N_3402);
nor U3720 (N_3720,N_3467,N_3368);
or U3721 (N_3721,N_3387,N_3252);
and U3722 (N_3722,N_3428,N_3322);
and U3723 (N_3723,N_3298,N_3365);
xor U3724 (N_3724,N_3269,N_3455);
nand U3725 (N_3725,N_3444,N_3368);
nor U3726 (N_3726,N_3452,N_3314);
nand U3727 (N_3727,N_3275,N_3437);
nand U3728 (N_3728,N_3375,N_3333);
xnor U3729 (N_3729,N_3318,N_3270);
or U3730 (N_3730,N_3372,N_3421);
and U3731 (N_3731,N_3491,N_3313);
xnor U3732 (N_3732,N_3421,N_3431);
nor U3733 (N_3733,N_3345,N_3443);
nand U3734 (N_3734,N_3283,N_3274);
xnor U3735 (N_3735,N_3391,N_3455);
xor U3736 (N_3736,N_3325,N_3262);
xor U3737 (N_3737,N_3325,N_3403);
xor U3738 (N_3738,N_3445,N_3438);
xor U3739 (N_3739,N_3495,N_3342);
xnor U3740 (N_3740,N_3295,N_3354);
nand U3741 (N_3741,N_3426,N_3390);
or U3742 (N_3742,N_3483,N_3339);
nor U3743 (N_3743,N_3276,N_3472);
and U3744 (N_3744,N_3412,N_3351);
nand U3745 (N_3745,N_3273,N_3458);
nor U3746 (N_3746,N_3460,N_3332);
xor U3747 (N_3747,N_3420,N_3320);
nand U3748 (N_3748,N_3353,N_3443);
and U3749 (N_3749,N_3428,N_3276);
xnor U3750 (N_3750,N_3730,N_3713);
or U3751 (N_3751,N_3646,N_3603);
or U3752 (N_3752,N_3611,N_3548);
or U3753 (N_3753,N_3536,N_3618);
and U3754 (N_3754,N_3591,N_3605);
nor U3755 (N_3755,N_3737,N_3742);
nor U3756 (N_3756,N_3564,N_3724);
or U3757 (N_3757,N_3575,N_3508);
or U3758 (N_3758,N_3720,N_3610);
xor U3759 (N_3759,N_3629,N_3597);
nor U3760 (N_3760,N_3745,N_3547);
xor U3761 (N_3761,N_3542,N_3643);
nand U3762 (N_3762,N_3543,N_3545);
or U3763 (N_3763,N_3577,N_3512);
xor U3764 (N_3764,N_3663,N_3540);
xnor U3765 (N_3765,N_3544,N_3516);
or U3766 (N_3766,N_3704,N_3722);
xor U3767 (N_3767,N_3641,N_3747);
and U3768 (N_3768,N_3652,N_3728);
or U3769 (N_3769,N_3683,N_3626);
and U3770 (N_3770,N_3589,N_3672);
xor U3771 (N_3771,N_3579,N_3656);
and U3772 (N_3772,N_3693,N_3550);
nor U3773 (N_3773,N_3584,N_3743);
nand U3774 (N_3774,N_3619,N_3677);
xnor U3775 (N_3775,N_3698,N_3710);
and U3776 (N_3776,N_3602,N_3740);
xor U3777 (N_3777,N_3563,N_3533);
nand U3778 (N_3778,N_3716,N_3669);
nand U3779 (N_3779,N_3608,N_3538);
or U3780 (N_3780,N_3732,N_3719);
or U3781 (N_3781,N_3668,N_3725);
nor U3782 (N_3782,N_3696,N_3522);
or U3783 (N_3783,N_3583,N_3681);
nand U3784 (N_3784,N_3746,N_3552);
xor U3785 (N_3785,N_3520,N_3505);
or U3786 (N_3786,N_3738,N_3596);
nor U3787 (N_3787,N_3501,N_3721);
xnor U3788 (N_3788,N_3606,N_3637);
or U3789 (N_3789,N_3506,N_3604);
nor U3790 (N_3790,N_3671,N_3650);
and U3791 (N_3791,N_3694,N_3749);
nor U3792 (N_3792,N_3703,N_3588);
nor U3793 (N_3793,N_3702,N_3562);
nand U3794 (N_3794,N_3572,N_3546);
and U3795 (N_3795,N_3503,N_3651);
nor U3796 (N_3796,N_3711,N_3507);
nand U3797 (N_3797,N_3735,N_3633);
nand U3798 (N_3798,N_3707,N_3624);
nand U3799 (N_3799,N_3685,N_3502);
xnor U3800 (N_3800,N_3565,N_3715);
and U3801 (N_3801,N_3593,N_3679);
xor U3802 (N_3802,N_3622,N_3535);
xnor U3803 (N_3803,N_3676,N_3662);
nand U3804 (N_3804,N_3609,N_3627);
nand U3805 (N_3805,N_3729,N_3714);
or U3806 (N_3806,N_3569,N_3748);
and U3807 (N_3807,N_3697,N_3660);
nand U3808 (N_3808,N_3553,N_3741);
xor U3809 (N_3809,N_3658,N_3708);
nor U3810 (N_3810,N_3576,N_3706);
nand U3811 (N_3811,N_3549,N_3689);
nor U3812 (N_3812,N_3541,N_3670);
and U3813 (N_3813,N_3511,N_3558);
xor U3814 (N_3814,N_3717,N_3574);
nor U3815 (N_3815,N_3688,N_3590);
xor U3816 (N_3816,N_3529,N_3709);
xor U3817 (N_3817,N_3649,N_3653);
nor U3818 (N_3818,N_3682,N_3645);
nor U3819 (N_3819,N_3638,N_3504);
xnor U3820 (N_3820,N_3517,N_3551);
xor U3821 (N_3821,N_3557,N_3699);
nor U3822 (N_3822,N_3586,N_3581);
or U3823 (N_3823,N_3570,N_3532);
xor U3824 (N_3824,N_3648,N_3515);
or U3825 (N_3825,N_3620,N_3647);
and U3826 (N_3826,N_3568,N_3518);
and U3827 (N_3827,N_3686,N_3733);
or U3828 (N_3828,N_3580,N_3661);
xor U3829 (N_3829,N_3734,N_3607);
nand U3830 (N_3830,N_3687,N_3665);
xnor U3831 (N_3831,N_3556,N_3560);
xor U3832 (N_3832,N_3617,N_3521);
or U3833 (N_3833,N_3573,N_3524);
nor U3834 (N_3834,N_3531,N_3684);
nor U3835 (N_3835,N_3640,N_3642);
and U3836 (N_3836,N_3635,N_3525);
and U3837 (N_3837,N_3659,N_3628);
nor U3838 (N_3838,N_3554,N_3527);
nor U3839 (N_3839,N_3598,N_3639);
or U3840 (N_3840,N_3625,N_3519);
nor U3841 (N_3841,N_3594,N_3530);
or U3842 (N_3842,N_3526,N_3666);
nand U3843 (N_3843,N_3634,N_3601);
nand U3844 (N_3844,N_3726,N_3630);
nor U3845 (N_3845,N_3644,N_3561);
nor U3846 (N_3846,N_3514,N_3655);
nor U3847 (N_3847,N_3528,N_3567);
and U3848 (N_3848,N_3509,N_3559);
nor U3849 (N_3849,N_3615,N_3595);
xor U3850 (N_3850,N_3571,N_3621);
nor U3851 (N_3851,N_3675,N_3667);
nor U3852 (N_3852,N_3700,N_3578);
xor U3853 (N_3853,N_3500,N_3736);
nand U3854 (N_3854,N_3701,N_3555);
and U3855 (N_3855,N_3537,N_3636);
xor U3856 (N_3856,N_3566,N_3585);
xor U3857 (N_3857,N_3678,N_3674);
nor U3858 (N_3858,N_3673,N_3523);
nor U3859 (N_3859,N_3616,N_3632);
nand U3860 (N_3860,N_3657,N_3631);
xor U3861 (N_3861,N_3513,N_3613);
xor U3862 (N_3862,N_3690,N_3718);
nor U3863 (N_3863,N_3510,N_3712);
nor U3864 (N_3864,N_3614,N_3705);
nor U3865 (N_3865,N_3592,N_3599);
or U3866 (N_3866,N_3539,N_3695);
xnor U3867 (N_3867,N_3534,N_3612);
nand U3868 (N_3868,N_3692,N_3727);
nor U3869 (N_3869,N_3623,N_3691);
or U3870 (N_3870,N_3654,N_3739);
xor U3871 (N_3871,N_3680,N_3731);
and U3872 (N_3872,N_3600,N_3744);
or U3873 (N_3873,N_3582,N_3587);
xnor U3874 (N_3874,N_3723,N_3664);
or U3875 (N_3875,N_3603,N_3678);
nand U3876 (N_3876,N_3619,N_3640);
or U3877 (N_3877,N_3576,N_3560);
and U3878 (N_3878,N_3551,N_3514);
nor U3879 (N_3879,N_3552,N_3567);
xor U3880 (N_3880,N_3686,N_3583);
nor U3881 (N_3881,N_3505,N_3642);
nor U3882 (N_3882,N_3745,N_3586);
and U3883 (N_3883,N_3611,N_3517);
xnor U3884 (N_3884,N_3697,N_3527);
xnor U3885 (N_3885,N_3684,N_3725);
nand U3886 (N_3886,N_3662,N_3531);
xor U3887 (N_3887,N_3721,N_3711);
or U3888 (N_3888,N_3692,N_3575);
nor U3889 (N_3889,N_3590,N_3702);
nor U3890 (N_3890,N_3727,N_3529);
nand U3891 (N_3891,N_3611,N_3684);
and U3892 (N_3892,N_3646,N_3580);
nand U3893 (N_3893,N_3507,N_3662);
nand U3894 (N_3894,N_3708,N_3633);
xnor U3895 (N_3895,N_3743,N_3640);
or U3896 (N_3896,N_3538,N_3518);
nand U3897 (N_3897,N_3520,N_3526);
or U3898 (N_3898,N_3725,N_3599);
xnor U3899 (N_3899,N_3571,N_3580);
or U3900 (N_3900,N_3656,N_3689);
nand U3901 (N_3901,N_3623,N_3610);
and U3902 (N_3902,N_3590,N_3693);
or U3903 (N_3903,N_3545,N_3522);
and U3904 (N_3904,N_3554,N_3702);
nor U3905 (N_3905,N_3728,N_3603);
or U3906 (N_3906,N_3737,N_3533);
xnor U3907 (N_3907,N_3619,N_3626);
and U3908 (N_3908,N_3704,N_3515);
and U3909 (N_3909,N_3585,N_3647);
xor U3910 (N_3910,N_3570,N_3576);
xor U3911 (N_3911,N_3501,N_3556);
or U3912 (N_3912,N_3537,N_3732);
nand U3913 (N_3913,N_3643,N_3580);
nand U3914 (N_3914,N_3525,N_3623);
nor U3915 (N_3915,N_3639,N_3733);
and U3916 (N_3916,N_3746,N_3502);
xor U3917 (N_3917,N_3516,N_3709);
and U3918 (N_3918,N_3595,N_3640);
and U3919 (N_3919,N_3723,N_3656);
nand U3920 (N_3920,N_3592,N_3627);
or U3921 (N_3921,N_3648,N_3538);
or U3922 (N_3922,N_3534,N_3510);
and U3923 (N_3923,N_3620,N_3720);
xnor U3924 (N_3924,N_3683,N_3615);
xnor U3925 (N_3925,N_3632,N_3553);
xnor U3926 (N_3926,N_3580,N_3739);
xnor U3927 (N_3927,N_3612,N_3678);
xnor U3928 (N_3928,N_3658,N_3559);
and U3929 (N_3929,N_3627,N_3666);
nand U3930 (N_3930,N_3586,N_3580);
nor U3931 (N_3931,N_3519,N_3665);
or U3932 (N_3932,N_3659,N_3634);
nor U3933 (N_3933,N_3500,N_3711);
nand U3934 (N_3934,N_3631,N_3692);
xnor U3935 (N_3935,N_3542,N_3676);
nor U3936 (N_3936,N_3628,N_3531);
nand U3937 (N_3937,N_3574,N_3739);
and U3938 (N_3938,N_3581,N_3738);
xor U3939 (N_3939,N_3690,N_3726);
xor U3940 (N_3940,N_3536,N_3608);
xnor U3941 (N_3941,N_3589,N_3613);
and U3942 (N_3942,N_3648,N_3705);
and U3943 (N_3943,N_3525,N_3550);
and U3944 (N_3944,N_3694,N_3589);
nor U3945 (N_3945,N_3524,N_3621);
or U3946 (N_3946,N_3714,N_3593);
nand U3947 (N_3947,N_3640,N_3707);
nor U3948 (N_3948,N_3651,N_3543);
and U3949 (N_3949,N_3686,N_3658);
and U3950 (N_3950,N_3710,N_3581);
and U3951 (N_3951,N_3666,N_3726);
nor U3952 (N_3952,N_3519,N_3598);
xnor U3953 (N_3953,N_3725,N_3647);
nor U3954 (N_3954,N_3655,N_3695);
nor U3955 (N_3955,N_3505,N_3740);
and U3956 (N_3956,N_3671,N_3591);
or U3957 (N_3957,N_3587,N_3708);
nor U3958 (N_3958,N_3689,N_3669);
or U3959 (N_3959,N_3691,N_3511);
and U3960 (N_3960,N_3728,N_3560);
nor U3961 (N_3961,N_3631,N_3530);
and U3962 (N_3962,N_3649,N_3569);
nor U3963 (N_3963,N_3635,N_3734);
xor U3964 (N_3964,N_3704,N_3577);
nand U3965 (N_3965,N_3631,N_3744);
and U3966 (N_3966,N_3653,N_3638);
nor U3967 (N_3967,N_3635,N_3580);
xnor U3968 (N_3968,N_3648,N_3630);
and U3969 (N_3969,N_3544,N_3597);
nand U3970 (N_3970,N_3739,N_3602);
or U3971 (N_3971,N_3672,N_3506);
xor U3972 (N_3972,N_3569,N_3664);
xnor U3973 (N_3973,N_3726,N_3735);
nor U3974 (N_3974,N_3716,N_3573);
or U3975 (N_3975,N_3603,N_3675);
nand U3976 (N_3976,N_3602,N_3748);
nor U3977 (N_3977,N_3611,N_3713);
nor U3978 (N_3978,N_3693,N_3572);
and U3979 (N_3979,N_3671,N_3598);
nor U3980 (N_3980,N_3500,N_3734);
and U3981 (N_3981,N_3612,N_3505);
nor U3982 (N_3982,N_3605,N_3637);
nand U3983 (N_3983,N_3518,N_3526);
or U3984 (N_3984,N_3526,N_3740);
and U3985 (N_3985,N_3735,N_3695);
nor U3986 (N_3986,N_3622,N_3744);
or U3987 (N_3987,N_3661,N_3557);
nand U3988 (N_3988,N_3652,N_3614);
or U3989 (N_3989,N_3722,N_3685);
and U3990 (N_3990,N_3556,N_3580);
nand U3991 (N_3991,N_3675,N_3610);
nor U3992 (N_3992,N_3687,N_3724);
nor U3993 (N_3993,N_3743,N_3745);
or U3994 (N_3994,N_3693,N_3501);
xnor U3995 (N_3995,N_3545,N_3708);
xnor U3996 (N_3996,N_3686,N_3645);
or U3997 (N_3997,N_3722,N_3537);
or U3998 (N_3998,N_3675,N_3733);
nor U3999 (N_3999,N_3740,N_3675);
nor U4000 (N_4000,N_3807,N_3793);
xnor U4001 (N_4001,N_3948,N_3763);
xor U4002 (N_4002,N_3936,N_3777);
nor U4003 (N_4003,N_3909,N_3843);
nor U4004 (N_4004,N_3769,N_3826);
and U4005 (N_4005,N_3782,N_3856);
nor U4006 (N_4006,N_3838,N_3832);
and U4007 (N_4007,N_3981,N_3894);
and U4008 (N_4008,N_3901,N_3995);
or U4009 (N_4009,N_3758,N_3905);
xor U4010 (N_4010,N_3929,N_3915);
xnor U4011 (N_4011,N_3932,N_3899);
or U4012 (N_4012,N_3892,N_3825);
nor U4013 (N_4013,N_3863,N_3865);
nand U4014 (N_4014,N_3784,N_3834);
nand U4015 (N_4015,N_3772,N_3795);
or U4016 (N_4016,N_3757,N_3873);
nand U4017 (N_4017,N_3878,N_3986);
xnor U4018 (N_4018,N_3766,N_3933);
nor U4019 (N_4019,N_3993,N_3831);
nor U4020 (N_4020,N_3774,N_3954);
xor U4021 (N_4021,N_3964,N_3781);
or U4022 (N_4022,N_3945,N_3851);
xor U4023 (N_4023,N_3762,N_3792);
nor U4024 (N_4024,N_3970,N_3980);
xnor U4025 (N_4025,N_3845,N_3950);
and U4026 (N_4026,N_3858,N_3778);
and U4027 (N_4027,N_3824,N_3926);
nand U4028 (N_4028,N_3849,N_3947);
xnor U4029 (N_4029,N_3846,N_3765);
and U4030 (N_4030,N_3850,N_3864);
and U4031 (N_4031,N_3903,N_3839);
and U4032 (N_4032,N_3988,N_3842);
nor U4033 (N_4033,N_3889,N_3885);
xnor U4034 (N_4034,N_3764,N_3989);
nor U4035 (N_4035,N_3770,N_3985);
nor U4036 (N_4036,N_3921,N_3877);
xor U4037 (N_4037,N_3771,N_3860);
or U4038 (N_4038,N_3794,N_3815);
and U4039 (N_4039,N_3943,N_3814);
nand U4040 (N_4040,N_3867,N_3797);
nor U4041 (N_4041,N_3890,N_3906);
or U4042 (N_4042,N_3934,N_3975);
and U4043 (N_4043,N_3907,N_3811);
xnor U4044 (N_4044,N_3830,N_3800);
xor U4045 (N_4045,N_3809,N_3802);
xor U4046 (N_4046,N_3820,N_3767);
nand U4047 (N_4047,N_3957,N_3895);
nand U4048 (N_4048,N_3941,N_3923);
or U4049 (N_4049,N_3768,N_3984);
or U4050 (N_4050,N_3871,N_3875);
nor U4051 (N_4051,N_3810,N_3952);
and U4052 (N_4052,N_3870,N_3783);
or U4053 (N_4053,N_3960,N_3847);
xor U4054 (N_4054,N_3869,N_3786);
xnor U4055 (N_4055,N_3791,N_3951);
and U4056 (N_4056,N_3968,N_3817);
and U4057 (N_4057,N_3829,N_3991);
nand U4058 (N_4058,N_3785,N_3854);
and U4059 (N_4059,N_3888,N_3937);
nor U4060 (N_4060,N_3812,N_3787);
xor U4061 (N_4061,N_3902,N_3799);
or U4062 (N_4062,N_3962,N_3898);
nor U4063 (N_4063,N_3884,N_3931);
and U4064 (N_4064,N_3977,N_3971);
xor U4065 (N_4065,N_3835,N_3868);
and U4066 (N_4066,N_3827,N_3761);
and U4067 (N_4067,N_3990,N_3788);
nor U4068 (N_4068,N_3917,N_3927);
nor U4069 (N_4069,N_3844,N_3818);
and U4070 (N_4070,N_3880,N_3779);
nand U4071 (N_4071,N_3806,N_3919);
xnor U4072 (N_4072,N_3756,N_3886);
xor U4073 (N_4073,N_3946,N_3904);
nand U4074 (N_4074,N_3857,N_3874);
nor U4075 (N_4075,N_3816,N_3808);
nand U4076 (N_4076,N_3956,N_3881);
and U4077 (N_4077,N_3925,N_3882);
nand U4078 (N_4078,N_3872,N_3805);
nand U4079 (N_4079,N_3979,N_3862);
xnor U4080 (N_4080,N_3823,N_3935);
nor U4081 (N_4081,N_3833,N_3966);
xor U4082 (N_4082,N_3879,N_3893);
nand U4083 (N_4083,N_3920,N_3914);
nand U4084 (N_4084,N_3776,N_3942);
or U4085 (N_4085,N_3949,N_3978);
and U4086 (N_4086,N_3753,N_3965);
or U4087 (N_4087,N_3855,N_3752);
xnor U4088 (N_4088,N_3959,N_3775);
nor U4089 (N_4089,N_3803,N_3883);
nand U4090 (N_4090,N_3940,N_3801);
xor U4091 (N_4091,N_3760,N_3755);
nand U4092 (N_4092,N_3840,N_3866);
xnor U4093 (N_4093,N_3998,N_3887);
or U4094 (N_4094,N_3804,N_3750);
and U4095 (N_4095,N_3780,N_3961);
or U4096 (N_4096,N_3754,N_3773);
nor U4097 (N_4097,N_3955,N_3911);
nand U4098 (N_4098,N_3972,N_3918);
nor U4099 (N_4099,N_3997,N_3759);
and U4100 (N_4100,N_3999,N_3994);
xor U4101 (N_4101,N_3908,N_3983);
xnor U4102 (N_4102,N_3922,N_3944);
or U4103 (N_4103,N_3992,N_3976);
nand U4104 (N_4104,N_3789,N_3828);
nor U4105 (N_4105,N_3900,N_3796);
nand U4106 (N_4106,N_3928,N_3987);
nand U4107 (N_4107,N_3859,N_3897);
nand U4108 (N_4108,N_3924,N_3953);
xor U4109 (N_4109,N_3848,N_3819);
nand U4110 (N_4110,N_3836,N_3813);
or U4111 (N_4111,N_3939,N_3963);
and U4112 (N_4112,N_3876,N_3852);
nand U4113 (N_4113,N_3938,N_3853);
nor U4114 (N_4114,N_3996,N_3896);
nor U4115 (N_4115,N_3751,N_3974);
or U4116 (N_4116,N_3958,N_3821);
or U4117 (N_4117,N_3861,N_3841);
xor U4118 (N_4118,N_3822,N_3912);
or U4119 (N_4119,N_3910,N_3969);
and U4120 (N_4120,N_3798,N_3913);
xnor U4121 (N_4121,N_3916,N_3973);
xor U4122 (N_4122,N_3790,N_3967);
xor U4123 (N_4123,N_3837,N_3982);
and U4124 (N_4124,N_3891,N_3930);
and U4125 (N_4125,N_3938,N_3856);
and U4126 (N_4126,N_3966,N_3853);
xnor U4127 (N_4127,N_3769,N_3856);
and U4128 (N_4128,N_3847,N_3957);
xor U4129 (N_4129,N_3829,N_3959);
nor U4130 (N_4130,N_3862,N_3969);
or U4131 (N_4131,N_3985,N_3923);
xnor U4132 (N_4132,N_3822,N_3927);
and U4133 (N_4133,N_3938,N_3787);
and U4134 (N_4134,N_3915,N_3910);
or U4135 (N_4135,N_3955,N_3931);
and U4136 (N_4136,N_3856,N_3829);
or U4137 (N_4137,N_3942,N_3867);
or U4138 (N_4138,N_3915,N_3992);
or U4139 (N_4139,N_3921,N_3993);
xor U4140 (N_4140,N_3861,N_3947);
nand U4141 (N_4141,N_3826,N_3860);
and U4142 (N_4142,N_3784,N_3766);
and U4143 (N_4143,N_3780,N_3772);
nor U4144 (N_4144,N_3884,N_3751);
xor U4145 (N_4145,N_3961,N_3936);
or U4146 (N_4146,N_3986,N_3800);
nand U4147 (N_4147,N_3847,N_3926);
nand U4148 (N_4148,N_3849,N_3896);
nand U4149 (N_4149,N_3871,N_3829);
and U4150 (N_4150,N_3788,N_3987);
nor U4151 (N_4151,N_3955,N_3882);
or U4152 (N_4152,N_3801,N_3923);
nor U4153 (N_4153,N_3792,N_3795);
or U4154 (N_4154,N_3848,N_3764);
nor U4155 (N_4155,N_3936,N_3771);
and U4156 (N_4156,N_3932,N_3765);
and U4157 (N_4157,N_3868,N_3768);
nor U4158 (N_4158,N_3993,N_3861);
nor U4159 (N_4159,N_3943,N_3954);
or U4160 (N_4160,N_3791,N_3840);
and U4161 (N_4161,N_3830,N_3948);
nand U4162 (N_4162,N_3829,N_3937);
xnor U4163 (N_4163,N_3963,N_3921);
xor U4164 (N_4164,N_3834,N_3852);
and U4165 (N_4165,N_3774,N_3817);
xnor U4166 (N_4166,N_3964,N_3959);
nor U4167 (N_4167,N_3775,N_3919);
xor U4168 (N_4168,N_3860,N_3875);
and U4169 (N_4169,N_3785,N_3815);
and U4170 (N_4170,N_3764,N_3776);
or U4171 (N_4171,N_3992,N_3906);
and U4172 (N_4172,N_3764,N_3981);
nand U4173 (N_4173,N_3845,N_3859);
or U4174 (N_4174,N_3760,N_3792);
nand U4175 (N_4175,N_3761,N_3869);
nand U4176 (N_4176,N_3874,N_3975);
nor U4177 (N_4177,N_3914,N_3763);
nand U4178 (N_4178,N_3992,N_3804);
or U4179 (N_4179,N_3943,N_3752);
xor U4180 (N_4180,N_3970,N_3990);
or U4181 (N_4181,N_3826,N_3990);
xnor U4182 (N_4182,N_3809,N_3855);
or U4183 (N_4183,N_3883,N_3828);
nand U4184 (N_4184,N_3883,N_3899);
nand U4185 (N_4185,N_3891,N_3919);
nor U4186 (N_4186,N_3771,N_3951);
and U4187 (N_4187,N_3990,N_3881);
and U4188 (N_4188,N_3904,N_3948);
or U4189 (N_4189,N_3991,N_3898);
and U4190 (N_4190,N_3771,N_3814);
or U4191 (N_4191,N_3890,N_3810);
nand U4192 (N_4192,N_3820,N_3788);
nand U4193 (N_4193,N_3827,N_3852);
nor U4194 (N_4194,N_3907,N_3756);
nor U4195 (N_4195,N_3995,N_3890);
nand U4196 (N_4196,N_3769,N_3781);
xor U4197 (N_4197,N_3925,N_3878);
nor U4198 (N_4198,N_3962,N_3836);
nand U4199 (N_4199,N_3762,N_3968);
nand U4200 (N_4200,N_3927,N_3877);
xnor U4201 (N_4201,N_3758,N_3827);
and U4202 (N_4202,N_3853,N_3780);
nand U4203 (N_4203,N_3937,N_3972);
nor U4204 (N_4204,N_3795,N_3851);
nor U4205 (N_4205,N_3901,N_3885);
nand U4206 (N_4206,N_3869,N_3997);
or U4207 (N_4207,N_3902,N_3964);
xor U4208 (N_4208,N_3819,N_3773);
or U4209 (N_4209,N_3892,N_3815);
and U4210 (N_4210,N_3781,N_3900);
nand U4211 (N_4211,N_3839,N_3924);
nand U4212 (N_4212,N_3836,N_3840);
xnor U4213 (N_4213,N_3779,N_3948);
nand U4214 (N_4214,N_3934,N_3922);
xor U4215 (N_4215,N_3801,N_3986);
and U4216 (N_4216,N_3886,N_3852);
and U4217 (N_4217,N_3763,N_3757);
nor U4218 (N_4218,N_3908,N_3875);
nor U4219 (N_4219,N_3900,N_3942);
xnor U4220 (N_4220,N_3933,N_3995);
xnor U4221 (N_4221,N_3876,N_3897);
nor U4222 (N_4222,N_3931,N_3817);
xnor U4223 (N_4223,N_3796,N_3850);
or U4224 (N_4224,N_3963,N_3855);
nor U4225 (N_4225,N_3804,N_3788);
or U4226 (N_4226,N_3855,N_3989);
nand U4227 (N_4227,N_3877,N_3890);
nand U4228 (N_4228,N_3898,N_3968);
xnor U4229 (N_4229,N_3838,N_3890);
or U4230 (N_4230,N_3960,N_3952);
nand U4231 (N_4231,N_3961,N_3760);
nor U4232 (N_4232,N_3982,N_3902);
xor U4233 (N_4233,N_3784,N_3968);
or U4234 (N_4234,N_3826,N_3928);
xnor U4235 (N_4235,N_3821,N_3767);
nand U4236 (N_4236,N_3795,N_3854);
or U4237 (N_4237,N_3889,N_3829);
nor U4238 (N_4238,N_3880,N_3860);
nand U4239 (N_4239,N_3955,N_3765);
nand U4240 (N_4240,N_3911,N_3944);
xor U4241 (N_4241,N_3778,N_3758);
nor U4242 (N_4242,N_3997,N_3828);
nor U4243 (N_4243,N_3821,N_3897);
nand U4244 (N_4244,N_3919,N_3811);
and U4245 (N_4245,N_3809,N_3949);
nor U4246 (N_4246,N_3935,N_3926);
nand U4247 (N_4247,N_3977,N_3879);
nor U4248 (N_4248,N_3984,N_3786);
xor U4249 (N_4249,N_3863,N_3859);
xnor U4250 (N_4250,N_4031,N_4182);
and U4251 (N_4251,N_4212,N_4044);
xor U4252 (N_4252,N_4187,N_4055);
nand U4253 (N_4253,N_4201,N_4092);
nor U4254 (N_4254,N_4150,N_4026);
or U4255 (N_4255,N_4239,N_4142);
nor U4256 (N_4256,N_4058,N_4101);
xnor U4257 (N_4257,N_4043,N_4116);
or U4258 (N_4258,N_4139,N_4246);
and U4259 (N_4259,N_4104,N_4036);
nor U4260 (N_4260,N_4033,N_4028);
or U4261 (N_4261,N_4180,N_4136);
or U4262 (N_4262,N_4048,N_4015);
or U4263 (N_4263,N_4222,N_4145);
or U4264 (N_4264,N_4225,N_4072);
nor U4265 (N_4265,N_4001,N_4042);
xnor U4266 (N_4266,N_4115,N_4087);
and U4267 (N_4267,N_4110,N_4007);
and U4268 (N_4268,N_4019,N_4181);
or U4269 (N_4269,N_4074,N_4069);
and U4270 (N_4270,N_4111,N_4119);
xor U4271 (N_4271,N_4062,N_4089);
xnor U4272 (N_4272,N_4234,N_4018);
and U4273 (N_4273,N_4020,N_4103);
or U4274 (N_4274,N_4146,N_4244);
xor U4275 (N_4275,N_4129,N_4094);
xnor U4276 (N_4276,N_4099,N_4170);
nor U4277 (N_4277,N_4236,N_4005);
and U4278 (N_4278,N_4230,N_4132);
nor U4279 (N_4279,N_4204,N_4191);
nand U4280 (N_4280,N_4071,N_4211);
and U4281 (N_4281,N_4137,N_4156);
and U4282 (N_4282,N_4004,N_4061);
nor U4283 (N_4283,N_4049,N_4199);
nand U4284 (N_4284,N_4093,N_4133);
or U4285 (N_4285,N_4091,N_4193);
nor U4286 (N_4286,N_4032,N_4034);
or U4287 (N_4287,N_4102,N_4192);
nor U4288 (N_4288,N_4154,N_4107);
nor U4289 (N_4289,N_4173,N_4175);
nand U4290 (N_4290,N_4114,N_4100);
and U4291 (N_4291,N_4027,N_4064);
nand U4292 (N_4292,N_4082,N_4118);
xor U4293 (N_4293,N_4214,N_4039);
xor U4294 (N_4294,N_4017,N_4210);
xor U4295 (N_4295,N_4079,N_4134);
and U4296 (N_4296,N_4120,N_4205);
or U4297 (N_4297,N_4000,N_4098);
xor U4298 (N_4298,N_4035,N_4096);
or U4299 (N_4299,N_4021,N_4179);
nand U4300 (N_4300,N_4127,N_4002);
nand U4301 (N_4301,N_4070,N_4147);
and U4302 (N_4302,N_4165,N_4029);
or U4303 (N_4303,N_4235,N_4190);
or U4304 (N_4304,N_4041,N_4090);
nand U4305 (N_4305,N_4149,N_4086);
nand U4306 (N_4306,N_4163,N_4243);
nand U4307 (N_4307,N_4059,N_4189);
and U4308 (N_4308,N_4112,N_4248);
and U4309 (N_4309,N_4057,N_4161);
or U4310 (N_4310,N_4078,N_4229);
nor U4311 (N_4311,N_4167,N_4196);
and U4312 (N_4312,N_4231,N_4172);
xnor U4313 (N_4313,N_4037,N_4218);
and U4314 (N_4314,N_4128,N_4108);
and U4315 (N_4315,N_4188,N_4085);
nor U4316 (N_4316,N_4171,N_4063);
and U4317 (N_4317,N_4117,N_4073);
and U4318 (N_4318,N_4008,N_4065);
and U4319 (N_4319,N_4077,N_4238);
or U4320 (N_4320,N_4138,N_4148);
and U4321 (N_4321,N_4153,N_4155);
nor U4322 (N_4322,N_4203,N_4249);
or U4323 (N_4323,N_4083,N_4232);
and U4324 (N_4324,N_4242,N_4075);
or U4325 (N_4325,N_4227,N_4054);
and U4326 (N_4326,N_4131,N_4162);
and U4327 (N_4327,N_4215,N_4095);
or U4328 (N_4328,N_4176,N_4228);
nand U4329 (N_4329,N_4233,N_4247);
nor U4330 (N_4330,N_4068,N_4053);
and U4331 (N_4331,N_4050,N_4030);
or U4332 (N_4332,N_4006,N_4224);
and U4333 (N_4333,N_4135,N_4194);
or U4334 (N_4334,N_4198,N_4076);
and U4335 (N_4335,N_4051,N_4144);
nand U4336 (N_4336,N_4217,N_4197);
and U4337 (N_4337,N_4124,N_4183);
or U4338 (N_4338,N_4024,N_4166);
or U4339 (N_4339,N_4056,N_4158);
nor U4340 (N_4340,N_4141,N_4003);
xor U4341 (N_4341,N_4178,N_4130);
nand U4342 (N_4342,N_4045,N_4174);
and U4343 (N_4343,N_4169,N_4164);
and U4344 (N_4344,N_4241,N_4200);
xor U4345 (N_4345,N_4226,N_4143);
or U4346 (N_4346,N_4184,N_4022);
nand U4347 (N_4347,N_4025,N_4195);
or U4348 (N_4348,N_4185,N_4223);
nor U4349 (N_4349,N_4207,N_4240);
nor U4350 (N_4350,N_4168,N_4152);
and U4351 (N_4351,N_4080,N_4220);
or U4352 (N_4352,N_4113,N_4109);
nand U4353 (N_4353,N_4216,N_4151);
xor U4354 (N_4354,N_4013,N_4010);
nor U4355 (N_4355,N_4206,N_4046);
nand U4356 (N_4356,N_4125,N_4213);
xor U4357 (N_4357,N_4081,N_4047);
xnor U4358 (N_4358,N_4084,N_4186);
nor U4359 (N_4359,N_4097,N_4038);
nand U4360 (N_4360,N_4123,N_4106);
nand U4361 (N_4361,N_4208,N_4209);
nand U4362 (N_4362,N_4011,N_4023);
or U4363 (N_4363,N_4012,N_4219);
nor U4364 (N_4364,N_4016,N_4014);
xor U4365 (N_4365,N_4009,N_4105);
or U4366 (N_4366,N_4067,N_4121);
or U4367 (N_4367,N_4088,N_4245);
nor U4368 (N_4368,N_4066,N_4237);
nor U4369 (N_4369,N_4202,N_4060);
nor U4370 (N_4370,N_4157,N_4159);
or U4371 (N_4371,N_4052,N_4140);
nand U4372 (N_4372,N_4221,N_4126);
or U4373 (N_4373,N_4177,N_4160);
or U4374 (N_4374,N_4122,N_4040);
and U4375 (N_4375,N_4170,N_4090);
or U4376 (N_4376,N_4205,N_4135);
or U4377 (N_4377,N_4164,N_4006);
and U4378 (N_4378,N_4131,N_4011);
and U4379 (N_4379,N_4116,N_4190);
and U4380 (N_4380,N_4025,N_4013);
nor U4381 (N_4381,N_4175,N_4180);
nor U4382 (N_4382,N_4204,N_4237);
nand U4383 (N_4383,N_4022,N_4220);
xor U4384 (N_4384,N_4081,N_4028);
or U4385 (N_4385,N_4105,N_4036);
nand U4386 (N_4386,N_4166,N_4100);
xnor U4387 (N_4387,N_4109,N_4048);
nand U4388 (N_4388,N_4022,N_4249);
nor U4389 (N_4389,N_4248,N_4071);
nor U4390 (N_4390,N_4135,N_4081);
xnor U4391 (N_4391,N_4210,N_4186);
nor U4392 (N_4392,N_4096,N_4117);
or U4393 (N_4393,N_4001,N_4241);
nor U4394 (N_4394,N_4214,N_4065);
nand U4395 (N_4395,N_4117,N_4052);
xor U4396 (N_4396,N_4154,N_4010);
and U4397 (N_4397,N_4247,N_4116);
or U4398 (N_4398,N_4234,N_4232);
nor U4399 (N_4399,N_4084,N_4106);
nor U4400 (N_4400,N_4145,N_4097);
nand U4401 (N_4401,N_4244,N_4072);
nand U4402 (N_4402,N_4016,N_4086);
and U4403 (N_4403,N_4042,N_4076);
nor U4404 (N_4404,N_4147,N_4148);
xnor U4405 (N_4405,N_4094,N_4188);
xor U4406 (N_4406,N_4185,N_4130);
xor U4407 (N_4407,N_4068,N_4025);
xnor U4408 (N_4408,N_4142,N_4167);
nand U4409 (N_4409,N_4156,N_4005);
or U4410 (N_4410,N_4115,N_4175);
and U4411 (N_4411,N_4170,N_4120);
and U4412 (N_4412,N_4213,N_4108);
and U4413 (N_4413,N_4242,N_4038);
and U4414 (N_4414,N_4054,N_4238);
nor U4415 (N_4415,N_4231,N_4100);
or U4416 (N_4416,N_4130,N_4108);
and U4417 (N_4417,N_4015,N_4067);
nand U4418 (N_4418,N_4178,N_4213);
xnor U4419 (N_4419,N_4050,N_4068);
and U4420 (N_4420,N_4173,N_4239);
xnor U4421 (N_4421,N_4217,N_4240);
xor U4422 (N_4422,N_4053,N_4028);
and U4423 (N_4423,N_4220,N_4082);
and U4424 (N_4424,N_4080,N_4111);
nor U4425 (N_4425,N_4223,N_4069);
nor U4426 (N_4426,N_4210,N_4085);
or U4427 (N_4427,N_4247,N_4081);
or U4428 (N_4428,N_4125,N_4031);
and U4429 (N_4429,N_4047,N_4208);
or U4430 (N_4430,N_4112,N_4081);
and U4431 (N_4431,N_4137,N_4050);
nand U4432 (N_4432,N_4217,N_4143);
and U4433 (N_4433,N_4093,N_4076);
nor U4434 (N_4434,N_4220,N_4065);
nand U4435 (N_4435,N_4219,N_4180);
and U4436 (N_4436,N_4022,N_4012);
nand U4437 (N_4437,N_4094,N_4242);
nor U4438 (N_4438,N_4171,N_4139);
xnor U4439 (N_4439,N_4122,N_4133);
and U4440 (N_4440,N_4218,N_4068);
or U4441 (N_4441,N_4082,N_4084);
or U4442 (N_4442,N_4195,N_4038);
xnor U4443 (N_4443,N_4193,N_4183);
or U4444 (N_4444,N_4138,N_4236);
nand U4445 (N_4445,N_4168,N_4199);
nor U4446 (N_4446,N_4114,N_4075);
xor U4447 (N_4447,N_4088,N_4093);
and U4448 (N_4448,N_4188,N_4114);
nor U4449 (N_4449,N_4203,N_4052);
xor U4450 (N_4450,N_4239,N_4032);
xnor U4451 (N_4451,N_4139,N_4127);
nor U4452 (N_4452,N_4066,N_4233);
or U4453 (N_4453,N_4133,N_4053);
nand U4454 (N_4454,N_4126,N_4100);
and U4455 (N_4455,N_4080,N_4212);
nor U4456 (N_4456,N_4196,N_4147);
and U4457 (N_4457,N_4118,N_4079);
nand U4458 (N_4458,N_4004,N_4046);
nor U4459 (N_4459,N_4246,N_4192);
and U4460 (N_4460,N_4025,N_4189);
or U4461 (N_4461,N_4004,N_4244);
and U4462 (N_4462,N_4135,N_4064);
nor U4463 (N_4463,N_4231,N_4105);
xor U4464 (N_4464,N_4188,N_4218);
nand U4465 (N_4465,N_4039,N_4072);
xnor U4466 (N_4466,N_4002,N_4209);
nor U4467 (N_4467,N_4230,N_4111);
nand U4468 (N_4468,N_4086,N_4063);
nor U4469 (N_4469,N_4051,N_4104);
and U4470 (N_4470,N_4004,N_4049);
and U4471 (N_4471,N_4100,N_4030);
and U4472 (N_4472,N_4196,N_4086);
nand U4473 (N_4473,N_4218,N_4179);
nand U4474 (N_4474,N_4209,N_4158);
or U4475 (N_4475,N_4046,N_4125);
and U4476 (N_4476,N_4012,N_4195);
xnor U4477 (N_4477,N_4078,N_4001);
or U4478 (N_4478,N_4195,N_4187);
and U4479 (N_4479,N_4137,N_4066);
nand U4480 (N_4480,N_4156,N_4239);
or U4481 (N_4481,N_4173,N_4231);
xnor U4482 (N_4482,N_4014,N_4092);
nand U4483 (N_4483,N_4216,N_4200);
nor U4484 (N_4484,N_4015,N_4068);
xnor U4485 (N_4485,N_4084,N_4051);
nand U4486 (N_4486,N_4177,N_4186);
nand U4487 (N_4487,N_4208,N_4110);
and U4488 (N_4488,N_4069,N_4022);
nor U4489 (N_4489,N_4080,N_4091);
or U4490 (N_4490,N_4013,N_4082);
nand U4491 (N_4491,N_4068,N_4216);
and U4492 (N_4492,N_4143,N_4047);
nand U4493 (N_4493,N_4034,N_4008);
nor U4494 (N_4494,N_4249,N_4027);
xnor U4495 (N_4495,N_4169,N_4181);
and U4496 (N_4496,N_4208,N_4019);
or U4497 (N_4497,N_4235,N_4194);
or U4498 (N_4498,N_4167,N_4249);
nand U4499 (N_4499,N_4198,N_4163);
nand U4500 (N_4500,N_4325,N_4395);
and U4501 (N_4501,N_4489,N_4288);
or U4502 (N_4502,N_4475,N_4353);
nand U4503 (N_4503,N_4410,N_4289);
and U4504 (N_4504,N_4321,N_4338);
nor U4505 (N_4505,N_4394,N_4432);
xor U4506 (N_4506,N_4258,N_4380);
and U4507 (N_4507,N_4402,N_4444);
xor U4508 (N_4508,N_4320,N_4460);
and U4509 (N_4509,N_4265,N_4332);
or U4510 (N_4510,N_4490,N_4401);
xor U4511 (N_4511,N_4278,N_4385);
or U4512 (N_4512,N_4326,N_4366);
and U4513 (N_4513,N_4373,N_4318);
or U4514 (N_4514,N_4340,N_4261);
nor U4515 (N_4515,N_4440,N_4372);
and U4516 (N_4516,N_4294,N_4364);
xor U4517 (N_4517,N_4419,N_4271);
and U4518 (N_4518,N_4491,N_4300);
nand U4519 (N_4519,N_4314,N_4267);
nor U4520 (N_4520,N_4350,N_4264);
and U4521 (N_4521,N_4421,N_4437);
xnor U4522 (N_4522,N_4290,N_4367);
or U4523 (N_4523,N_4461,N_4442);
xor U4524 (N_4524,N_4428,N_4420);
nor U4525 (N_4525,N_4487,N_4315);
or U4526 (N_4526,N_4473,N_4287);
nor U4527 (N_4527,N_4447,N_4497);
xnor U4528 (N_4528,N_4336,N_4406);
nand U4529 (N_4529,N_4416,N_4408);
nand U4530 (N_4530,N_4352,N_4455);
nand U4531 (N_4531,N_4369,N_4431);
nor U4532 (N_4532,N_4349,N_4306);
xnor U4533 (N_4533,N_4342,N_4302);
and U4534 (N_4534,N_4310,N_4371);
nand U4535 (N_4535,N_4331,N_4355);
nand U4536 (N_4536,N_4422,N_4313);
xnor U4537 (N_4537,N_4301,N_4478);
and U4538 (N_4538,N_4370,N_4260);
nor U4539 (N_4539,N_4480,N_4386);
or U4540 (N_4540,N_4347,N_4275);
nand U4541 (N_4541,N_4304,N_4412);
or U4542 (N_4542,N_4327,N_4383);
and U4543 (N_4543,N_4413,N_4345);
xor U4544 (N_4544,N_4441,N_4333);
nand U4545 (N_4545,N_4423,N_4256);
and U4546 (N_4546,N_4493,N_4456);
and U4547 (N_4547,N_4449,N_4293);
nor U4548 (N_4548,N_4439,N_4409);
nor U4549 (N_4549,N_4329,N_4381);
nor U4550 (N_4550,N_4341,N_4463);
xnor U4551 (N_4551,N_4479,N_4376);
xnor U4552 (N_4552,N_4317,N_4282);
nor U4553 (N_4553,N_4362,N_4468);
or U4554 (N_4554,N_4330,N_4450);
or U4555 (N_4555,N_4356,N_4360);
and U4556 (N_4556,N_4426,N_4397);
xor U4557 (N_4557,N_4443,N_4251);
and U4558 (N_4558,N_4472,N_4492);
or U4559 (N_4559,N_4453,N_4465);
nand U4560 (N_4560,N_4281,N_4375);
or U4561 (N_4561,N_4476,N_4398);
and U4562 (N_4562,N_4291,N_4407);
xor U4563 (N_4563,N_4430,N_4494);
nor U4564 (N_4564,N_4404,N_4266);
nand U4565 (N_4565,N_4400,N_4448);
or U4566 (N_4566,N_4252,N_4484);
xnor U4567 (N_4567,N_4257,N_4393);
or U4568 (N_4568,N_4469,N_4378);
nand U4569 (N_4569,N_4481,N_4295);
nand U4570 (N_4570,N_4464,N_4477);
nand U4571 (N_4571,N_4496,N_4319);
nand U4572 (N_4572,N_4284,N_4458);
or U4573 (N_4573,N_4296,N_4414);
or U4574 (N_4574,N_4312,N_4466);
nor U4575 (N_4575,N_4399,N_4499);
nor U4576 (N_4576,N_4322,N_4274);
nor U4577 (N_4577,N_4280,N_4323);
nor U4578 (N_4578,N_4417,N_4311);
xnor U4579 (N_4579,N_4299,N_4368);
and U4580 (N_4580,N_4396,N_4451);
and U4581 (N_4581,N_4390,N_4357);
nand U4582 (N_4582,N_4348,N_4298);
xnor U4583 (N_4583,N_4337,N_4305);
and U4584 (N_4584,N_4415,N_4474);
or U4585 (N_4585,N_4259,N_4485);
nor U4586 (N_4586,N_4498,N_4316);
nor U4587 (N_4587,N_4339,N_4433);
nor U4588 (N_4588,N_4405,N_4324);
and U4589 (N_4589,N_4403,N_4361);
nand U4590 (N_4590,N_4384,N_4268);
nand U4591 (N_4591,N_4358,N_4262);
nor U4592 (N_4592,N_4425,N_4411);
nand U4593 (N_4593,N_4292,N_4276);
or U4594 (N_4594,N_4270,N_4436);
nor U4595 (N_4595,N_4427,N_4363);
nand U4596 (N_4596,N_4269,N_4354);
xnor U4597 (N_4597,N_4454,N_4263);
or U4598 (N_4598,N_4471,N_4277);
nand U4599 (N_4599,N_4346,N_4470);
nand U4600 (N_4600,N_4374,N_4389);
or U4601 (N_4601,N_4387,N_4344);
and U4602 (N_4602,N_4379,N_4273);
and U4603 (N_4603,N_4377,N_4285);
nor U4604 (N_4604,N_4392,N_4459);
nand U4605 (N_4605,N_4334,N_4457);
xnor U4606 (N_4606,N_4254,N_4438);
or U4607 (N_4607,N_4359,N_4435);
nor U4608 (N_4608,N_4418,N_4482);
nor U4609 (N_4609,N_4328,N_4297);
xor U4610 (N_4610,N_4343,N_4382);
or U4611 (N_4611,N_4445,N_4452);
nand U4612 (N_4612,N_4488,N_4365);
nor U4613 (N_4613,N_4303,N_4467);
xor U4614 (N_4614,N_4351,N_4308);
xnor U4615 (N_4615,N_4253,N_4283);
nor U4616 (N_4616,N_4309,N_4307);
nor U4617 (N_4617,N_4434,N_4486);
and U4618 (N_4618,N_4286,N_4279);
xnor U4619 (N_4619,N_4391,N_4424);
nor U4620 (N_4620,N_4255,N_4446);
xnor U4621 (N_4621,N_4483,N_4429);
nor U4622 (N_4622,N_4250,N_4388);
nand U4623 (N_4623,N_4462,N_4272);
and U4624 (N_4624,N_4335,N_4495);
and U4625 (N_4625,N_4432,N_4487);
xor U4626 (N_4626,N_4333,N_4477);
and U4627 (N_4627,N_4390,N_4476);
and U4628 (N_4628,N_4382,N_4394);
xor U4629 (N_4629,N_4350,N_4464);
xnor U4630 (N_4630,N_4256,N_4419);
nor U4631 (N_4631,N_4307,N_4435);
xnor U4632 (N_4632,N_4473,N_4325);
nor U4633 (N_4633,N_4427,N_4473);
nand U4634 (N_4634,N_4415,N_4427);
nand U4635 (N_4635,N_4336,N_4408);
and U4636 (N_4636,N_4270,N_4262);
nor U4637 (N_4637,N_4495,N_4442);
nand U4638 (N_4638,N_4444,N_4470);
or U4639 (N_4639,N_4260,N_4459);
nor U4640 (N_4640,N_4283,N_4491);
and U4641 (N_4641,N_4391,N_4261);
nand U4642 (N_4642,N_4310,N_4397);
nor U4643 (N_4643,N_4378,N_4451);
nand U4644 (N_4644,N_4455,N_4339);
or U4645 (N_4645,N_4437,N_4379);
nand U4646 (N_4646,N_4378,N_4300);
xor U4647 (N_4647,N_4401,N_4271);
or U4648 (N_4648,N_4491,N_4353);
and U4649 (N_4649,N_4461,N_4275);
nand U4650 (N_4650,N_4280,N_4343);
nand U4651 (N_4651,N_4352,N_4468);
and U4652 (N_4652,N_4337,N_4296);
and U4653 (N_4653,N_4499,N_4256);
nor U4654 (N_4654,N_4455,N_4399);
and U4655 (N_4655,N_4424,N_4253);
nor U4656 (N_4656,N_4399,N_4344);
and U4657 (N_4657,N_4455,N_4416);
nor U4658 (N_4658,N_4272,N_4282);
or U4659 (N_4659,N_4473,N_4464);
xor U4660 (N_4660,N_4454,N_4492);
nand U4661 (N_4661,N_4328,N_4318);
and U4662 (N_4662,N_4389,N_4288);
or U4663 (N_4663,N_4402,N_4460);
or U4664 (N_4664,N_4372,N_4272);
and U4665 (N_4665,N_4378,N_4430);
or U4666 (N_4666,N_4490,N_4290);
xor U4667 (N_4667,N_4437,N_4468);
nor U4668 (N_4668,N_4276,N_4278);
nor U4669 (N_4669,N_4378,N_4477);
or U4670 (N_4670,N_4462,N_4354);
xor U4671 (N_4671,N_4403,N_4418);
nand U4672 (N_4672,N_4363,N_4469);
and U4673 (N_4673,N_4423,N_4445);
xor U4674 (N_4674,N_4332,N_4382);
and U4675 (N_4675,N_4406,N_4453);
nor U4676 (N_4676,N_4399,N_4347);
xnor U4677 (N_4677,N_4428,N_4449);
and U4678 (N_4678,N_4433,N_4408);
and U4679 (N_4679,N_4271,N_4277);
and U4680 (N_4680,N_4378,N_4474);
and U4681 (N_4681,N_4272,N_4294);
and U4682 (N_4682,N_4308,N_4266);
nor U4683 (N_4683,N_4278,N_4491);
xor U4684 (N_4684,N_4363,N_4488);
and U4685 (N_4685,N_4306,N_4284);
and U4686 (N_4686,N_4375,N_4383);
and U4687 (N_4687,N_4352,N_4347);
nand U4688 (N_4688,N_4274,N_4302);
and U4689 (N_4689,N_4302,N_4446);
xnor U4690 (N_4690,N_4498,N_4429);
nor U4691 (N_4691,N_4424,N_4410);
nand U4692 (N_4692,N_4302,N_4267);
nand U4693 (N_4693,N_4271,N_4457);
nand U4694 (N_4694,N_4464,N_4495);
or U4695 (N_4695,N_4320,N_4372);
and U4696 (N_4696,N_4417,N_4462);
nand U4697 (N_4697,N_4486,N_4389);
nand U4698 (N_4698,N_4276,N_4311);
and U4699 (N_4699,N_4335,N_4390);
xnor U4700 (N_4700,N_4448,N_4352);
and U4701 (N_4701,N_4492,N_4326);
and U4702 (N_4702,N_4291,N_4416);
nand U4703 (N_4703,N_4340,N_4275);
nor U4704 (N_4704,N_4434,N_4482);
xnor U4705 (N_4705,N_4493,N_4483);
nand U4706 (N_4706,N_4365,N_4342);
or U4707 (N_4707,N_4269,N_4487);
nand U4708 (N_4708,N_4463,N_4447);
or U4709 (N_4709,N_4328,N_4443);
or U4710 (N_4710,N_4371,N_4395);
or U4711 (N_4711,N_4312,N_4428);
nand U4712 (N_4712,N_4475,N_4320);
xor U4713 (N_4713,N_4468,N_4341);
nor U4714 (N_4714,N_4390,N_4318);
nor U4715 (N_4715,N_4356,N_4275);
nand U4716 (N_4716,N_4326,N_4333);
nand U4717 (N_4717,N_4343,N_4411);
or U4718 (N_4718,N_4469,N_4362);
nand U4719 (N_4719,N_4359,N_4363);
nand U4720 (N_4720,N_4494,N_4282);
nand U4721 (N_4721,N_4480,N_4430);
nor U4722 (N_4722,N_4254,N_4402);
xnor U4723 (N_4723,N_4444,N_4483);
and U4724 (N_4724,N_4345,N_4492);
xor U4725 (N_4725,N_4282,N_4316);
nand U4726 (N_4726,N_4367,N_4300);
xnor U4727 (N_4727,N_4409,N_4416);
xnor U4728 (N_4728,N_4479,N_4427);
xor U4729 (N_4729,N_4297,N_4448);
nand U4730 (N_4730,N_4429,N_4318);
or U4731 (N_4731,N_4270,N_4280);
and U4732 (N_4732,N_4483,N_4469);
nor U4733 (N_4733,N_4469,N_4422);
xnor U4734 (N_4734,N_4355,N_4372);
nand U4735 (N_4735,N_4498,N_4306);
or U4736 (N_4736,N_4308,N_4424);
nor U4737 (N_4737,N_4347,N_4445);
xor U4738 (N_4738,N_4396,N_4341);
nor U4739 (N_4739,N_4499,N_4443);
or U4740 (N_4740,N_4318,N_4496);
nand U4741 (N_4741,N_4360,N_4490);
and U4742 (N_4742,N_4489,N_4490);
nand U4743 (N_4743,N_4294,N_4250);
nor U4744 (N_4744,N_4276,N_4350);
nor U4745 (N_4745,N_4261,N_4304);
xnor U4746 (N_4746,N_4444,N_4255);
nor U4747 (N_4747,N_4397,N_4285);
xor U4748 (N_4748,N_4363,N_4327);
nand U4749 (N_4749,N_4288,N_4305);
and U4750 (N_4750,N_4739,N_4536);
nand U4751 (N_4751,N_4563,N_4551);
nor U4752 (N_4752,N_4597,N_4560);
nand U4753 (N_4753,N_4729,N_4727);
and U4754 (N_4754,N_4590,N_4733);
nand U4755 (N_4755,N_4662,N_4743);
and U4756 (N_4756,N_4701,N_4591);
xor U4757 (N_4757,N_4648,N_4512);
nor U4758 (N_4758,N_4587,N_4691);
xnor U4759 (N_4759,N_4737,N_4695);
or U4760 (N_4760,N_4593,N_4725);
and U4761 (N_4761,N_4564,N_4717);
nor U4762 (N_4762,N_4653,N_4632);
xor U4763 (N_4763,N_4613,N_4507);
xor U4764 (N_4764,N_4710,N_4672);
xnor U4765 (N_4765,N_4579,N_4630);
and U4766 (N_4766,N_4555,N_4643);
nand U4767 (N_4767,N_4712,N_4610);
and U4768 (N_4768,N_4547,N_4523);
nand U4769 (N_4769,N_4618,N_4520);
nand U4770 (N_4770,N_4627,N_4576);
nor U4771 (N_4771,N_4654,N_4562);
and U4772 (N_4772,N_4708,N_4616);
nor U4773 (N_4773,N_4641,N_4696);
nand U4774 (N_4774,N_4693,N_4736);
and U4775 (N_4775,N_4516,N_4598);
xor U4776 (N_4776,N_4561,N_4675);
nor U4777 (N_4777,N_4645,N_4676);
or U4778 (N_4778,N_4521,N_4724);
xor U4779 (N_4779,N_4678,N_4522);
xnor U4780 (N_4780,N_4570,N_4742);
xor U4781 (N_4781,N_4651,N_4673);
or U4782 (N_4782,N_4625,N_4646);
xnor U4783 (N_4783,N_4619,N_4671);
xor U4784 (N_4784,N_4661,N_4720);
nor U4785 (N_4785,N_4663,N_4502);
xnor U4786 (N_4786,N_4689,N_4549);
or U4787 (N_4787,N_4510,N_4674);
nand U4788 (N_4788,N_4734,N_4707);
nand U4789 (N_4789,N_4596,N_4740);
and U4790 (N_4790,N_4548,N_4706);
xor U4791 (N_4791,N_4670,N_4732);
nor U4792 (N_4792,N_4554,N_4668);
or U4793 (N_4793,N_4718,N_4532);
nand U4794 (N_4794,N_4544,N_4639);
nand U4795 (N_4795,N_4543,N_4575);
or U4796 (N_4796,N_4601,N_4665);
nor U4797 (N_4797,N_4711,N_4682);
nor U4798 (N_4798,N_4650,N_4621);
xor U4799 (N_4799,N_4571,N_4624);
nand U4800 (N_4800,N_4538,N_4716);
nand U4801 (N_4801,N_4633,N_4715);
nor U4802 (N_4802,N_4531,N_4735);
nand U4803 (N_4803,N_4514,N_4588);
nand U4804 (N_4804,N_4535,N_4684);
xor U4805 (N_4805,N_4638,N_4617);
xnor U4806 (N_4806,N_4569,N_4629);
xor U4807 (N_4807,N_4541,N_4647);
or U4808 (N_4808,N_4685,N_4565);
and U4809 (N_4809,N_4745,N_4608);
or U4810 (N_4810,N_4686,N_4605);
nor U4811 (N_4811,N_4524,N_4726);
or U4812 (N_4812,N_4628,N_4603);
nand U4813 (N_4813,N_4594,N_4635);
nand U4814 (N_4814,N_4609,N_4660);
xnor U4815 (N_4815,N_4595,N_4679);
nand U4816 (N_4816,N_4604,N_4700);
nor U4817 (N_4817,N_4713,N_4704);
nand U4818 (N_4818,N_4583,N_4688);
and U4819 (N_4819,N_4659,N_4527);
or U4820 (N_4820,N_4748,N_4620);
and U4821 (N_4821,N_4586,N_4644);
and U4822 (N_4822,N_4500,N_4669);
and U4823 (N_4823,N_4505,N_4584);
nand U4824 (N_4824,N_4506,N_4656);
nor U4825 (N_4825,N_4622,N_4600);
or U4826 (N_4826,N_4657,N_4690);
and U4827 (N_4827,N_4746,N_4658);
and U4828 (N_4828,N_4687,N_4714);
nor U4829 (N_4829,N_4612,N_4655);
or U4830 (N_4830,N_4649,N_4517);
nor U4831 (N_4831,N_4666,N_4537);
and U4832 (N_4832,N_4580,N_4703);
or U4833 (N_4833,N_4556,N_4529);
nand U4834 (N_4834,N_4722,N_4738);
and U4835 (N_4835,N_4747,N_4567);
or U4836 (N_4836,N_4615,N_4592);
and U4837 (N_4837,N_4744,N_4719);
and U4838 (N_4838,N_4721,N_4542);
or U4839 (N_4839,N_4557,N_4636);
or U4840 (N_4840,N_4545,N_4574);
nor U4841 (N_4841,N_4578,N_4585);
nand U4842 (N_4842,N_4741,N_4642);
or U4843 (N_4843,N_4681,N_4634);
or U4844 (N_4844,N_4640,N_4515);
xnor U4845 (N_4845,N_4581,N_4589);
nand U4846 (N_4846,N_4683,N_4553);
or U4847 (N_4847,N_4749,N_4568);
nor U4848 (N_4848,N_4623,N_4731);
nor U4849 (N_4849,N_4677,N_4508);
and U4850 (N_4850,N_4631,N_4680);
nor U4851 (N_4851,N_4552,N_4540);
xor U4852 (N_4852,N_4559,N_4511);
and U4853 (N_4853,N_4546,N_4652);
nand U4854 (N_4854,N_4599,N_4558);
and U4855 (N_4855,N_4582,N_4528);
or U4856 (N_4856,N_4534,N_4503);
xnor U4857 (N_4857,N_4539,N_4667);
nand U4858 (N_4858,N_4637,N_4504);
nor U4859 (N_4859,N_4728,N_4602);
and U4860 (N_4860,N_4519,N_4730);
nor U4861 (N_4861,N_4611,N_4626);
and U4862 (N_4862,N_4509,N_4723);
and U4863 (N_4863,N_4606,N_4577);
or U4864 (N_4864,N_4566,N_4501);
nor U4865 (N_4865,N_4692,N_4614);
nand U4866 (N_4866,N_4518,N_4573);
nand U4867 (N_4867,N_4697,N_4530);
or U4868 (N_4868,N_4525,N_4664);
and U4869 (N_4869,N_4513,N_4705);
and U4870 (N_4870,N_4533,N_4550);
and U4871 (N_4871,N_4699,N_4698);
or U4872 (N_4872,N_4702,N_4607);
nor U4873 (N_4873,N_4572,N_4526);
xnor U4874 (N_4874,N_4694,N_4709);
or U4875 (N_4875,N_4548,N_4680);
and U4876 (N_4876,N_4552,N_4649);
or U4877 (N_4877,N_4699,N_4611);
nand U4878 (N_4878,N_4574,N_4692);
or U4879 (N_4879,N_4712,N_4558);
or U4880 (N_4880,N_4651,N_4717);
nand U4881 (N_4881,N_4695,N_4717);
and U4882 (N_4882,N_4684,N_4729);
or U4883 (N_4883,N_4600,N_4627);
nor U4884 (N_4884,N_4738,N_4664);
and U4885 (N_4885,N_4606,N_4674);
or U4886 (N_4886,N_4721,N_4511);
nand U4887 (N_4887,N_4510,N_4550);
nor U4888 (N_4888,N_4560,N_4626);
or U4889 (N_4889,N_4590,N_4564);
and U4890 (N_4890,N_4589,N_4502);
xor U4891 (N_4891,N_4704,N_4555);
or U4892 (N_4892,N_4554,N_4733);
nor U4893 (N_4893,N_4624,N_4593);
or U4894 (N_4894,N_4644,N_4680);
xor U4895 (N_4895,N_4653,N_4635);
and U4896 (N_4896,N_4693,N_4579);
nand U4897 (N_4897,N_4718,N_4651);
xor U4898 (N_4898,N_4506,N_4636);
nor U4899 (N_4899,N_4644,N_4739);
and U4900 (N_4900,N_4718,N_4674);
and U4901 (N_4901,N_4687,N_4710);
or U4902 (N_4902,N_4682,N_4506);
nand U4903 (N_4903,N_4551,N_4512);
xnor U4904 (N_4904,N_4526,N_4680);
and U4905 (N_4905,N_4677,N_4520);
and U4906 (N_4906,N_4574,N_4562);
or U4907 (N_4907,N_4667,N_4744);
nor U4908 (N_4908,N_4698,N_4548);
and U4909 (N_4909,N_4674,N_4723);
or U4910 (N_4910,N_4583,N_4685);
or U4911 (N_4911,N_4545,N_4679);
nand U4912 (N_4912,N_4563,N_4721);
nor U4913 (N_4913,N_4620,N_4688);
nor U4914 (N_4914,N_4727,N_4519);
nor U4915 (N_4915,N_4706,N_4735);
xnor U4916 (N_4916,N_4669,N_4610);
and U4917 (N_4917,N_4654,N_4571);
or U4918 (N_4918,N_4514,N_4508);
xor U4919 (N_4919,N_4589,N_4573);
xnor U4920 (N_4920,N_4610,N_4595);
nor U4921 (N_4921,N_4542,N_4575);
and U4922 (N_4922,N_4617,N_4631);
or U4923 (N_4923,N_4622,N_4675);
nand U4924 (N_4924,N_4515,N_4670);
xnor U4925 (N_4925,N_4574,N_4525);
xor U4926 (N_4926,N_4632,N_4503);
xor U4927 (N_4927,N_4711,N_4744);
and U4928 (N_4928,N_4732,N_4735);
nor U4929 (N_4929,N_4706,N_4724);
nand U4930 (N_4930,N_4559,N_4732);
xor U4931 (N_4931,N_4519,N_4514);
and U4932 (N_4932,N_4665,N_4598);
nand U4933 (N_4933,N_4526,N_4610);
xor U4934 (N_4934,N_4572,N_4604);
and U4935 (N_4935,N_4647,N_4726);
and U4936 (N_4936,N_4597,N_4701);
nor U4937 (N_4937,N_4520,N_4700);
and U4938 (N_4938,N_4548,N_4525);
and U4939 (N_4939,N_4555,N_4610);
xor U4940 (N_4940,N_4513,N_4637);
or U4941 (N_4941,N_4625,N_4670);
nor U4942 (N_4942,N_4556,N_4672);
nand U4943 (N_4943,N_4611,N_4583);
nand U4944 (N_4944,N_4586,N_4599);
nand U4945 (N_4945,N_4508,N_4576);
or U4946 (N_4946,N_4528,N_4615);
and U4947 (N_4947,N_4649,N_4740);
nand U4948 (N_4948,N_4608,N_4531);
or U4949 (N_4949,N_4617,N_4722);
nand U4950 (N_4950,N_4727,N_4521);
xor U4951 (N_4951,N_4557,N_4730);
nor U4952 (N_4952,N_4719,N_4549);
xnor U4953 (N_4953,N_4733,N_4654);
or U4954 (N_4954,N_4604,N_4609);
nand U4955 (N_4955,N_4655,N_4664);
nand U4956 (N_4956,N_4597,N_4669);
xnor U4957 (N_4957,N_4731,N_4537);
nor U4958 (N_4958,N_4688,N_4578);
or U4959 (N_4959,N_4519,N_4578);
and U4960 (N_4960,N_4514,N_4653);
and U4961 (N_4961,N_4561,N_4571);
nor U4962 (N_4962,N_4642,N_4706);
or U4963 (N_4963,N_4581,N_4732);
nand U4964 (N_4964,N_4592,N_4523);
and U4965 (N_4965,N_4733,N_4501);
or U4966 (N_4966,N_4538,N_4586);
and U4967 (N_4967,N_4710,N_4569);
or U4968 (N_4968,N_4653,N_4640);
or U4969 (N_4969,N_4663,N_4565);
xor U4970 (N_4970,N_4688,N_4682);
or U4971 (N_4971,N_4540,N_4725);
nand U4972 (N_4972,N_4733,N_4638);
xnor U4973 (N_4973,N_4707,N_4681);
or U4974 (N_4974,N_4604,N_4695);
nor U4975 (N_4975,N_4687,N_4688);
and U4976 (N_4976,N_4549,N_4735);
or U4977 (N_4977,N_4541,N_4633);
and U4978 (N_4978,N_4624,N_4607);
nor U4979 (N_4979,N_4651,N_4746);
or U4980 (N_4980,N_4644,N_4723);
and U4981 (N_4981,N_4509,N_4556);
nand U4982 (N_4982,N_4662,N_4728);
nand U4983 (N_4983,N_4570,N_4704);
and U4984 (N_4984,N_4737,N_4636);
xnor U4985 (N_4985,N_4683,N_4530);
nand U4986 (N_4986,N_4555,N_4646);
xnor U4987 (N_4987,N_4634,N_4604);
nand U4988 (N_4988,N_4661,N_4674);
xor U4989 (N_4989,N_4665,N_4597);
or U4990 (N_4990,N_4596,N_4598);
xor U4991 (N_4991,N_4568,N_4535);
nor U4992 (N_4992,N_4657,N_4716);
nand U4993 (N_4993,N_4639,N_4518);
or U4994 (N_4994,N_4546,N_4670);
or U4995 (N_4995,N_4631,N_4607);
nand U4996 (N_4996,N_4652,N_4737);
nand U4997 (N_4997,N_4585,N_4501);
nand U4998 (N_4998,N_4523,N_4651);
nand U4999 (N_4999,N_4559,N_4598);
and U5000 (N_5000,N_4974,N_4851);
nand U5001 (N_5001,N_4752,N_4891);
nand U5002 (N_5002,N_4826,N_4967);
nand U5003 (N_5003,N_4757,N_4866);
xnor U5004 (N_5004,N_4846,N_4875);
nand U5005 (N_5005,N_4986,N_4801);
and U5006 (N_5006,N_4840,N_4820);
xor U5007 (N_5007,N_4992,N_4969);
nand U5008 (N_5008,N_4936,N_4965);
and U5009 (N_5009,N_4937,N_4772);
xor U5010 (N_5010,N_4802,N_4951);
or U5011 (N_5011,N_4862,N_4913);
or U5012 (N_5012,N_4993,N_4779);
or U5013 (N_5013,N_4943,N_4878);
xnor U5014 (N_5014,N_4976,N_4865);
or U5015 (N_5015,N_4977,N_4784);
nand U5016 (N_5016,N_4896,N_4956);
and U5017 (N_5017,N_4983,N_4910);
or U5018 (N_5018,N_4980,N_4822);
xnor U5019 (N_5019,N_4829,N_4867);
xor U5020 (N_5020,N_4817,N_4796);
and U5021 (N_5021,N_4984,N_4894);
and U5022 (N_5022,N_4985,N_4755);
nand U5023 (N_5023,N_4856,N_4957);
xor U5024 (N_5024,N_4893,N_4958);
xor U5025 (N_5025,N_4869,N_4847);
xnor U5026 (N_5026,N_4860,N_4898);
or U5027 (N_5027,N_4837,N_4979);
and U5028 (N_5028,N_4803,N_4787);
xnor U5029 (N_5029,N_4835,N_4874);
or U5030 (N_5030,N_4827,N_4991);
nand U5031 (N_5031,N_4909,N_4999);
or U5032 (N_5032,N_4816,N_4794);
nand U5033 (N_5033,N_4906,N_4915);
xor U5034 (N_5034,N_4836,N_4804);
nor U5035 (N_5035,N_4927,N_4844);
or U5036 (N_5036,N_4806,N_4933);
nor U5037 (N_5037,N_4814,N_4810);
nand U5038 (N_5038,N_4761,N_4883);
nor U5039 (N_5039,N_4899,N_4811);
xnor U5040 (N_5040,N_4885,N_4750);
nor U5041 (N_5041,N_4934,N_4897);
and U5042 (N_5042,N_4978,N_4926);
or U5043 (N_5043,N_4948,N_4981);
or U5044 (N_5044,N_4854,N_4920);
and U5045 (N_5045,N_4873,N_4895);
nor U5046 (N_5046,N_4905,N_4950);
xnor U5047 (N_5047,N_4903,N_4925);
xor U5048 (N_5048,N_4962,N_4793);
and U5049 (N_5049,N_4799,N_4959);
xnor U5050 (N_5050,N_4759,N_4975);
and U5051 (N_5051,N_4908,N_4767);
or U5052 (N_5052,N_4795,N_4886);
and U5053 (N_5053,N_4941,N_4988);
or U5054 (N_5054,N_4788,N_4760);
nand U5055 (N_5055,N_4855,N_4863);
nor U5056 (N_5056,N_4997,N_4889);
nand U5057 (N_5057,N_4924,N_4852);
nor U5058 (N_5058,N_4754,N_4850);
nor U5059 (N_5059,N_4868,N_4756);
nor U5060 (N_5060,N_4914,N_4982);
or U5061 (N_5061,N_4890,N_4901);
and U5062 (N_5062,N_4824,N_4764);
and U5063 (N_5063,N_4768,N_4871);
or U5064 (N_5064,N_4766,N_4809);
nor U5065 (N_5065,N_4825,N_4938);
or U5066 (N_5066,N_4808,N_4907);
xor U5067 (N_5067,N_4805,N_4830);
xnor U5068 (N_5068,N_4918,N_4944);
and U5069 (N_5069,N_4770,N_4940);
nor U5070 (N_5070,N_4845,N_4785);
nor U5071 (N_5071,N_4987,N_4797);
or U5072 (N_5072,N_4904,N_4776);
nor U5073 (N_5073,N_4902,N_4877);
nand U5074 (N_5074,N_4819,N_4880);
xor U5075 (N_5075,N_4769,N_4912);
and U5076 (N_5076,N_4762,N_4841);
and U5077 (N_5077,N_4931,N_4998);
nand U5078 (N_5078,N_4953,N_4839);
xnor U5079 (N_5079,N_4900,N_4765);
xnor U5080 (N_5080,N_4884,N_4831);
nor U5081 (N_5081,N_4857,N_4946);
nand U5082 (N_5082,N_4876,N_4939);
or U5083 (N_5083,N_4995,N_4786);
xnor U5084 (N_5084,N_4791,N_4882);
and U5085 (N_5085,N_4949,N_4963);
or U5086 (N_5086,N_4947,N_4888);
xnor U5087 (N_5087,N_4838,N_4848);
or U5088 (N_5088,N_4881,N_4782);
and U5089 (N_5089,N_4821,N_4872);
xor U5090 (N_5090,N_4968,N_4778);
or U5091 (N_5091,N_4773,N_4961);
nor U5092 (N_5092,N_4813,N_4753);
nor U5093 (N_5093,N_4922,N_4973);
or U5094 (N_5094,N_4989,N_4887);
nor U5095 (N_5095,N_4777,N_4932);
xnor U5096 (N_5096,N_4921,N_4781);
and U5097 (N_5097,N_4792,N_4930);
and U5098 (N_5098,N_4843,N_4774);
xnor U5099 (N_5099,N_4763,N_4800);
or U5100 (N_5100,N_4923,N_4970);
xor U5101 (N_5101,N_4919,N_4853);
nand U5102 (N_5102,N_4864,N_4858);
and U5103 (N_5103,N_4960,N_4916);
or U5104 (N_5104,N_4952,N_4828);
nor U5105 (N_5105,N_4928,N_4945);
or U5106 (N_5106,N_4954,N_4990);
or U5107 (N_5107,N_4818,N_4861);
and U5108 (N_5108,N_4879,N_4789);
nand U5109 (N_5109,N_4832,N_4917);
nand U5110 (N_5110,N_4790,N_4758);
nor U5111 (N_5111,N_4964,N_4849);
or U5112 (N_5112,N_4994,N_4834);
nor U5113 (N_5113,N_4771,N_4859);
nand U5114 (N_5114,N_4870,N_4780);
nor U5115 (N_5115,N_4972,N_4833);
nor U5116 (N_5116,N_4911,N_4966);
xor U5117 (N_5117,N_4807,N_4798);
xnor U5118 (N_5118,N_4842,N_4812);
and U5119 (N_5119,N_4942,N_4929);
nor U5120 (N_5120,N_4783,N_4955);
xor U5121 (N_5121,N_4775,N_4996);
nor U5122 (N_5122,N_4815,N_4751);
nor U5123 (N_5123,N_4892,N_4935);
nand U5124 (N_5124,N_4971,N_4823);
nand U5125 (N_5125,N_4789,N_4755);
xor U5126 (N_5126,N_4947,N_4830);
and U5127 (N_5127,N_4981,N_4972);
xor U5128 (N_5128,N_4808,N_4968);
nor U5129 (N_5129,N_4890,N_4866);
xor U5130 (N_5130,N_4898,N_4768);
nand U5131 (N_5131,N_4913,N_4944);
and U5132 (N_5132,N_4853,N_4992);
xnor U5133 (N_5133,N_4826,N_4754);
nor U5134 (N_5134,N_4970,N_4878);
nor U5135 (N_5135,N_4792,N_4822);
nor U5136 (N_5136,N_4788,N_4903);
nor U5137 (N_5137,N_4880,N_4758);
xnor U5138 (N_5138,N_4911,N_4957);
nor U5139 (N_5139,N_4947,N_4768);
nor U5140 (N_5140,N_4950,N_4974);
or U5141 (N_5141,N_4916,N_4769);
or U5142 (N_5142,N_4753,N_4870);
or U5143 (N_5143,N_4869,N_4890);
xnor U5144 (N_5144,N_4784,N_4972);
or U5145 (N_5145,N_4971,N_4814);
nand U5146 (N_5146,N_4961,N_4866);
nand U5147 (N_5147,N_4998,N_4838);
or U5148 (N_5148,N_4892,N_4989);
xor U5149 (N_5149,N_4793,N_4951);
nor U5150 (N_5150,N_4794,N_4914);
nand U5151 (N_5151,N_4753,N_4911);
xor U5152 (N_5152,N_4797,N_4929);
nand U5153 (N_5153,N_4867,N_4857);
or U5154 (N_5154,N_4981,N_4865);
or U5155 (N_5155,N_4817,N_4934);
and U5156 (N_5156,N_4944,N_4805);
xnor U5157 (N_5157,N_4928,N_4806);
or U5158 (N_5158,N_4975,N_4869);
nand U5159 (N_5159,N_4838,N_4975);
and U5160 (N_5160,N_4880,N_4784);
nand U5161 (N_5161,N_4806,N_4906);
xor U5162 (N_5162,N_4899,N_4886);
nor U5163 (N_5163,N_4914,N_4770);
nand U5164 (N_5164,N_4764,N_4816);
nand U5165 (N_5165,N_4834,N_4783);
and U5166 (N_5166,N_4871,N_4904);
and U5167 (N_5167,N_4946,N_4922);
nand U5168 (N_5168,N_4828,N_4964);
and U5169 (N_5169,N_4754,N_4894);
nand U5170 (N_5170,N_4839,N_4815);
nor U5171 (N_5171,N_4952,N_4764);
nand U5172 (N_5172,N_4868,N_4971);
or U5173 (N_5173,N_4804,N_4813);
and U5174 (N_5174,N_4781,N_4946);
nor U5175 (N_5175,N_4977,N_4887);
or U5176 (N_5176,N_4870,N_4899);
xnor U5177 (N_5177,N_4777,N_4782);
xor U5178 (N_5178,N_4851,N_4858);
nor U5179 (N_5179,N_4953,N_4975);
nand U5180 (N_5180,N_4917,N_4856);
or U5181 (N_5181,N_4882,N_4840);
nor U5182 (N_5182,N_4934,N_4767);
xor U5183 (N_5183,N_4770,N_4811);
xnor U5184 (N_5184,N_4948,N_4929);
nand U5185 (N_5185,N_4797,N_4847);
nand U5186 (N_5186,N_4914,N_4845);
nor U5187 (N_5187,N_4931,N_4758);
nor U5188 (N_5188,N_4885,N_4772);
xnor U5189 (N_5189,N_4793,N_4913);
nand U5190 (N_5190,N_4770,N_4845);
and U5191 (N_5191,N_4903,N_4815);
and U5192 (N_5192,N_4816,N_4904);
or U5193 (N_5193,N_4795,N_4939);
or U5194 (N_5194,N_4924,N_4820);
nor U5195 (N_5195,N_4989,N_4770);
xor U5196 (N_5196,N_4838,N_4809);
nor U5197 (N_5197,N_4763,N_4993);
nand U5198 (N_5198,N_4800,N_4798);
and U5199 (N_5199,N_4830,N_4900);
nor U5200 (N_5200,N_4759,N_4816);
nand U5201 (N_5201,N_4853,N_4831);
or U5202 (N_5202,N_4994,N_4972);
nand U5203 (N_5203,N_4923,N_4925);
and U5204 (N_5204,N_4873,N_4770);
or U5205 (N_5205,N_4991,N_4895);
and U5206 (N_5206,N_4974,N_4924);
nor U5207 (N_5207,N_4823,N_4923);
and U5208 (N_5208,N_4995,N_4970);
or U5209 (N_5209,N_4797,N_4867);
and U5210 (N_5210,N_4875,N_4861);
nor U5211 (N_5211,N_4827,N_4980);
nand U5212 (N_5212,N_4781,N_4750);
or U5213 (N_5213,N_4987,N_4888);
nor U5214 (N_5214,N_4792,N_4760);
nor U5215 (N_5215,N_4787,N_4756);
or U5216 (N_5216,N_4788,N_4849);
nor U5217 (N_5217,N_4960,N_4971);
nor U5218 (N_5218,N_4765,N_4882);
xnor U5219 (N_5219,N_4762,N_4887);
nand U5220 (N_5220,N_4787,N_4874);
xnor U5221 (N_5221,N_4764,N_4957);
and U5222 (N_5222,N_4846,N_4957);
xor U5223 (N_5223,N_4816,N_4875);
nand U5224 (N_5224,N_4917,N_4958);
nand U5225 (N_5225,N_4763,N_4903);
xor U5226 (N_5226,N_4770,N_4789);
or U5227 (N_5227,N_4955,N_4863);
and U5228 (N_5228,N_4830,N_4873);
xor U5229 (N_5229,N_4778,N_4762);
and U5230 (N_5230,N_4763,N_4780);
nor U5231 (N_5231,N_4892,N_4802);
nor U5232 (N_5232,N_4840,N_4855);
or U5233 (N_5233,N_4854,N_4960);
xnor U5234 (N_5234,N_4939,N_4873);
or U5235 (N_5235,N_4973,N_4858);
nor U5236 (N_5236,N_4840,N_4998);
nand U5237 (N_5237,N_4803,N_4987);
xnor U5238 (N_5238,N_4993,N_4830);
nand U5239 (N_5239,N_4783,N_4885);
or U5240 (N_5240,N_4790,N_4907);
nand U5241 (N_5241,N_4965,N_4836);
nor U5242 (N_5242,N_4966,N_4756);
and U5243 (N_5243,N_4988,N_4944);
nor U5244 (N_5244,N_4949,N_4814);
xnor U5245 (N_5245,N_4920,N_4832);
or U5246 (N_5246,N_4856,N_4976);
or U5247 (N_5247,N_4849,N_4879);
or U5248 (N_5248,N_4912,N_4964);
and U5249 (N_5249,N_4858,N_4826);
or U5250 (N_5250,N_5214,N_5061);
nand U5251 (N_5251,N_5217,N_5154);
nand U5252 (N_5252,N_5241,N_5219);
nand U5253 (N_5253,N_5118,N_5147);
nor U5254 (N_5254,N_5062,N_5234);
xnor U5255 (N_5255,N_5198,N_5164);
or U5256 (N_5256,N_5189,N_5005);
and U5257 (N_5257,N_5203,N_5179);
or U5258 (N_5258,N_5215,N_5195);
or U5259 (N_5259,N_5029,N_5191);
nand U5260 (N_5260,N_5123,N_5160);
xor U5261 (N_5261,N_5020,N_5199);
or U5262 (N_5262,N_5175,N_5000);
or U5263 (N_5263,N_5222,N_5110);
nor U5264 (N_5264,N_5065,N_5078);
xor U5265 (N_5265,N_5059,N_5091);
xor U5266 (N_5266,N_5151,N_5157);
xnor U5267 (N_5267,N_5122,N_5224);
nand U5268 (N_5268,N_5206,N_5071);
nor U5269 (N_5269,N_5039,N_5133);
and U5270 (N_5270,N_5009,N_5054);
nand U5271 (N_5271,N_5193,N_5001);
or U5272 (N_5272,N_5004,N_5096);
and U5273 (N_5273,N_5050,N_5087);
nand U5274 (N_5274,N_5130,N_5233);
and U5275 (N_5275,N_5144,N_5044);
and U5276 (N_5276,N_5173,N_5053);
nor U5277 (N_5277,N_5247,N_5121);
or U5278 (N_5278,N_5126,N_5155);
nor U5279 (N_5279,N_5011,N_5064);
xnor U5280 (N_5280,N_5162,N_5094);
and U5281 (N_5281,N_5161,N_5131);
or U5282 (N_5282,N_5142,N_5235);
xor U5283 (N_5283,N_5066,N_5055);
and U5284 (N_5284,N_5143,N_5242);
xnor U5285 (N_5285,N_5098,N_5223);
and U5286 (N_5286,N_5231,N_5220);
and U5287 (N_5287,N_5041,N_5014);
nand U5288 (N_5288,N_5080,N_5112);
nor U5289 (N_5289,N_5145,N_5141);
and U5290 (N_5290,N_5106,N_5172);
nand U5291 (N_5291,N_5017,N_5188);
nor U5292 (N_5292,N_5230,N_5031);
and U5293 (N_5293,N_5019,N_5072);
nor U5294 (N_5294,N_5115,N_5006);
nor U5295 (N_5295,N_5148,N_5132);
nand U5296 (N_5296,N_5084,N_5114);
and U5297 (N_5297,N_5090,N_5119);
nor U5298 (N_5298,N_5025,N_5074);
nand U5299 (N_5299,N_5149,N_5137);
xnor U5300 (N_5300,N_5184,N_5170);
xor U5301 (N_5301,N_5192,N_5152);
nor U5302 (N_5302,N_5129,N_5018);
or U5303 (N_5303,N_5205,N_5245);
and U5304 (N_5304,N_5088,N_5165);
nor U5305 (N_5305,N_5047,N_5086);
nand U5306 (N_5306,N_5225,N_5239);
or U5307 (N_5307,N_5196,N_5043);
or U5308 (N_5308,N_5040,N_5183);
or U5309 (N_5309,N_5034,N_5153);
xor U5310 (N_5310,N_5128,N_5120);
or U5311 (N_5311,N_5216,N_5246);
nand U5312 (N_5312,N_5048,N_5167);
or U5313 (N_5313,N_5060,N_5063);
nand U5314 (N_5314,N_5238,N_5102);
xor U5315 (N_5315,N_5159,N_5049);
and U5316 (N_5316,N_5103,N_5135);
and U5317 (N_5317,N_5136,N_5227);
nor U5318 (N_5318,N_5036,N_5056);
nand U5319 (N_5319,N_5076,N_5028);
and U5320 (N_5320,N_5185,N_5013);
nand U5321 (N_5321,N_5107,N_5008);
and U5322 (N_5322,N_5075,N_5211);
and U5323 (N_5323,N_5010,N_5002);
nand U5324 (N_5324,N_5140,N_5201);
or U5325 (N_5325,N_5204,N_5139);
xnor U5326 (N_5326,N_5111,N_5081);
xnor U5327 (N_5327,N_5101,N_5244);
xor U5328 (N_5328,N_5038,N_5026);
and U5329 (N_5329,N_5213,N_5229);
or U5330 (N_5330,N_5124,N_5085);
and U5331 (N_5331,N_5146,N_5035);
and U5332 (N_5332,N_5032,N_5207);
and U5333 (N_5333,N_5202,N_5209);
nor U5334 (N_5334,N_5007,N_5127);
or U5335 (N_5335,N_5022,N_5237);
and U5336 (N_5336,N_5200,N_5095);
and U5337 (N_5337,N_5150,N_5092);
xnor U5338 (N_5338,N_5181,N_5099);
xor U5339 (N_5339,N_5194,N_5228);
and U5340 (N_5340,N_5109,N_5057);
nor U5341 (N_5341,N_5218,N_5174);
or U5342 (N_5342,N_5226,N_5024);
xor U5343 (N_5343,N_5180,N_5003);
nor U5344 (N_5344,N_5125,N_5030);
xnor U5345 (N_5345,N_5012,N_5212);
and U5346 (N_5346,N_5163,N_5077);
xor U5347 (N_5347,N_5116,N_5051);
xor U5348 (N_5348,N_5221,N_5079);
nor U5349 (N_5349,N_5037,N_5083);
and U5350 (N_5350,N_5182,N_5104);
or U5351 (N_5351,N_5243,N_5023);
xnor U5352 (N_5352,N_5176,N_5069);
xnor U5353 (N_5353,N_5187,N_5158);
nand U5354 (N_5354,N_5156,N_5236);
nand U5355 (N_5355,N_5046,N_5058);
nand U5356 (N_5356,N_5210,N_5138);
nor U5357 (N_5357,N_5240,N_5033);
nor U5358 (N_5358,N_5168,N_5186);
and U5359 (N_5359,N_5016,N_5100);
or U5360 (N_5360,N_5042,N_5070);
xnor U5361 (N_5361,N_5178,N_5052);
nor U5362 (N_5362,N_5232,N_5108);
and U5363 (N_5363,N_5249,N_5067);
xnor U5364 (N_5364,N_5097,N_5093);
xnor U5365 (N_5365,N_5248,N_5197);
nand U5366 (N_5366,N_5068,N_5190);
nor U5367 (N_5367,N_5027,N_5045);
nand U5368 (N_5368,N_5166,N_5169);
nor U5369 (N_5369,N_5171,N_5082);
and U5370 (N_5370,N_5208,N_5073);
and U5371 (N_5371,N_5021,N_5015);
nor U5372 (N_5372,N_5089,N_5134);
nand U5373 (N_5373,N_5117,N_5177);
nand U5374 (N_5374,N_5105,N_5113);
or U5375 (N_5375,N_5170,N_5210);
or U5376 (N_5376,N_5071,N_5086);
or U5377 (N_5377,N_5195,N_5122);
xor U5378 (N_5378,N_5169,N_5157);
and U5379 (N_5379,N_5099,N_5009);
nor U5380 (N_5380,N_5186,N_5067);
or U5381 (N_5381,N_5210,N_5073);
and U5382 (N_5382,N_5214,N_5166);
nand U5383 (N_5383,N_5234,N_5226);
nor U5384 (N_5384,N_5153,N_5128);
or U5385 (N_5385,N_5001,N_5118);
xor U5386 (N_5386,N_5155,N_5112);
and U5387 (N_5387,N_5006,N_5182);
xnor U5388 (N_5388,N_5107,N_5105);
xor U5389 (N_5389,N_5078,N_5230);
xor U5390 (N_5390,N_5009,N_5194);
nor U5391 (N_5391,N_5014,N_5155);
nor U5392 (N_5392,N_5009,N_5097);
xor U5393 (N_5393,N_5042,N_5093);
nor U5394 (N_5394,N_5056,N_5100);
nand U5395 (N_5395,N_5239,N_5230);
and U5396 (N_5396,N_5187,N_5194);
xnor U5397 (N_5397,N_5005,N_5239);
nor U5398 (N_5398,N_5176,N_5109);
or U5399 (N_5399,N_5163,N_5075);
or U5400 (N_5400,N_5239,N_5211);
nor U5401 (N_5401,N_5008,N_5116);
nor U5402 (N_5402,N_5246,N_5100);
xor U5403 (N_5403,N_5019,N_5023);
or U5404 (N_5404,N_5159,N_5077);
nand U5405 (N_5405,N_5239,N_5185);
nand U5406 (N_5406,N_5038,N_5191);
nand U5407 (N_5407,N_5005,N_5177);
nand U5408 (N_5408,N_5009,N_5146);
and U5409 (N_5409,N_5194,N_5248);
nor U5410 (N_5410,N_5136,N_5089);
and U5411 (N_5411,N_5193,N_5093);
and U5412 (N_5412,N_5042,N_5139);
or U5413 (N_5413,N_5200,N_5008);
nand U5414 (N_5414,N_5060,N_5020);
xor U5415 (N_5415,N_5066,N_5187);
or U5416 (N_5416,N_5175,N_5227);
nor U5417 (N_5417,N_5052,N_5011);
nor U5418 (N_5418,N_5191,N_5248);
nor U5419 (N_5419,N_5052,N_5015);
xnor U5420 (N_5420,N_5051,N_5162);
nand U5421 (N_5421,N_5092,N_5207);
or U5422 (N_5422,N_5208,N_5099);
xor U5423 (N_5423,N_5017,N_5101);
xnor U5424 (N_5424,N_5228,N_5233);
nor U5425 (N_5425,N_5037,N_5000);
nor U5426 (N_5426,N_5170,N_5000);
nor U5427 (N_5427,N_5161,N_5232);
nand U5428 (N_5428,N_5173,N_5221);
xnor U5429 (N_5429,N_5020,N_5198);
nand U5430 (N_5430,N_5121,N_5067);
and U5431 (N_5431,N_5092,N_5101);
nand U5432 (N_5432,N_5051,N_5001);
nand U5433 (N_5433,N_5008,N_5167);
nor U5434 (N_5434,N_5168,N_5093);
nor U5435 (N_5435,N_5029,N_5213);
nand U5436 (N_5436,N_5184,N_5154);
or U5437 (N_5437,N_5097,N_5249);
and U5438 (N_5438,N_5044,N_5156);
or U5439 (N_5439,N_5157,N_5038);
nor U5440 (N_5440,N_5228,N_5225);
xor U5441 (N_5441,N_5113,N_5156);
nor U5442 (N_5442,N_5184,N_5139);
xor U5443 (N_5443,N_5036,N_5197);
xor U5444 (N_5444,N_5045,N_5064);
or U5445 (N_5445,N_5143,N_5218);
nand U5446 (N_5446,N_5213,N_5010);
and U5447 (N_5447,N_5086,N_5187);
nand U5448 (N_5448,N_5116,N_5075);
nor U5449 (N_5449,N_5128,N_5103);
nor U5450 (N_5450,N_5042,N_5095);
and U5451 (N_5451,N_5031,N_5144);
xnor U5452 (N_5452,N_5096,N_5201);
or U5453 (N_5453,N_5117,N_5124);
nand U5454 (N_5454,N_5171,N_5053);
or U5455 (N_5455,N_5204,N_5183);
nand U5456 (N_5456,N_5194,N_5161);
nor U5457 (N_5457,N_5149,N_5197);
nand U5458 (N_5458,N_5028,N_5110);
nor U5459 (N_5459,N_5002,N_5060);
or U5460 (N_5460,N_5064,N_5208);
nand U5461 (N_5461,N_5238,N_5245);
xnor U5462 (N_5462,N_5108,N_5118);
and U5463 (N_5463,N_5019,N_5084);
nand U5464 (N_5464,N_5019,N_5229);
nor U5465 (N_5465,N_5249,N_5087);
or U5466 (N_5466,N_5216,N_5056);
or U5467 (N_5467,N_5068,N_5011);
nor U5468 (N_5468,N_5101,N_5069);
nand U5469 (N_5469,N_5111,N_5242);
or U5470 (N_5470,N_5115,N_5065);
nor U5471 (N_5471,N_5106,N_5206);
and U5472 (N_5472,N_5014,N_5114);
and U5473 (N_5473,N_5104,N_5064);
or U5474 (N_5474,N_5077,N_5046);
xor U5475 (N_5475,N_5084,N_5186);
or U5476 (N_5476,N_5170,N_5187);
or U5477 (N_5477,N_5054,N_5187);
or U5478 (N_5478,N_5142,N_5211);
nor U5479 (N_5479,N_5043,N_5183);
and U5480 (N_5480,N_5233,N_5080);
nand U5481 (N_5481,N_5002,N_5139);
nand U5482 (N_5482,N_5196,N_5201);
or U5483 (N_5483,N_5201,N_5073);
xor U5484 (N_5484,N_5000,N_5110);
and U5485 (N_5485,N_5119,N_5117);
or U5486 (N_5486,N_5242,N_5229);
or U5487 (N_5487,N_5169,N_5041);
nand U5488 (N_5488,N_5011,N_5026);
and U5489 (N_5489,N_5188,N_5057);
or U5490 (N_5490,N_5011,N_5047);
or U5491 (N_5491,N_5246,N_5170);
and U5492 (N_5492,N_5133,N_5196);
xor U5493 (N_5493,N_5010,N_5099);
nand U5494 (N_5494,N_5081,N_5035);
nand U5495 (N_5495,N_5122,N_5055);
xnor U5496 (N_5496,N_5162,N_5015);
nand U5497 (N_5497,N_5139,N_5009);
nand U5498 (N_5498,N_5039,N_5057);
and U5499 (N_5499,N_5115,N_5013);
or U5500 (N_5500,N_5255,N_5492);
nor U5501 (N_5501,N_5461,N_5374);
or U5502 (N_5502,N_5455,N_5252);
nor U5503 (N_5503,N_5346,N_5298);
or U5504 (N_5504,N_5266,N_5413);
and U5505 (N_5505,N_5475,N_5474);
or U5506 (N_5506,N_5478,N_5420);
xor U5507 (N_5507,N_5408,N_5250);
and U5508 (N_5508,N_5378,N_5306);
nand U5509 (N_5509,N_5385,N_5407);
and U5510 (N_5510,N_5270,N_5359);
nand U5511 (N_5511,N_5389,N_5457);
nand U5512 (N_5512,N_5263,N_5327);
xnor U5513 (N_5513,N_5358,N_5326);
or U5514 (N_5514,N_5421,N_5318);
nor U5515 (N_5515,N_5332,N_5394);
nand U5516 (N_5516,N_5280,N_5459);
or U5517 (N_5517,N_5290,N_5456);
nor U5518 (N_5518,N_5291,N_5440);
or U5519 (N_5519,N_5341,N_5350);
xnor U5520 (N_5520,N_5432,N_5330);
nand U5521 (N_5521,N_5364,N_5393);
or U5522 (N_5522,N_5452,N_5495);
or U5523 (N_5523,N_5286,N_5314);
and U5524 (N_5524,N_5347,N_5409);
nand U5525 (N_5525,N_5377,N_5472);
and U5526 (N_5526,N_5372,N_5426);
and U5527 (N_5527,N_5483,N_5337);
or U5528 (N_5528,N_5484,N_5397);
nand U5529 (N_5529,N_5391,N_5296);
nand U5530 (N_5530,N_5438,N_5311);
nand U5531 (N_5531,N_5422,N_5256);
nor U5532 (N_5532,N_5329,N_5417);
nor U5533 (N_5533,N_5373,N_5390);
xnor U5534 (N_5534,N_5260,N_5328);
and U5535 (N_5535,N_5331,N_5261);
or U5536 (N_5536,N_5376,N_5448);
and U5537 (N_5537,N_5424,N_5464);
nor U5538 (N_5538,N_5349,N_5313);
nor U5539 (N_5539,N_5499,N_5405);
and U5540 (N_5540,N_5361,N_5398);
and U5541 (N_5541,N_5251,N_5253);
or U5542 (N_5542,N_5435,N_5354);
nand U5543 (N_5543,N_5356,N_5302);
nor U5544 (N_5544,N_5319,N_5275);
and U5545 (N_5545,N_5324,N_5315);
and U5546 (N_5546,N_5375,N_5282);
and U5547 (N_5547,N_5363,N_5272);
nor U5548 (N_5548,N_5352,N_5418);
nor U5549 (N_5549,N_5355,N_5439);
nor U5550 (N_5550,N_5279,N_5254);
nor U5551 (N_5551,N_5369,N_5437);
nand U5552 (N_5552,N_5292,N_5485);
xor U5553 (N_5553,N_5382,N_5338);
nor U5554 (N_5554,N_5415,N_5258);
and U5555 (N_5555,N_5316,N_5379);
nor U5556 (N_5556,N_5479,N_5477);
and U5557 (N_5557,N_5486,N_5274);
nand U5558 (N_5558,N_5339,N_5257);
xnor U5559 (N_5559,N_5396,N_5293);
or U5560 (N_5560,N_5433,N_5404);
or U5561 (N_5561,N_5366,N_5493);
nand U5562 (N_5562,N_5269,N_5265);
nand U5563 (N_5563,N_5446,N_5262);
or U5564 (N_5564,N_5383,N_5368);
and U5565 (N_5565,N_5277,N_5476);
and U5566 (N_5566,N_5289,N_5410);
xor U5567 (N_5567,N_5287,N_5310);
or U5568 (N_5568,N_5288,N_5268);
and U5569 (N_5569,N_5336,N_5321);
or U5570 (N_5570,N_5348,N_5304);
and U5571 (N_5571,N_5462,N_5412);
nand U5572 (N_5572,N_5294,N_5299);
and U5573 (N_5573,N_5480,N_5362);
xor U5574 (N_5574,N_5365,N_5283);
and U5575 (N_5575,N_5490,N_5482);
or U5576 (N_5576,N_5301,N_5465);
or U5577 (N_5577,N_5453,N_5449);
nor U5578 (N_5578,N_5307,N_5323);
xor U5579 (N_5579,N_5463,N_5343);
nor U5580 (N_5580,N_5458,N_5491);
and U5581 (N_5581,N_5371,N_5384);
and U5582 (N_5582,N_5345,N_5344);
xor U5583 (N_5583,N_5488,N_5427);
and U5584 (N_5584,N_5494,N_5357);
nand U5585 (N_5585,N_5429,N_5317);
or U5586 (N_5586,N_5447,N_5498);
and U5587 (N_5587,N_5395,N_5325);
nor U5588 (N_5588,N_5406,N_5454);
or U5589 (N_5589,N_5419,N_5387);
and U5590 (N_5590,N_5481,N_5468);
nand U5591 (N_5591,N_5308,N_5416);
xnor U5592 (N_5592,N_5443,N_5467);
or U5593 (N_5593,N_5436,N_5403);
nand U5594 (N_5594,N_5450,N_5473);
nand U5595 (N_5595,N_5466,N_5333);
xnor U5596 (N_5596,N_5281,N_5425);
and U5597 (N_5597,N_5400,N_5312);
and U5598 (N_5598,N_5381,N_5303);
nand U5599 (N_5599,N_5411,N_5444);
nand U5600 (N_5600,N_5305,N_5285);
nor U5601 (N_5601,N_5273,N_5367);
or U5602 (N_5602,N_5267,N_5423);
and U5603 (N_5603,N_5445,N_5297);
nand U5604 (N_5604,N_5271,N_5386);
nor U5605 (N_5605,N_5442,N_5434);
and U5606 (N_5606,N_5370,N_5489);
or U5607 (N_5607,N_5497,N_5470);
xnor U5608 (N_5608,N_5496,N_5431);
nand U5609 (N_5609,N_5320,N_5351);
xor U5610 (N_5610,N_5264,N_5401);
xnor U5611 (N_5611,N_5334,N_5399);
nor U5612 (N_5612,N_5295,N_5460);
and U5613 (N_5613,N_5380,N_5388);
or U5614 (N_5614,N_5278,N_5441);
or U5615 (N_5615,N_5469,N_5284);
and U5616 (N_5616,N_5402,N_5342);
or U5617 (N_5617,N_5300,N_5309);
xnor U5618 (N_5618,N_5471,N_5353);
or U5619 (N_5619,N_5360,N_5487);
and U5620 (N_5620,N_5335,N_5451);
and U5621 (N_5621,N_5430,N_5392);
nor U5622 (N_5622,N_5276,N_5414);
nor U5623 (N_5623,N_5428,N_5259);
xor U5624 (N_5624,N_5340,N_5322);
and U5625 (N_5625,N_5262,N_5344);
xor U5626 (N_5626,N_5429,N_5435);
nor U5627 (N_5627,N_5452,N_5349);
xor U5628 (N_5628,N_5256,N_5427);
nor U5629 (N_5629,N_5347,N_5486);
xnor U5630 (N_5630,N_5389,N_5298);
or U5631 (N_5631,N_5352,N_5435);
and U5632 (N_5632,N_5395,N_5354);
or U5633 (N_5633,N_5370,N_5377);
xnor U5634 (N_5634,N_5468,N_5440);
xor U5635 (N_5635,N_5420,N_5431);
xor U5636 (N_5636,N_5499,N_5264);
xor U5637 (N_5637,N_5308,N_5425);
and U5638 (N_5638,N_5390,N_5426);
or U5639 (N_5639,N_5428,N_5368);
and U5640 (N_5640,N_5493,N_5401);
nor U5641 (N_5641,N_5280,N_5336);
xnor U5642 (N_5642,N_5264,N_5388);
nor U5643 (N_5643,N_5389,N_5260);
nand U5644 (N_5644,N_5483,N_5276);
or U5645 (N_5645,N_5272,N_5325);
or U5646 (N_5646,N_5433,N_5441);
nand U5647 (N_5647,N_5335,N_5284);
xnor U5648 (N_5648,N_5339,N_5313);
or U5649 (N_5649,N_5359,N_5457);
or U5650 (N_5650,N_5360,N_5298);
and U5651 (N_5651,N_5400,N_5453);
xnor U5652 (N_5652,N_5317,N_5342);
xor U5653 (N_5653,N_5274,N_5469);
nor U5654 (N_5654,N_5471,N_5463);
nand U5655 (N_5655,N_5304,N_5340);
and U5656 (N_5656,N_5374,N_5445);
nor U5657 (N_5657,N_5398,N_5408);
and U5658 (N_5658,N_5285,N_5272);
nor U5659 (N_5659,N_5264,N_5458);
nand U5660 (N_5660,N_5398,N_5268);
nor U5661 (N_5661,N_5312,N_5335);
nor U5662 (N_5662,N_5389,N_5422);
or U5663 (N_5663,N_5317,N_5259);
or U5664 (N_5664,N_5335,N_5383);
nand U5665 (N_5665,N_5496,N_5493);
xnor U5666 (N_5666,N_5283,N_5285);
nor U5667 (N_5667,N_5321,N_5460);
xnor U5668 (N_5668,N_5343,N_5459);
or U5669 (N_5669,N_5387,N_5471);
and U5670 (N_5670,N_5462,N_5398);
xor U5671 (N_5671,N_5390,N_5499);
and U5672 (N_5672,N_5259,N_5401);
and U5673 (N_5673,N_5428,N_5299);
nand U5674 (N_5674,N_5406,N_5479);
and U5675 (N_5675,N_5433,N_5333);
xnor U5676 (N_5676,N_5392,N_5407);
and U5677 (N_5677,N_5440,N_5483);
or U5678 (N_5678,N_5400,N_5484);
and U5679 (N_5679,N_5451,N_5341);
or U5680 (N_5680,N_5495,N_5277);
xnor U5681 (N_5681,N_5440,N_5340);
nand U5682 (N_5682,N_5274,N_5320);
or U5683 (N_5683,N_5404,N_5415);
nand U5684 (N_5684,N_5329,N_5286);
and U5685 (N_5685,N_5263,N_5314);
xor U5686 (N_5686,N_5462,N_5456);
nor U5687 (N_5687,N_5415,N_5390);
nand U5688 (N_5688,N_5424,N_5374);
xnor U5689 (N_5689,N_5281,N_5426);
nor U5690 (N_5690,N_5469,N_5278);
or U5691 (N_5691,N_5481,N_5310);
and U5692 (N_5692,N_5284,N_5347);
or U5693 (N_5693,N_5343,N_5424);
and U5694 (N_5694,N_5343,N_5347);
or U5695 (N_5695,N_5421,N_5348);
or U5696 (N_5696,N_5469,N_5481);
nand U5697 (N_5697,N_5414,N_5480);
and U5698 (N_5698,N_5301,N_5345);
or U5699 (N_5699,N_5334,N_5341);
nand U5700 (N_5700,N_5400,N_5344);
nor U5701 (N_5701,N_5349,N_5437);
xor U5702 (N_5702,N_5303,N_5334);
nor U5703 (N_5703,N_5250,N_5331);
nor U5704 (N_5704,N_5416,N_5306);
xor U5705 (N_5705,N_5435,N_5455);
nand U5706 (N_5706,N_5296,N_5428);
nor U5707 (N_5707,N_5259,N_5338);
nand U5708 (N_5708,N_5447,N_5448);
and U5709 (N_5709,N_5309,N_5432);
nand U5710 (N_5710,N_5430,N_5489);
or U5711 (N_5711,N_5494,N_5349);
or U5712 (N_5712,N_5384,N_5313);
nand U5713 (N_5713,N_5287,N_5368);
or U5714 (N_5714,N_5451,N_5426);
and U5715 (N_5715,N_5424,N_5382);
and U5716 (N_5716,N_5435,N_5437);
xor U5717 (N_5717,N_5299,N_5253);
nor U5718 (N_5718,N_5259,N_5290);
or U5719 (N_5719,N_5382,N_5393);
nand U5720 (N_5720,N_5264,N_5323);
or U5721 (N_5721,N_5282,N_5318);
nor U5722 (N_5722,N_5379,N_5401);
nor U5723 (N_5723,N_5313,N_5411);
xnor U5724 (N_5724,N_5267,N_5319);
and U5725 (N_5725,N_5267,N_5337);
or U5726 (N_5726,N_5461,N_5480);
nor U5727 (N_5727,N_5350,N_5254);
or U5728 (N_5728,N_5423,N_5410);
or U5729 (N_5729,N_5311,N_5365);
or U5730 (N_5730,N_5278,N_5323);
and U5731 (N_5731,N_5377,N_5492);
and U5732 (N_5732,N_5337,N_5378);
and U5733 (N_5733,N_5280,N_5307);
or U5734 (N_5734,N_5330,N_5373);
nor U5735 (N_5735,N_5293,N_5349);
and U5736 (N_5736,N_5382,N_5345);
nand U5737 (N_5737,N_5323,N_5324);
or U5738 (N_5738,N_5444,N_5319);
xnor U5739 (N_5739,N_5474,N_5345);
and U5740 (N_5740,N_5380,N_5295);
and U5741 (N_5741,N_5397,N_5319);
xor U5742 (N_5742,N_5339,N_5496);
nand U5743 (N_5743,N_5462,N_5409);
and U5744 (N_5744,N_5414,N_5259);
nand U5745 (N_5745,N_5267,N_5482);
xnor U5746 (N_5746,N_5362,N_5460);
nor U5747 (N_5747,N_5471,N_5355);
nor U5748 (N_5748,N_5290,N_5276);
nor U5749 (N_5749,N_5302,N_5461);
nor U5750 (N_5750,N_5591,N_5544);
nor U5751 (N_5751,N_5546,N_5727);
and U5752 (N_5752,N_5539,N_5534);
and U5753 (N_5753,N_5631,N_5717);
nor U5754 (N_5754,N_5592,N_5731);
xnor U5755 (N_5755,N_5506,N_5582);
xnor U5756 (N_5756,N_5668,N_5739);
or U5757 (N_5757,N_5703,N_5681);
xnor U5758 (N_5758,N_5562,N_5527);
or U5759 (N_5759,N_5699,N_5677);
and U5760 (N_5760,N_5533,N_5589);
nor U5761 (N_5761,N_5580,N_5667);
xnor U5762 (N_5762,N_5720,N_5537);
nand U5763 (N_5763,N_5623,N_5569);
nor U5764 (N_5764,N_5637,N_5556);
and U5765 (N_5765,N_5672,N_5605);
or U5766 (N_5766,N_5726,N_5545);
xnor U5767 (N_5767,N_5614,N_5653);
nand U5768 (N_5768,N_5721,N_5564);
and U5769 (N_5769,N_5612,N_5593);
or U5770 (N_5770,N_5509,N_5704);
nand U5771 (N_5771,N_5708,N_5738);
xor U5772 (N_5772,N_5629,N_5741);
or U5773 (N_5773,N_5647,N_5692);
xnor U5774 (N_5774,N_5554,N_5662);
nor U5775 (N_5775,N_5526,N_5743);
nor U5776 (N_5776,N_5665,N_5548);
and U5777 (N_5777,N_5635,N_5638);
xnor U5778 (N_5778,N_5748,N_5684);
nand U5779 (N_5779,N_5568,N_5552);
nand U5780 (N_5780,N_5573,N_5728);
nand U5781 (N_5781,N_5734,N_5510);
or U5782 (N_5782,N_5599,N_5620);
xor U5783 (N_5783,N_5567,N_5598);
nor U5784 (N_5784,N_5633,N_5735);
xor U5785 (N_5785,N_5651,N_5695);
nor U5786 (N_5786,N_5641,N_5710);
or U5787 (N_5787,N_5659,N_5516);
and U5788 (N_5788,N_5724,N_5602);
and U5789 (N_5789,N_5634,N_5682);
nand U5790 (N_5790,N_5557,N_5640);
nand U5791 (N_5791,N_5660,N_5687);
nand U5792 (N_5792,N_5521,N_5585);
and U5793 (N_5793,N_5555,N_5590);
or U5794 (N_5794,N_5697,N_5518);
nand U5795 (N_5795,N_5504,N_5693);
or U5796 (N_5796,N_5581,N_5654);
nor U5797 (N_5797,N_5563,N_5577);
and U5798 (N_5798,N_5719,N_5532);
xnor U5799 (N_5799,N_5642,N_5649);
xnor U5800 (N_5800,N_5500,N_5702);
and U5801 (N_5801,N_5630,N_5528);
nor U5802 (N_5802,N_5571,N_5747);
and U5803 (N_5803,N_5689,N_5503);
and U5804 (N_5804,N_5514,N_5566);
nor U5805 (N_5805,N_5676,N_5597);
xnor U5806 (N_5806,N_5587,N_5715);
or U5807 (N_5807,N_5522,N_5547);
and U5808 (N_5808,N_5520,N_5565);
nand U5809 (N_5809,N_5744,N_5669);
xor U5810 (N_5810,N_5683,N_5502);
xor U5811 (N_5811,N_5586,N_5524);
nor U5812 (N_5812,N_5658,N_5746);
and U5813 (N_5813,N_5621,N_5732);
and U5814 (N_5814,N_5505,N_5679);
xnor U5815 (N_5815,N_5745,N_5517);
nand U5816 (N_5816,N_5722,N_5671);
and U5817 (N_5817,N_5696,N_5561);
nand U5818 (N_5818,N_5616,N_5711);
xor U5819 (N_5819,N_5604,N_5627);
or U5820 (N_5820,N_5558,N_5579);
xor U5821 (N_5821,N_5601,N_5622);
or U5822 (N_5822,N_5639,N_5523);
and U5823 (N_5823,N_5570,N_5511);
nand U5824 (N_5824,N_5663,N_5729);
and U5825 (N_5825,N_5636,N_5650);
and U5826 (N_5826,N_5553,N_5512);
or U5827 (N_5827,N_5560,N_5559);
and U5828 (N_5828,N_5619,N_5628);
and U5829 (N_5829,N_5594,N_5576);
nand U5830 (N_5830,N_5714,N_5698);
nor U5831 (N_5831,N_5740,N_5705);
nor U5832 (N_5832,N_5678,N_5575);
and U5833 (N_5833,N_5644,N_5685);
nor U5834 (N_5834,N_5691,N_5736);
nand U5835 (N_5835,N_5615,N_5723);
and U5836 (N_5836,N_5656,N_5513);
and U5837 (N_5837,N_5648,N_5595);
nor U5838 (N_5838,N_5655,N_5536);
or U5839 (N_5839,N_5608,N_5670);
nor U5840 (N_5840,N_5657,N_5501);
and U5841 (N_5841,N_5673,N_5632);
nor U5842 (N_5842,N_5700,N_5543);
nor U5843 (N_5843,N_5611,N_5733);
or U5844 (N_5844,N_5645,N_5730);
nand U5845 (N_5845,N_5609,N_5690);
xor U5846 (N_5846,N_5701,N_5515);
xor U5847 (N_5847,N_5674,N_5713);
and U5848 (N_5848,N_5574,N_5742);
and U5849 (N_5849,N_5709,N_5718);
or U5850 (N_5850,N_5507,N_5531);
or U5851 (N_5851,N_5578,N_5618);
nor U5852 (N_5852,N_5652,N_5661);
and U5853 (N_5853,N_5706,N_5588);
xnor U5854 (N_5854,N_5749,N_5646);
xnor U5855 (N_5855,N_5529,N_5626);
or U5856 (N_5856,N_5600,N_5716);
and U5857 (N_5857,N_5538,N_5643);
and U5858 (N_5858,N_5550,N_5613);
nor U5859 (N_5859,N_5680,N_5624);
nand U5860 (N_5860,N_5519,N_5596);
xnor U5861 (N_5861,N_5617,N_5712);
nand U5862 (N_5862,N_5551,N_5686);
and U5863 (N_5863,N_5666,N_5549);
and U5864 (N_5864,N_5572,N_5535);
nor U5865 (N_5865,N_5664,N_5737);
and U5866 (N_5866,N_5606,N_5694);
nor U5867 (N_5867,N_5607,N_5610);
nand U5868 (N_5868,N_5525,N_5725);
or U5869 (N_5869,N_5541,N_5583);
xor U5870 (N_5870,N_5542,N_5688);
nor U5871 (N_5871,N_5625,N_5707);
xor U5872 (N_5872,N_5540,N_5603);
or U5873 (N_5873,N_5584,N_5508);
nand U5874 (N_5874,N_5675,N_5530);
nor U5875 (N_5875,N_5709,N_5595);
nand U5876 (N_5876,N_5624,N_5732);
xnor U5877 (N_5877,N_5626,N_5715);
nand U5878 (N_5878,N_5732,N_5693);
nor U5879 (N_5879,N_5701,N_5608);
and U5880 (N_5880,N_5702,N_5596);
and U5881 (N_5881,N_5574,N_5746);
xor U5882 (N_5882,N_5594,N_5727);
and U5883 (N_5883,N_5749,N_5548);
nand U5884 (N_5884,N_5549,N_5522);
nor U5885 (N_5885,N_5638,N_5688);
or U5886 (N_5886,N_5581,N_5727);
and U5887 (N_5887,N_5559,N_5558);
nand U5888 (N_5888,N_5732,N_5728);
or U5889 (N_5889,N_5648,N_5511);
or U5890 (N_5890,N_5571,N_5727);
nor U5891 (N_5891,N_5582,N_5500);
or U5892 (N_5892,N_5656,N_5660);
nor U5893 (N_5893,N_5506,N_5711);
xor U5894 (N_5894,N_5745,N_5654);
nor U5895 (N_5895,N_5691,N_5557);
and U5896 (N_5896,N_5647,N_5563);
or U5897 (N_5897,N_5690,N_5603);
nand U5898 (N_5898,N_5729,N_5575);
nor U5899 (N_5899,N_5676,N_5543);
or U5900 (N_5900,N_5537,N_5663);
nand U5901 (N_5901,N_5712,N_5626);
nor U5902 (N_5902,N_5664,N_5683);
xnor U5903 (N_5903,N_5649,N_5584);
nor U5904 (N_5904,N_5651,N_5648);
xor U5905 (N_5905,N_5697,N_5551);
nor U5906 (N_5906,N_5744,N_5593);
nor U5907 (N_5907,N_5614,N_5700);
and U5908 (N_5908,N_5720,N_5513);
and U5909 (N_5909,N_5545,N_5617);
xor U5910 (N_5910,N_5658,N_5555);
nor U5911 (N_5911,N_5610,N_5586);
nor U5912 (N_5912,N_5675,N_5685);
xor U5913 (N_5913,N_5660,N_5585);
nor U5914 (N_5914,N_5730,N_5692);
and U5915 (N_5915,N_5717,N_5636);
or U5916 (N_5916,N_5681,N_5633);
nor U5917 (N_5917,N_5724,N_5650);
or U5918 (N_5918,N_5727,N_5654);
xnor U5919 (N_5919,N_5516,N_5546);
and U5920 (N_5920,N_5559,N_5648);
nor U5921 (N_5921,N_5555,N_5672);
nor U5922 (N_5922,N_5693,N_5735);
xor U5923 (N_5923,N_5548,N_5645);
nor U5924 (N_5924,N_5645,N_5652);
xnor U5925 (N_5925,N_5519,N_5738);
nor U5926 (N_5926,N_5603,N_5677);
xor U5927 (N_5927,N_5513,N_5516);
or U5928 (N_5928,N_5693,N_5551);
nand U5929 (N_5929,N_5519,N_5610);
or U5930 (N_5930,N_5621,N_5565);
nand U5931 (N_5931,N_5590,N_5601);
nor U5932 (N_5932,N_5644,N_5532);
or U5933 (N_5933,N_5648,N_5731);
nor U5934 (N_5934,N_5698,N_5521);
and U5935 (N_5935,N_5686,N_5734);
or U5936 (N_5936,N_5567,N_5656);
or U5937 (N_5937,N_5591,N_5628);
xnor U5938 (N_5938,N_5611,N_5651);
or U5939 (N_5939,N_5672,N_5603);
or U5940 (N_5940,N_5543,N_5501);
xor U5941 (N_5941,N_5593,N_5549);
or U5942 (N_5942,N_5576,N_5681);
or U5943 (N_5943,N_5644,N_5546);
nor U5944 (N_5944,N_5585,N_5559);
nor U5945 (N_5945,N_5513,N_5735);
or U5946 (N_5946,N_5688,N_5609);
xnor U5947 (N_5947,N_5507,N_5720);
or U5948 (N_5948,N_5554,N_5732);
xnor U5949 (N_5949,N_5725,N_5625);
nor U5950 (N_5950,N_5638,N_5576);
nor U5951 (N_5951,N_5747,N_5575);
nor U5952 (N_5952,N_5528,N_5571);
or U5953 (N_5953,N_5721,N_5714);
xor U5954 (N_5954,N_5741,N_5665);
xor U5955 (N_5955,N_5673,N_5564);
and U5956 (N_5956,N_5592,N_5715);
nand U5957 (N_5957,N_5592,N_5603);
nand U5958 (N_5958,N_5695,N_5714);
and U5959 (N_5959,N_5723,N_5730);
or U5960 (N_5960,N_5745,N_5630);
and U5961 (N_5961,N_5593,N_5721);
nor U5962 (N_5962,N_5584,N_5515);
xor U5963 (N_5963,N_5521,N_5523);
and U5964 (N_5964,N_5604,N_5580);
nor U5965 (N_5965,N_5584,N_5619);
or U5966 (N_5966,N_5653,N_5595);
or U5967 (N_5967,N_5692,N_5720);
nand U5968 (N_5968,N_5561,N_5679);
nor U5969 (N_5969,N_5530,N_5507);
xnor U5970 (N_5970,N_5565,N_5612);
xnor U5971 (N_5971,N_5526,N_5532);
nand U5972 (N_5972,N_5747,N_5691);
nor U5973 (N_5973,N_5695,N_5600);
or U5974 (N_5974,N_5735,N_5658);
and U5975 (N_5975,N_5705,N_5587);
and U5976 (N_5976,N_5511,N_5608);
or U5977 (N_5977,N_5541,N_5537);
and U5978 (N_5978,N_5544,N_5733);
xor U5979 (N_5979,N_5742,N_5613);
nand U5980 (N_5980,N_5722,N_5515);
nor U5981 (N_5981,N_5640,N_5675);
or U5982 (N_5982,N_5563,N_5678);
xor U5983 (N_5983,N_5659,N_5699);
nor U5984 (N_5984,N_5532,N_5663);
or U5985 (N_5985,N_5633,N_5609);
nand U5986 (N_5986,N_5509,N_5524);
nand U5987 (N_5987,N_5508,N_5677);
and U5988 (N_5988,N_5740,N_5695);
and U5989 (N_5989,N_5556,N_5544);
nand U5990 (N_5990,N_5563,N_5576);
or U5991 (N_5991,N_5671,N_5653);
nand U5992 (N_5992,N_5656,N_5538);
xnor U5993 (N_5993,N_5530,N_5520);
and U5994 (N_5994,N_5599,N_5586);
xor U5995 (N_5995,N_5518,N_5696);
and U5996 (N_5996,N_5609,N_5628);
and U5997 (N_5997,N_5514,N_5666);
nor U5998 (N_5998,N_5643,N_5559);
xnor U5999 (N_5999,N_5507,N_5641);
or U6000 (N_6000,N_5797,N_5922);
or U6001 (N_6001,N_5760,N_5875);
nor U6002 (N_6002,N_5755,N_5946);
or U6003 (N_6003,N_5910,N_5756);
xor U6004 (N_6004,N_5983,N_5856);
nand U6005 (N_6005,N_5976,N_5991);
xor U6006 (N_6006,N_5994,N_5768);
and U6007 (N_6007,N_5827,N_5980);
and U6008 (N_6008,N_5885,N_5759);
and U6009 (N_6009,N_5934,N_5761);
nor U6010 (N_6010,N_5883,N_5811);
and U6011 (N_6011,N_5825,N_5804);
nand U6012 (N_6012,N_5935,N_5771);
nand U6013 (N_6013,N_5920,N_5834);
nand U6014 (N_6014,N_5995,N_5766);
nor U6015 (N_6015,N_5943,N_5785);
xnor U6016 (N_6016,N_5780,N_5906);
nor U6017 (N_6017,N_5950,N_5996);
xor U6018 (N_6018,N_5919,N_5973);
xnor U6019 (N_6019,N_5762,N_5803);
xnor U6020 (N_6020,N_5902,N_5765);
xnor U6021 (N_6021,N_5982,N_5763);
xnor U6022 (N_6022,N_5789,N_5817);
and U6023 (N_6023,N_5928,N_5860);
and U6024 (N_6024,N_5904,N_5849);
nor U6025 (N_6025,N_5862,N_5940);
and U6026 (N_6026,N_5964,N_5819);
and U6027 (N_6027,N_5897,N_5957);
nor U6028 (N_6028,N_5911,N_5882);
xnor U6029 (N_6029,N_5975,N_5857);
xnor U6030 (N_6030,N_5848,N_5843);
nand U6031 (N_6031,N_5779,N_5784);
and U6032 (N_6032,N_5824,N_5839);
nand U6033 (N_6033,N_5853,N_5774);
and U6034 (N_6034,N_5974,N_5826);
or U6035 (N_6035,N_5778,N_5847);
nor U6036 (N_6036,N_5786,N_5787);
xnor U6037 (N_6037,N_5988,N_5870);
nand U6038 (N_6038,N_5970,N_5969);
or U6039 (N_6039,N_5753,N_5927);
nand U6040 (N_6040,N_5990,N_5966);
and U6041 (N_6041,N_5893,N_5767);
and U6042 (N_6042,N_5796,N_5872);
xnor U6043 (N_6043,N_5793,N_5801);
and U6044 (N_6044,N_5931,N_5782);
nor U6045 (N_6045,N_5813,N_5963);
nor U6046 (N_6046,N_5790,N_5757);
xnor U6047 (N_6047,N_5799,N_5947);
nor U6048 (N_6048,N_5908,N_5865);
nor U6049 (N_6049,N_5907,N_5816);
nor U6050 (N_6050,N_5806,N_5751);
xnor U6051 (N_6051,N_5833,N_5924);
nor U6052 (N_6052,N_5769,N_5840);
or U6053 (N_6053,N_5829,N_5820);
and U6054 (N_6054,N_5845,N_5913);
or U6055 (N_6055,N_5754,N_5890);
and U6056 (N_6056,N_5818,N_5773);
or U6057 (N_6057,N_5854,N_5989);
nand U6058 (N_6058,N_5841,N_5798);
nor U6059 (N_6059,N_5901,N_5836);
or U6060 (N_6060,N_5936,N_5823);
and U6061 (N_6061,N_5933,N_5955);
or U6062 (N_6062,N_5838,N_5909);
nand U6063 (N_6063,N_5832,N_5859);
xor U6064 (N_6064,N_5891,N_5858);
nand U6065 (N_6065,N_5929,N_5821);
nor U6066 (N_6066,N_5772,N_5867);
or U6067 (N_6067,N_5894,N_5886);
xor U6068 (N_6068,N_5861,N_5900);
xor U6069 (N_6069,N_5977,N_5878);
xor U6070 (N_6070,N_5948,N_5792);
nor U6071 (N_6071,N_5831,N_5959);
and U6072 (N_6072,N_5998,N_5997);
xor U6073 (N_6073,N_5846,N_5815);
nor U6074 (N_6074,N_5889,N_5944);
nand U6075 (N_6075,N_5863,N_5981);
xnor U6076 (N_6076,N_5992,N_5932);
xnor U6077 (N_6077,N_5949,N_5962);
nor U6078 (N_6078,N_5956,N_5937);
and U6079 (N_6079,N_5809,N_5835);
nor U6080 (N_6080,N_5979,N_5921);
or U6081 (N_6081,N_5898,N_5884);
or U6082 (N_6082,N_5930,N_5952);
and U6083 (N_6083,N_5783,N_5942);
or U6084 (N_6084,N_5776,N_5800);
nor U6085 (N_6085,N_5939,N_5864);
nor U6086 (N_6086,N_5781,N_5877);
or U6087 (N_6087,N_5874,N_5805);
xnor U6088 (N_6088,N_5968,N_5895);
nand U6089 (N_6089,N_5986,N_5752);
nor U6090 (N_6090,N_5802,N_5868);
xor U6091 (N_6091,N_5915,N_5999);
nand U6092 (N_6092,N_5916,N_5866);
xnor U6093 (N_6093,N_5794,N_5855);
nor U6094 (N_6094,N_5770,N_5830);
nor U6095 (N_6095,N_5961,N_5795);
xor U6096 (N_6096,N_5828,N_5958);
or U6097 (N_6097,N_5871,N_5810);
and U6098 (N_6098,N_5852,N_5844);
nand U6099 (N_6099,N_5941,N_5750);
or U6100 (N_6100,N_5873,N_5788);
nor U6101 (N_6101,N_5881,N_5960);
xor U6102 (N_6102,N_5791,N_5869);
or U6103 (N_6103,N_5965,N_5967);
nand U6104 (N_6104,N_5987,N_5837);
nor U6105 (N_6105,N_5917,N_5775);
nor U6106 (N_6106,N_5945,N_5896);
or U6107 (N_6107,N_5842,N_5876);
and U6108 (N_6108,N_5912,N_5880);
nand U6109 (N_6109,N_5985,N_5925);
and U6110 (N_6110,N_5814,N_5777);
nand U6111 (N_6111,N_5905,N_5807);
and U6112 (N_6112,N_5808,N_5954);
xnor U6113 (N_6113,N_5822,N_5892);
nor U6114 (N_6114,N_5758,N_5914);
and U6115 (N_6115,N_5978,N_5971);
nor U6116 (N_6116,N_5951,N_5888);
nand U6117 (N_6117,N_5764,N_5879);
xnor U6118 (N_6118,N_5993,N_5918);
nand U6119 (N_6119,N_5812,N_5850);
nor U6120 (N_6120,N_5903,N_5972);
nand U6121 (N_6121,N_5926,N_5899);
xnor U6122 (N_6122,N_5938,N_5887);
nor U6123 (N_6123,N_5851,N_5953);
xnor U6124 (N_6124,N_5923,N_5984);
xnor U6125 (N_6125,N_5963,N_5894);
xnor U6126 (N_6126,N_5755,N_5773);
nand U6127 (N_6127,N_5997,N_5782);
or U6128 (N_6128,N_5918,N_5750);
xnor U6129 (N_6129,N_5754,N_5990);
nand U6130 (N_6130,N_5893,N_5848);
nand U6131 (N_6131,N_5766,N_5945);
xor U6132 (N_6132,N_5984,N_5910);
nor U6133 (N_6133,N_5949,N_5819);
and U6134 (N_6134,N_5837,N_5819);
and U6135 (N_6135,N_5916,N_5827);
and U6136 (N_6136,N_5836,N_5770);
nand U6137 (N_6137,N_5833,N_5776);
and U6138 (N_6138,N_5872,N_5928);
nand U6139 (N_6139,N_5976,N_5826);
or U6140 (N_6140,N_5907,N_5848);
nand U6141 (N_6141,N_5775,N_5874);
and U6142 (N_6142,N_5913,N_5768);
nor U6143 (N_6143,N_5831,N_5980);
and U6144 (N_6144,N_5898,N_5752);
xnor U6145 (N_6145,N_5804,N_5820);
or U6146 (N_6146,N_5758,N_5848);
and U6147 (N_6147,N_5987,N_5767);
and U6148 (N_6148,N_5954,N_5834);
nand U6149 (N_6149,N_5770,N_5845);
xnor U6150 (N_6150,N_5814,N_5979);
xnor U6151 (N_6151,N_5948,N_5795);
xnor U6152 (N_6152,N_5877,N_5997);
nand U6153 (N_6153,N_5925,N_5891);
and U6154 (N_6154,N_5817,N_5930);
or U6155 (N_6155,N_5759,N_5954);
or U6156 (N_6156,N_5867,N_5892);
nor U6157 (N_6157,N_5839,N_5914);
and U6158 (N_6158,N_5840,N_5854);
and U6159 (N_6159,N_5971,N_5772);
or U6160 (N_6160,N_5758,N_5802);
nor U6161 (N_6161,N_5801,N_5991);
nand U6162 (N_6162,N_5817,N_5763);
and U6163 (N_6163,N_5865,N_5757);
or U6164 (N_6164,N_5949,N_5927);
and U6165 (N_6165,N_5750,N_5991);
and U6166 (N_6166,N_5973,N_5860);
or U6167 (N_6167,N_5884,N_5752);
xor U6168 (N_6168,N_5995,N_5815);
nor U6169 (N_6169,N_5932,N_5753);
nand U6170 (N_6170,N_5966,N_5960);
nor U6171 (N_6171,N_5786,N_5831);
or U6172 (N_6172,N_5925,N_5913);
xnor U6173 (N_6173,N_5905,N_5980);
nor U6174 (N_6174,N_5945,N_5847);
xor U6175 (N_6175,N_5844,N_5993);
and U6176 (N_6176,N_5915,N_5821);
xnor U6177 (N_6177,N_5773,N_5943);
and U6178 (N_6178,N_5768,N_5857);
and U6179 (N_6179,N_5903,N_5766);
nor U6180 (N_6180,N_5810,N_5814);
nor U6181 (N_6181,N_5782,N_5816);
xnor U6182 (N_6182,N_5895,N_5928);
nand U6183 (N_6183,N_5750,N_5776);
nor U6184 (N_6184,N_5948,N_5796);
nor U6185 (N_6185,N_5993,N_5851);
nand U6186 (N_6186,N_5850,N_5942);
or U6187 (N_6187,N_5967,N_5854);
nor U6188 (N_6188,N_5897,N_5951);
nor U6189 (N_6189,N_5939,N_5787);
or U6190 (N_6190,N_5790,N_5777);
and U6191 (N_6191,N_5908,N_5786);
and U6192 (N_6192,N_5860,N_5811);
xnor U6193 (N_6193,N_5857,N_5887);
or U6194 (N_6194,N_5938,N_5967);
or U6195 (N_6195,N_5818,N_5783);
nand U6196 (N_6196,N_5826,N_5803);
or U6197 (N_6197,N_5881,N_5941);
xnor U6198 (N_6198,N_5795,N_5857);
or U6199 (N_6199,N_5766,N_5862);
nor U6200 (N_6200,N_5888,N_5885);
nand U6201 (N_6201,N_5939,N_5812);
nand U6202 (N_6202,N_5868,N_5949);
nand U6203 (N_6203,N_5901,N_5830);
and U6204 (N_6204,N_5958,N_5971);
and U6205 (N_6205,N_5932,N_5822);
nor U6206 (N_6206,N_5966,N_5840);
nor U6207 (N_6207,N_5922,N_5981);
nor U6208 (N_6208,N_5908,N_5811);
nand U6209 (N_6209,N_5765,N_5769);
xnor U6210 (N_6210,N_5932,N_5808);
xnor U6211 (N_6211,N_5867,N_5938);
xor U6212 (N_6212,N_5815,N_5764);
and U6213 (N_6213,N_5776,N_5895);
xor U6214 (N_6214,N_5816,N_5850);
xnor U6215 (N_6215,N_5900,N_5795);
xnor U6216 (N_6216,N_5962,N_5977);
nand U6217 (N_6217,N_5814,N_5825);
nor U6218 (N_6218,N_5848,N_5791);
nor U6219 (N_6219,N_5845,N_5946);
nor U6220 (N_6220,N_5946,N_5829);
nor U6221 (N_6221,N_5819,N_5786);
or U6222 (N_6222,N_5845,N_5932);
nor U6223 (N_6223,N_5995,N_5921);
nor U6224 (N_6224,N_5776,N_5945);
nand U6225 (N_6225,N_5831,N_5930);
and U6226 (N_6226,N_5951,N_5882);
xor U6227 (N_6227,N_5957,N_5890);
nand U6228 (N_6228,N_5754,N_5908);
or U6229 (N_6229,N_5979,N_5942);
and U6230 (N_6230,N_5805,N_5981);
and U6231 (N_6231,N_5960,N_5855);
or U6232 (N_6232,N_5959,N_5780);
xor U6233 (N_6233,N_5818,N_5811);
or U6234 (N_6234,N_5922,N_5931);
nand U6235 (N_6235,N_5896,N_5768);
or U6236 (N_6236,N_5949,N_5899);
nor U6237 (N_6237,N_5825,N_5873);
or U6238 (N_6238,N_5998,N_5890);
and U6239 (N_6239,N_5803,N_5867);
or U6240 (N_6240,N_5908,N_5977);
xnor U6241 (N_6241,N_5863,N_5919);
xnor U6242 (N_6242,N_5985,N_5780);
nand U6243 (N_6243,N_5971,N_5954);
xnor U6244 (N_6244,N_5937,N_5935);
xor U6245 (N_6245,N_5936,N_5859);
or U6246 (N_6246,N_5914,N_5818);
xor U6247 (N_6247,N_5977,N_5987);
xnor U6248 (N_6248,N_5943,N_5827);
nor U6249 (N_6249,N_5947,N_5963);
nand U6250 (N_6250,N_6124,N_6010);
nor U6251 (N_6251,N_6141,N_6059);
xnor U6252 (N_6252,N_6173,N_6171);
nand U6253 (N_6253,N_6092,N_6053);
and U6254 (N_6254,N_6148,N_6196);
or U6255 (N_6255,N_6075,N_6052);
or U6256 (N_6256,N_6071,N_6137);
or U6257 (N_6257,N_6076,N_6208);
and U6258 (N_6258,N_6100,N_6147);
or U6259 (N_6259,N_6027,N_6248);
xnor U6260 (N_6260,N_6226,N_6180);
nor U6261 (N_6261,N_6082,N_6049);
xnor U6262 (N_6262,N_6058,N_6087);
and U6263 (N_6263,N_6077,N_6078);
nand U6264 (N_6264,N_6031,N_6228);
nand U6265 (N_6265,N_6002,N_6184);
nor U6266 (N_6266,N_6190,N_6215);
nor U6267 (N_6267,N_6094,N_6070);
and U6268 (N_6268,N_6174,N_6073);
xnor U6269 (N_6269,N_6111,N_6225);
nand U6270 (N_6270,N_6041,N_6212);
xor U6271 (N_6271,N_6001,N_6000);
xor U6272 (N_6272,N_6139,N_6121);
nor U6273 (N_6273,N_6216,N_6181);
nor U6274 (N_6274,N_6193,N_6242);
xor U6275 (N_6275,N_6102,N_6224);
nand U6276 (N_6276,N_6074,N_6104);
xnor U6277 (N_6277,N_6129,N_6038);
xor U6278 (N_6278,N_6083,N_6126);
or U6279 (N_6279,N_6179,N_6182);
nand U6280 (N_6280,N_6195,N_6048);
or U6281 (N_6281,N_6192,N_6172);
nor U6282 (N_6282,N_6061,N_6239);
and U6283 (N_6283,N_6188,N_6134);
nand U6284 (N_6284,N_6037,N_6057);
nor U6285 (N_6285,N_6085,N_6163);
xnor U6286 (N_6286,N_6206,N_6130);
nor U6287 (N_6287,N_6161,N_6185);
or U6288 (N_6288,N_6003,N_6122);
nand U6289 (N_6289,N_6213,N_6211);
nand U6290 (N_6290,N_6245,N_6160);
or U6291 (N_6291,N_6066,N_6136);
nor U6292 (N_6292,N_6116,N_6011);
xnor U6293 (N_6293,N_6125,N_6247);
or U6294 (N_6294,N_6145,N_6246);
xor U6295 (N_6295,N_6197,N_6089);
and U6296 (N_6296,N_6205,N_6149);
nor U6297 (N_6297,N_6103,N_6217);
and U6298 (N_6298,N_6112,N_6007);
or U6299 (N_6299,N_6093,N_6158);
nor U6300 (N_6300,N_6146,N_6118);
nand U6301 (N_6301,N_6209,N_6015);
nand U6302 (N_6302,N_6095,N_6183);
and U6303 (N_6303,N_6028,N_6025);
nand U6304 (N_6304,N_6120,N_6156);
or U6305 (N_6305,N_6065,N_6203);
nand U6306 (N_6306,N_6099,N_6243);
nand U6307 (N_6307,N_6133,N_6198);
or U6308 (N_6308,N_6119,N_6056);
and U6309 (N_6309,N_6016,N_6244);
and U6310 (N_6310,N_6021,N_6020);
nand U6311 (N_6311,N_6067,N_6050);
and U6312 (N_6312,N_6151,N_6108);
nand U6313 (N_6313,N_6159,N_6237);
nor U6314 (N_6314,N_6032,N_6034);
nor U6315 (N_6315,N_6040,N_6046);
nand U6316 (N_6316,N_6227,N_6200);
and U6317 (N_6317,N_6017,N_6138);
xor U6318 (N_6318,N_6096,N_6101);
nor U6319 (N_6319,N_6229,N_6154);
and U6320 (N_6320,N_6230,N_6091);
nor U6321 (N_6321,N_6202,N_6231);
or U6322 (N_6322,N_6191,N_6098);
nand U6323 (N_6323,N_6047,N_6249);
xnor U6324 (N_6324,N_6238,N_6113);
nand U6325 (N_6325,N_6039,N_6033);
and U6326 (N_6326,N_6081,N_6187);
or U6327 (N_6327,N_6170,N_6150);
nor U6328 (N_6328,N_6201,N_6029);
and U6329 (N_6329,N_6064,N_6063);
nor U6330 (N_6330,N_6169,N_6090);
xnor U6331 (N_6331,N_6107,N_6194);
or U6332 (N_6332,N_6117,N_6152);
or U6333 (N_6333,N_6175,N_6055);
or U6334 (N_6334,N_6210,N_6036);
nand U6335 (N_6335,N_6026,N_6164);
xor U6336 (N_6336,N_6043,N_6080);
xnor U6337 (N_6337,N_6013,N_6018);
nor U6338 (N_6338,N_6223,N_6123);
and U6339 (N_6339,N_6218,N_6135);
xnor U6340 (N_6340,N_6084,N_6004);
nand U6341 (N_6341,N_6186,N_6177);
nand U6342 (N_6342,N_6005,N_6166);
and U6343 (N_6343,N_6221,N_6051);
and U6344 (N_6344,N_6023,N_6044);
nor U6345 (N_6345,N_6233,N_6054);
and U6346 (N_6346,N_6199,N_6240);
or U6347 (N_6347,N_6178,N_6035);
nand U6348 (N_6348,N_6167,N_6222);
xnor U6349 (N_6349,N_6006,N_6128);
nand U6350 (N_6350,N_6144,N_6072);
and U6351 (N_6351,N_6069,N_6131);
and U6352 (N_6352,N_6068,N_6109);
nand U6353 (N_6353,N_6012,N_6132);
or U6354 (N_6354,N_6142,N_6008);
xnor U6355 (N_6355,N_6204,N_6042);
or U6356 (N_6356,N_6079,N_6060);
nand U6357 (N_6357,N_6014,N_6106);
or U6358 (N_6358,N_6153,N_6127);
xnor U6359 (N_6359,N_6140,N_6143);
nor U6360 (N_6360,N_6241,N_6162);
nand U6361 (N_6361,N_6234,N_6207);
and U6362 (N_6362,N_6176,N_6214);
nor U6363 (N_6363,N_6155,N_6097);
xor U6364 (N_6364,N_6024,N_6105);
nand U6365 (N_6365,N_6009,N_6086);
xnor U6366 (N_6366,N_6115,N_6165);
xnor U6367 (N_6367,N_6110,N_6045);
or U6368 (N_6368,N_6114,N_6022);
nor U6369 (N_6369,N_6062,N_6235);
and U6370 (N_6370,N_6232,N_6189);
or U6371 (N_6371,N_6236,N_6220);
nor U6372 (N_6372,N_6157,N_6168);
xnor U6373 (N_6373,N_6219,N_6088);
and U6374 (N_6374,N_6030,N_6019);
xnor U6375 (N_6375,N_6147,N_6041);
nand U6376 (N_6376,N_6122,N_6063);
nor U6377 (N_6377,N_6095,N_6157);
or U6378 (N_6378,N_6200,N_6191);
nand U6379 (N_6379,N_6121,N_6031);
nor U6380 (N_6380,N_6149,N_6036);
and U6381 (N_6381,N_6175,N_6095);
xor U6382 (N_6382,N_6049,N_6084);
xor U6383 (N_6383,N_6021,N_6214);
nand U6384 (N_6384,N_6151,N_6127);
nor U6385 (N_6385,N_6007,N_6236);
and U6386 (N_6386,N_6097,N_6175);
xor U6387 (N_6387,N_6216,N_6131);
or U6388 (N_6388,N_6209,N_6244);
and U6389 (N_6389,N_6115,N_6111);
nand U6390 (N_6390,N_6228,N_6191);
xor U6391 (N_6391,N_6174,N_6065);
and U6392 (N_6392,N_6237,N_6043);
or U6393 (N_6393,N_6238,N_6024);
or U6394 (N_6394,N_6005,N_6207);
xnor U6395 (N_6395,N_6037,N_6226);
and U6396 (N_6396,N_6104,N_6167);
nand U6397 (N_6397,N_6052,N_6078);
nor U6398 (N_6398,N_6026,N_6153);
xnor U6399 (N_6399,N_6011,N_6244);
xor U6400 (N_6400,N_6201,N_6154);
and U6401 (N_6401,N_6118,N_6066);
and U6402 (N_6402,N_6216,N_6162);
or U6403 (N_6403,N_6078,N_6200);
nor U6404 (N_6404,N_6059,N_6190);
or U6405 (N_6405,N_6165,N_6122);
nor U6406 (N_6406,N_6033,N_6120);
nor U6407 (N_6407,N_6049,N_6237);
xor U6408 (N_6408,N_6105,N_6084);
nor U6409 (N_6409,N_6038,N_6240);
xnor U6410 (N_6410,N_6167,N_6143);
and U6411 (N_6411,N_6187,N_6150);
or U6412 (N_6412,N_6162,N_6101);
and U6413 (N_6413,N_6043,N_6087);
nand U6414 (N_6414,N_6196,N_6035);
and U6415 (N_6415,N_6068,N_6039);
xor U6416 (N_6416,N_6204,N_6039);
xnor U6417 (N_6417,N_6229,N_6145);
or U6418 (N_6418,N_6185,N_6194);
xor U6419 (N_6419,N_6219,N_6065);
nor U6420 (N_6420,N_6013,N_6149);
or U6421 (N_6421,N_6145,N_6159);
or U6422 (N_6422,N_6065,N_6141);
nor U6423 (N_6423,N_6097,N_6164);
nand U6424 (N_6424,N_6118,N_6051);
xnor U6425 (N_6425,N_6189,N_6142);
xor U6426 (N_6426,N_6087,N_6030);
nand U6427 (N_6427,N_6066,N_6194);
xnor U6428 (N_6428,N_6003,N_6070);
or U6429 (N_6429,N_6228,N_6016);
nor U6430 (N_6430,N_6046,N_6053);
nand U6431 (N_6431,N_6099,N_6022);
nand U6432 (N_6432,N_6176,N_6178);
and U6433 (N_6433,N_6161,N_6141);
or U6434 (N_6434,N_6059,N_6026);
or U6435 (N_6435,N_6153,N_6193);
or U6436 (N_6436,N_6223,N_6099);
and U6437 (N_6437,N_6224,N_6163);
or U6438 (N_6438,N_6153,N_6246);
or U6439 (N_6439,N_6137,N_6098);
nand U6440 (N_6440,N_6241,N_6244);
and U6441 (N_6441,N_6064,N_6176);
and U6442 (N_6442,N_6229,N_6227);
and U6443 (N_6443,N_6152,N_6171);
nor U6444 (N_6444,N_6156,N_6218);
and U6445 (N_6445,N_6134,N_6198);
xor U6446 (N_6446,N_6181,N_6004);
and U6447 (N_6447,N_6009,N_6184);
or U6448 (N_6448,N_6209,N_6012);
and U6449 (N_6449,N_6219,N_6033);
nand U6450 (N_6450,N_6197,N_6056);
and U6451 (N_6451,N_6095,N_6073);
xor U6452 (N_6452,N_6137,N_6187);
xor U6453 (N_6453,N_6009,N_6249);
nand U6454 (N_6454,N_6113,N_6183);
nor U6455 (N_6455,N_6160,N_6053);
nand U6456 (N_6456,N_6200,N_6010);
and U6457 (N_6457,N_6192,N_6068);
xnor U6458 (N_6458,N_6243,N_6053);
nand U6459 (N_6459,N_6025,N_6152);
nand U6460 (N_6460,N_6239,N_6044);
xnor U6461 (N_6461,N_6046,N_6027);
and U6462 (N_6462,N_6142,N_6249);
nor U6463 (N_6463,N_6196,N_6063);
nor U6464 (N_6464,N_6012,N_6065);
nand U6465 (N_6465,N_6144,N_6065);
nand U6466 (N_6466,N_6046,N_6247);
and U6467 (N_6467,N_6120,N_6129);
nor U6468 (N_6468,N_6083,N_6060);
and U6469 (N_6469,N_6166,N_6027);
nand U6470 (N_6470,N_6019,N_6144);
or U6471 (N_6471,N_6159,N_6028);
xnor U6472 (N_6472,N_6166,N_6173);
or U6473 (N_6473,N_6153,N_6219);
nand U6474 (N_6474,N_6205,N_6008);
nor U6475 (N_6475,N_6024,N_6183);
nor U6476 (N_6476,N_6036,N_6131);
and U6477 (N_6477,N_6238,N_6180);
nand U6478 (N_6478,N_6135,N_6219);
and U6479 (N_6479,N_6063,N_6229);
or U6480 (N_6480,N_6149,N_6240);
or U6481 (N_6481,N_6033,N_6036);
or U6482 (N_6482,N_6187,N_6057);
or U6483 (N_6483,N_6014,N_6072);
nor U6484 (N_6484,N_6213,N_6180);
nor U6485 (N_6485,N_6067,N_6227);
xnor U6486 (N_6486,N_6208,N_6007);
and U6487 (N_6487,N_6183,N_6101);
or U6488 (N_6488,N_6055,N_6213);
and U6489 (N_6489,N_6105,N_6026);
xor U6490 (N_6490,N_6120,N_6110);
xor U6491 (N_6491,N_6069,N_6006);
nor U6492 (N_6492,N_6044,N_6175);
or U6493 (N_6493,N_6241,N_6075);
and U6494 (N_6494,N_6035,N_6242);
xor U6495 (N_6495,N_6160,N_6158);
or U6496 (N_6496,N_6075,N_6015);
and U6497 (N_6497,N_6179,N_6116);
xor U6498 (N_6498,N_6081,N_6198);
and U6499 (N_6499,N_6071,N_6124);
nor U6500 (N_6500,N_6477,N_6298);
and U6501 (N_6501,N_6423,N_6401);
nand U6502 (N_6502,N_6262,N_6466);
xnor U6503 (N_6503,N_6250,N_6337);
nor U6504 (N_6504,N_6411,N_6448);
or U6505 (N_6505,N_6436,N_6288);
nand U6506 (N_6506,N_6270,N_6278);
and U6507 (N_6507,N_6344,N_6398);
xor U6508 (N_6508,N_6264,N_6340);
or U6509 (N_6509,N_6263,N_6357);
nand U6510 (N_6510,N_6486,N_6474);
xnor U6511 (N_6511,N_6495,N_6472);
or U6512 (N_6512,N_6476,N_6451);
xor U6513 (N_6513,N_6343,N_6353);
and U6514 (N_6514,N_6299,N_6428);
xor U6515 (N_6515,N_6279,N_6351);
and U6516 (N_6516,N_6433,N_6471);
nor U6517 (N_6517,N_6404,N_6373);
nor U6518 (N_6518,N_6386,N_6393);
and U6519 (N_6519,N_6267,N_6341);
nand U6520 (N_6520,N_6331,N_6256);
nand U6521 (N_6521,N_6350,N_6284);
or U6522 (N_6522,N_6335,N_6292);
nor U6523 (N_6523,N_6385,N_6300);
nor U6524 (N_6524,N_6437,N_6326);
nor U6525 (N_6525,N_6376,N_6355);
nand U6526 (N_6526,N_6384,N_6443);
or U6527 (N_6527,N_6266,N_6372);
and U6528 (N_6528,N_6321,N_6460);
or U6529 (N_6529,N_6441,N_6402);
nor U6530 (N_6530,N_6457,N_6309);
and U6531 (N_6531,N_6452,N_6367);
or U6532 (N_6532,N_6491,N_6287);
or U6533 (N_6533,N_6275,N_6489);
nand U6534 (N_6534,N_6318,N_6362);
nand U6535 (N_6535,N_6308,N_6317);
or U6536 (N_6536,N_6358,N_6368);
nor U6537 (N_6537,N_6462,N_6281);
xnor U6538 (N_6538,N_6446,N_6383);
or U6539 (N_6539,N_6498,N_6432);
or U6540 (N_6540,N_6253,N_6359);
and U6541 (N_6541,N_6255,N_6315);
nor U6542 (N_6542,N_6382,N_6492);
xnor U6543 (N_6543,N_6449,N_6403);
xnor U6544 (N_6544,N_6306,N_6416);
and U6545 (N_6545,N_6470,N_6328);
or U6546 (N_6546,N_6282,N_6319);
nor U6547 (N_6547,N_6469,N_6394);
and U6548 (N_6548,N_6320,N_6271);
and U6549 (N_6549,N_6378,N_6377);
nor U6550 (N_6550,N_6496,N_6289);
nand U6551 (N_6551,N_6396,N_6369);
nor U6552 (N_6552,N_6258,N_6295);
or U6553 (N_6553,N_6338,N_6464);
xor U6554 (N_6554,N_6493,N_6487);
and U6555 (N_6555,N_6490,N_6483);
or U6556 (N_6556,N_6479,N_6458);
xor U6557 (N_6557,N_6388,N_6347);
and U6558 (N_6558,N_6283,N_6430);
nand U6559 (N_6559,N_6294,N_6391);
or U6560 (N_6560,N_6374,N_6467);
nor U6561 (N_6561,N_6334,N_6375);
and U6562 (N_6562,N_6395,N_6349);
xor U6563 (N_6563,N_6332,N_6265);
xor U6564 (N_6564,N_6456,N_6342);
and U6565 (N_6565,N_6463,N_6442);
nor U6566 (N_6566,N_6307,N_6371);
and U6567 (N_6567,N_6336,N_6325);
nor U6568 (N_6568,N_6468,N_6354);
or U6569 (N_6569,N_6484,N_6329);
and U6570 (N_6570,N_6459,N_6274);
and U6571 (N_6571,N_6435,N_6389);
or U6572 (N_6572,N_6346,N_6421);
and U6573 (N_6573,N_6333,N_6409);
nand U6574 (N_6574,N_6313,N_6494);
nor U6575 (N_6575,N_6444,N_6420);
nand U6576 (N_6576,N_6426,N_6414);
nor U6577 (N_6577,N_6445,N_6364);
xnor U6578 (N_6578,N_6361,N_6392);
or U6579 (N_6579,N_6497,N_6390);
or U6580 (N_6580,N_6381,N_6400);
or U6581 (N_6581,N_6480,N_6418);
nor U6582 (N_6582,N_6296,N_6254);
nor U6583 (N_6583,N_6410,N_6252);
nor U6584 (N_6584,N_6434,N_6251);
nand U6585 (N_6585,N_6380,N_6293);
and U6586 (N_6586,N_6356,N_6297);
or U6587 (N_6587,N_6304,N_6379);
or U6588 (N_6588,N_6269,N_6482);
nand U6589 (N_6589,N_6429,N_6323);
nor U6590 (N_6590,N_6310,N_6327);
nand U6591 (N_6591,N_6365,N_6285);
and U6592 (N_6592,N_6415,N_6303);
or U6593 (N_6593,N_6465,N_6424);
or U6594 (N_6594,N_6290,N_6478);
nand U6595 (N_6595,N_6425,N_6454);
or U6596 (N_6596,N_6360,N_6268);
nor U6597 (N_6597,N_6461,N_6276);
nor U6598 (N_6598,N_6431,N_6387);
and U6599 (N_6599,N_6286,N_6273);
nand U6600 (N_6600,N_6450,N_6257);
xor U6601 (N_6601,N_6427,N_6440);
and U6602 (N_6602,N_6301,N_6422);
xnor U6603 (N_6603,N_6322,N_6408);
nor U6604 (N_6604,N_6302,N_6419);
nand U6605 (N_6605,N_6339,N_6314);
nor U6606 (N_6606,N_6370,N_6447);
xor U6607 (N_6607,N_6399,N_6311);
nand U6608 (N_6608,N_6324,N_6330);
nor U6609 (N_6609,N_6352,N_6407);
xor U6610 (N_6610,N_6488,N_6439);
nand U6611 (N_6611,N_6499,N_6312);
and U6612 (N_6612,N_6397,N_6305);
or U6613 (N_6613,N_6277,N_6366);
nand U6614 (N_6614,N_6261,N_6272);
or U6615 (N_6615,N_6363,N_6453);
nor U6616 (N_6616,N_6455,N_6316);
nand U6617 (N_6617,N_6438,N_6406);
or U6618 (N_6618,N_6473,N_6345);
nand U6619 (N_6619,N_6291,N_6481);
and U6620 (N_6620,N_6348,N_6485);
nand U6621 (N_6621,N_6412,N_6259);
or U6622 (N_6622,N_6280,N_6417);
nand U6623 (N_6623,N_6475,N_6405);
or U6624 (N_6624,N_6260,N_6413);
and U6625 (N_6625,N_6351,N_6256);
nand U6626 (N_6626,N_6329,N_6494);
xnor U6627 (N_6627,N_6301,N_6313);
or U6628 (N_6628,N_6305,N_6266);
or U6629 (N_6629,N_6425,N_6346);
or U6630 (N_6630,N_6361,N_6401);
nand U6631 (N_6631,N_6258,N_6484);
nand U6632 (N_6632,N_6450,N_6492);
and U6633 (N_6633,N_6257,N_6334);
xnor U6634 (N_6634,N_6440,N_6434);
nor U6635 (N_6635,N_6266,N_6298);
nor U6636 (N_6636,N_6291,N_6313);
xor U6637 (N_6637,N_6472,N_6367);
xnor U6638 (N_6638,N_6443,N_6474);
nor U6639 (N_6639,N_6385,N_6491);
and U6640 (N_6640,N_6448,N_6488);
nand U6641 (N_6641,N_6469,N_6417);
and U6642 (N_6642,N_6469,N_6377);
nor U6643 (N_6643,N_6424,N_6293);
nand U6644 (N_6644,N_6291,N_6441);
and U6645 (N_6645,N_6372,N_6486);
xnor U6646 (N_6646,N_6305,N_6454);
xor U6647 (N_6647,N_6434,N_6497);
nor U6648 (N_6648,N_6371,N_6398);
nor U6649 (N_6649,N_6499,N_6390);
or U6650 (N_6650,N_6367,N_6454);
nor U6651 (N_6651,N_6486,N_6281);
or U6652 (N_6652,N_6335,N_6355);
xor U6653 (N_6653,N_6370,N_6349);
or U6654 (N_6654,N_6295,N_6293);
or U6655 (N_6655,N_6496,N_6321);
nor U6656 (N_6656,N_6457,N_6429);
or U6657 (N_6657,N_6316,N_6456);
xor U6658 (N_6658,N_6282,N_6450);
nand U6659 (N_6659,N_6433,N_6320);
nand U6660 (N_6660,N_6422,N_6415);
and U6661 (N_6661,N_6306,N_6390);
or U6662 (N_6662,N_6354,N_6297);
or U6663 (N_6663,N_6422,N_6443);
xnor U6664 (N_6664,N_6352,N_6323);
and U6665 (N_6665,N_6396,N_6255);
and U6666 (N_6666,N_6280,N_6366);
and U6667 (N_6667,N_6336,N_6252);
nor U6668 (N_6668,N_6344,N_6336);
xnor U6669 (N_6669,N_6335,N_6312);
or U6670 (N_6670,N_6264,N_6324);
xor U6671 (N_6671,N_6353,N_6254);
nor U6672 (N_6672,N_6410,N_6388);
or U6673 (N_6673,N_6428,N_6414);
xor U6674 (N_6674,N_6382,N_6301);
xnor U6675 (N_6675,N_6254,N_6334);
xnor U6676 (N_6676,N_6458,N_6441);
or U6677 (N_6677,N_6448,N_6285);
and U6678 (N_6678,N_6255,N_6335);
xnor U6679 (N_6679,N_6494,N_6476);
nand U6680 (N_6680,N_6332,N_6441);
nand U6681 (N_6681,N_6264,N_6306);
nor U6682 (N_6682,N_6466,N_6381);
nor U6683 (N_6683,N_6430,N_6469);
nand U6684 (N_6684,N_6270,N_6392);
nor U6685 (N_6685,N_6479,N_6422);
nand U6686 (N_6686,N_6324,N_6445);
nand U6687 (N_6687,N_6270,N_6264);
xnor U6688 (N_6688,N_6413,N_6481);
or U6689 (N_6689,N_6298,N_6299);
xor U6690 (N_6690,N_6489,N_6404);
nand U6691 (N_6691,N_6282,N_6357);
nor U6692 (N_6692,N_6428,N_6391);
or U6693 (N_6693,N_6468,N_6442);
or U6694 (N_6694,N_6288,N_6401);
or U6695 (N_6695,N_6379,N_6346);
and U6696 (N_6696,N_6482,N_6410);
nand U6697 (N_6697,N_6475,N_6332);
or U6698 (N_6698,N_6289,N_6304);
nand U6699 (N_6699,N_6445,N_6314);
nor U6700 (N_6700,N_6374,N_6496);
or U6701 (N_6701,N_6284,N_6400);
nand U6702 (N_6702,N_6457,N_6324);
nand U6703 (N_6703,N_6374,N_6359);
nor U6704 (N_6704,N_6488,N_6395);
or U6705 (N_6705,N_6451,N_6453);
nor U6706 (N_6706,N_6384,N_6282);
or U6707 (N_6707,N_6333,N_6491);
nand U6708 (N_6708,N_6458,N_6373);
and U6709 (N_6709,N_6423,N_6328);
nand U6710 (N_6710,N_6305,N_6317);
nand U6711 (N_6711,N_6398,N_6350);
nor U6712 (N_6712,N_6391,N_6377);
xnor U6713 (N_6713,N_6273,N_6438);
xor U6714 (N_6714,N_6395,N_6385);
xor U6715 (N_6715,N_6485,N_6481);
and U6716 (N_6716,N_6410,N_6290);
nor U6717 (N_6717,N_6379,N_6320);
or U6718 (N_6718,N_6272,N_6394);
and U6719 (N_6719,N_6304,N_6490);
nand U6720 (N_6720,N_6348,N_6271);
or U6721 (N_6721,N_6435,N_6464);
nor U6722 (N_6722,N_6478,N_6411);
nor U6723 (N_6723,N_6395,N_6458);
nand U6724 (N_6724,N_6312,N_6497);
and U6725 (N_6725,N_6455,N_6484);
or U6726 (N_6726,N_6266,N_6272);
nor U6727 (N_6727,N_6383,N_6488);
or U6728 (N_6728,N_6413,N_6320);
nand U6729 (N_6729,N_6376,N_6481);
nand U6730 (N_6730,N_6278,N_6494);
nand U6731 (N_6731,N_6310,N_6401);
nor U6732 (N_6732,N_6367,N_6325);
nand U6733 (N_6733,N_6425,N_6321);
and U6734 (N_6734,N_6400,N_6259);
nor U6735 (N_6735,N_6405,N_6315);
nor U6736 (N_6736,N_6343,N_6499);
nand U6737 (N_6737,N_6472,N_6498);
xnor U6738 (N_6738,N_6391,N_6317);
xor U6739 (N_6739,N_6295,N_6426);
or U6740 (N_6740,N_6362,N_6497);
or U6741 (N_6741,N_6313,N_6282);
xor U6742 (N_6742,N_6278,N_6289);
xor U6743 (N_6743,N_6454,N_6490);
or U6744 (N_6744,N_6276,N_6332);
nand U6745 (N_6745,N_6384,N_6354);
or U6746 (N_6746,N_6460,N_6311);
xnor U6747 (N_6747,N_6393,N_6466);
or U6748 (N_6748,N_6436,N_6306);
and U6749 (N_6749,N_6267,N_6398);
xnor U6750 (N_6750,N_6682,N_6638);
xnor U6751 (N_6751,N_6514,N_6701);
xor U6752 (N_6752,N_6606,N_6575);
nand U6753 (N_6753,N_6567,N_6600);
nor U6754 (N_6754,N_6627,N_6536);
xnor U6755 (N_6755,N_6705,N_6747);
xnor U6756 (N_6756,N_6692,N_6640);
and U6757 (N_6757,N_6535,N_6667);
and U6758 (N_6758,N_6681,N_6566);
and U6759 (N_6759,N_6612,N_6516);
and U6760 (N_6760,N_6576,N_6617);
xnor U6761 (N_6761,N_6557,N_6501);
or U6762 (N_6762,N_6581,N_6620);
or U6763 (N_6763,N_6744,N_6673);
and U6764 (N_6764,N_6707,N_6724);
and U6765 (N_6765,N_6716,N_6730);
or U6766 (N_6766,N_6732,N_6528);
and U6767 (N_6767,N_6597,N_6723);
or U6768 (N_6768,N_6718,N_6533);
xnor U6769 (N_6769,N_6689,N_6662);
and U6770 (N_6770,N_6683,N_6670);
nand U6771 (N_6771,N_6595,N_6582);
nor U6772 (N_6772,N_6526,N_6562);
or U6773 (N_6773,N_6635,N_6548);
nor U6774 (N_6774,N_6537,N_6655);
or U6775 (N_6775,N_6672,N_6529);
nand U6776 (N_6776,N_6502,N_6608);
nand U6777 (N_6777,N_6740,N_6573);
and U6778 (N_6778,N_6527,N_6614);
or U6779 (N_6779,N_6518,N_6715);
nor U6780 (N_6780,N_6733,N_6645);
and U6781 (N_6781,N_6714,N_6569);
or U6782 (N_6782,N_6632,N_6719);
xor U6783 (N_6783,N_6579,N_6694);
or U6784 (N_6784,N_6626,N_6742);
and U6785 (N_6785,N_6663,N_6686);
xor U6786 (N_6786,N_6578,N_6570);
nand U6787 (N_6787,N_6674,N_6648);
and U6788 (N_6788,N_6589,N_6622);
and U6789 (N_6789,N_6583,N_6746);
xnor U6790 (N_6790,N_6649,N_6659);
and U6791 (N_6791,N_6734,N_6748);
nor U6792 (N_6792,N_6717,N_6611);
xor U6793 (N_6793,N_6675,N_6669);
nand U6794 (N_6794,N_6510,N_6610);
nand U6795 (N_6795,N_6621,N_6619);
xnor U6796 (N_6796,N_6712,N_6731);
xor U6797 (N_6797,N_6658,N_6603);
nor U6798 (N_6798,N_6656,N_6738);
nand U6799 (N_6799,N_6531,N_6704);
nor U6800 (N_6800,N_6546,N_6699);
and U6801 (N_6801,N_6591,N_6698);
and U6802 (N_6802,N_6678,N_6585);
and U6803 (N_6803,N_6513,N_6671);
nor U6804 (N_6804,N_6685,N_6602);
and U6805 (N_6805,N_6598,N_6605);
nand U6806 (N_6806,N_6511,N_6521);
and U6807 (N_6807,N_6630,N_6625);
nand U6808 (N_6808,N_6563,N_6596);
xor U6809 (N_6809,N_6559,N_6544);
nand U6810 (N_6810,N_6697,N_6515);
or U6811 (N_6811,N_6572,N_6539);
nand U6812 (N_6812,N_6644,N_6580);
xnor U6813 (N_6813,N_6609,N_6534);
xor U6814 (N_6814,N_6532,N_6636);
xor U6815 (N_6815,N_6652,N_6711);
nor U6816 (N_6816,N_6651,N_6509);
xnor U6817 (N_6817,N_6618,N_6550);
nor U6818 (N_6818,N_6650,N_6592);
nor U6819 (N_6819,N_6604,N_6696);
nand U6820 (N_6820,N_6590,N_6506);
xnor U6821 (N_6821,N_6646,N_6586);
nor U6822 (N_6822,N_6708,N_6519);
xor U6823 (N_6823,N_6588,N_6637);
nand U6824 (N_6824,N_6739,N_6577);
nor U6825 (N_6825,N_6735,N_6549);
and U6826 (N_6826,N_6709,N_6525);
xor U6827 (N_6827,N_6512,N_6561);
nor U6828 (N_6828,N_6547,N_6553);
and U6829 (N_6829,N_6693,N_6555);
and U6830 (N_6830,N_6593,N_6503);
nand U6831 (N_6831,N_6607,N_6721);
or U6832 (N_6832,N_6727,N_6530);
nand U6833 (N_6833,N_6599,N_6538);
nand U6834 (N_6834,N_6560,N_6710);
or U6835 (N_6835,N_6700,N_6584);
xnor U6836 (N_6836,N_6676,N_6737);
and U6837 (N_6837,N_6556,N_6641);
and U6838 (N_6838,N_6545,N_6691);
or U6839 (N_6839,N_6541,N_6729);
nor U6840 (N_6840,N_6647,N_6660);
nand U6841 (N_6841,N_6664,N_6633);
and U6842 (N_6842,N_6615,N_6571);
and U6843 (N_6843,N_6568,N_6564);
nand U6844 (N_6844,N_6639,N_6507);
or U6845 (N_6845,N_6749,N_6679);
xnor U6846 (N_6846,N_6624,N_6594);
and U6847 (N_6847,N_6720,N_6628);
or U6848 (N_6848,N_6543,N_6623);
and U6849 (N_6849,N_6695,N_6680);
or U6850 (N_6850,N_6517,N_6574);
or U6851 (N_6851,N_6523,N_6587);
nand U6852 (N_6852,N_6702,N_6690);
nand U6853 (N_6853,N_6554,N_6558);
xor U6854 (N_6854,N_6653,N_6524);
nand U6855 (N_6855,N_6668,N_6520);
or U6856 (N_6856,N_6741,N_6684);
nand U6857 (N_6857,N_6736,N_6631);
or U6858 (N_6858,N_6706,N_6505);
nand U6859 (N_6859,N_6522,N_6500);
nand U6860 (N_6860,N_6542,N_6642);
nand U6861 (N_6861,N_6687,N_6728);
and U6862 (N_6862,N_6657,N_6613);
or U6863 (N_6863,N_6677,N_6661);
or U6864 (N_6864,N_6634,N_6743);
or U6865 (N_6865,N_6616,N_6703);
nand U6866 (N_6866,N_6551,N_6722);
xor U6867 (N_6867,N_6504,N_6629);
and U6868 (N_6868,N_6713,N_6725);
nand U6869 (N_6869,N_6552,N_6540);
xnor U6870 (N_6870,N_6601,N_6688);
nor U6871 (N_6871,N_6508,N_6666);
and U6872 (N_6872,N_6745,N_6726);
and U6873 (N_6873,N_6654,N_6565);
nand U6874 (N_6874,N_6643,N_6665);
and U6875 (N_6875,N_6630,N_6609);
or U6876 (N_6876,N_6633,N_6647);
nor U6877 (N_6877,N_6689,N_6726);
nor U6878 (N_6878,N_6638,N_6512);
nand U6879 (N_6879,N_6680,N_6741);
xnor U6880 (N_6880,N_6678,N_6542);
and U6881 (N_6881,N_6617,N_6722);
and U6882 (N_6882,N_6505,N_6519);
or U6883 (N_6883,N_6507,N_6549);
nor U6884 (N_6884,N_6534,N_6670);
or U6885 (N_6885,N_6718,N_6610);
and U6886 (N_6886,N_6640,N_6739);
and U6887 (N_6887,N_6735,N_6604);
and U6888 (N_6888,N_6672,N_6506);
nor U6889 (N_6889,N_6586,N_6502);
and U6890 (N_6890,N_6722,N_6674);
nor U6891 (N_6891,N_6588,N_6670);
nand U6892 (N_6892,N_6621,N_6651);
xnor U6893 (N_6893,N_6542,N_6673);
nor U6894 (N_6894,N_6722,N_6626);
nor U6895 (N_6895,N_6678,N_6747);
or U6896 (N_6896,N_6707,N_6698);
and U6897 (N_6897,N_6523,N_6722);
nor U6898 (N_6898,N_6736,N_6639);
nor U6899 (N_6899,N_6591,N_6516);
nand U6900 (N_6900,N_6651,N_6743);
and U6901 (N_6901,N_6635,N_6708);
or U6902 (N_6902,N_6540,N_6675);
xor U6903 (N_6903,N_6501,N_6505);
nand U6904 (N_6904,N_6617,N_6520);
nand U6905 (N_6905,N_6644,N_6632);
or U6906 (N_6906,N_6669,N_6569);
or U6907 (N_6907,N_6691,N_6540);
and U6908 (N_6908,N_6568,N_6658);
nand U6909 (N_6909,N_6515,N_6629);
nor U6910 (N_6910,N_6707,N_6607);
xnor U6911 (N_6911,N_6629,N_6609);
xnor U6912 (N_6912,N_6514,N_6741);
or U6913 (N_6913,N_6568,N_6695);
nor U6914 (N_6914,N_6684,N_6519);
xnor U6915 (N_6915,N_6515,N_6582);
or U6916 (N_6916,N_6554,N_6654);
and U6917 (N_6917,N_6606,N_6690);
nor U6918 (N_6918,N_6654,N_6664);
nand U6919 (N_6919,N_6701,N_6558);
xnor U6920 (N_6920,N_6715,N_6571);
or U6921 (N_6921,N_6633,N_6593);
nand U6922 (N_6922,N_6531,N_6547);
and U6923 (N_6923,N_6740,N_6500);
nand U6924 (N_6924,N_6693,N_6673);
nand U6925 (N_6925,N_6723,N_6518);
nor U6926 (N_6926,N_6585,N_6711);
or U6927 (N_6927,N_6612,N_6674);
nand U6928 (N_6928,N_6732,N_6684);
nand U6929 (N_6929,N_6738,N_6632);
xor U6930 (N_6930,N_6657,N_6673);
and U6931 (N_6931,N_6522,N_6647);
nand U6932 (N_6932,N_6636,N_6603);
nand U6933 (N_6933,N_6618,N_6595);
xor U6934 (N_6934,N_6613,N_6660);
nor U6935 (N_6935,N_6512,N_6563);
xor U6936 (N_6936,N_6508,N_6682);
nor U6937 (N_6937,N_6663,N_6619);
nor U6938 (N_6938,N_6609,N_6720);
xor U6939 (N_6939,N_6746,N_6684);
nor U6940 (N_6940,N_6591,N_6737);
nand U6941 (N_6941,N_6619,N_6607);
xnor U6942 (N_6942,N_6703,N_6620);
or U6943 (N_6943,N_6732,N_6512);
xnor U6944 (N_6944,N_6502,N_6601);
or U6945 (N_6945,N_6672,N_6640);
nor U6946 (N_6946,N_6647,N_6585);
nor U6947 (N_6947,N_6502,N_6678);
and U6948 (N_6948,N_6670,N_6529);
xnor U6949 (N_6949,N_6511,N_6587);
or U6950 (N_6950,N_6590,N_6511);
nor U6951 (N_6951,N_6677,N_6646);
xnor U6952 (N_6952,N_6658,N_6719);
nand U6953 (N_6953,N_6576,N_6543);
and U6954 (N_6954,N_6560,N_6661);
nand U6955 (N_6955,N_6681,N_6704);
nor U6956 (N_6956,N_6533,N_6517);
and U6957 (N_6957,N_6510,N_6598);
nor U6958 (N_6958,N_6660,N_6626);
nand U6959 (N_6959,N_6574,N_6683);
nor U6960 (N_6960,N_6572,N_6609);
nand U6961 (N_6961,N_6509,N_6646);
xnor U6962 (N_6962,N_6726,N_6744);
nor U6963 (N_6963,N_6626,N_6624);
or U6964 (N_6964,N_6644,N_6712);
nor U6965 (N_6965,N_6677,N_6746);
nor U6966 (N_6966,N_6629,N_6523);
nand U6967 (N_6967,N_6658,N_6745);
and U6968 (N_6968,N_6582,N_6517);
xor U6969 (N_6969,N_6675,N_6744);
nand U6970 (N_6970,N_6648,N_6536);
or U6971 (N_6971,N_6522,N_6689);
xor U6972 (N_6972,N_6672,N_6636);
nand U6973 (N_6973,N_6629,N_6730);
xnor U6974 (N_6974,N_6623,N_6664);
nand U6975 (N_6975,N_6503,N_6736);
nand U6976 (N_6976,N_6709,N_6667);
nand U6977 (N_6977,N_6609,N_6587);
and U6978 (N_6978,N_6504,N_6694);
xor U6979 (N_6979,N_6627,N_6746);
nor U6980 (N_6980,N_6650,N_6554);
xor U6981 (N_6981,N_6747,N_6738);
or U6982 (N_6982,N_6579,N_6525);
and U6983 (N_6983,N_6545,N_6542);
nand U6984 (N_6984,N_6666,N_6728);
nor U6985 (N_6985,N_6606,N_6625);
nand U6986 (N_6986,N_6648,N_6689);
xor U6987 (N_6987,N_6609,N_6731);
and U6988 (N_6988,N_6688,N_6504);
and U6989 (N_6989,N_6650,N_6525);
xnor U6990 (N_6990,N_6629,N_6616);
xnor U6991 (N_6991,N_6522,N_6747);
nand U6992 (N_6992,N_6533,N_6700);
or U6993 (N_6993,N_6548,N_6601);
nand U6994 (N_6994,N_6610,N_6724);
and U6995 (N_6995,N_6671,N_6519);
xnor U6996 (N_6996,N_6502,N_6736);
and U6997 (N_6997,N_6734,N_6605);
or U6998 (N_6998,N_6726,N_6567);
nor U6999 (N_6999,N_6628,N_6546);
and U7000 (N_7000,N_6937,N_6835);
and U7001 (N_7001,N_6766,N_6880);
nor U7002 (N_7002,N_6867,N_6815);
and U7003 (N_7003,N_6758,N_6898);
and U7004 (N_7004,N_6764,N_6863);
xnor U7005 (N_7005,N_6926,N_6939);
nand U7006 (N_7006,N_6813,N_6922);
xnor U7007 (N_7007,N_6824,N_6757);
and U7008 (N_7008,N_6808,N_6977);
nor U7009 (N_7009,N_6802,N_6969);
nand U7010 (N_7010,N_6872,N_6991);
xnor U7011 (N_7011,N_6938,N_6933);
nor U7012 (N_7012,N_6804,N_6777);
nand U7013 (N_7013,N_6942,N_6838);
or U7014 (N_7014,N_6828,N_6853);
nor U7015 (N_7015,N_6826,N_6791);
and U7016 (N_7016,N_6751,N_6906);
or U7017 (N_7017,N_6836,N_6874);
or U7018 (N_7018,N_6752,N_6899);
xor U7019 (N_7019,N_6805,N_6830);
nand U7020 (N_7020,N_6958,N_6785);
and U7021 (N_7021,N_6895,N_6810);
xnor U7022 (N_7022,N_6784,N_6888);
nand U7023 (N_7023,N_6782,N_6847);
xor U7024 (N_7024,N_6894,N_6846);
and U7025 (N_7025,N_6797,N_6765);
or U7026 (N_7026,N_6796,N_6893);
nor U7027 (N_7027,N_6916,N_6961);
xor U7028 (N_7028,N_6923,N_6754);
or U7029 (N_7029,N_6806,N_6914);
nor U7030 (N_7030,N_6783,N_6882);
and U7031 (N_7031,N_6845,N_6989);
or U7032 (N_7032,N_6908,N_6809);
nand U7033 (N_7033,N_6935,N_6983);
or U7034 (N_7034,N_6753,N_6781);
and U7035 (N_7035,N_6965,N_6931);
or U7036 (N_7036,N_6994,N_6865);
xor U7037 (N_7037,N_6812,N_6801);
xor U7038 (N_7038,N_6952,N_6869);
nor U7039 (N_7039,N_6966,N_6875);
nor U7040 (N_7040,N_6901,N_6821);
nand U7041 (N_7041,N_6920,N_6822);
nor U7042 (N_7042,N_6771,N_6978);
nor U7043 (N_7043,N_6930,N_6998);
nor U7044 (N_7044,N_6775,N_6790);
or U7045 (N_7045,N_6891,N_6780);
and U7046 (N_7046,N_6951,N_6981);
and U7047 (N_7047,N_6912,N_6940);
nand U7048 (N_7048,N_6871,N_6843);
nor U7049 (N_7049,N_6964,N_6968);
xnor U7050 (N_7050,N_6928,N_6884);
or U7051 (N_7051,N_6918,N_6852);
and U7052 (N_7052,N_6772,N_6941);
or U7053 (N_7053,N_6924,N_6995);
or U7054 (N_7054,N_6881,N_6756);
or U7055 (N_7055,N_6949,N_6996);
or U7056 (N_7056,N_6857,N_6788);
nand U7057 (N_7057,N_6768,N_6792);
xnor U7058 (N_7058,N_6892,N_6816);
and U7059 (N_7059,N_6900,N_6982);
nor U7060 (N_7060,N_6887,N_6832);
nor U7061 (N_7061,N_6825,N_6851);
and U7062 (N_7062,N_6963,N_6763);
nand U7063 (N_7063,N_6819,N_6903);
and U7064 (N_7064,N_6913,N_6955);
nor U7065 (N_7065,N_6929,N_6936);
and U7066 (N_7066,N_6798,N_6962);
nor U7067 (N_7067,N_6840,N_6823);
or U7068 (N_7068,N_6879,N_6957);
nand U7069 (N_7069,N_6934,N_6868);
and U7070 (N_7070,N_6886,N_6786);
nor U7071 (N_7071,N_6870,N_6876);
xor U7072 (N_7072,N_6945,N_6859);
or U7073 (N_7073,N_6946,N_6837);
nand U7074 (N_7074,N_6789,N_6890);
nor U7075 (N_7075,N_6988,N_6755);
and U7076 (N_7076,N_6985,N_6959);
xor U7077 (N_7077,N_6814,N_6896);
and U7078 (N_7078,N_6855,N_6807);
or U7079 (N_7079,N_6762,N_6904);
xor U7080 (N_7080,N_6820,N_6774);
xnor U7081 (N_7081,N_6944,N_6787);
and U7082 (N_7082,N_6910,N_6844);
or U7083 (N_7083,N_6954,N_6987);
xor U7084 (N_7084,N_6866,N_6834);
and U7085 (N_7085,N_6776,N_6921);
nor U7086 (N_7086,N_6850,N_6839);
xor U7087 (N_7087,N_6778,N_6833);
and U7088 (N_7088,N_6897,N_6948);
and U7089 (N_7089,N_6905,N_6990);
nor U7090 (N_7090,N_6975,N_6769);
xor U7091 (N_7091,N_6759,N_6818);
nor U7092 (N_7092,N_6971,N_6993);
nor U7093 (N_7093,N_6750,N_6760);
nand U7094 (N_7094,N_6947,N_6793);
or U7095 (N_7095,N_6858,N_6799);
or U7096 (N_7096,N_6761,N_6883);
xnor U7097 (N_7097,N_6967,N_6885);
nand U7098 (N_7098,N_6770,N_6767);
xnor U7099 (N_7099,N_6972,N_6779);
and U7100 (N_7100,N_6795,N_6950);
and U7101 (N_7101,N_6829,N_6862);
and U7102 (N_7102,N_6800,N_6878);
nor U7103 (N_7103,N_6943,N_6831);
and U7104 (N_7104,N_6873,N_6849);
nand U7105 (N_7105,N_6803,N_6980);
nand U7106 (N_7106,N_6842,N_6999);
and U7107 (N_7107,N_6976,N_6877);
nor U7108 (N_7108,N_6992,N_6889);
or U7109 (N_7109,N_6960,N_6925);
nor U7110 (N_7110,N_6953,N_6979);
and U7111 (N_7111,N_6854,N_6856);
nor U7112 (N_7112,N_6919,N_6811);
xnor U7113 (N_7113,N_6794,N_6970);
nand U7114 (N_7114,N_6927,N_6841);
or U7115 (N_7115,N_6956,N_6911);
or U7116 (N_7116,N_6932,N_6917);
xor U7117 (N_7117,N_6773,N_6860);
or U7118 (N_7118,N_6861,N_6902);
or U7119 (N_7119,N_6974,N_6827);
or U7120 (N_7120,N_6915,N_6907);
nand U7121 (N_7121,N_6864,N_6986);
or U7122 (N_7122,N_6848,N_6909);
and U7123 (N_7123,N_6817,N_6997);
nor U7124 (N_7124,N_6973,N_6984);
nand U7125 (N_7125,N_6961,N_6931);
and U7126 (N_7126,N_6754,N_6910);
nand U7127 (N_7127,N_6892,N_6862);
nor U7128 (N_7128,N_6769,N_6955);
or U7129 (N_7129,N_6783,N_6832);
xnor U7130 (N_7130,N_6954,N_6939);
nor U7131 (N_7131,N_6908,N_6881);
and U7132 (N_7132,N_6940,N_6756);
or U7133 (N_7133,N_6820,N_6842);
nand U7134 (N_7134,N_6893,N_6990);
nand U7135 (N_7135,N_6871,N_6784);
nor U7136 (N_7136,N_6843,N_6929);
nor U7137 (N_7137,N_6835,N_6919);
xnor U7138 (N_7138,N_6898,N_6794);
or U7139 (N_7139,N_6997,N_6766);
nor U7140 (N_7140,N_6903,N_6859);
or U7141 (N_7141,N_6944,N_6774);
nand U7142 (N_7142,N_6986,N_6948);
or U7143 (N_7143,N_6843,N_6859);
nor U7144 (N_7144,N_6763,N_6818);
xor U7145 (N_7145,N_6800,N_6972);
or U7146 (N_7146,N_6998,N_6888);
nor U7147 (N_7147,N_6870,N_6758);
and U7148 (N_7148,N_6767,N_6825);
or U7149 (N_7149,N_6912,N_6870);
or U7150 (N_7150,N_6867,N_6892);
or U7151 (N_7151,N_6796,N_6896);
and U7152 (N_7152,N_6989,N_6821);
nor U7153 (N_7153,N_6883,N_6818);
nand U7154 (N_7154,N_6884,N_6794);
nand U7155 (N_7155,N_6893,N_6787);
nor U7156 (N_7156,N_6952,N_6789);
or U7157 (N_7157,N_6875,N_6996);
xnor U7158 (N_7158,N_6863,N_6954);
xnor U7159 (N_7159,N_6785,N_6914);
nor U7160 (N_7160,N_6842,N_6806);
or U7161 (N_7161,N_6999,N_6839);
and U7162 (N_7162,N_6998,N_6958);
and U7163 (N_7163,N_6823,N_6964);
xnor U7164 (N_7164,N_6918,N_6919);
nor U7165 (N_7165,N_6963,N_6862);
and U7166 (N_7166,N_6937,N_6943);
and U7167 (N_7167,N_6911,N_6998);
nand U7168 (N_7168,N_6759,N_6986);
nor U7169 (N_7169,N_6803,N_6877);
xnor U7170 (N_7170,N_6760,N_6772);
or U7171 (N_7171,N_6834,N_6871);
nand U7172 (N_7172,N_6841,N_6943);
or U7173 (N_7173,N_6986,N_6867);
and U7174 (N_7174,N_6845,N_6774);
nor U7175 (N_7175,N_6910,N_6926);
xor U7176 (N_7176,N_6868,N_6886);
xor U7177 (N_7177,N_6759,N_6826);
or U7178 (N_7178,N_6848,N_6808);
nand U7179 (N_7179,N_6949,N_6784);
nand U7180 (N_7180,N_6769,N_6889);
xnor U7181 (N_7181,N_6920,N_6852);
xor U7182 (N_7182,N_6813,N_6987);
nor U7183 (N_7183,N_6838,N_6949);
xor U7184 (N_7184,N_6765,N_6937);
nor U7185 (N_7185,N_6772,N_6839);
and U7186 (N_7186,N_6910,N_6957);
nor U7187 (N_7187,N_6960,N_6911);
and U7188 (N_7188,N_6767,N_6827);
xnor U7189 (N_7189,N_6770,N_6774);
nor U7190 (N_7190,N_6834,N_6770);
nand U7191 (N_7191,N_6962,N_6922);
or U7192 (N_7192,N_6895,N_6801);
xor U7193 (N_7193,N_6787,N_6795);
nand U7194 (N_7194,N_6948,N_6889);
or U7195 (N_7195,N_6792,N_6835);
nor U7196 (N_7196,N_6841,N_6762);
xnor U7197 (N_7197,N_6970,N_6842);
or U7198 (N_7198,N_6818,N_6997);
nor U7199 (N_7199,N_6961,N_6815);
or U7200 (N_7200,N_6789,N_6867);
nand U7201 (N_7201,N_6996,N_6916);
and U7202 (N_7202,N_6889,N_6929);
nor U7203 (N_7203,N_6796,N_6979);
nor U7204 (N_7204,N_6990,N_6954);
nor U7205 (N_7205,N_6937,N_6995);
and U7206 (N_7206,N_6919,N_6938);
xor U7207 (N_7207,N_6822,N_6825);
nand U7208 (N_7208,N_6772,N_6949);
nand U7209 (N_7209,N_6890,N_6832);
and U7210 (N_7210,N_6995,N_6803);
xnor U7211 (N_7211,N_6852,N_6989);
nor U7212 (N_7212,N_6891,N_6902);
xor U7213 (N_7213,N_6943,N_6944);
xnor U7214 (N_7214,N_6876,N_6829);
or U7215 (N_7215,N_6927,N_6810);
or U7216 (N_7216,N_6947,N_6886);
xor U7217 (N_7217,N_6861,N_6860);
xor U7218 (N_7218,N_6816,N_6977);
or U7219 (N_7219,N_6758,N_6833);
and U7220 (N_7220,N_6997,N_6764);
nand U7221 (N_7221,N_6789,N_6764);
and U7222 (N_7222,N_6836,N_6868);
xor U7223 (N_7223,N_6977,N_6772);
nor U7224 (N_7224,N_6976,N_6805);
nand U7225 (N_7225,N_6802,N_6976);
nor U7226 (N_7226,N_6753,N_6973);
or U7227 (N_7227,N_6852,N_6859);
and U7228 (N_7228,N_6920,N_6770);
xor U7229 (N_7229,N_6819,N_6843);
xnor U7230 (N_7230,N_6800,N_6913);
xnor U7231 (N_7231,N_6762,N_6805);
xnor U7232 (N_7232,N_6975,N_6994);
and U7233 (N_7233,N_6920,N_6781);
or U7234 (N_7234,N_6912,N_6888);
nor U7235 (N_7235,N_6961,N_6918);
or U7236 (N_7236,N_6839,N_6946);
xnor U7237 (N_7237,N_6776,N_6804);
xnor U7238 (N_7238,N_6871,N_6966);
nand U7239 (N_7239,N_6919,N_6871);
nor U7240 (N_7240,N_6801,N_6844);
nor U7241 (N_7241,N_6983,N_6912);
or U7242 (N_7242,N_6983,N_6750);
xor U7243 (N_7243,N_6785,N_6772);
nand U7244 (N_7244,N_6900,N_6968);
xnor U7245 (N_7245,N_6978,N_6879);
xnor U7246 (N_7246,N_6977,N_6953);
and U7247 (N_7247,N_6919,N_6846);
xnor U7248 (N_7248,N_6855,N_6929);
or U7249 (N_7249,N_6865,N_6928);
xnor U7250 (N_7250,N_7034,N_7015);
xor U7251 (N_7251,N_7041,N_7045);
or U7252 (N_7252,N_7101,N_7179);
or U7253 (N_7253,N_7175,N_7168);
nor U7254 (N_7254,N_7003,N_7167);
nand U7255 (N_7255,N_7114,N_7176);
and U7256 (N_7256,N_7171,N_7042);
nor U7257 (N_7257,N_7187,N_7018);
or U7258 (N_7258,N_7150,N_7007);
or U7259 (N_7259,N_7155,N_7038);
nor U7260 (N_7260,N_7013,N_7203);
and U7261 (N_7261,N_7239,N_7165);
and U7262 (N_7262,N_7095,N_7115);
or U7263 (N_7263,N_7202,N_7166);
and U7264 (N_7264,N_7149,N_7244);
and U7265 (N_7265,N_7213,N_7146);
nor U7266 (N_7266,N_7241,N_7248);
and U7267 (N_7267,N_7033,N_7172);
xor U7268 (N_7268,N_7208,N_7199);
and U7269 (N_7269,N_7064,N_7097);
or U7270 (N_7270,N_7092,N_7243);
xnor U7271 (N_7271,N_7242,N_7031);
xor U7272 (N_7272,N_7132,N_7020);
and U7273 (N_7273,N_7117,N_7052);
nand U7274 (N_7274,N_7198,N_7140);
xor U7275 (N_7275,N_7035,N_7044);
xor U7276 (N_7276,N_7185,N_7159);
nor U7277 (N_7277,N_7008,N_7192);
nand U7278 (N_7278,N_7037,N_7107);
nand U7279 (N_7279,N_7133,N_7222);
nand U7280 (N_7280,N_7011,N_7170);
and U7281 (N_7281,N_7094,N_7012);
and U7282 (N_7282,N_7090,N_7209);
xnor U7283 (N_7283,N_7189,N_7183);
and U7284 (N_7284,N_7205,N_7125);
nor U7285 (N_7285,N_7067,N_7195);
nor U7286 (N_7286,N_7105,N_7046);
xor U7287 (N_7287,N_7194,N_7002);
nand U7288 (N_7288,N_7173,N_7188);
nor U7289 (N_7289,N_7048,N_7130);
or U7290 (N_7290,N_7049,N_7106);
nor U7291 (N_7291,N_7026,N_7224);
nand U7292 (N_7292,N_7055,N_7053);
xnor U7293 (N_7293,N_7004,N_7060);
and U7294 (N_7294,N_7093,N_7072);
xor U7295 (N_7295,N_7163,N_7063);
xor U7296 (N_7296,N_7074,N_7223);
nor U7297 (N_7297,N_7153,N_7010);
xor U7298 (N_7298,N_7186,N_7120);
nand U7299 (N_7299,N_7103,N_7204);
and U7300 (N_7300,N_7191,N_7231);
nand U7301 (N_7301,N_7190,N_7025);
or U7302 (N_7302,N_7099,N_7169);
xnor U7303 (N_7303,N_7238,N_7108);
or U7304 (N_7304,N_7181,N_7220);
xor U7305 (N_7305,N_7073,N_7193);
nand U7306 (N_7306,N_7214,N_7024);
or U7307 (N_7307,N_7138,N_7098);
nor U7308 (N_7308,N_7017,N_7177);
xnor U7309 (N_7309,N_7069,N_7030);
or U7310 (N_7310,N_7182,N_7080);
xor U7311 (N_7311,N_7174,N_7112);
nor U7312 (N_7312,N_7200,N_7068);
or U7313 (N_7313,N_7144,N_7040);
nand U7314 (N_7314,N_7139,N_7000);
or U7315 (N_7315,N_7128,N_7104);
xnor U7316 (N_7316,N_7152,N_7201);
or U7317 (N_7317,N_7233,N_7021);
and U7318 (N_7318,N_7219,N_7086);
nor U7319 (N_7319,N_7089,N_7210);
nor U7320 (N_7320,N_7197,N_7229);
xnor U7321 (N_7321,N_7043,N_7221);
xor U7322 (N_7322,N_7148,N_7160);
xor U7323 (N_7323,N_7102,N_7161);
nor U7324 (N_7324,N_7158,N_7116);
xor U7325 (N_7325,N_7058,N_7084);
nor U7326 (N_7326,N_7096,N_7156);
nor U7327 (N_7327,N_7065,N_7247);
xnor U7328 (N_7328,N_7057,N_7076);
nand U7329 (N_7329,N_7136,N_7022);
or U7330 (N_7330,N_7180,N_7051);
and U7331 (N_7331,N_7083,N_7014);
xnor U7332 (N_7332,N_7109,N_7211);
nand U7333 (N_7333,N_7054,N_7028);
or U7334 (N_7334,N_7126,N_7147);
xor U7335 (N_7335,N_7145,N_7056);
and U7336 (N_7336,N_7164,N_7245);
nand U7337 (N_7337,N_7062,N_7135);
nand U7338 (N_7338,N_7023,N_7079);
xnor U7339 (N_7339,N_7228,N_7151);
and U7340 (N_7340,N_7006,N_7218);
nand U7341 (N_7341,N_7077,N_7016);
xor U7342 (N_7342,N_7206,N_7082);
nor U7343 (N_7343,N_7131,N_7081);
nand U7344 (N_7344,N_7196,N_7087);
nor U7345 (N_7345,N_7111,N_7119);
nand U7346 (N_7346,N_7127,N_7240);
xnor U7347 (N_7347,N_7207,N_7184);
or U7348 (N_7348,N_7134,N_7078);
xnor U7349 (N_7349,N_7143,N_7088);
or U7350 (N_7350,N_7032,N_7039);
or U7351 (N_7351,N_7178,N_7059);
nand U7352 (N_7352,N_7009,N_7029);
nand U7353 (N_7353,N_7212,N_7124);
or U7354 (N_7354,N_7071,N_7235);
and U7355 (N_7355,N_7123,N_7110);
or U7356 (N_7356,N_7154,N_7230);
nand U7357 (N_7357,N_7227,N_7215);
nor U7358 (N_7358,N_7061,N_7137);
or U7359 (N_7359,N_7237,N_7122);
and U7360 (N_7360,N_7249,N_7236);
xor U7361 (N_7361,N_7226,N_7047);
nand U7362 (N_7362,N_7075,N_7162);
nor U7363 (N_7363,N_7019,N_7005);
xor U7364 (N_7364,N_7036,N_7070);
nor U7365 (N_7365,N_7246,N_7027);
xor U7366 (N_7366,N_7118,N_7216);
or U7367 (N_7367,N_7129,N_7232);
nand U7368 (N_7368,N_7066,N_7121);
xor U7369 (N_7369,N_7050,N_7234);
nand U7370 (N_7370,N_7217,N_7141);
nor U7371 (N_7371,N_7225,N_7001);
or U7372 (N_7372,N_7142,N_7085);
xnor U7373 (N_7373,N_7100,N_7157);
or U7374 (N_7374,N_7113,N_7091);
nor U7375 (N_7375,N_7048,N_7201);
xor U7376 (N_7376,N_7197,N_7027);
or U7377 (N_7377,N_7227,N_7196);
nor U7378 (N_7378,N_7091,N_7033);
nor U7379 (N_7379,N_7113,N_7107);
nor U7380 (N_7380,N_7078,N_7131);
and U7381 (N_7381,N_7084,N_7047);
nand U7382 (N_7382,N_7088,N_7108);
or U7383 (N_7383,N_7176,N_7137);
xnor U7384 (N_7384,N_7152,N_7093);
nand U7385 (N_7385,N_7151,N_7061);
nand U7386 (N_7386,N_7023,N_7028);
and U7387 (N_7387,N_7023,N_7082);
and U7388 (N_7388,N_7216,N_7222);
nand U7389 (N_7389,N_7054,N_7127);
xnor U7390 (N_7390,N_7164,N_7248);
and U7391 (N_7391,N_7187,N_7040);
and U7392 (N_7392,N_7183,N_7059);
nand U7393 (N_7393,N_7053,N_7240);
or U7394 (N_7394,N_7147,N_7150);
nand U7395 (N_7395,N_7004,N_7151);
nand U7396 (N_7396,N_7150,N_7178);
nand U7397 (N_7397,N_7166,N_7046);
nor U7398 (N_7398,N_7165,N_7036);
or U7399 (N_7399,N_7071,N_7094);
xor U7400 (N_7400,N_7200,N_7039);
nor U7401 (N_7401,N_7205,N_7214);
nand U7402 (N_7402,N_7202,N_7229);
nand U7403 (N_7403,N_7011,N_7066);
and U7404 (N_7404,N_7091,N_7046);
nand U7405 (N_7405,N_7042,N_7103);
nor U7406 (N_7406,N_7007,N_7194);
or U7407 (N_7407,N_7201,N_7127);
nor U7408 (N_7408,N_7209,N_7012);
xnor U7409 (N_7409,N_7110,N_7098);
or U7410 (N_7410,N_7064,N_7074);
nand U7411 (N_7411,N_7160,N_7061);
nor U7412 (N_7412,N_7212,N_7132);
or U7413 (N_7413,N_7181,N_7238);
nor U7414 (N_7414,N_7069,N_7022);
nand U7415 (N_7415,N_7148,N_7223);
nor U7416 (N_7416,N_7008,N_7073);
or U7417 (N_7417,N_7128,N_7109);
xor U7418 (N_7418,N_7000,N_7181);
and U7419 (N_7419,N_7098,N_7168);
xor U7420 (N_7420,N_7189,N_7024);
xnor U7421 (N_7421,N_7042,N_7172);
nor U7422 (N_7422,N_7153,N_7048);
xnor U7423 (N_7423,N_7217,N_7025);
nor U7424 (N_7424,N_7115,N_7247);
xnor U7425 (N_7425,N_7108,N_7082);
xor U7426 (N_7426,N_7184,N_7066);
nand U7427 (N_7427,N_7219,N_7034);
xnor U7428 (N_7428,N_7175,N_7188);
and U7429 (N_7429,N_7133,N_7024);
xnor U7430 (N_7430,N_7004,N_7223);
nand U7431 (N_7431,N_7092,N_7043);
and U7432 (N_7432,N_7054,N_7102);
nand U7433 (N_7433,N_7071,N_7236);
nor U7434 (N_7434,N_7235,N_7025);
nand U7435 (N_7435,N_7165,N_7066);
or U7436 (N_7436,N_7043,N_7005);
and U7437 (N_7437,N_7133,N_7127);
or U7438 (N_7438,N_7101,N_7175);
nor U7439 (N_7439,N_7144,N_7152);
xnor U7440 (N_7440,N_7198,N_7223);
nand U7441 (N_7441,N_7010,N_7089);
xnor U7442 (N_7442,N_7021,N_7109);
xor U7443 (N_7443,N_7035,N_7147);
xnor U7444 (N_7444,N_7022,N_7000);
or U7445 (N_7445,N_7197,N_7119);
xnor U7446 (N_7446,N_7016,N_7078);
or U7447 (N_7447,N_7129,N_7113);
nor U7448 (N_7448,N_7096,N_7203);
nor U7449 (N_7449,N_7219,N_7100);
nand U7450 (N_7450,N_7177,N_7138);
nand U7451 (N_7451,N_7224,N_7030);
nand U7452 (N_7452,N_7242,N_7219);
xnor U7453 (N_7453,N_7224,N_7209);
nor U7454 (N_7454,N_7124,N_7103);
and U7455 (N_7455,N_7046,N_7021);
nor U7456 (N_7456,N_7127,N_7155);
nor U7457 (N_7457,N_7073,N_7231);
or U7458 (N_7458,N_7157,N_7125);
or U7459 (N_7459,N_7153,N_7018);
and U7460 (N_7460,N_7183,N_7214);
xor U7461 (N_7461,N_7030,N_7057);
xor U7462 (N_7462,N_7194,N_7068);
nor U7463 (N_7463,N_7028,N_7096);
xor U7464 (N_7464,N_7015,N_7049);
nor U7465 (N_7465,N_7196,N_7032);
or U7466 (N_7466,N_7077,N_7029);
xor U7467 (N_7467,N_7112,N_7217);
and U7468 (N_7468,N_7040,N_7086);
or U7469 (N_7469,N_7027,N_7217);
nor U7470 (N_7470,N_7226,N_7118);
or U7471 (N_7471,N_7200,N_7181);
or U7472 (N_7472,N_7058,N_7203);
or U7473 (N_7473,N_7157,N_7086);
or U7474 (N_7474,N_7002,N_7134);
nand U7475 (N_7475,N_7064,N_7180);
and U7476 (N_7476,N_7102,N_7201);
nor U7477 (N_7477,N_7112,N_7064);
nor U7478 (N_7478,N_7106,N_7235);
nor U7479 (N_7479,N_7068,N_7066);
nand U7480 (N_7480,N_7011,N_7107);
and U7481 (N_7481,N_7162,N_7195);
xor U7482 (N_7482,N_7012,N_7030);
and U7483 (N_7483,N_7082,N_7085);
nor U7484 (N_7484,N_7110,N_7225);
xor U7485 (N_7485,N_7097,N_7173);
or U7486 (N_7486,N_7178,N_7172);
xor U7487 (N_7487,N_7090,N_7179);
and U7488 (N_7488,N_7245,N_7002);
and U7489 (N_7489,N_7101,N_7233);
xor U7490 (N_7490,N_7066,N_7034);
nand U7491 (N_7491,N_7075,N_7187);
nor U7492 (N_7492,N_7164,N_7078);
nor U7493 (N_7493,N_7010,N_7008);
xnor U7494 (N_7494,N_7151,N_7229);
nor U7495 (N_7495,N_7041,N_7141);
xnor U7496 (N_7496,N_7101,N_7095);
or U7497 (N_7497,N_7233,N_7106);
nand U7498 (N_7498,N_7099,N_7243);
xor U7499 (N_7499,N_7103,N_7018);
nor U7500 (N_7500,N_7413,N_7443);
or U7501 (N_7501,N_7282,N_7490);
nand U7502 (N_7502,N_7366,N_7392);
and U7503 (N_7503,N_7381,N_7293);
or U7504 (N_7504,N_7271,N_7478);
and U7505 (N_7505,N_7396,N_7441);
and U7506 (N_7506,N_7477,N_7493);
nand U7507 (N_7507,N_7264,N_7439);
nand U7508 (N_7508,N_7328,N_7495);
xnor U7509 (N_7509,N_7305,N_7465);
or U7510 (N_7510,N_7445,N_7474);
or U7511 (N_7511,N_7352,N_7317);
and U7512 (N_7512,N_7321,N_7268);
nand U7513 (N_7513,N_7440,N_7260);
and U7514 (N_7514,N_7491,N_7284);
xor U7515 (N_7515,N_7342,N_7404);
or U7516 (N_7516,N_7452,N_7279);
xnor U7517 (N_7517,N_7315,N_7471);
nor U7518 (N_7518,N_7298,N_7416);
nor U7519 (N_7519,N_7330,N_7411);
xor U7520 (N_7520,N_7361,N_7395);
or U7521 (N_7521,N_7384,N_7270);
or U7522 (N_7522,N_7438,N_7360);
and U7523 (N_7523,N_7364,N_7374);
xor U7524 (N_7524,N_7437,N_7300);
nand U7525 (N_7525,N_7383,N_7281);
nor U7526 (N_7526,N_7464,N_7424);
nor U7527 (N_7527,N_7409,N_7292);
nand U7528 (N_7528,N_7322,N_7336);
nand U7529 (N_7529,N_7388,N_7355);
nand U7530 (N_7530,N_7475,N_7299);
and U7531 (N_7531,N_7459,N_7362);
nand U7532 (N_7532,N_7447,N_7309);
xnor U7533 (N_7533,N_7435,N_7291);
nand U7534 (N_7534,N_7423,N_7346);
nor U7535 (N_7535,N_7399,N_7324);
and U7536 (N_7536,N_7455,N_7433);
nand U7537 (N_7537,N_7348,N_7486);
and U7538 (N_7538,N_7430,N_7469);
or U7539 (N_7539,N_7481,N_7320);
xnor U7540 (N_7540,N_7269,N_7426);
and U7541 (N_7541,N_7273,N_7325);
xnor U7542 (N_7542,N_7255,N_7254);
nor U7543 (N_7543,N_7393,N_7276);
nand U7544 (N_7544,N_7473,N_7340);
nand U7545 (N_7545,N_7417,N_7451);
nor U7546 (N_7546,N_7462,N_7334);
nand U7547 (N_7547,N_7405,N_7333);
and U7548 (N_7548,N_7419,N_7310);
nand U7549 (N_7549,N_7446,N_7327);
or U7550 (N_7550,N_7376,N_7338);
xnor U7551 (N_7551,N_7302,N_7422);
and U7552 (N_7552,N_7484,N_7341);
and U7553 (N_7553,N_7468,N_7343);
and U7554 (N_7554,N_7347,N_7373);
nand U7555 (N_7555,N_7483,N_7421);
nor U7556 (N_7556,N_7326,N_7354);
nor U7557 (N_7557,N_7467,N_7287);
and U7558 (N_7558,N_7337,N_7391);
xor U7559 (N_7559,N_7267,N_7407);
nand U7560 (N_7560,N_7259,N_7288);
and U7561 (N_7561,N_7345,N_7410);
xor U7562 (N_7562,N_7363,N_7494);
nor U7563 (N_7563,N_7262,N_7369);
nor U7564 (N_7564,N_7290,N_7316);
xor U7565 (N_7565,N_7349,N_7379);
or U7566 (N_7566,N_7296,N_7263);
or U7567 (N_7567,N_7250,N_7266);
nand U7568 (N_7568,N_7278,N_7353);
and U7569 (N_7569,N_7331,N_7257);
nor U7570 (N_7570,N_7377,N_7442);
and U7571 (N_7571,N_7251,N_7496);
xor U7572 (N_7572,N_7371,N_7488);
xnor U7573 (N_7573,N_7357,N_7400);
or U7574 (N_7574,N_7265,N_7294);
and U7575 (N_7575,N_7286,N_7301);
nor U7576 (N_7576,N_7358,N_7303);
nand U7577 (N_7577,N_7311,N_7444);
nand U7578 (N_7578,N_7323,N_7431);
and U7579 (N_7579,N_7428,N_7482);
or U7580 (N_7580,N_7314,N_7487);
or U7581 (N_7581,N_7449,N_7472);
nor U7582 (N_7582,N_7350,N_7356);
or U7583 (N_7583,N_7339,N_7274);
nor U7584 (N_7584,N_7318,N_7253);
nand U7585 (N_7585,N_7418,N_7402);
nor U7586 (N_7586,N_7401,N_7272);
nor U7587 (N_7587,N_7319,N_7485);
nor U7588 (N_7588,N_7463,N_7461);
and U7589 (N_7589,N_7436,N_7460);
nand U7590 (N_7590,N_7387,N_7492);
or U7591 (N_7591,N_7365,N_7261);
nand U7592 (N_7592,N_7499,N_7456);
nand U7593 (N_7593,N_7372,N_7458);
xor U7594 (N_7594,N_7295,N_7307);
nor U7595 (N_7595,N_7386,N_7308);
nor U7596 (N_7596,N_7252,N_7277);
nor U7597 (N_7597,N_7448,N_7258);
xor U7598 (N_7598,N_7432,N_7329);
and U7599 (N_7599,N_7427,N_7312);
nand U7600 (N_7600,N_7389,N_7313);
xnor U7601 (N_7601,N_7297,N_7497);
nor U7602 (N_7602,N_7479,N_7332);
and U7603 (N_7603,N_7476,N_7398);
xor U7604 (N_7604,N_7466,N_7367);
nor U7605 (N_7605,N_7498,N_7380);
xor U7606 (N_7606,N_7275,N_7480);
nand U7607 (N_7607,N_7370,N_7453);
or U7608 (N_7608,N_7256,N_7344);
xor U7609 (N_7609,N_7429,N_7457);
nor U7610 (N_7610,N_7306,N_7425);
and U7611 (N_7611,N_7415,N_7403);
nor U7612 (N_7612,N_7394,N_7280);
xor U7613 (N_7613,N_7335,N_7382);
nor U7614 (N_7614,N_7368,N_7397);
or U7615 (N_7615,N_7283,N_7390);
nor U7616 (N_7616,N_7414,N_7450);
and U7617 (N_7617,N_7408,N_7470);
nor U7618 (N_7618,N_7434,N_7406);
xor U7619 (N_7619,N_7289,N_7454);
and U7620 (N_7620,N_7385,N_7285);
or U7621 (N_7621,N_7351,N_7359);
xor U7622 (N_7622,N_7412,N_7378);
or U7623 (N_7623,N_7489,N_7304);
nand U7624 (N_7624,N_7375,N_7420);
nand U7625 (N_7625,N_7270,N_7473);
nor U7626 (N_7626,N_7471,N_7360);
and U7627 (N_7627,N_7362,N_7440);
and U7628 (N_7628,N_7264,N_7332);
xor U7629 (N_7629,N_7496,N_7308);
and U7630 (N_7630,N_7272,N_7342);
nor U7631 (N_7631,N_7280,N_7365);
xor U7632 (N_7632,N_7466,N_7492);
xnor U7633 (N_7633,N_7403,N_7373);
nand U7634 (N_7634,N_7257,N_7264);
nand U7635 (N_7635,N_7407,N_7369);
or U7636 (N_7636,N_7472,N_7468);
nand U7637 (N_7637,N_7276,N_7252);
nor U7638 (N_7638,N_7423,N_7428);
and U7639 (N_7639,N_7455,N_7462);
xnor U7640 (N_7640,N_7297,N_7419);
xnor U7641 (N_7641,N_7401,N_7350);
nand U7642 (N_7642,N_7417,N_7374);
nor U7643 (N_7643,N_7481,N_7441);
and U7644 (N_7644,N_7407,N_7289);
nor U7645 (N_7645,N_7397,N_7296);
nand U7646 (N_7646,N_7408,N_7466);
nor U7647 (N_7647,N_7418,N_7357);
and U7648 (N_7648,N_7437,N_7315);
xnor U7649 (N_7649,N_7491,N_7378);
nand U7650 (N_7650,N_7265,N_7318);
and U7651 (N_7651,N_7464,N_7316);
or U7652 (N_7652,N_7299,N_7458);
or U7653 (N_7653,N_7312,N_7392);
nand U7654 (N_7654,N_7268,N_7251);
xor U7655 (N_7655,N_7421,N_7278);
and U7656 (N_7656,N_7448,N_7329);
and U7657 (N_7657,N_7463,N_7343);
nand U7658 (N_7658,N_7492,N_7352);
xor U7659 (N_7659,N_7284,N_7305);
nand U7660 (N_7660,N_7348,N_7312);
xor U7661 (N_7661,N_7497,N_7411);
and U7662 (N_7662,N_7474,N_7421);
nor U7663 (N_7663,N_7309,N_7427);
nor U7664 (N_7664,N_7477,N_7429);
nand U7665 (N_7665,N_7395,N_7333);
nor U7666 (N_7666,N_7313,N_7369);
xnor U7667 (N_7667,N_7473,N_7256);
and U7668 (N_7668,N_7255,N_7312);
nand U7669 (N_7669,N_7455,N_7277);
nand U7670 (N_7670,N_7263,N_7299);
nand U7671 (N_7671,N_7271,N_7444);
or U7672 (N_7672,N_7405,N_7481);
nor U7673 (N_7673,N_7444,N_7381);
nand U7674 (N_7674,N_7301,N_7330);
nand U7675 (N_7675,N_7349,N_7411);
nor U7676 (N_7676,N_7255,N_7314);
nor U7677 (N_7677,N_7276,N_7480);
nand U7678 (N_7678,N_7297,N_7421);
xnor U7679 (N_7679,N_7299,N_7440);
and U7680 (N_7680,N_7327,N_7431);
xor U7681 (N_7681,N_7289,N_7394);
and U7682 (N_7682,N_7396,N_7300);
xnor U7683 (N_7683,N_7264,N_7489);
nand U7684 (N_7684,N_7419,N_7333);
xnor U7685 (N_7685,N_7329,N_7461);
and U7686 (N_7686,N_7274,N_7487);
or U7687 (N_7687,N_7446,N_7278);
nor U7688 (N_7688,N_7475,N_7469);
xnor U7689 (N_7689,N_7323,N_7391);
or U7690 (N_7690,N_7258,N_7369);
and U7691 (N_7691,N_7260,N_7364);
nand U7692 (N_7692,N_7441,N_7378);
xor U7693 (N_7693,N_7276,N_7322);
nor U7694 (N_7694,N_7421,N_7250);
or U7695 (N_7695,N_7260,N_7468);
or U7696 (N_7696,N_7356,N_7452);
and U7697 (N_7697,N_7278,N_7401);
or U7698 (N_7698,N_7303,N_7447);
nand U7699 (N_7699,N_7427,N_7319);
nand U7700 (N_7700,N_7386,N_7331);
or U7701 (N_7701,N_7299,N_7309);
nand U7702 (N_7702,N_7375,N_7493);
xor U7703 (N_7703,N_7432,N_7262);
and U7704 (N_7704,N_7438,N_7466);
or U7705 (N_7705,N_7397,N_7335);
xor U7706 (N_7706,N_7307,N_7277);
nand U7707 (N_7707,N_7469,N_7476);
and U7708 (N_7708,N_7280,N_7291);
nand U7709 (N_7709,N_7279,N_7490);
xor U7710 (N_7710,N_7334,N_7331);
xnor U7711 (N_7711,N_7482,N_7265);
xnor U7712 (N_7712,N_7362,N_7467);
nor U7713 (N_7713,N_7270,N_7263);
and U7714 (N_7714,N_7400,N_7314);
nand U7715 (N_7715,N_7415,N_7333);
and U7716 (N_7716,N_7262,N_7346);
and U7717 (N_7717,N_7379,N_7466);
nor U7718 (N_7718,N_7489,N_7434);
nor U7719 (N_7719,N_7299,N_7498);
and U7720 (N_7720,N_7299,N_7300);
or U7721 (N_7721,N_7344,N_7477);
nor U7722 (N_7722,N_7453,N_7473);
xor U7723 (N_7723,N_7351,N_7445);
nor U7724 (N_7724,N_7380,N_7276);
nand U7725 (N_7725,N_7357,N_7390);
nand U7726 (N_7726,N_7451,N_7384);
or U7727 (N_7727,N_7381,N_7454);
and U7728 (N_7728,N_7290,N_7435);
xor U7729 (N_7729,N_7251,N_7299);
xor U7730 (N_7730,N_7490,N_7257);
nand U7731 (N_7731,N_7474,N_7306);
xor U7732 (N_7732,N_7348,N_7309);
nand U7733 (N_7733,N_7374,N_7276);
and U7734 (N_7734,N_7448,N_7433);
xnor U7735 (N_7735,N_7478,N_7364);
xnor U7736 (N_7736,N_7292,N_7322);
or U7737 (N_7737,N_7271,N_7336);
nand U7738 (N_7738,N_7327,N_7445);
or U7739 (N_7739,N_7307,N_7292);
nor U7740 (N_7740,N_7479,N_7314);
and U7741 (N_7741,N_7467,N_7253);
xor U7742 (N_7742,N_7273,N_7323);
xnor U7743 (N_7743,N_7363,N_7298);
nand U7744 (N_7744,N_7420,N_7401);
or U7745 (N_7745,N_7423,N_7255);
nor U7746 (N_7746,N_7391,N_7258);
or U7747 (N_7747,N_7495,N_7408);
nor U7748 (N_7748,N_7300,N_7328);
xor U7749 (N_7749,N_7413,N_7467);
xnor U7750 (N_7750,N_7709,N_7734);
or U7751 (N_7751,N_7612,N_7701);
and U7752 (N_7752,N_7685,N_7746);
xor U7753 (N_7753,N_7660,N_7652);
nor U7754 (N_7754,N_7742,N_7663);
and U7755 (N_7755,N_7716,N_7538);
xnor U7756 (N_7756,N_7715,N_7659);
and U7757 (N_7757,N_7729,N_7597);
nand U7758 (N_7758,N_7618,N_7605);
nand U7759 (N_7759,N_7599,N_7667);
xor U7760 (N_7760,N_7521,N_7523);
nor U7761 (N_7761,N_7625,N_7519);
and U7762 (N_7762,N_7745,N_7693);
nand U7763 (N_7763,N_7551,N_7526);
nand U7764 (N_7764,N_7589,N_7641);
nand U7765 (N_7765,N_7545,N_7524);
nor U7766 (N_7766,N_7689,N_7723);
nand U7767 (N_7767,N_7520,N_7593);
xnor U7768 (N_7768,N_7635,N_7570);
nor U7769 (N_7769,N_7596,N_7602);
or U7770 (N_7770,N_7557,N_7740);
and U7771 (N_7771,N_7555,N_7670);
nor U7772 (N_7772,N_7540,N_7686);
or U7773 (N_7773,N_7529,N_7654);
or U7774 (N_7774,N_7661,N_7512);
xor U7775 (N_7775,N_7518,N_7676);
or U7776 (N_7776,N_7731,N_7564);
nor U7777 (N_7777,N_7682,N_7724);
nand U7778 (N_7778,N_7633,N_7665);
and U7779 (N_7779,N_7580,N_7616);
and U7780 (N_7780,N_7515,N_7705);
and U7781 (N_7781,N_7629,N_7717);
nand U7782 (N_7782,N_7584,N_7531);
and U7783 (N_7783,N_7643,N_7547);
or U7784 (N_7784,N_7714,N_7588);
or U7785 (N_7785,N_7636,N_7650);
xnor U7786 (N_7786,N_7696,N_7614);
nand U7787 (N_7787,N_7658,N_7749);
and U7788 (N_7788,N_7514,N_7632);
nand U7789 (N_7789,N_7510,N_7536);
or U7790 (N_7790,N_7702,N_7563);
or U7791 (N_7791,N_7725,N_7624);
xor U7792 (N_7792,N_7528,N_7527);
nand U7793 (N_7793,N_7592,N_7577);
nand U7794 (N_7794,N_7594,N_7657);
and U7795 (N_7795,N_7543,N_7720);
or U7796 (N_7796,N_7626,N_7640);
and U7797 (N_7797,N_7506,N_7573);
xnor U7798 (N_7798,N_7671,N_7733);
or U7799 (N_7799,N_7735,N_7642);
nand U7800 (N_7800,N_7673,N_7628);
and U7801 (N_7801,N_7569,N_7645);
nor U7802 (N_7802,N_7620,N_7732);
or U7803 (N_7803,N_7544,N_7613);
nor U7804 (N_7804,N_7537,N_7741);
or U7805 (N_7805,N_7722,N_7743);
and U7806 (N_7806,N_7662,N_7503);
xnor U7807 (N_7807,N_7611,N_7559);
or U7808 (N_7808,N_7617,N_7678);
nor U7809 (N_7809,N_7598,N_7508);
or U7810 (N_7810,N_7517,N_7530);
xnor U7811 (N_7811,N_7627,N_7695);
and U7812 (N_7812,N_7585,N_7623);
nor U7813 (N_7813,N_7542,N_7560);
nand U7814 (N_7814,N_7718,N_7595);
nand U7815 (N_7815,N_7558,N_7567);
nor U7816 (N_7816,N_7549,N_7600);
xnor U7817 (N_7817,N_7677,N_7691);
nor U7818 (N_7818,N_7622,N_7728);
or U7819 (N_7819,N_7601,N_7698);
nand U7820 (N_7820,N_7699,N_7694);
xor U7821 (N_7821,N_7575,N_7681);
and U7822 (N_7822,N_7513,N_7587);
or U7823 (N_7823,N_7744,N_7552);
nand U7824 (N_7824,N_7683,N_7648);
nand U7825 (N_7825,N_7738,N_7501);
xnor U7826 (N_7826,N_7631,N_7535);
and U7827 (N_7827,N_7668,N_7591);
and U7828 (N_7828,N_7649,N_7730);
nand U7829 (N_7829,N_7692,N_7646);
xor U7830 (N_7830,N_7562,N_7644);
and U7831 (N_7831,N_7609,N_7516);
or U7832 (N_7832,N_7727,N_7711);
nand U7833 (N_7833,N_7606,N_7687);
and U7834 (N_7834,N_7697,N_7556);
or U7835 (N_7835,N_7736,N_7619);
and U7836 (N_7836,N_7533,N_7706);
xnor U7837 (N_7837,N_7532,N_7553);
nor U7838 (N_7838,N_7704,N_7656);
and U7839 (N_7839,N_7726,N_7546);
and U7840 (N_7840,N_7747,N_7548);
and U7841 (N_7841,N_7615,N_7621);
xor U7842 (N_7842,N_7653,N_7688);
nor U7843 (N_7843,N_7630,N_7737);
or U7844 (N_7844,N_7578,N_7566);
xor U7845 (N_7845,N_7590,N_7690);
and U7846 (N_7846,N_7541,N_7582);
and U7847 (N_7847,N_7581,N_7586);
nor U7848 (N_7848,N_7707,N_7708);
nor U7849 (N_7849,N_7739,N_7509);
nor U7850 (N_7850,N_7669,N_7554);
nand U7851 (N_7851,N_7525,N_7607);
xnor U7852 (N_7852,N_7684,N_7505);
nor U7853 (N_7853,N_7672,N_7583);
nand U7854 (N_7854,N_7713,N_7748);
nand U7855 (N_7855,N_7664,N_7550);
or U7856 (N_7856,N_7712,N_7647);
nand U7857 (N_7857,N_7561,N_7638);
or U7858 (N_7858,N_7655,N_7507);
nor U7859 (N_7859,N_7680,N_7666);
nor U7860 (N_7860,N_7568,N_7700);
nand U7861 (N_7861,N_7679,N_7710);
or U7862 (N_7862,N_7571,N_7604);
or U7863 (N_7863,N_7539,N_7703);
and U7864 (N_7864,N_7610,N_7576);
nand U7865 (N_7865,N_7500,N_7574);
or U7866 (N_7866,N_7603,N_7674);
nor U7867 (N_7867,N_7634,N_7511);
and U7868 (N_7868,N_7719,N_7721);
nand U7869 (N_7869,N_7565,N_7675);
and U7870 (N_7870,N_7651,N_7639);
nand U7871 (N_7871,N_7608,N_7637);
and U7872 (N_7872,N_7534,N_7504);
nor U7873 (N_7873,N_7572,N_7522);
or U7874 (N_7874,N_7579,N_7502);
or U7875 (N_7875,N_7525,N_7540);
or U7876 (N_7876,N_7636,N_7509);
and U7877 (N_7877,N_7579,N_7626);
xnor U7878 (N_7878,N_7551,N_7518);
and U7879 (N_7879,N_7669,N_7507);
nand U7880 (N_7880,N_7603,N_7671);
or U7881 (N_7881,N_7650,N_7621);
nor U7882 (N_7882,N_7698,N_7625);
or U7883 (N_7883,N_7541,N_7599);
or U7884 (N_7884,N_7719,N_7516);
xnor U7885 (N_7885,N_7658,N_7613);
or U7886 (N_7886,N_7604,N_7676);
and U7887 (N_7887,N_7679,N_7736);
and U7888 (N_7888,N_7593,N_7568);
xnor U7889 (N_7889,N_7620,N_7705);
nor U7890 (N_7890,N_7507,N_7653);
xnor U7891 (N_7891,N_7666,N_7603);
nor U7892 (N_7892,N_7524,N_7584);
nor U7893 (N_7893,N_7614,N_7577);
or U7894 (N_7894,N_7743,N_7588);
nand U7895 (N_7895,N_7596,N_7694);
nor U7896 (N_7896,N_7692,N_7706);
or U7897 (N_7897,N_7714,N_7581);
and U7898 (N_7898,N_7712,N_7516);
nor U7899 (N_7899,N_7554,N_7610);
nand U7900 (N_7900,N_7669,N_7728);
nand U7901 (N_7901,N_7747,N_7685);
nand U7902 (N_7902,N_7512,N_7599);
or U7903 (N_7903,N_7665,N_7546);
xor U7904 (N_7904,N_7665,N_7632);
xnor U7905 (N_7905,N_7606,N_7546);
or U7906 (N_7906,N_7526,N_7701);
and U7907 (N_7907,N_7545,N_7705);
nor U7908 (N_7908,N_7736,N_7512);
or U7909 (N_7909,N_7570,N_7748);
xnor U7910 (N_7910,N_7625,N_7689);
nor U7911 (N_7911,N_7577,N_7685);
xor U7912 (N_7912,N_7512,N_7728);
nor U7913 (N_7913,N_7509,N_7622);
nand U7914 (N_7914,N_7737,N_7748);
xor U7915 (N_7915,N_7691,N_7745);
or U7916 (N_7916,N_7610,N_7627);
and U7917 (N_7917,N_7510,N_7731);
and U7918 (N_7918,N_7514,N_7668);
nor U7919 (N_7919,N_7687,N_7587);
or U7920 (N_7920,N_7607,N_7709);
xor U7921 (N_7921,N_7618,N_7540);
or U7922 (N_7922,N_7639,N_7551);
xnor U7923 (N_7923,N_7525,N_7558);
and U7924 (N_7924,N_7738,N_7631);
nand U7925 (N_7925,N_7622,N_7652);
nand U7926 (N_7926,N_7711,N_7530);
and U7927 (N_7927,N_7526,N_7672);
xor U7928 (N_7928,N_7648,N_7669);
or U7929 (N_7929,N_7575,N_7592);
or U7930 (N_7930,N_7651,N_7595);
xor U7931 (N_7931,N_7580,N_7561);
nor U7932 (N_7932,N_7660,N_7524);
xor U7933 (N_7933,N_7575,N_7503);
xor U7934 (N_7934,N_7723,N_7639);
xnor U7935 (N_7935,N_7618,N_7648);
nand U7936 (N_7936,N_7508,N_7561);
nand U7937 (N_7937,N_7573,N_7695);
or U7938 (N_7938,N_7745,N_7550);
xnor U7939 (N_7939,N_7568,N_7613);
nor U7940 (N_7940,N_7650,N_7692);
or U7941 (N_7941,N_7743,N_7715);
nand U7942 (N_7942,N_7747,N_7686);
and U7943 (N_7943,N_7601,N_7749);
nand U7944 (N_7944,N_7568,N_7543);
or U7945 (N_7945,N_7540,N_7701);
and U7946 (N_7946,N_7622,N_7695);
nor U7947 (N_7947,N_7665,N_7513);
nor U7948 (N_7948,N_7661,N_7674);
nor U7949 (N_7949,N_7693,N_7661);
and U7950 (N_7950,N_7602,N_7598);
and U7951 (N_7951,N_7612,N_7603);
nor U7952 (N_7952,N_7564,N_7554);
and U7953 (N_7953,N_7503,N_7602);
and U7954 (N_7954,N_7613,N_7701);
nand U7955 (N_7955,N_7643,N_7528);
or U7956 (N_7956,N_7579,N_7538);
and U7957 (N_7957,N_7641,N_7567);
or U7958 (N_7958,N_7544,N_7721);
or U7959 (N_7959,N_7731,N_7588);
nor U7960 (N_7960,N_7689,N_7690);
or U7961 (N_7961,N_7529,N_7660);
xor U7962 (N_7962,N_7515,N_7514);
nand U7963 (N_7963,N_7583,N_7641);
xor U7964 (N_7964,N_7736,N_7606);
and U7965 (N_7965,N_7548,N_7620);
nor U7966 (N_7966,N_7684,N_7530);
nor U7967 (N_7967,N_7527,N_7529);
or U7968 (N_7968,N_7639,N_7629);
and U7969 (N_7969,N_7610,N_7670);
or U7970 (N_7970,N_7683,N_7550);
nand U7971 (N_7971,N_7729,N_7633);
xor U7972 (N_7972,N_7591,N_7664);
and U7973 (N_7973,N_7680,N_7749);
or U7974 (N_7974,N_7558,N_7529);
nand U7975 (N_7975,N_7589,N_7719);
nand U7976 (N_7976,N_7689,N_7704);
nor U7977 (N_7977,N_7521,N_7511);
nand U7978 (N_7978,N_7504,N_7700);
xor U7979 (N_7979,N_7682,N_7606);
nor U7980 (N_7980,N_7691,N_7627);
xnor U7981 (N_7981,N_7506,N_7684);
nand U7982 (N_7982,N_7520,N_7744);
or U7983 (N_7983,N_7535,N_7532);
xor U7984 (N_7984,N_7679,N_7558);
xor U7985 (N_7985,N_7510,N_7732);
and U7986 (N_7986,N_7744,N_7506);
nor U7987 (N_7987,N_7730,N_7742);
xnor U7988 (N_7988,N_7559,N_7514);
nor U7989 (N_7989,N_7740,N_7505);
nand U7990 (N_7990,N_7511,N_7516);
xor U7991 (N_7991,N_7590,N_7639);
nand U7992 (N_7992,N_7619,N_7616);
nand U7993 (N_7993,N_7741,N_7681);
nand U7994 (N_7994,N_7727,N_7616);
nor U7995 (N_7995,N_7516,N_7549);
nand U7996 (N_7996,N_7535,N_7618);
nor U7997 (N_7997,N_7585,N_7650);
and U7998 (N_7998,N_7585,N_7669);
xor U7999 (N_7999,N_7659,N_7692);
nor U8000 (N_8000,N_7753,N_7961);
nor U8001 (N_8001,N_7801,N_7885);
nor U8002 (N_8002,N_7756,N_7758);
nor U8003 (N_8003,N_7828,N_7760);
nand U8004 (N_8004,N_7965,N_7912);
xor U8005 (N_8005,N_7779,N_7794);
nand U8006 (N_8006,N_7963,N_7977);
xor U8007 (N_8007,N_7791,N_7861);
nand U8008 (N_8008,N_7800,N_7902);
nand U8009 (N_8009,N_7838,N_7754);
nand U8010 (N_8010,N_7813,N_7875);
or U8011 (N_8011,N_7859,N_7968);
nand U8012 (N_8012,N_7825,N_7814);
and U8013 (N_8013,N_7880,N_7820);
nand U8014 (N_8014,N_7877,N_7909);
nand U8015 (N_8015,N_7763,N_7768);
or U8016 (N_8016,N_7958,N_7911);
or U8017 (N_8017,N_7752,N_7987);
nand U8018 (N_8018,N_7864,N_7766);
and U8019 (N_8019,N_7849,N_7933);
nand U8020 (N_8020,N_7939,N_7765);
and U8021 (N_8021,N_7901,N_7917);
or U8022 (N_8022,N_7954,N_7767);
nand U8023 (N_8023,N_7974,N_7918);
nand U8024 (N_8024,N_7850,N_7876);
and U8025 (N_8025,N_7986,N_7793);
nand U8026 (N_8026,N_7936,N_7955);
and U8027 (N_8027,N_7797,N_7834);
or U8028 (N_8028,N_7915,N_7823);
nand U8029 (N_8029,N_7950,N_7996);
and U8030 (N_8030,N_7809,N_7985);
and U8031 (N_8031,N_7998,N_7982);
nand U8032 (N_8032,N_7817,N_7951);
or U8033 (N_8033,N_7935,N_7931);
nor U8034 (N_8034,N_7962,N_7932);
nand U8035 (N_8035,N_7926,N_7827);
nand U8036 (N_8036,N_7837,N_7870);
or U8037 (N_8037,N_7947,N_7882);
or U8038 (N_8038,N_7881,N_7810);
or U8039 (N_8039,N_7841,N_7854);
xnor U8040 (N_8040,N_7789,N_7921);
nand U8041 (N_8041,N_7908,N_7769);
and U8042 (N_8042,N_7920,N_7957);
nor U8043 (N_8043,N_7816,N_7824);
and U8044 (N_8044,N_7750,N_7896);
and U8045 (N_8045,N_7929,N_7862);
nor U8046 (N_8046,N_7970,N_7860);
nand U8047 (N_8047,N_7845,N_7757);
or U8048 (N_8048,N_7840,N_7784);
xnor U8049 (N_8049,N_7821,N_7806);
xor U8050 (N_8050,N_7966,N_7833);
xnor U8051 (N_8051,N_7983,N_7778);
nor U8052 (N_8052,N_7969,N_7780);
and U8053 (N_8053,N_7964,N_7761);
or U8054 (N_8054,N_7960,N_7853);
nand U8055 (N_8055,N_7990,N_7873);
xnor U8056 (N_8056,N_7847,N_7904);
nand U8057 (N_8057,N_7907,N_7952);
xor U8058 (N_8058,N_7762,N_7826);
and U8059 (N_8059,N_7925,N_7771);
or U8060 (N_8060,N_7792,N_7916);
nand U8061 (N_8061,N_7946,N_7796);
xnor U8062 (N_8062,N_7997,N_7973);
or U8063 (N_8063,N_7900,N_7804);
and U8064 (N_8064,N_7895,N_7874);
nand U8065 (N_8065,N_7790,N_7959);
xor U8066 (N_8066,N_7891,N_7795);
xnor U8067 (N_8067,N_7914,N_7991);
nand U8068 (N_8068,N_7910,N_7811);
nor U8069 (N_8069,N_7822,N_7787);
xor U8070 (N_8070,N_7759,N_7906);
nor U8071 (N_8071,N_7905,N_7989);
or U8072 (N_8072,N_7812,N_7981);
and U8073 (N_8073,N_7843,N_7869);
xor U8074 (N_8074,N_7818,N_7781);
xnor U8075 (N_8075,N_7903,N_7856);
nand U8076 (N_8076,N_7819,N_7770);
and U8077 (N_8077,N_7894,N_7831);
xnor U8078 (N_8078,N_7956,N_7949);
and U8079 (N_8079,N_7978,N_7993);
nor U8080 (N_8080,N_7971,N_7967);
nand U8081 (N_8081,N_7937,N_7898);
or U8082 (N_8082,N_7930,N_7865);
xnor U8083 (N_8083,N_7774,N_7887);
nor U8084 (N_8084,N_7830,N_7984);
and U8085 (N_8085,N_7858,N_7808);
or U8086 (N_8086,N_7888,N_7934);
or U8087 (N_8087,N_7940,N_7923);
nand U8088 (N_8088,N_7892,N_7976);
nand U8089 (N_8089,N_7863,N_7884);
nor U8090 (N_8090,N_7785,N_7879);
and U8091 (N_8091,N_7835,N_7979);
or U8092 (N_8092,N_7868,N_7913);
and U8093 (N_8093,N_7871,N_7803);
and U8094 (N_8094,N_7815,N_7855);
xnor U8095 (N_8095,N_7878,N_7846);
and U8096 (N_8096,N_7943,N_7953);
or U8097 (N_8097,N_7786,N_7999);
nand U8098 (N_8098,N_7805,N_7751);
and U8099 (N_8099,N_7848,N_7948);
and U8100 (N_8100,N_7941,N_7839);
nor U8101 (N_8101,N_7852,N_7944);
and U8102 (N_8102,N_7938,N_7844);
nand U8103 (N_8103,N_7857,N_7886);
and U8104 (N_8104,N_7802,N_7783);
and U8105 (N_8105,N_7807,N_7872);
xor U8106 (N_8106,N_7788,N_7893);
or U8107 (N_8107,N_7992,N_7897);
nor U8108 (N_8108,N_7777,N_7975);
or U8109 (N_8109,N_7773,N_7832);
nand U8110 (N_8110,N_7782,N_7772);
or U8111 (N_8111,N_7883,N_7988);
nor U8112 (N_8112,N_7776,N_7866);
nand U8113 (N_8113,N_7799,N_7945);
nand U8114 (N_8114,N_7899,N_7972);
nor U8115 (N_8115,N_7994,N_7851);
xnor U8116 (N_8116,N_7755,N_7836);
nand U8117 (N_8117,N_7995,N_7942);
and U8118 (N_8118,N_7775,N_7890);
nor U8119 (N_8119,N_7829,N_7927);
and U8120 (N_8120,N_7889,N_7922);
and U8121 (N_8121,N_7919,N_7764);
xor U8122 (N_8122,N_7867,N_7980);
or U8123 (N_8123,N_7798,N_7924);
or U8124 (N_8124,N_7928,N_7842);
nand U8125 (N_8125,N_7847,N_7757);
xnor U8126 (N_8126,N_7830,N_7879);
xnor U8127 (N_8127,N_7889,N_7957);
and U8128 (N_8128,N_7998,N_7851);
and U8129 (N_8129,N_7826,N_7854);
nor U8130 (N_8130,N_7756,N_7812);
nand U8131 (N_8131,N_7864,N_7778);
xor U8132 (N_8132,N_7878,N_7896);
and U8133 (N_8133,N_7864,N_7825);
or U8134 (N_8134,N_7954,N_7816);
nand U8135 (N_8135,N_7859,N_7996);
nand U8136 (N_8136,N_7766,N_7859);
xor U8137 (N_8137,N_7970,N_7947);
xor U8138 (N_8138,N_7860,N_7753);
nor U8139 (N_8139,N_7999,N_7858);
or U8140 (N_8140,N_7987,N_7972);
nor U8141 (N_8141,N_7817,N_7906);
nand U8142 (N_8142,N_7750,N_7977);
xor U8143 (N_8143,N_7776,N_7933);
and U8144 (N_8144,N_7866,N_7833);
or U8145 (N_8145,N_7772,N_7867);
or U8146 (N_8146,N_7993,N_7906);
and U8147 (N_8147,N_7947,N_7949);
or U8148 (N_8148,N_7994,N_7910);
or U8149 (N_8149,N_7912,N_7757);
xor U8150 (N_8150,N_7875,N_7952);
or U8151 (N_8151,N_7913,N_7912);
or U8152 (N_8152,N_7760,N_7806);
nor U8153 (N_8153,N_7963,N_7809);
nor U8154 (N_8154,N_7989,N_7840);
xnor U8155 (N_8155,N_7762,N_7968);
xor U8156 (N_8156,N_7787,N_7812);
or U8157 (N_8157,N_7850,N_7881);
nor U8158 (N_8158,N_7864,N_7937);
xnor U8159 (N_8159,N_7815,N_7980);
nor U8160 (N_8160,N_7987,N_7893);
and U8161 (N_8161,N_7949,N_7778);
xor U8162 (N_8162,N_7948,N_7796);
or U8163 (N_8163,N_7894,N_7968);
nor U8164 (N_8164,N_7869,N_7963);
nand U8165 (N_8165,N_7908,N_7786);
nand U8166 (N_8166,N_7955,N_7999);
or U8167 (N_8167,N_7942,N_7785);
or U8168 (N_8168,N_7973,N_7805);
or U8169 (N_8169,N_7926,N_7909);
xor U8170 (N_8170,N_7885,N_7998);
xnor U8171 (N_8171,N_7873,N_7959);
nor U8172 (N_8172,N_7902,N_7943);
and U8173 (N_8173,N_7787,N_7883);
xnor U8174 (N_8174,N_7909,N_7775);
or U8175 (N_8175,N_7961,N_7969);
and U8176 (N_8176,N_7811,N_7791);
nor U8177 (N_8177,N_7751,N_7852);
or U8178 (N_8178,N_7758,N_7910);
or U8179 (N_8179,N_7809,N_7965);
nor U8180 (N_8180,N_7892,N_7942);
or U8181 (N_8181,N_7860,N_7822);
nand U8182 (N_8182,N_7974,N_7987);
nand U8183 (N_8183,N_7764,N_7806);
or U8184 (N_8184,N_7890,N_7974);
or U8185 (N_8185,N_7806,N_7796);
nand U8186 (N_8186,N_7981,N_7999);
nand U8187 (N_8187,N_7974,N_7915);
or U8188 (N_8188,N_7944,N_7883);
and U8189 (N_8189,N_7968,N_7917);
nor U8190 (N_8190,N_7816,N_7841);
and U8191 (N_8191,N_7997,N_7802);
nor U8192 (N_8192,N_7997,N_7961);
nand U8193 (N_8193,N_7871,N_7926);
and U8194 (N_8194,N_7825,N_7972);
xor U8195 (N_8195,N_7758,N_7823);
xor U8196 (N_8196,N_7776,N_7837);
and U8197 (N_8197,N_7858,N_7860);
and U8198 (N_8198,N_7939,N_7884);
xor U8199 (N_8199,N_7828,N_7920);
and U8200 (N_8200,N_7794,N_7963);
and U8201 (N_8201,N_7913,N_7818);
nand U8202 (N_8202,N_7774,N_7805);
xnor U8203 (N_8203,N_7894,N_7807);
or U8204 (N_8204,N_7820,N_7993);
nor U8205 (N_8205,N_7874,N_7980);
xor U8206 (N_8206,N_7923,N_7758);
xor U8207 (N_8207,N_7921,N_7956);
and U8208 (N_8208,N_7897,N_7990);
nand U8209 (N_8209,N_7923,N_7792);
xnor U8210 (N_8210,N_7967,N_7980);
xor U8211 (N_8211,N_7859,N_7765);
or U8212 (N_8212,N_7991,N_7767);
xnor U8213 (N_8213,N_7856,N_7904);
nand U8214 (N_8214,N_7782,N_7760);
and U8215 (N_8215,N_7966,N_7947);
nand U8216 (N_8216,N_7756,N_7778);
or U8217 (N_8217,N_7833,N_7976);
xnor U8218 (N_8218,N_7820,N_7767);
nor U8219 (N_8219,N_7768,N_7954);
nand U8220 (N_8220,N_7777,N_7993);
nor U8221 (N_8221,N_7969,N_7860);
nor U8222 (N_8222,N_7933,N_7923);
nor U8223 (N_8223,N_7970,N_7820);
or U8224 (N_8224,N_7896,N_7897);
nand U8225 (N_8225,N_7784,N_7977);
and U8226 (N_8226,N_7918,N_7935);
xor U8227 (N_8227,N_7751,N_7918);
nor U8228 (N_8228,N_7817,N_7839);
and U8229 (N_8229,N_7960,N_7834);
and U8230 (N_8230,N_7800,N_7997);
xor U8231 (N_8231,N_7966,N_7848);
nand U8232 (N_8232,N_7957,N_7941);
nand U8233 (N_8233,N_7794,N_7822);
nor U8234 (N_8234,N_7870,N_7926);
and U8235 (N_8235,N_7859,N_7869);
or U8236 (N_8236,N_7942,N_7809);
or U8237 (N_8237,N_7864,N_7906);
xor U8238 (N_8238,N_7798,N_7838);
nand U8239 (N_8239,N_7898,N_7884);
or U8240 (N_8240,N_7801,N_7835);
xor U8241 (N_8241,N_7892,N_7805);
nor U8242 (N_8242,N_7956,N_7751);
or U8243 (N_8243,N_7838,N_7967);
nand U8244 (N_8244,N_7779,N_7869);
nor U8245 (N_8245,N_7780,N_7952);
and U8246 (N_8246,N_7878,N_7774);
and U8247 (N_8247,N_7892,N_7863);
nor U8248 (N_8248,N_7755,N_7982);
nand U8249 (N_8249,N_7811,N_7980);
or U8250 (N_8250,N_8007,N_8118);
nand U8251 (N_8251,N_8194,N_8162);
and U8252 (N_8252,N_8011,N_8179);
nand U8253 (N_8253,N_8019,N_8200);
or U8254 (N_8254,N_8097,N_8117);
or U8255 (N_8255,N_8204,N_8103);
nor U8256 (N_8256,N_8074,N_8091);
nand U8257 (N_8257,N_8021,N_8025);
nor U8258 (N_8258,N_8243,N_8207);
xnor U8259 (N_8259,N_8053,N_8170);
nor U8260 (N_8260,N_8056,N_8107);
and U8261 (N_8261,N_8130,N_8211);
nor U8262 (N_8262,N_8168,N_8049);
or U8263 (N_8263,N_8101,N_8045);
nor U8264 (N_8264,N_8147,N_8212);
or U8265 (N_8265,N_8129,N_8219);
or U8266 (N_8266,N_8041,N_8137);
or U8267 (N_8267,N_8163,N_8171);
nand U8268 (N_8268,N_8023,N_8027);
or U8269 (N_8269,N_8038,N_8225);
xnor U8270 (N_8270,N_8010,N_8191);
xor U8271 (N_8271,N_8052,N_8017);
or U8272 (N_8272,N_8150,N_8061);
or U8273 (N_8273,N_8132,N_8001);
nand U8274 (N_8274,N_8154,N_8223);
xor U8275 (N_8275,N_8085,N_8188);
nand U8276 (N_8276,N_8002,N_8175);
nand U8277 (N_8277,N_8192,N_8231);
nand U8278 (N_8278,N_8151,N_8140);
nand U8279 (N_8279,N_8184,N_8218);
nor U8280 (N_8280,N_8088,N_8022);
nand U8281 (N_8281,N_8159,N_8018);
and U8282 (N_8282,N_8115,N_8189);
nor U8283 (N_8283,N_8051,N_8127);
nor U8284 (N_8284,N_8028,N_8148);
nand U8285 (N_8285,N_8063,N_8165);
nand U8286 (N_8286,N_8145,N_8226);
or U8287 (N_8287,N_8201,N_8213);
nand U8288 (N_8288,N_8004,N_8076);
xor U8289 (N_8289,N_8238,N_8026);
xnor U8290 (N_8290,N_8065,N_8020);
and U8291 (N_8291,N_8072,N_8032);
xnor U8292 (N_8292,N_8105,N_8146);
and U8293 (N_8293,N_8141,N_8067);
and U8294 (N_8294,N_8234,N_8214);
nand U8295 (N_8295,N_8157,N_8087);
xnor U8296 (N_8296,N_8081,N_8120);
xnor U8297 (N_8297,N_8128,N_8078);
and U8298 (N_8298,N_8060,N_8003);
nand U8299 (N_8299,N_8153,N_8094);
nor U8300 (N_8300,N_8031,N_8245);
xnor U8301 (N_8301,N_8066,N_8124);
nor U8302 (N_8302,N_8138,N_8116);
or U8303 (N_8303,N_8182,N_8244);
xor U8304 (N_8304,N_8156,N_8142);
nor U8305 (N_8305,N_8177,N_8106);
and U8306 (N_8306,N_8195,N_8050);
or U8307 (N_8307,N_8108,N_8073);
nor U8308 (N_8308,N_8064,N_8099);
nand U8309 (N_8309,N_8100,N_8048);
or U8310 (N_8310,N_8178,N_8209);
and U8311 (N_8311,N_8241,N_8233);
nand U8312 (N_8312,N_8172,N_8229);
nand U8313 (N_8313,N_8126,N_8113);
nor U8314 (N_8314,N_8196,N_8055);
nor U8315 (N_8315,N_8034,N_8139);
nand U8316 (N_8316,N_8110,N_8033);
xnor U8317 (N_8317,N_8143,N_8059);
or U8318 (N_8318,N_8198,N_8062);
or U8319 (N_8319,N_8000,N_8239);
nand U8320 (N_8320,N_8144,N_8246);
nand U8321 (N_8321,N_8221,N_8047);
nand U8322 (N_8322,N_8069,N_8125);
and U8323 (N_8323,N_8216,N_8095);
and U8324 (N_8324,N_8084,N_8230);
nand U8325 (N_8325,N_8024,N_8096);
nor U8326 (N_8326,N_8043,N_8035);
xor U8327 (N_8327,N_8111,N_8135);
nand U8328 (N_8328,N_8122,N_8228);
nor U8329 (N_8329,N_8015,N_8220);
nand U8330 (N_8330,N_8236,N_8005);
nand U8331 (N_8331,N_8012,N_8104);
xnor U8332 (N_8332,N_8131,N_8112);
nand U8333 (N_8333,N_8016,N_8217);
and U8334 (N_8334,N_8039,N_8190);
or U8335 (N_8335,N_8173,N_8071);
nor U8336 (N_8336,N_8199,N_8240);
or U8337 (N_8337,N_8161,N_8235);
and U8338 (N_8338,N_8242,N_8222);
nor U8339 (N_8339,N_8058,N_8044);
and U8340 (N_8340,N_8187,N_8183);
or U8341 (N_8341,N_8167,N_8068);
and U8342 (N_8342,N_8070,N_8114);
or U8343 (N_8343,N_8208,N_8227);
nand U8344 (N_8344,N_8098,N_8089);
or U8345 (N_8345,N_8040,N_8119);
nor U8346 (N_8346,N_8176,N_8037);
xnor U8347 (N_8347,N_8164,N_8158);
nor U8348 (N_8348,N_8042,N_8152);
nand U8349 (N_8349,N_8036,N_8121);
nand U8350 (N_8350,N_8014,N_8030);
nor U8351 (N_8351,N_8210,N_8029);
or U8352 (N_8352,N_8193,N_8197);
xor U8353 (N_8353,N_8232,N_8093);
and U8354 (N_8354,N_8248,N_8009);
nand U8355 (N_8355,N_8185,N_8169);
nand U8356 (N_8356,N_8075,N_8123);
or U8357 (N_8357,N_8006,N_8054);
nor U8358 (N_8358,N_8149,N_8077);
or U8359 (N_8359,N_8237,N_8057);
nor U8360 (N_8360,N_8013,N_8203);
or U8361 (N_8361,N_8090,N_8134);
nand U8362 (N_8362,N_8186,N_8079);
xor U8363 (N_8363,N_8109,N_8247);
xnor U8364 (N_8364,N_8136,N_8215);
nor U8365 (N_8365,N_8202,N_8206);
xor U8366 (N_8366,N_8086,N_8160);
nand U8367 (N_8367,N_8102,N_8224);
xnor U8368 (N_8368,N_8166,N_8174);
nor U8369 (N_8369,N_8082,N_8249);
and U8370 (N_8370,N_8181,N_8092);
nor U8371 (N_8371,N_8155,N_8008);
xor U8372 (N_8372,N_8180,N_8133);
xnor U8373 (N_8373,N_8046,N_8205);
nor U8374 (N_8374,N_8083,N_8080);
nor U8375 (N_8375,N_8242,N_8134);
xnor U8376 (N_8376,N_8167,N_8048);
xor U8377 (N_8377,N_8038,N_8223);
or U8378 (N_8378,N_8067,N_8148);
or U8379 (N_8379,N_8150,N_8108);
and U8380 (N_8380,N_8249,N_8121);
xor U8381 (N_8381,N_8133,N_8088);
and U8382 (N_8382,N_8047,N_8044);
nand U8383 (N_8383,N_8240,N_8108);
nor U8384 (N_8384,N_8111,N_8089);
nand U8385 (N_8385,N_8102,N_8062);
and U8386 (N_8386,N_8150,N_8035);
and U8387 (N_8387,N_8095,N_8087);
or U8388 (N_8388,N_8224,N_8232);
and U8389 (N_8389,N_8116,N_8171);
and U8390 (N_8390,N_8096,N_8245);
xnor U8391 (N_8391,N_8032,N_8172);
nand U8392 (N_8392,N_8003,N_8068);
nor U8393 (N_8393,N_8179,N_8052);
nand U8394 (N_8394,N_8206,N_8017);
xnor U8395 (N_8395,N_8213,N_8071);
nor U8396 (N_8396,N_8186,N_8013);
nor U8397 (N_8397,N_8079,N_8132);
xnor U8398 (N_8398,N_8040,N_8163);
nand U8399 (N_8399,N_8239,N_8011);
nand U8400 (N_8400,N_8059,N_8238);
nand U8401 (N_8401,N_8064,N_8140);
nor U8402 (N_8402,N_8236,N_8011);
and U8403 (N_8403,N_8055,N_8178);
xor U8404 (N_8404,N_8194,N_8210);
and U8405 (N_8405,N_8039,N_8194);
and U8406 (N_8406,N_8214,N_8179);
nor U8407 (N_8407,N_8169,N_8047);
xnor U8408 (N_8408,N_8180,N_8215);
or U8409 (N_8409,N_8067,N_8236);
or U8410 (N_8410,N_8139,N_8058);
nand U8411 (N_8411,N_8159,N_8161);
and U8412 (N_8412,N_8152,N_8205);
or U8413 (N_8413,N_8203,N_8086);
nor U8414 (N_8414,N_8079,N_8048);
and U8415 (N_8415,N_8049,N_8229);
nand U8416 (N_8416,N_8110,N_8070);
nand U8417 (N_8417,N_8172,N_8174);
and U8418 (N_8418,N_8219,N_8003);
or U8419 (N_8419,N_8063,N_8098);
nor U8420 (N_8420,N_8120,N_8188);
nor U8421 (N_8421,N_8052,N_8146);
and U8422 (N_8422,N_8072,N_8099);
or U8423 (N_8423,N_8132,N_8179);
and U8424 (N_8424,N_8010,N_8093);
or U8425 (N_8425,N_8130,N_8172);
nand U8426 (N_8426,N_8054,N_8212);
and U8427 (N_8427,N_8222,N_8010);
nor U8428 (N_8428,N_8107,N_8036);
nand U8429 (N_8429,N_8201,N_8190);
and U8430 (N_8430,N_8172,N_8190);
or U8431 (N_8431,N_8048,N_8131);
or U8432 (N_8432,N_8115,N_8063);
or U8433 (N_8433,N_8041,N_8157);
nand U8434 (N_8434,N_8197,N_8218);
nor U8435 (N_8435,N_8084,N_8082);
or U8436 (N_8436,N_8200,N_8061);
xnor U8437 (N_8437,N_8031,N_8153);
nand U8438 (N_8438,N_8211,N_8039);
and U8439 (N_8439,N_8165,N_8241);
nor U8440 (N_8440,N_8044,N_8084);
and U8441 (N_8441,N_8128,N_8087);
xnor U8442 (N_8442,N_8208,N_8159);
xor U8443 (N_8443,N_8181,N_8227);
and U8444 (N_8444,N_8076,N_8006);
and U8445 (N_8445,N_8074,N_8176);
nor U8446 (N_8446,N_8004,N_8117);
nor U8447 (N_8447,N_8126,N_8033);
xnor U8448 (N_8448,N_8065,N_8238);
or U8449 (N_8449,N_8040,N_8209);
nor U8450 (N_8450,N_8018,N_8088);
nand U8451 (N_8451,N_8040,N_8221);
and U8452 (N_8452,N_8099,N_8022);
nor U8453 (N_8453,N_8136,N_8183);
and U8454 (N_8454,N_8063,N_8096);
nand U8455 (N_8455,N_8143,N_8099);
or U8456 (N_8456,N_8249,N_8112);
nor U8457 (N_8457,N_8063,N_8222);
and U8458 (N_8458,N_8047,N_8032);
or U8459 (N_8459,N_8219,N_8173);
xor U8460 (N_8460,N_8189,N_8044);
nor U8461 (N_8461,N_8005,N_8162);
and U8462 (N_8462,N_8096,N_8098);
nor U8463 (N_8463,N_8240,N_8059);
nand U8464 (N_8464,N_8021,N_8072);
xor U8465 (N_8465,N_8068,N_8237);
nor U8466 (N_8466,N_8108,N_8084);
and U8467 (N_8467,N_8206,N_8116);
or U8468 (N_8468,N_8075,N_8225);
and U8469 (N_8469,N_8239,N_8209);
nand U8470 (N_8470,N_8220,N_8243);
nand U8471 (N_8471,N_8013,N_8118);
and U8472 (N_8472,N_8060,N_8068);
xnor U8473 (N_8473,N_8244,N_8123);
nor U8474 (N_8474,N_8117,N_8212);
nand U8475 (N_8475,N_8088,N_8033);
nand U8476 (N_8476,N_8083,N_8054);
xnor U8477 (N_8477,N_8123,N_8240);
nand U8478 (N_8478,N_8221,N_8062);
xnor U8479 (N_8479,N_8162,N_8196);
nor U8480 (N_8480,N_8174,N_8011);
nand U8481 (N_8481,N_8165,N_8191);
xor U8482 (N_8482,N_8058,N_8230);
or U8483 (N_8483,N_8182,N_8042);
nor U8484 (N_8484,N_8199,N_8156);
nor U8485 (N_8485,N_8039,N_8086);
nand U8486 (N_8486,N_8121,N_8016);
or U8487 (N_8487,N_8132,N_8134);
nor U8488 (N_8488,N_8138,N_8243);
and U8489 (N_8489,N_8119,N_8144);
nand U8490 (N_8490,N_8044,N_8033);
nor U8491 (N_8491,N_8187,N_8196);
xor U8492 (N_8492,N_8093,N_8020);
nand U8493 (N_8493,N_8046,N_8038);
nor U8494 (N_8494,N_8071,N_8245);
and U8495 (N_8495,N_8244,N_8079);
nand U8496 (N_8496,N_8009,N_8219);
xor U8497 (N_8497,N_8174,N_8234);
xnor U8498 (N_8498,N_8018,N_8171);
nand U8499 (N_8499,N_8009,N_8159);
xnor U8500 (N_8500,N_8322,N_8371);
nand U8501 (N_8501,N_8261,N_8443);
xnor U8502 (N_8502,N_8453,N_8484);
nand U8503 (N_8503,N_8394,N_8479);
or U8504 (N_8504,N_8387,N_8364);
and U8505 (N_8505,N_8478,N_8349);
nand U8506 (N_8506,N_8458,N_8469);
xnor U8507 (N_8507,N_8282,N_8471);
or U8508 (N_8508,N_8417,N_8369);
and U8509 (N_8509,N_8444,N_8385);
xor U8510 (N_8510,N_8375,N_8320);
or U8511 (N_8511,N_8348,N_8337);
nand U8512 (N_8512,N_8275,N_8428);
or U8513 (N_8513,N_8495,N_8376);
nor U8514 (N_8514,N_8475,N_8476);
nor U8515 (N_8515,N_8388,N_8323);
or U8516 (N_8516,N_8398,N_8499);
xor U8517 (N_8517,N_8255,N_8461);
and U8518 (N_8518,N_8473,N_8276);
nand U8519 (N_8519,N_8271,N_8436);
xnor U8520 (N_8520,N_8415,N_8277);
and U8521 (N_8521,N_8358,N_8268);
or U8522 (N_8522,N_8332,N_8407);
xnor U8523 (N_8523,N_8267,N_8284);
nor U8524 (N_8524,N_8381,N_8346);
nor U8525 (N_8525,N_8370,N_8402);
or U8526 (N_8526,N_8359,N_8451);
xnor U8527 (N_8527,N_8382,N_8338);
xor U8528 (N_8528,N_8343,N_8327);
nor U8529 (N_8529,N_8286,N_8367);
nor U8530 (N_8530,N_8449,N_8424);
and U8531 (N_8531,N_8279,N_8290);
nor U8532 (N_8532,N_8485,N_8254);
and U8533 (N_8533,N_8314,N_8361);
nand U8534 (N_8534,N_8465,N_8468);
or U8535 (N_8535,N_8391,N_8347);
nor U8536 (N_8536,N_8423,N_8426);
or U8537 (N_8537,N_8374,N_8351);
or U8538 (N_8538,N_8410,N_8306);
xor U8539 (N_8539,N_8345,N_8368);
and U8540 (N_8540,N_8389,N_8263);
or U8541 (N_8541,N_8422,N_8312);
and U8542 (N_8542,N_8420,N_8435);
nand U8543 (N_8543,N_8496,N_8294);
nor U8544 (N_8544,N_8299,N_8377);
or U8545 (N_8545,N_8488,N_8397);
nor U8546 (N_8546,N_8437,N_8304);
nor U8547 (N_8547,N_8403,N_8427);
nand U8548 (N_8548,N_8464,N_8431);
and U8549 (N_8549,N_8406,N_8409);
and U8550 (N_8550,N_8411,N_8378);
nand U8551 (N_8551,N_8497,N_8356);
nor U8552 (N_8552,N_8430,N_8316);
nor U8553 (N_8553,N_8467,N_8425);
xor U8554 (N_8554,N_8298,N_8326);
nor U8555 (N_8555,N_8335,N_8419);
nor U8556 (N_8556,N_8405,N_8357);
nor U8557 (N_8557,N_8413,N_8315);
or U8558 (N_8558,N_8283,N_8390);
xor U8559 (N_8559,N_8281,N_8384);
and U8560 (N_8560,N_8456,N_8330);
and U8561 (N_8561,N_8309,N_8416);
nand U8562 (N_8562,N_8455,N_8393);
nand U8563 (N_8563,N_8438,N_8273);
and U8564 (N_8564,N_8295,N_8310);
nand U8565 (N_8565,N_8480,N_8264);
or U8566 (N_8566,N_8448,N_8311);
xor U8567 (N_8567,N_8472,N_8439);
nor U8568 (N_8568,N_8462,N_8445);
xnor U8569 (N_8569,N_8318,N_8412);
and U8570 (N_8570,N_8252,N_8256);
nor U8571 (N_8571,N_8395,N_8313);
and U8572 (N_8572,N_8486,N_8251);
or U8573 (N_8573,N_8257,N_8296);
nor U8574 (N_8574,N_8408,N_8308);
nand U8575 (N_8575,N_8432,N_8386);
or U8576 (N_8576,N_8272,N_8399);
xnor U8577 (N_8577,N_8289,N_8492);
and U8578 (N_8578,N_8334,N_8440);
and U8579 (N_8579,N_8396,N_8270);
or U8580 (N_8580,N_8447,N_8260);
or U8581 (N_8581,N_8482,N_8250);
nand U8582 (N_8582,N_8360,N_8434);
and U8583 (N_8583,N_8477,N_8342);
and U8584 (N_8584,N_8328,N_8404);
xor U8585 (N_8585,N_8494,N_8373);
xnor U8586 (N_8586,N_8452,N_8344);
xor U8587 (N_8587,N_8383,N_8450);
nand U8588 (N_8588,N_8291,N_8274);
nand U8589 (N_8589,N_8331,N_8259);
and U8590 (N_8590,N_8305,N_8421);
nor U8591 (N_8591,N_8262,N_8329);
xor U8592 (N_8592,N_8303,N_8340);
nor U8593 (N_8593,N_8302,N_8363);
nand U8594 (N_8594,N_8372,N_8483);
nor U8595 (N_8595,N_8463,N_8429);
nand U8596 (N_8596,N_8339,N_8442);
or U8597 (N_8597,N_8285,N_8280);
nand U8598 (N_8598,N_8418,N_8352);
or U8599 (N_8599,N_8300,N_8481);
or U8600 (N_8600,N_8498,N_8446);
or U8601 (N_8601,N_8355,N_8454);
nand U8602 (N_8602,N_8474,N_8489);
nor U8603 (N_8603,N_8433,N_8297);
and U8604 (N_8604,N_8400,N_8287);
nand U8605 (N_8605,N_8379,N_8401);
nand U8606 (N_8606,N_8354,N_8278);
and U8607 (N_8607,N_8301,N_8380);
nand U8608 (N_8608,N_8466,N_8266);
and U8609 (N_8609,N_8317,N_8258);
nor U8610 (N_8610,N_8333,N_8414);
nand U8611 (N_8611,N_8321,N_8362);
or U8612 (N_8612,N_8307,N_8441);
and U8613 (N_8613,N_8319,N_8365);
nand U8614 (N_8614,N_8490,N_8341);
or U8615 (N_8615,N_8353,N_8253);
or U8616 (N_8616,N_8336,N_8265);
nand U8617 (N_8617,N_8491,N_8487);
nor U8618 (N_8618,N_8324,N_8392);
nor U8619 (N_8619,N_8457,N_8470);
xnor U8620 (N_8620,N_8459,N_8493);
xor U8621 (N_8621,N_8269,N_8366);
and U8622 (N_8622,N_8288,N_8293);
and U8623 (N_8623,N_8325,N_8460);
xor U8624 (N_8624,N_8350,N_8292);
nor U8625 (N_8625,N_8447,N_8405);
xnor U8626 (N_8626,N_8352,N_8310);
nand U8627 (N_8627,N_8295,N_8426);
or U8628 (N_8628,N_8469,N_8297);
or U8629 (N_8629,N_8384,N_8360);
or U8630 (N_8630,N_8302,N_8469);
and U8631 (N_8631,N_8253,N_8325);
nand U8632 (N_8632,N_8341,N_8295);
xnor U8633 (N_8633,N_8496,N_8394);
and U8634 (N_8634,N_8310,N_8492);
xor U8635 (N_8635,N_8320,N_8288);
nand U8636 (N_8636,N_8412,N_8271);
or U8637 (N_8637,N_8499,N_8489);
nor U8638 (N_8638,N_8255,N_8349);
or U8639 (N_8639,N_8396,N_8363);
or U8640 (N_8640,N_8288,N_8347);
nor U8641 (N_8641,N_8433,N_8469);
xnor U8642 (N_8642,N_8400,N_8291);
or U8643 (N_8643,N_8407,N_8276);
xor U8644 (N_8644,N_8330,N_8324);
nor U8645 (N_8645,N_8434,N_8264);
nor U8646 (N_8646,N_8370,N_8413);
xor U8647 (N_8647,N_8453,N_8472);
nand U8648 (N_8648,N_8486,N_8374);
and U8649 (N_8649,N_8407,N_8322);
nor U8650 (N_8650,N_8406,N_8309);
xnor U8651 (N_8651,N_8379,N_8356);
xnor U8652 (N_8652,N_8356,N_8459);
xor U8653 (N_8653,N_8413,N_8363);
xor U8654 (N_8654,N_8469,N_8499);
nand U8655 (N_8655,N_8455,N_8490);
or U8656 (N_8656,N_8417,N_8395);
nand U8657 (N_8657,N_8407,N_8490);
or U8658 (N_8658,N_8374,N_8381);
and U8659 (N_8659,N_8388,N_8267);
nor U8660 (N_8660,N_8268,N_8315);
xor U8661 (N_8661,N_8458,N_8436);
and U8662 (N_8662,N_8439,N_8288);
nor U8663 (N_8663,N_8496,N_8437);
nor U8664 (N_8664,N_8429,N_8342);
nand U8665 (N_8665,N_8410,N_8336);
nor U8666 (N_8666,N_8319,N_8253);
nor U8667 (N_8667,N_8408,N_8311);
xor U8668 (N_8668,N_8370,N_8397);
and U8669 (N_8669,N_8293,N_8339);
nor U8670 (N_8670,N_8388,N_8293);
and U8671 (N_8671,N_8399,N_8463);
or U8672 (N_8672,N_8404,N_8250);
xnor U8673 (N_8673,N_8390,N_8352);
xnor U8674 (N_8674,N_8345,N_8258);
nand U8675 (N_8675,N_8290,N_8347);
nand U8676 (N_8676,N_8265,N_8310);
xor U8677 (N_8677,N_8434,N_8259);
nand U8678 (N_8678,N_8339,N_8305);
nand U8679 (N_8679,N_8375,N_8357);
nor U8680 (N_8680,N_8452,N_8329);
or U8681 (N_8681,N_8329,N_8413);
nor U8682 (N_8682,N_8354,N_8332);
or U8683 (N_8683,N_8380,N_8317);
xnor U8684 (N_8684,N_8424,N_8488);
nand U8685 (N_8685,N_8250,N_8411);
nand U8686 (N_8686,N_8271,N_8295);
xnor U8687 (N_8687,N_8285,N_8250);
nand U8688 (N_8688,N_8450,N_8471);
nor U8689 (N_8689,N_8438,N_8271);
xnor U8690 (N_8690,N_8312,N_8364);
xor U8691 (N_8691,N_8294,N_8386);
nor U8692 (N_8692,N_8396,N_8443);
or U8693 (N_8693,N_8300,N_8366);
nor U8694 (N_8694,N_8327,N_8350);
or U8695 (N_8695,N_8388,N_8415);
and U8696 (N_8696,N_8417,N_8434);
or U8697 (N_8697,N_8310,N_8369);
or U8698 (N_8698,N_8285,N_8370);
nand U8699 (N_8699,N_8379,N_8435);
xnor U8700 (N_8700,N_8418,N_8334);
and U8701 (N_8701,N_8408,N_8272);
xnor U8702 (N_8702,N_8420,N_8365);
and U8703 (N_8703,N_8411,N_8496);
or U8704 (N_8704,N_8445,N_8428);
nor U8705 (N_8705,N_8479,N_8486);
nand U8706 (N_8706,N_8287,N_8468);
nor U8707 (N_8707,N_8252,N_8257);
nor U8708 (N_8708,N_8402,N_8319);
and U8709 (N_8709,N_8254,N_8344);
and U8710 (N_8710,N_8289,N_8481);
xnor U8711 (N_8711,N_8418,N_8299);
xnor U8712 (N_8712,N_8406,N_8470);
nor U8713 (N_8713,N_8450,N_8263);
and U8714 (N_8714,N_8290,N_8383);
nor U8715 (N_8715,N_8307,N_8447);
nor U8716 (N_8716,N_8330,N_8371);
or U8717 (N_8717,N_8347,N_8250);
xor U8718 (N_8718,N_8296,N_8338);
and U8719 (N_8719,N_8493,N_8289);
and U8720 (N_8720,N_8441,N_8290);
xor U8721 (N_8721,N_8390,N_8446);
xor U8722 (N_8722,N_8409,N_8384);
nand U8723 (N_8723,N_8492,N_8464);
nand U8724 (N_8724,N_8263,N_8281);
nand U8725 (N_8725,N_8295,N_8350);
nor U8726 (N_8726,N_8497,N_8422);
nor U8727 (N_8727,N_8497,N_8345);
and U8728 (N_8728,N_8463,N_8252);
nor U8729 (N_8729,N_8467,N_8270);
nand U8730 (N_8730,N_8490,N_8471);
nor U8731 (N_8731,N_8307,N_8476);
xnor U8732 (N_8732,N_8295,N_8293);
and U8733 (N_8733,N_8482,N_8464);
nand U8734 (N_8734,N_8354,N_8312);
or U8735 (N_8735,N_8429,N_8424);
nor U8736 (N_8736,N_8494,N_8346);
nor U8737 (N_8737,N_8336,N_8255);
and U8738 (N_8738,N_8370,N_8401);
xor U8739 (N_8739,N_8353,N_8255);
or U8740 (N_8740,N_8260,N_8390);
nand U8741 (N_8741,N_8306,N_8418);
or U8742 (N_8742,N_8264,N_8411);
nand U8743 (N_8743,N_8400,N_8450);
xnor U8744 (N_8744,N_8258,N_8259);
and U8745 (N_8745,N_8483,N_8496);
nand U8746 (N_8746,N_8327,N_8352);
and U8747 (N_8747,N_8308,N_8418);
nand U8748 (N_8748,N_8252,N_8347);
nand U8749 (N_8749,N_8382,N_8261);
nor U8750 (N_8750,N_8544,N_8694);
and U8751 (N_8751,N_8714,N_8618);
nor U8752 (N_8752,N_8506,N_8573);
or U8753 (N_8753,N_8681,N_8530);
nand U8754 (N_8754,N_8624,N_8523);
and U8755 (N_8755,N_8522,N_8712);
and U8756 (N_8756,N_8602,N_8627);
and U8757 (N_8757,N_8713,N_8722);
nand U8758 (N_8758,N_8519,N_8543);
xnor U8759 (N_8759,N_8696,N_8661);
and U8760 (N_8760,N_8656,N_8630);
nor U8761 (N_8761,N_8725,N_8621);
nor U8762 (N_8762,N_8553,N_8562);
xnor U8763 (N_8763,N_8625,N_8643);
nor U8764 (N_8764,N_8699,N_8646);
nor U8765 (N_8765,N_8668,N_8509);
or U8766 (N_8766,N_8613,N_8547);
nor U8767 (N_8767,N_8595,N_8549);
or U8768 (N_8768,N_8555,N_8729);
and U8769 (N_8769,N_8749,N_8538);
or U8770 (N_8770,N_8503,N_8690);
nand U8771 (N_8771,N_8675,N_8708);
and U8772 (N_8772,N_8706,N_8651);
xor U8773 (N_8773,N_8679,N_8589);
nor U8774 (N_8774,N_8584,N_8680);
or U8775 (N_8775,N_8501,N_8537);
and U8776 (N_8776,N_8609,N_8684);
or U8777 (N_8777,N_8603,N_8719);
nor U8778 (N_8778,N_8510,N_8600);
xor U8779 (N_8779,N_8535,N_8673);
and U8780 (N_8780,N_8735,N_8724);
and U8781 (N_8781,N_8515,N_8727);
xor U8782 (N_8782,N_8581,N_8610);
and U8783 (N_8783,N_8570,N_8676);
nor U8784 (N_8784,N_8660,N_8578);
nand U8785 (N_8785,N_8663,N_8601);
or U8786 (N_8786,N_8507,N_8733);
or U8787 (N_8787,N_8718,N_8742);
nor U8788 (N_8788,N_8648,N_8731);
xnor U8789 (N_8789,N_8697,N_8560);
xor U8790 (N_8790,N_8649,N_8730);
or U8791 (N_8791,N_8521,N_8534);
or U8792 (N_8792,N_8616,N_8520);
and U8793 (N_8793,N_8586,N_8606);
nand U8794 (N_8794,N_8726,N_8700);
and U8795 (N_8795,N_8524,N_8525);
nand U8796 (N_8796,N_8505,N_8596);
xnor U8797 (N_8797,N_8662,N_8612);
xor U8798 (N_8798,N_8559,N_8633);
nand U8799 (N_8799,N_8667,N_8682);
nor U8800 (N_8800,N_8611,N_8644);
or U8801 (N_8801,N_8640,N_8631);
nor U8802 (N_8802,N_8736,N_8585);
nor U8803 (N_8803,N_8691,N_8715);
and U8804 (N_8804,N_8591,N_8634);
nand U8805 (N_8805,N_8737,N_8598);
or U8806 (N_8806,N_8568,N_8615);
or U8807 (N_8807,N_8693,N_8658);
nor U8808 (N_8808,N_8707,N_8744);
or U8809 (N_8809,N_8593,N_8604);
xor U8810 (N_8810,N_8532,N_8641);
and U8811 (N_8811,N_8677,N_8716);
xnor U8812 (N_8812,N_8659,N_8687);
nand U8813 (N_8813,N_8626,N_8747);
and U8814 (N_8814,N_8709,N_8587);
nor U8815 (N_8815,N_8550,N_8545);
nor U8816 (N_8816,N_8539,N_8664);
or U8817 (N_8817,N_8678,N_8685);
and U8818 (N_8818,N_8642,N_8527);
and U8819 (N_8819,N_8552,N_8701);
or U8820 (N_8820,N_8582,N_8579);
nor U8821 (N_8821,N_8597,N_8617);
xnor U8822 (N_8822,N_8548,N_8689);
nand U8823 (N_8823,N_8732,N_8575);
xor U8824 (N_8824,N_8569,N_8526);
nand U8825 (N_8825,N_8635,N_8551);
xor U8826 (N_8826,N_8739,N_8720);
and U8827 (N_8827,N_8705,N_8745);
and U8828 (N_8828,N_8723,N_8511);
nor U8829 (N_8829,N_8546,N_8672);
or U8830 (N_8830,N_8688,N_8698);
and U8831 (N_8831,N_8567,N_8728);
nand U8832 (N_8832,N_8518,N_8541);
xor U8833 (N_8833,N_8704,N_8666);
and U8834 (N_8834,N_8607,N_8557);
and U8835 (N_8835,N_8528,N_8536);
or U8836 (N_8836,N_8623,N_8734);
or U8837 (N_8837,N_8533,N_8746);
or U8838 (N_8838,N_8517,N_8558);
nor U8839 (N_8839,N_8592,N_8703);
nand U8840 (N_8840,N_8695,N_8628);
xor U8841 (N_8841,N_8561,N_8638);
or U8842 (N_8842,N_8669,N_8653);
or U8843 (N_8843,N_8599,N_8529);
or U8844 (N_8844,N_8683,N_8508);
or U8845 (N_8845,N_8500,N_8563);
nor U8846 (N_8846,N_8702,N_8590);
nor U8847 (N_8847,N_8571,N_8608);
or U8848 (N_8848,N_8622,N_8512);
nor U8849 (N_8849,N_8556,N_8652);
xnor U8850 (N_8850,N_8632,N_8605);
or U8851 (N_8851,N_8513,N_8721);
nor U8852 (N_8852,N_8636,N_8576);
nand U8853 (N_8853,N_8674,N_8614);
nor U8854 (N_8854,N_8514,N_8637);
or U8855 (N_8855,N_8738,N_8647);
and U8856 (N_8856,N_8577,N_8619);
xnor U8857 (N_8857,N_8502,N_8743);
nor U8858 (N_8858,N_8542,N_8692);
nor U8859 (N_8859,N_8741,N_8504);
nand U8860 (N_8860,N_8540,N_8670);
nand U8861 (N_8861,N_8531,N_8665);
or U8862 (N_8862,N_8657,N_8565);
and U8863 (N_8863,N_8583,N_8574);
and U8864 (N_8864,N_8748,N_8566);
or U8865 (N_8865,N_8594,N_8686);
and U8866 (N_8866,N_8645,N_8654);
and U8867 (N_8867,N_8629,N_8516);
or U8868 (N_8868,N_8572,N_8717);
nand U8869 (N_8869,N_8655,N_8639);
nand U8870 (N_8870,N_8740,N_8620);
nor U8871 (N_8871,N_8554,N_8671);
or U8872 (N_8872,N_8580,N_8711);
or U8873 (N_8873,N_8564,N_8588);
or U8874 (N_8874,N_8650,N_8710);
xnor U8875 (N_8875,N_8519,N_8698);
nand U8876 (N_8876,N_8555,N_8722);
nor U8877 (N_8877,N_8642,N_8510);
and U8878 (N_8878,N_8734,N_8702);
nand U8879 (N_8879,N_8540,N_8558);
and U8880 (N_8880,N_8538,N_8746);
xnor U8881 (N_8881,N_8662,N_8507);
and U8882 (N_8882,N_8510,N_8612);
nand U8883 (N_8883,N_8642,N_8740);
xnor U8884 (N_8884,N_8512,N_8727);
or U8885 (N_8885,N_8597,N_8708);
xor U8886 (N_8886,N_8747,N_8726);
nand U8887 (N_8887,N_8599,N_8635);
and U8888 (N_8888,N_8518,N_8564);
xor U8889 (N_8889,N_8724,N_8581);
nor U8890 (N_8890,N_8598,N_8507);
xor U8891 (N_8891,N_8688,N_8740);
nand U8892 (N_8892,N_8712,N_8715);
nor U8893 (N_8893,N_8690,N_8745);
or U8894 (N_8894,N_8505,N_8688);
or U8895 (N_8895,N_8502,N_8746);
and U8896 (N_8896,N_8565,N_8630);
xor U8897 (N_8897,N_8539,N_8677);
or U8898 (N_8898,N_8697,N_8671);
xnor U8899 (N_8899,N_8726,N_8695);
nor U8900 (N_8900,N_8667,N_8530);
xnor U8901 (N_8901,N_8668,N_8502);
and U8902 (N_8902,N_8651,N_8620);
or U8903 (N_8903,N_8698,N_8704);
or U8904 (N_8904,N_8736,N_8732);
nor U8905 (N_8905,N_8516,N_8550);
nand U8906 (N_8906,N_8593,N_8725);
nand U8907 (N_8907,N_8651,N_8714);
xor U8908 (N_8908,N_8587,N_8726);
and U8909 (N_8909,N_8668,N_8591);
xor U8910 (N_8910,N_8543,N_8634);
xor U8911 (N_8911,N_8614,N_8714);
and U8912 (N_8912,N_8723,N_8660);
and U8913 (N_8913,N_8588,N_8531);
and U8914 (N_8914,N_8727,N_8598);
nor U8915 (N_8915,N_8523,N_8633);
or U8916 (N_8916,N_8561,N_8537);
xor U8917 (N_8917,N_8568,N_8648);
nor U8918 (N_8918,N_8574,N_8509);
or U8919 (N_8919,N_8619,N_8739);
or U8920 (N_8920,N_8694,N_8599);
and U8921 (N_8921,N_8691,N_8571);
xnor U8922 (N_8922,N_8641,N_8640);
nand U8923 (N_8923,N_8743,N_8626);
xnor U8924 (N_8924,N_8666,N_8708);
or U8925 (N_8925,N_8557,N_8513);
nand U8926 (N_8926,N_8581,N_8737);
and U8927 (N_8927,N_8588,N_8590);
xnor U8928 (N_8928,N_8626,N_8585);
or U8929 (N_8929,N_8664,N_8676);
and U8930 (N_8930,N_8696,N_8573);
and U8931 (N_8931,N_8711,N_8745);
xnor U8932 (N_8932,N_8622,N_8687);
nor U8933 (N_8933,N_8721,N_8726);
or U8934 (N_8934,N_8606,N_8697);
or U8935 (N_8935,N_8584,N_8691);
nand U8936 (N_8936,N_8689,N_8590);
nor U8937 (N_8937,N_8691,N_8551);
nor U8938 (N_8938,N_8514,N_8668);
nor U8939 (N_8939,N_8505,N_8695);
xor U8940 (N_8940,N_8633,N_8710);
xnor U8941 (N_8941,N_8656,N_8717);
nor U8942 (N_8942,N_8721,N_8732);
or U8943 (N_8943,N_8552,N_8677);
nand U8944 (N_8944,N_8600,N_8699);
nor U8945 (N_8945,N_8673,N_8501);
and U8946 (N_8946,N_8643,N_8617);
or U8947 (N_8947,N_8623,N_8657);
xnor U8948 (N_8948,N_8674,N_8568);
nand U8949 (N_8949,N_8599,N_8536);
nor U8950 (N_8950,N_8629,N_8502);
and U8951 (N_8951,N_8523,N_8669);
or U8952 (N_8952,N_8727,N_8510);
nand U8953 (N_8953,N_8586,N_8611);
nor U8954 (N_8954,N_8643,N_8515);
and U8955 (N_8955,N_8504,N_8509);
and U8956 (N_8956,N_8510,N_8647);
nand U8957 (N_8957,N_8669,N_8637);
nor U8958 (N_8958,N_8688,N_8598);
xnor U8959 (N_8959,N_8740,N_8508);
or U8960 (N_8960,N_8528,N_8561);
nand U8961 (N_8961,N_8672,N_8599);
nand U8962 (N_8962,N_8714,N_8679);
xor U8963 (N_8963,N_8690,N_8609);
xnor U8964 (N_8964,N_8630,N_8729);
nor U8965 (N_8965,N_8617,N_8672);
nor U8966 (N_8966,N_8546,N_8589);
and U8967 (N_8967,N_8637,N_8684);
or U8968 (N_8968,N_8581,N_8535);
nor U8969 (N_8969,N_8606,N_8642);
and U8970 (N_8970,N_8648,N_8524);
and U8971 (N_8971,N_8701,N_8558);
nand U8972 (N_8972,N_8732,N_8670);
nor U8973 (N_8973,N_8671,N_8744);
nor U8974 (N_8974,N_8718,N_8564);
xor U8975 (N_8975,N_8554,N_8597);
xnor U8976 (N_8976,N_8666,N_8624);
nand U8977 (N_8977,N_8601,N_8507);
xor U8978 (N_8978,N_8501,N_8522);
or U8979 (N_8979,N_8690,N_8593);
and U8980 (N_8980,N_8527,N_8608);
or U8981 (N_8981,N_8508,N_8659);
and U8982 (N_8982,N_8560,N_8711);
and U8983 (N_8983,N_8585,N_8665);
and U8984 (N_8984,N_8631,N_8528);
nand U8985 (N_8985,N_8697,N_8702);
or U8986 (N_8986,N_8523,N_8648);
nand U8987 (N_8987,N_8644,N_8592);
xor U8988 (N_8988,N_8572,N_8569);
nor U8989 (N_8989,N_8686,N_8556);
nor U8990 (N_8990,N_8638,N_8692);
nand U8991 (N_8991,N_8610,N_8604);
and U8992 (N_8992,N_8705,N_8649);
or U8993 (N_8993,N_8522,N_8508);
xor U8994 (N_8994,N_8661,N_8663);
or U8995 (N_8995,N_8686,N_8614);
xor U8996 (N_8996,N_8599,N_8593);
or U8997 (N_8997,N_8728,N_8740);
or U8998 (N_8998,N_8501,N_8606);
and U8999 (N_8999,N_8732,N_8531);
or U9000 (N_9000,N_8937,N_8844);
or U9001 (N_9001,N_8908,N_8752);
nand U9002 (N_9002,N_8809,N_8893);
and U9003 (N_9003,N_8952,N_8961);
xnor U9004 (N_9004,N_8972,N_8969);
or U9005 (N_9005,N_8878,N_8933);
xor U9006 (N_9006,N_8996,N_8928);
nor U9007 (N_9007,N_8785,N_8847);
and U9008 (N_9008,N_8850,N_8976);
and U9009 (N_9009,N_8962,N_8794);
xor U9010 (N_9010,N_8966,N_8776);
nand U9011 (N_9011,N_8762,N_8832);
xnor U9012 (N_9012,N_8868,N_8894);
xnor U9013 (N_9013,N_8859,N_8754);
xnor U9014 (N_9014,N_8964,N_8842);
and U9015 (N_9015,N_8796,N_8958);
xor U9016 (N_9016,N_8770,N_8947);
xor U9017 (N_9017,N_8769,N_8863);
nand U9018 (N_9018,N_8824,N_8880);
nand U9019 (N_9019,N_8887,N_8916);
nand U9020 (N_9020,N_8789,N_8956);
xor U9021 (N_9021,N_8860,N_8876);
xor U9022 (N_9022,N_8786,N_8765);
and U9023 (N_9023,N_8873,N_8861);
nor U9024 (N_9024,N_8780,N_8926);
nand U9025 (N_9025,N_8831,N_8979);
nor U9026 (N_9026,N_8772,N_8800);
or U9027 (N_9027,N_8803,N_8934);
and U9028 (N_9028,N_8750,N_8892);
nor U9029 (N_9029,N_8829,N_8825);
and U9030 (N_9030,N_8913,N_8977);
nor U9031 (N_9031,N_8806,N_8995);
nor U9032 (N_9032,N_8938,N_8848);
nor U9033 (N_9033,N_8862,N_8918);
nor U9034 (N_9034,N_8759,N_8895);
or U9035 (N_9035,N_8897,N_8965);
and U9036 (N_9036,N_8915,N_8778);
nor U9037 (N_9037,N_8812,N_8753);
or U9038 (N_9038,N_8925,N_8851);
nor U9039 (N_9039,N_8874,N_8830);
and U9040 (N_9040,N_8982,N_8857);
xor U9041 (N_9041,N_8886,N_8950);
xnor U9042 (N_9042,N_8828,N_8801);
or U9043 (N_9043,N_8811,N_8784);
xnor U9044 (N_9044,N_8764,N_8758);
xor U9045 (N_9045,N_8920,N_8902);
or U9046 (N_9046,N_8767,N_8757);
nand U9047 (N_9047,N_8927,N_8833);
nand U9048 (N_9048,N_8974,N_8804);
nand U9049 (N_9049,N_8912,N_8990);
nor U9050 (N_9050,N_8881,N_8838);
or U9051 (N_9051,N_8883,N_8791);
or U9052 (N_9052,N_8852,N_8779);
nand U9053 (N_9053,N_8932,N_8756);
xnor U9054 (N_9054,N_8808,N_8890);
nor U9055 (N_9055,N_8827,N_8948);
nor U9056 (N_9056,N_8807,N_8781);
or U9057 (N_9057,N_8967,N_8849);
and U9058 (N_9058,N_8960,N_8760);
nand U9059 (N_9059,N_8896,N_8782);
and U9060 (N_9060,N_8855,N_8986);
nor U9061 (N_9061,N_8904,N_8929);
nor U9062 (N_9062,N_8983,N_8815);
nor U9063 (N_9063,N_8888,N_8816);
nand U9064 (N_9064,N_8936,N_8840);
xor U9065 (N_9065,N_8981,N_8856);
xnor U9066 (N_9066,N_8841,N_8884);
or U9067 (N_9067,N_8865,N_8775);
nor U9068 (N_9068,N_8994,N_8975);
or U9069 (N_9069,N_8768,N_8853);
xor U9070 (N_9070,N_8795,N_8957);
nor U9071 (N_9071,N_8858,N_8879);
nor U9072 (N_9072,N_8835,N_8817);
xor U9073 (N_9073,N_8845,N_8820);
xnor U9074 (N_9074,N_8954,N_8872);
and U9075 (N_9075,N_8875,N_8940);
or U9076 (N_9076,N_8930,N_8959);
xor U9077 (N_9077,N_8923,N_8899);
nand U9078 (N_9078,N_8905,N_8792);
nor U9079 (N_9079,N_8991,N_8968);
or U9080 (N_9080,N_8971,N_8846);
or U9081 (N_9081,N_8942,N_8989);
or U9082 (N_9082,N_8935,N_8955);
or U9083 (N_9083,N_8919,N_8854);
xor U9084 (N_9084,N_8805,N_8882);
and U9085 (N_9085,N_8924,N_8783);
xnor U9086 (N_9086,N_8963,N_8889);
xnor U9087 (N_9087,N_8870,N_8907);
xnor U9088 (N_9088,N_8931,N_8793);
and U9089 (N_9089,N_8980,N_8777);
and U9090 (N_9090,N_8911,N_8939);
nor U9091 (N_9091,N_8946,N_8798);
xor U9092 (N_9092,N_8987,N_8891);
and U9093 (N_9093,N_8790,N_8843);
or U9094 (N_9094,N_8951,N_8993);
xnor U9095 (N_9095,N_8802,N_8985);
xor U9096 (N_9096,N_8944,N_8978);
xor U9097 (N_9097,N_8837,N_8799);
nand U9098 (N_9098,N_8766,N_8751);
nand U9099 (N_9099,N_8909,N_8819);
nor U9100 (N_9100,N_8885,N_8821);
nand U9101 (N_9101,N_8877,N_8943);
nor U9102 (N_9102,N_8823,N_8898);
nand U9103 (N_9103,N_8997,N_8866);
or U9104 (N_9104,N_8864,N_8761);
or U9105 (N_9105,N_8834,N_8988);
xnor U9106 (N_9106,N_8901,N_8953);
or U9107 (N_9107,N_8970,N_8900);
nand U9108 (N_9108,N_8839,N_8771);
nand U9109 (N_9109,N_8945,N_8992);
or U9110 (N_9110,N_8867,N_8818);
xnor U9111 (N_9111,N_8788,N_8973);
xnor U9112 (N_9112,N_8814,N_8822);
nor U9113 (N_9113,N_8755,N_8906);
and U9114 (N_9114,N_8914,N_8773);
nand U9115 (N_9115,N_8813,N_8836);
or U9116 (N_9116,N_8787,N_8999);
xor U9117 (N_9117,N_8941,N_8949);
and U9118 (N_9118,N_8917,N_8774);
nor U9119 (N_9119,N_8763,N_8910);
and U9120 (N_9120,N_8922,N_8826);
xnor U9121 (N_9121,N_8871,N_8869);
nor U9122 (N_9122,N_8810,N_8998);
nor U9123 (N_9123,N_8903,N_8921);
or U9124 (N_9124,N_8797,N_8984);
or U9125 (N_9125,N_8853,N_8980);
nand U9126 (N_9126,N_8799,N_8890);
nor U9127 (N_9127,N_8986,N_8754);
nor U9128 (N_9128,N_8841,N_8972);
nand U9129 (N_9129,N_8930,N_8975);
nor U9130 (N_9130,N_8817,N_8872);
nor U9131 (N_9131,N_8945,N_8937);
or U9132 (N_9132,N_8927,N_8801);
xor U9133 (N_9133,N_8852,N_8878);
xor U9134 (N_9134,N_8826,N_8756);
nor U9135 (N_9135,N_8759,N_8979);
and U9136 (N_9136,N_8761,N_8808);
nor U9137 (N_9137,N_8895,N_8978);
nand U9138 (N_9138,N_8838,N_8899);
and U9139 (N_9139,N_8821,N_8921);
or U9140 (N_9140,N_8993,N_8771);
nor U9141 (N_9141,N_8952,N_8761);
nand U9142 (N_9142,N_8979,N_8766);
nand U9143 (N_9143,N_8970,N_8869);
and U9144 (N_9144,N_8843,N_8846);
xor U9145 (N_9145,N_8853,N_8933);
or U9146 (N_9146,N_8940,N_8794);
nand U9147 (N_9147,N_8752,N_8936);
and U9148 (N_9148,N_8923,N_8971);
and U9149 (N_9149,N_8988,N_8966);
and U9150 (N_9150,N_8962,N_8980);
and U9151 (N_9151,N_8867,N_8956);
and U9152 (N_9152,N_8814,N_8937);
and U9153 (N_9153,N_8875,N_8786);
or U9154 (N_9154,N_8904,N_8992);
nand U9155 (N_9155,N_8768,N_8756);
nand U9156 (N_9156,N_8793,N_8985);
and U9157 (N_9157,N_8872,N_8974);
or U9158 (N_9158,N_8865,N_8874);
xnor U9159 (N_9159,N_8765,N_8920);
xor U9160 (N_9160,N_8852,N_8835);
xor U9161 (N_9161,N_8912,N_8775);
and U9162 (N_9162,N_8883,N_8878);
nand U9163 (N_9163,N_8883,N_8808);
nand U9164 (N_9164,N_8774,N_8951);
nor U9165 (N_9165,N_8779,N_8927);
nand U9166 (N_9166,N_8780,N_8918);
or U9167 (N_9167,N_8872,N_8981);
and U9168 (N_9168,N_8962,N_8968);
and U9169 (N_9169,N_8801,N_8943);
and U9170 (N_9170,N_8845,N_8752);
nand U9171 (N_9171,N_8923,N_8940);
nand U9172 (N_9172,N_8765,N_8946);
nor U9173 (N_9173,N_8912,N_8948);
nor U9174 (N_9174,N_8760,N_8955);
and U9175 (N_9175,N_8978,N_8842);
and U9176 (N_9176,N_8893,N_8967);
nand U9177 (N_9177,N_8784,N_8868);
xnor U9178 (N_9178,N_8865,N_8779);
or U9179 (N_9179,N_8915,N_8846);
xor U9180 (N_9180,N_8944,N_8801);
and U9181 (N_9181,N_8783,N_8832);
nand U9182 (N_9182,N_8814,N_8847);
nor U9183 (N_9183,N_8969,N_8943);
nand U9184 (N_9184,N_8772,N_8836);
and U9185 (N_9185,N_8755,N_8852);
or U9186 (N_9186,N_8774,N_8998);
or U9187 (N_9187,N_8954,N_8985);
xnor U9188 (N_9188,N_8978,N_8931);
nor U9189 (N_9189,N_8927,N_8772);
nor U9190 (N_9190,N_8976,N_8776);
nor U9191 (N_9191,N_8833,N_8998);
nand U9192 (N_9192,N_8904,N_8888);
and U9193 (N_9193,N_8878,N_8978);
xor U9194 (N_9194,N_8971,N_8796);
xnor U9195 (N_9195,N_8964,N_8888);
nand U9196 (N_9196,N_8759,N_8788);
xnor U9197 (N_9197,N_8866,N_8813);
nand U9198 (N_9198,N_8858,N_8894);
xnor U9199 (N_9199,N_8818,N_8879);
nor U9200 (N_9200,N_8966,N_8807);
nand U9201 (N_9201,N_8927,N_8832);
xor U9202 (N_9202,N_8937,N_8910);
xnor U9203 (N_9203,N_8826,N_8917);
xor U9204 (N_9204,N_8852,N_8924);
xor U9205 (N_9205,N_8806,N_8883);
xor U9206 (N_9206,N_8958,N_8942);
or U9207 (N_9207,N_8982,N_8762);
or U9208 (N_9208,N_8762,N_8899);
and U9209 (N_9209,N_8847,N_8780);
xnor U9210 (N_9210,N_8943,N_8859);
nor U9211 (N_9211,N_8761,N_8981);
nand U9212 (N_9212,N_8874,N_8848);
or U9213 (N_9213,N_8759,N_8781);
and U9214 (N_9214,N_8757,N_8825);
xnor U9215 (N_9215,N_8823,N_8811);
nand U9216 (N_9216,N_8815,N_8962);
or U9217 (N_9217,N_8901,N_8982);
nor U9218 (N_9218,N_8844,N_8829);
and U9219 (N_9219,N_8884,N_8959);
nor U9220 (N_9220,N_8847,N_8774);
nor U9221 (N_9221,N_8983,N_8762);
xnor U9222 (N_9222,N_8973,N_8813);
nand U9223 (N_9223,N_8773,N_8808);
or U9224 (N_9224,N_8933,N_8921);
and U9225 (N_9225,N_8798,N_8927);
nand U9226 (N_9226,N_8920,N_8791);
and U9227 (N_9227,N_8786,N_8979);
xor U9228 (N_9228,N_8862,N_8752);
nand U9229 (N_9229,N_8908,N_8950);
and U9230 (N_9230,N_8944,N_8997);
nand U9231 (N_9231,N_8981,N_8860);
and U9232 (N_9232,N_8779,N_8853);
and U9233 (N_9233,N_8792,N_8810);
or U9234 (N_9234,N_8923,N_8941);
and U9235 (N_9235,N_8797,N_8900);
nor U9236 (N_9236,N_8771,N_8911);
nand U9237 (N_9237,N_8993,N_8881);
nand U9238 (N_9238,N_8757,N_8917);
nand U9239 (N_9239,N_8899,N_8976);
and U9240 (N_9240,N_8809,N_8750);
nor U9241 (N_9241,N_8897,N_8921);
nor U9242 (N_9242,N_8795,N_8990);
or U9243 (N_9243,N_8969,N_8806);
xnor U9244 (N_9244,N_8922,N_8944);
nand U9245 (N_9245,N_8948,N_8960);
xor U9246 (N_9246,N_8768,N_8781);
and U9247 (N_9247,N_8752,N_8880);
or U9248 (N_9248,N_8843,N_8912);
or U9249 (N_9249,N_8763,N_8907);
or U9250 (N_9250,N_9109,N_9120);
nand U9251 (N_9251,N_9065,N_9168);
or U9252 (N_9252,N_9089,N_9228);
nand U9253 (N_9253,N_9125,N_9210);
nor U9254 (N_9254,N_9003,N_9181);
xnor U9255 (N_9255,N_9000,N_9019);
nor U9256 (N_9256,N_9209,N_9198);
xor U9257 (N_9257,N_9025,N_9174);
or U9258 (N_9258,N_9024,N_9161);
nor U9259 (N_9259,N_9203,N_9190);
nor U9260 (N_9260,N_9068,N_9159);
and U9261 (N_9261,N_9141,N_9213);
and U9262 (N_9262,N_9239,N_9149);
xor U9263 (N_9263,N_9045,N_9046);
or U9264 (N_9264,N_9047,N_9195);
xor U9265 (N_9265,N_9212,N_9129);
xnor U9266 (N_9266,N_9083,N_9085);
xor U9267 (N_9267,N_9075,N_9111);
xor U9268 (N_9268,N_9116,N_9041);
nor U9269 (N_9269,N_9147,N_9172);
nor U9270 (N_9270,N_9022,N_9169);
nor U9271 (N_9271,N_9215,N_9063);
nor U9272 (N_9272,N_9069,N_9217);
and U9273 (N_9273,N_9031,N_9013);
xor U9274 (N_9274,N_9021,N_9052);
nor U9275 (N_9275,N_9238,N_9163);
nor U9276 (N_9276,N_9035,N_9178);
or U9277 (N_9277,N_9206,N_9173);
nand U9278 (N_9278,N_9225,N_9230);
xor U9279 (N_9279,N_9102,N_9182);
nor U9280 (N_9280,N_9002,N_9216);
nand U9281 (N_9281,N_9023,N_9026);
xor U9282 (N_9282,N_9134,N_9082);
nand U9283 (N_9283,N_9144,N_9097);
nand U9284 (N_9284,N_9152,N_9167);
or U9285 (N_9285,N_9148,N_9233);
nor U9286 (N_9286,N_9014,N_9008);
nand U9287 (N_9287,N_9186,N_9027);
nor U9288 (N_9288,N_9162,N_9249);
nand U9289 (N_9289,N_9241,N_9077);
or U9290 (N_9290,N_9177,N_9179);
nor U9291 (N_9291,N_9101,N_9086);
nand U9292 (N_9292,N_9191,N_9006);
and U9293 (N_9293,N_9048,N_9007);
xnor U9294 (N_9294,N_9017,N_9115);
or U9295 (N_9295,N_9166,N_9033);
and U9296 (N_9296,N_9151,N_9237);
or U9297 (N_9297,N_9087,N_9124);
or U9298 (N_9298,N_9088,N_9245);
nor U9299 (N_9299,N_9098,N_9070);
nor U9300 (N_9300,N_9053,N_9030);
xor U9301 (N_9301,N_9180,N_9090);
nor U9302 (N_9302,N_9011,N_9200);
nand U9303 (N_9303,N_9040,N_9114);
and U9304 (N_9304,N_9153,N_9223);
nand U9305 (N_9305,N_9096,N_9062);
or U9306 (N_9306,N_9232,N_9135);
and U9307 (N_9307,N_9234,N_9059);
nor U9308 (N_9308,N_9220,N_9012);
and U9309 (N_9309,N_9073,N_9242);
xnor U9310 (N_9310,N_9100,N_9103);
and U9311 (N_9311,N_9156,N_9074);
nor U9312 (N_9312,N_9154,N_9229);
or U9313 (N_9313,N_9187,N_9044);
xnor U9314 (N_9314,N_9104,N_9171);
xor U9315 (N_9315,N_9043,N_9132);
or U9316 (N_9316,N_9054,N_9139);
nand U9317 (N_9317,N_9176,N_9165);
xnor U9318 (N_9318,N_9184,N_9080);
and U9319 (N_9319,N_9146,N_9016);
nand U9320 (N_9320,N_9227,N_9049);
nand U9321 (N_9321,N_9060,N_9004);
nor U9322 (N_9322,N_9057,N_9076);
and U9323 (N_9323,N_9244,N_9218);
nand U9324 (N_9324,N_9038,N_9020);
nor U9325 (N_9325,N_9034,N_9028);
nand U9326 (N_9326,N_9126,N_9235);
xnor U9327 (N_9327,N_9160,N_9246);
nand U9328 (N_9328,N_9106,N_9064);
and U9329 (N_9329,N_9183,N_9155);
nand U9330 (N_9330,N_9099,N_9196);
and U9331 (N_9331,N_9066,N_9042);
nor U9332 (N_9332,N_9197,N_9015);
and U9333 (N_9333,N_9123,N_9010);
nand U9334 (N_9334,N_9072,N_9001);
nor U9335 (N_9335,N_9071,N_9204);
xor U9336 (N_9336,N_9158,N_9029);
and U9337 (N_9337,N_9092,N_9058);
nor U9338 (N_9338,N_9145,N_9248);
xnor U9339 (N_9339,N_9136,N_9036);
nor U9340 (N_9340,N_9084,N_9110);
xnor U9341 (N_9341,N_9224,N_9222);
nor U9342 (N_9342,N_9009,N_9193);
and U9343 (N_9343,N_9189,N_9055);
xnor U9344 (N_9344,N_9137,N_9091);
xor U9345 (N_9345,N_9039,N_9175);
or U9346 (N_9346,N_9240,N_9170);
nand U9347 (N_9347,N_9208,N_9079);
or U9348 (N_9348,N_9108,N_9051);
or U9349 (N_9349,N_9150,N_9105);
nor U9350 (N_9350,N_9067,N_9112);
xor U9351 (N_9351,N_9018,N_9050);
xnor U9352 (N_9352,N_9118,N_9093);
nand U9353 (N_9353,N_9219,N_9202);
xnor U9354 (N_9354,N_9133,N_9226);
nor U9355 (N_9355,N_9128,N_9127);
xnor U9356 (N_9356,N_9113,N_9243);
nor U9357 (N_9357,N_9130,N_9140);
xor U9358 (N_9358,N_9157,N_9231);
nand U9359 (N_9359,N_9081,N_9005);
nand U9360 (N_9360,N_9078,N_9061);
nor U9361 (N_9361,N_9121,N_9143);
nor U9362 (N_9362,N_9107,N_9199);
and U9363 (N_9363,N_9211,N_9236);
nand U9364 (N_9364,N_9207,N_9185);
or U9365 (N_9365,N_9119,N_9201);
nand U9366 (N_9366,N_9117,N_9138);
nor U9367 (N_9367,N_9164,N_9122);
nand U9368 (N_9368,N_9194,N_9037);
nand U9369 (N_9369,N_9032,N_9056);
nor U9370 (N_9370,N_9094,N_9214);
nand U9371 (N_9371,N_9221,N_9142);
xnor U9372 (N_9372,N_9205,N_9192);
and U9373 (N_9373,N_9188,N_9095);
and U9374 (N_9374,N_9131,N_9247);
or U9375 (N_9375,N_9171,N_9147);
nor U9376 (N_9376,N_9087,N_9140);
and U9377 (N_9377,N_9161,N_9149);
and U9378 (N_9378,N_9049,N_9055);
or U9379 (N_9379,N_9222,N_9158);
or U9380 (N_9380,N_9101,N_9046);
or U9381 (N_9381,N_9172,N_9101);
nor U9382 (N_9382,N_9188,N_9232);
or U9383 (N_9383,N_9179,N_9000);
or U9384 (N_9384,N_9109,N_9042);
nor U9385 (N_9385,N_9246,N_9081);
and U9386 (N_9386,N_9150,N_9100);
or U9387 (N_9387,N_9078,N_9221);
or U9388 (N_9388,N_9015,N_9246);
nor U9389 (N_9389,N_9028,N_9123);
nand U9390 (N_9390,N_9155,N_9021);
xor U9391 (N_9391,N_9093,N_9016);
xnor U9392 (N_9392,N_9223,N_9241);
or U9393 (N_9393,N_9144,N_9127);
nor U9394 (N_9394,N_9094,N_9150);
nand U9395 (N_9395,N_9041,N_9136);
nand U9396 (N_9396,N_9220,N_9202);
and U9397 (N_9397,N_9152,N_9193);
xor U9398 (N_9398,N_9142,N_9106);
nand U9399 (N_9399,N_9129,N_9187);
and U9400 (N_9400,N_9112,N_9117);
nor U9401 (N_9401,N_9033,N_9151);
or U9402 (N_9402,N_9055,N_9214);
xor U9403 (N_9403,N_9233,N_9135);
and U9404 (N_9404,N_9045,N_9191);
nor U9405 (N_9405,N_9019,N_9004);
nor U9406 (N_9406,N_9068,N_9155);
and U9407 (N_9407,N_9039,N_9213);
or U9408 (N_9408,N_9134,N_9090);
nor U9409 (N_9409,N_9150,N_9225);
xnor U9410 (N_9410,N_9083,N_9074);
and U9411 (N_9411,N_9078,N_9077);
xor U9412 (N_9412,N_9244,N_9045);
nand U9413 (N_9413,N_9134,N_9236);
and U9414 (N_9414,N_9206,N_9210);
and U9415 (N_9415,N_9187,N_9123);
nor U9416 (N_9416,N_9091,N_9145);
and U9417 (N_9417,N_9183,N_9010);
nand U9418 (N_9418,N_9121,N_9244);
xnor U9419 (N_9419,N_9008,N_9049);
or U9420 (N_9420,N_9109,N_9239);
or U9421 (N_9421,N_9172,N_9214);
or U9422 (N_9422,N_9159,N_9098);
and U9423 (N_9423,N_9248,N_9226);
xnor U9424 (N_9424,N_9124,N_9033);
xnor U9425 (N_9425,N_9106,N_9062);
nor U9426 (N_9426,N_9066,N_9198);
nor U9427 (N_9427,N_9015,N_9081);
nor U9428 (N_9428,N_9042,N_9052);
xnor U9429 (N_9429,N_9087,N_9032);
nor U9430 (N_9430,N_9129,N_9110);
nor U9431 (N_9431,N_9102,N_9091);
xor U9432 (N_9432,N_9047,N_9149);
or U9433 (N_9433,N_9106,N_9100);
nand U9434 (N_9434,N_9148,N_9097);
nor U9435 (N_9435,N_9137,N_9196);
nor U9436 (N_9436,N_9006,N_9148);
or U9437 (N_9437,N_9037,N_9176);
nand U9438 (N_9438,N_9186,N_9185);
and U9439 (N_9439,N_9033,N_9117);
xor U9440 (N_9440,N_9055,N_9241);
or U9441 (N_9441,N_9157,N_9061);
and U9442 (N_9442,N_9015,N_9002);
nor U9443 (N_9443,N_9228,N_9008);
nand U9444 (N_9444,N_9029,N_9149);
xnor U9445 (N_9445,N_9116,N_9038);
or U9446 (N_9446,N_9168,N_9060);
or U9447 (N_9447,N_9247,N_9220);
or U9448 (N_9448,N_9233,N_9196);
nor U9449 (N_9449,N_9038,N_9196);
nand U9450 (N_9450,N_9054,N_9070);
nor U9451 (N_9451,N_9060,N_9222);
nand U9452 (N_9452,N_9214,N_9068);
and U9453 (N_9453,N_9195,N_9027);
nand U9454 (N_9454,N_9069,N_9219);
or U9455 (N_9455,N_9057,N_9032);
xnor U9456 (N_9456,N_9017,N_9018);
nor U9457 (N_9457,N_9115,N_9025);
xor U9458 (N_9458,N_9205,N_9128);
xnor U9459 (N_9459,N_9114,N_9159);
or U9460 (N_9460,N_9179,N_9003);
or U9461 (N_9461,N_9175,N_9180);
and U9462 (N_9462,N_9046,N_9184);
xnor U9463 (N_9463,N_9019,N_9134);
xnor U9464 (N_9464,N_9162,N_9142);
xnor U9465 (N_9465,N_9003,N_9001);
or U9466 (N_9466,N_9023,N_9160);
nor U9467 (N_9467,N_9234,N_9052);
or U9468 (N_9468,N_9206,N_9132);
nand U9469 (N_9469,N_9168,N_9114);
xnor U9470 (N_9470,N_9172,N_9131);
nor U9471 (N_9471,N_9121,N_9105);
or U9472 (N_9472,N_9080,N_9141);
nand U9473 (N_9473,N_9113,N_9013);
nor U9474 (N_9474,N_9048,N_9200);
xnor U9475 (N_9475,N_9056,N_9029);
xnor U9476 (N_9476,N_9059,N_9171);
nor U9477 (N_9477,N_9224,N_9210);
or U9478 (N_9478,N_9209,N_9233);
nor U9479 (N_9479,N_9105,N_9019);
and U9480 (N_9480,N_9021,N_9080);
and U9481 (N_9481,N_9184,N_9022);
nor U9482 (N_9482,N_9163,N_9174);
or U9483 (N_9483,N_9241,N_9164);
nand U9484 (N_9484,N_9169,N_9199);
nor U9485 (N_9485,N_9226,N_9121);
and U9486 (N_9486,N_9144,N_9011);
nand U9487 (N_9487,N_9007,N_9164);
xnor U9488 (N_9488,N_9028,N_9246);
or U9489 (N_9489,N_9194,N_9116);
xnor U9490 (N_9490,N_9065,N_9061);
xor U9491 (N_9491,N_9020,N_9013);
xnor U9492 (N_9492,N_9035,N_9132);
nand U9493 (N_9493,N_9131,N_9074);
and U9494 (N_9494,N_9069,N_9008);
xor U9495 (N_9495,N_9106,N_9099);
nand U9496 (N_9496,N_9122,N_9169);
nand U9497 (N_9497,N_9058,N_9134);
xor U9498 (N_9498,N_9121,N_9024);
or U9499 (N_9499,N_9027,N_9040);
or U9500 (N_9500,N_9299,N_9465);
nor U9501 (N_9501,N_9311,N_9288);
nand U9502 (N_9502,N_9477,N_9374);
or U9503 (N_9503,N_9432,N_9423);
nand U9504 (N_9504,N_9467,N_9487);
xnor U9505 (N_9505,N_9348,N_9356);
and U9506 (N_9506,N_9407,N_9491);
and U9507 (N_9507,N_9425,N_9268);
and U9508 (N_9508,N_9284,N_9424);
xor U9509 (N_9509,N_9305,N_9285);
or U9510 (N_9510,N_9361,N_9283);
xor U9511 (N_9511,N_9486,N_9275);
or U9512 (N_9512,N_9406,N_9346);
nand U9513 (N_9513,N_9418,N_9381);
xor U9514 (N_9514,N_9294,N_9302);
and U9515 (N_9515,N_9250,N_9429);
or U9516 (N_9516,N_9449,N_9321);
nor U9517 (N_9517,N_9456,N_9323);
nor U9518 (N_9518,N_9427,N_9493);
xor U9519 (N_9519,N_9415,N_9396);
xnor U9520 (N_9520,N_9363,N_9395);
nor U9521 (N_9521,N_9278,N_9386);
and U9522 (N_9522,N_9495,N_9496);
and U9523 (N_9523,N_9382,N_9409);
nor U9524 (N_9524,N_9375,N_9295);
nand U9525 (N_9525,N_9410,N_9251);
xor U9526 (N_9526,N_9324,N_9454);
nand U9527 (N_9527,N_9282,N_9271);
or U9528 (N_9528,N_9314,N_9378);
and U9529 (N_9529,N_9292,N_9408);
and U9530 (N_9530,N_9400,N_9475);
and U9531 (N_9531,N_9428,N_9266);
and U9532 (N_9532,N_9254,N_9379);
nor U9533 (N_9533,N_9264,N_9277);
and U9534 (N_9534,N_9478,N_9335);
xnor U9535 (N_9535,N_9322,N_9347);
and U9536 (N_9536,N_9404,N_9256);
and U9537 (N_9537,N_9485,N_9473);
nor U9538 (N_9538,N_9460,N_9304);
and U9539 (N_9539,N_9480,N_9492);
or U9540 (N_9540,N_9483,N_9336);
nor U9541 (N_9541,N_9482,N_9479);
nand U9542 (N_9542,N_9355,N_9393);
nand U9543 (N_9543,N_9330,N_9466);
nor U9544 (N_9544,N_9376,N_9463);
nor U9545 (N_9545,N_9436,N_9269);
or U9546 (N_9546,N_9366,N_9403);
xor U9547 (N_9547,N_9272,N_9385);
and U9548 (N_9548,N_9354,N_9344);
and U9549 (N_9549,N_9293,N_9319);
nor U9550 (N_9550,N_9416,N_9301);
nor U9551 (N_9551,N_9367,N_9325);
nor U9552 (N_9552,N_9434,N_9498);
and U9553 (N_9553,N_9419,N_9274);
or U9554 (N_9554,N_9469,N_9497);
and U9555 (N_9555,N_9459,N_9370);
nand U9556 (N_9556,N_9279,N_9387);
nor U9557 (N_9557,N_9281,N_9368);
xnor U9558 (N_9558,N_9364,N_9448);
or U9559 (N_9559,N_9345,N_9340);
xor U9560 (N_9560,N_9398,N_9414);
nand U9561 (N_9561,N_9280,N_9310);
and U9562 (N_9562,N_9391,N_9470);
and U9563 (N_9563,N_9358,N_9405);
nor U9564 (N_9564,N_9444,N_9259);
nand U9565 (N_9565,N_9258,N_9339);
nor U9566 (N_9566,N_9341,N_9372);
or U9567 (N_9567,N_9326,N_9494);
nand U9568 (N_9568,N_9377,N_9342);
or U9569 (N_9569,N_9445,N_9362);
and U9570 (N_9570,N_9457,N_9472);
xor U9571 (N_9571,N_9420,N_9422);
xnor U9572 (N_9572,N_9318,N_9352);
or U9573 (N_9573,N_9300,N_9296);
nor U9574 (N_9574,N_9307,N_9402);
nor U9575 (N_9575,N_9431,N_9462);
nand U9576 (N_9576,N_9262,N_9389);
nand U9577 (N_9577,N_9265,N_9388);
nor U9578 (N_9578,N_9317,N_9430);
nor U9579 (N_9579,N_9455,N_9290);
xor U9580 (N_9580,N_9426,N_9412);
nand U9581 (N_9581,N_9488,N_9312);
or U9582 (N_9582,N_9333,N_9371);
and U9583 (N_9583,N_9287,N_9357);
nor U9584 (N_9584,N_9452,N_9257);
nand U9585 (N_9585,N_9446,N_9337);
xor U9586 (N_9586,N_9468,N_9440);
or U9587 (N_9587,N_9474,N_9451);
nor U9588 (N_9588,N_9252,N_9328);
nor U9589 (N_9589,N_9447,N_9298);
nor U9590 (N_9590,N_9499,N_9349);
nand U9591 (N_9591,N_9306,N_9450);
or U9592 (N_9592,N_9413,N_9438);
nand U9593 (N_9593,N_9332,N_9289);
or U9594 (N_9594,N_9353,N_9421);
nand U9595 (N_9595,N_9481,N_9399);
xnor U9596 (N_9596,N_9327,N_9343);
nand U9597 (N_9597,N_9490,N_9442);
nand U9598 (N_9598,N_9484,N_9369);
and U9599 (N_9599,N_9458,N_9394);
or U9600 (N_9600,N_9267,N_9263);
xor U9601 (N_9601,N_9433,N_9411);
or U9602 (N_9602,N_9315,N_9313);
nor U9603 (N_9603,N_9331,N_9461);
and U9604 (N_9604,N_9308,N_9334);
xnor U9605 (N_9605,N_9286,N_9297);
or U9606 (N_9606,N_9384,N_9273);
nor U9607 (N_9607,N_9276,N_9360);
nor U9608 (N_9608,N_9350,N_9320);
nand U9609 (N_9609,N_9260,N_9435);
or U9610 (N_9610,N_9365,N_9329);
nand U9611 (N_9611,N_9261,N_9437);
and U9612 (N_9612,N_9316,N_9303);
nand U9613 (N_9613,N_9439,N_9471);
xor U9614 (N_9614,N_9441,N_9291);
or U9615 (N_9615,N_9390,N_9453);
xnor U9616 (N_9616,N_9443,N_9373);
nand U9617 (N_9617,N_9401,N_9359);
nand U9618 (N_9618,N_9464,N_9309);
nand U9619 (N_9619,N_9351,N_9397);
nor U9620 (N_9620,N_9338,N_9383);
xor U9621 (N_9621,N_9417,N_9253);
xnor U9622 (N_9622,N_9255,N_9392);
xnor U9623 (N_9623,N_9489,N_9380);
or U9624 (N_9624,N_9476,N_9270);
or U9625 (N_9625,N_9329,N_9369);
xnor U9626 (N_9626,N_9390,N_9287);
nand U9627 (N_9627,N_9275,N_9470);
and U9628 (N_9628,N_9300,N_9478);
and U9629 (N_9629,N_9495,N_9446);
nor U9630 (N_9630,N_9294,N_9326);
nand U9631 (N_9631,N_9452,N_9281);
nand U9632 (N_9632,N_9376,N_9256);
and U9633 (N_9633,N_9376,N_9277);
xnor U9634 (N_9634,N_9377,N_9346);
nor U9635 (N_9635,N_9267,N_9431);
xor U9636 (N_9636,N_9356,N_9487);
and U9637 (N_9637,N_9299,N_9443);
xnor U9638 (N_9638,N_9478,N_9281);
or U9639 (N_9639,N_9442,N_9279);
xnor U9640 (N_9640,N_9347,N_9429);
xnor U9641 (N_9641,N_9272,N_9480);
xor U9642 (N_9642,N_9276,N_9451);
nor U9643 (N_9643,N_9407,N_9263);
nand U9644 (N_9644,N_9404,N_9381);
nand U9645 (N_9645,N_9261,N_9341);
xor U9646 (N_9646,N_9351,N_9389);
or U9647 (N_9647,N_9432,N_9437);
xor U9648 (N_9648,N_9419,N_9362);
or U9649 (N_9649,N_9452,N_9337);
and U9650 (N_9650,N_9499,N_9478);
or U9651 (N_9651,N_9362,N_9327);
or U9652 (N_9652,N_9252,N_9329);
nand U9653 (N_9653,N_9283,N_9380);
nand U9654 (N_9654,N_9390,N_9297);
nand U9655 (N_9655,N_9420,N_9305);
xnor U9656 (N_9656,N_9353,N_9329);
and U9657 (N_9657,N_9349,N_9450);
nor U9658 (N_9658,N_9390,N_9285);
xnor U9659 (N_9659,N_9301,N_9338);
nor U9660 (N_9660,N_9489,N_9326);
xnor U9661 (N_9661,N_9341,N_9451);
nor U9662 (N_9662,N_9463,N_9343);
nand U9663 (N_9663,N_9408,N_9344);
xor U9664 (N_9664,N_9316,N_9428);
or U9665 (N_9665,N_9493,N_9486);
nand U9666 (N_9666,N_9439,N_9290);
and U9667 (N_9667,N_9364,N_9438);
and U9668 (N_9668,N_9294,N_9312);
nand U9669 (N_9669,N_9383,N_9391);
nand U9670 (N_9670,N_9416,N_9320);
and U9671 (N_9671,N_9318,N_9260);
nand U9672 (N_9672,N_9415,N_9301);
and U9673 (N_9673,N_9477,N_9410);
or U9674 (N_9674,N_9292,N_9409);
or U9675 (N_9675,N_9473,N_9392);
xnor U9676 (N_9676,N_9375,N_9361);
nand U9677 (N_9677,N_9359,N_9280);
xnor U9678 (N_9678,N_9263,N_9313);
and U9679 (N_9679,N_9333,N_9453);
nor U9680 (N_9680,N_9335,N_9352);
xor U9681 (N_9681,N_9296,N_9343);
or U9682 (N_9682,N_9434,N_9302);
nor U9683 (N_9683,N_9343,N_9419);
or U9684 (N_9684,N_9254,N_9495);
or U9685 (N_9685,N_9397,N_9409);
nand U9686 (N_9686,N_9459,N_9408);
xnor U9687 (N_9687,N_9386,N_9492);
or U9688 (N_9688,N_9367,N_9467);
nor U9689 (N_9689,N_9260,N_9467);
and U9690 (N_9690,N_9431,N_9348);
nor U9691 (N_9691,N_9481,N_9272);
nand U9692 (N_9692,N_9403,N_9455);
and U9693 (N_9693,N_9318,N_9462);
nand U9694 (N_9694,N_9251,N_9451);
xor U9695 (N_9695,N_9340,N_9402);
nor U9696 (N_9696,N_9454,N_9447);
nor U9697 (N_9697,N_9306,N_9409);
nand U9698 (N_9698,N_9256,N_9281);
and U9699 (N_9699,N_9273,N_9442);
nor U9700 (N_9700,N_9382,N_9258);
and U9701 (N_9701,N_9326,N_9315);
and U9702 (N_9702,N_9399,N_9439);
or U9703 (N_9703,N_9345,N_9495);
nand U9704 (N_9704,N_9487,N_9337);
nor U9705 (N_9705,N_9365,N_9478);
xnor U9706 (N_9706,N_9479,N_9262);
xor U9707 (N_9707,N_9488,N_9365);
nand U9708 (N_9708,N_9474,N_9443);
or U9709 (N_9709,N_9343,N_9368);
xor U9710 (N_9710,N_9409,N_9442);
and U9711 (N_9711,N_9251,N_9349);
xor U9712 (N_9712,N_9261,N_9272);
nor U9713 (N_9713,N_9325,N_9301);
xnor U9714 (N_9714,N_9320,N_9281);
and U9715 (N_9715,N_9281,N_9473);
or U9716 (N_9716,N_9451,N_9310);
nor U9717 (N_9717,N_9413,N_9400);
xor U9718 (N_9718,N_9312,N_9347);
nand U9719 (N_9719,N_9435,N_9252);
nor U9720 (N_9720,N_9363,N_9265);
nand U9721 (N_9721,N_9429,N_9489);
nor U9722 (N_9722,N_9348,N_9364);
xnor U9723 (N_9723,N_9429,N_9342);
nand U9724 (N_9724,N_9444,N_9458);
or U9725 (N_9725,N_9492,N_9486);
nor U9726 (N_9726,N_9321,N_9377);
nand U9727 (N_9727,N_9381,N_9396);
and U9728 (N_9728,N_9352,N_9268);
nor U9729 (N_9729,N_9419,N_9291);
nand U9730 (N_9730,N_9255,N_9313);
xor U9731 (N_9731,N_9330,N_9258);
xor U9732 (N_9732,N_9351,N_9444);
nor U9733 (N_9733,N_9324,N_9405);
and U9734 (N_9734,N_9254,N_9262);
and U9735 (N_9735,N_9408,N_9433);
nand U9736 (N_9736,N_9467,N_9375);
nor U9737 (N_9737,N_9360,N_9441);
nand U9738 (N_9738,N_9357,N_9412);
and U9739 (N_9739,N_9393,N_9286);
nand U9740 (N_9740,N_9387,N_9261);
nor U9741 (N_9741,N_9494,N_9261);
or U9742 (N_9742,N_9283,N_9365);
or U9743 (N_9743,N_9294,N_9443);
nor U9744 (N_9744,N_9461,N_9450);
nor U9745 (N_9745,N_9450,N_9279);
nor U9746 (N_9746,N_9489,N_9311);
and U9747 (N_9747,N_9498,N_9333);
or U9748 (N_9748,N_9276,N_9416);
and U9749 (N_9749,N_9358,N_9335);
or U9750 (N_9750,N_9719,N_9640);
and U9751 (N_9751,N_9637,N_9550);
and U9752 (N_9752,N_9518,N_9681);
xnor U9753 (N_9753,N_9739,N_9656);
or U9754 (N_9754,N_9695,N_9747);
xnor U9755 (N_9755,N_9743,N_9737);
nand U9756 (N_9756,N_9588,N_9506);
and U9757 (N_9757,N_9597,N_9668);
and U9758 (N_9758,N_9636,N_9539);
xor U9759 (N_9759,N_9674,N_9714);
xor U9760 (N_9760,N_9523,N_9628);
xnor U9761 (N_9761,N_9593,N_9621);
or U9762 (N_9762,N_9586,N_9577);
xor U9763 (N_9763,N_9678,N_9730);
or U9764 (N_9764,N_9665,N_9648);
and U9765 (N_9765,N_9531,N_9547);
or U9766 (N_9766,N_9643,N_9604);
nand U9767 (N_9767,N_9653,N_9603);
nor U9768 (N_9768,N_9677,N_9611);
and U9769 (N_9769,N_9572,N_9585);
or U9770 (N_9770,N_9693,N_9736);
and U9771 (N_9771,N_9587,N_9559);
nand U9772 (N_9772,N_9619,N_9646);
nor U9773 (N_9773,N_9654,N_9745);
nor U9774 (N_9774,N_9712,N_9694);
nand U9775 (N_9775,N_9617,N_9669);
nor U9776 (N_9776,N_9749,N_9647);
nor U9777 (N_9777,N_9689,N_9558);
xnor U9778 (N_9778,N_9717,N_9715);
nand U9779 (N_9779,N_9673,N_9684);
and U9780 (N_9780,N_9546,N_9567);
or U9781 (N_9781,N_9501,N_9671);
nand U9782 (N_9782,N_9610,N_9716);
nor U9783 (N_9783,N_9513,N_9562);
xnor U9784 (N_9784,N_9578,N_9720);
or U9785 (N_9785,N_9700,N_9598);
and U9786 (N_9786,N_9505,N_9521);
or U9787 (N_9787,N_9589,N_9741);
xor U9788 (N_9788,N_9528,N_9670);
and U9789 (N_9789,N_9551,N_9516);
nand U9790 (N_9790,N_9721,N_9691);
xor U9791 (N_9791,N_9740,N_9500);
xnor U9792 (N_9792,N_9725,N_9744);
and U9793 (N_9793,N_9512,N_9595);
and U9794 (N_9794,N_9625,N_9552);
or U9795 (N_9795,N_9727,N_9627);
nor U9796 (N_9796,N_9662,N_9606);
xor U9797 (N_9797,N_9591,N_9599);
nand U9798 (N_9798,N_9549,N_9746);
xor U9799 (N_9799,N_9652,N_9520);
or U9800 (N_9800,N_9532,N_9545);
nand U9801 (N_9801,N_9663,N_9602);
nand U9802 (N_9802,N_9639,N_9675);
nand U9803 (N_9803,N_9540,N_9633);
and U9804 (N_9804,N_9536,N_9735);
xnor U9805 (N_9805,N_9748,N_9724);
xnor U9806 (N_9806,N_9679,N_9583);
xnor U9807 (N_9807,N_9680,N_9711);
or U9808 (N_9808,N_9657,N_9732);
xor U9809 (N_9809,N_9605,N_9527);
and U9810 (N_9810,N_9601,N_9519);
nor U9811 (N_9811,N_9514,N_9733);
xnor U9812 (N_9812,N_9542,N_9707);
or U9813 (N_9813,N_9544,N_9710);
nand U9814 (N_9814,N_9722,N_9563);
nand U9815 (N_9815,N_9502,N_9533);
xnor U9816 (N_9816,N_9568,N_9510);
nor U9817 (N_9817,N_9509,N_9703);
nand U9818 (N_9818,N_9615,N_9729);
xor U9819 (N_9819,N_9742,N_9581);
or U9820 (N_9820,N_9503,N_9534);
and U9821 (N_9821,N_9655,N_9687);
or U9822 (N_9822,N_9709,N_9697);
and U9823 (N_9823,N_9706,N_9543);
nand U9824 (N_9824,N_9728,N_9580);
and U9825 (N_9825,N_9576,N_9696);
xnor U9826 (N_9826,N_9609,N_9734);
nor U9827 (N_9827,N_9530,N_9570);
and U9828 (N_9828,N_9651,N_9612);
xor U9829 (N_9829,N_9659,N_9624);
and U9830 (N_9830,N_9666,N_9555);
or U9831 (N_9831,N_9731,N_9644);
xor U9832 (N_9832,N_9569,N_9626);
xor U9833 (N_9833,N_9708,N_9688);
xor U9834 (N_9834,N_9629,N_9515);
xnor U9835 (N_9835,N_9692,N_9660);
or U9836 (N_9836,N_9616,N_9623);
xor U9837 (N_9837,N_9635,N_9682);
nor U9838 (N_9838,N_9672,N_9592);
xnor U9839 (N_9839,N_9522,N_9590);
nand U9840 (N_9840,N_9560,N_9538);
xor U9841 (N_9841,N_9594,N_9596);
and U9842 (N_9842,N_9622,N_9683);
and U9843 (N_9843,N_9630,N_9632);
nand U9844 (N_9844,N_9579,N_9614);
and U9845 (N_9845,N_9548,N_9575);
xor U9846 (N_9846,N_9667,N_9649);
and U9847 (N_9847,N_9613,N_9704);
or U9848 (N_9848,N_9525,N_9517);
xor U9849 (N_9849,N_9641,N_9698);
or U9850 (N_9850,N_9600,N_9566);
xor U9851 (N_9851,N_9650,N_9573);
or U9852 (N_9852,N_9608,N_9584);
or U9853 (N_9853,N_9658,N_9723);
nand U9854 (N_9854,N_9699,N_9537);
or U9855 (N_9855,N_9564,N_9557);
xnor U9856 (N_9856,N_9634,N_9690);
nor U9857 (N_9857,N_9738,N_9620);
xor U9858 (N_9858,N_9676,N_9718);
nor U9859 (N_9859,N_9524,N_9511);
nor U9860 (N_9860,N_9686,N_9582);
xnor U9861 (N_9861,N_9504,N_9553);
and U9862 (N_9862,N_9705,N_9618);
and U9863 (N_9863,N_9561,N_9565);
and U9864 (N_9864,N_9645,N_9571);
and U9865 (N_9865,N_9631,N_9541);
xnor U9866 (N_9866,N_9554,N_9574);
nand U9867 (N_9867,N_9507,N_9642);
or U9868 (N_9868,N_9529,N_9713);
nand U9869 (N_9869,N_9701,N_9535);
or U9870 (N_9870,N_9664,N_9726);
or U9871 (N_9871,N_9661,N_9526);
or U9872 (N_9872,N_9556,N_9702);
nand U9873 (N_9873,N_9607,N_9508);
or U9874 (N_9874,N_9685,N_9638);
nor U9875 (N_9875,N_9702,N_9519);
and U9876 (N_9876,N_9657,N_9563);
nand U9877 (N_9877,N_9673,N_9748);
xor U9878 (N_9878,N_9599,N_9549);
nand U9879 (N_9879,N_9640,N_9729);
and U9880 (N_9880,N_9697,N_9624);
and U9881 (N_9881,N_9511,N_9664);
xor U9882 (N_9882,N_9585,N_9727);
nor U9883 (N_9883,N_9700,N_9690);
nor U9884 (N_9884,N_9602,N_9713);
nand U9885 (N_9885,N_9586,N_9610);
or U9886 (N_9886,N_9700,N_9623);
nand U9887 (N_9887,N_9595,N_9569);
or U9888 (N_9888,N_9627,N_9645);
nand U9889 (N_9889,N_9741,N_9636);
nor U9890 (N_9890,N_9640,N_9580);
and U9891 (N_9891,N_9660,N_9666);
and U9892 (N_9892,N_9586,N_9569);
nand U9893 (N_9893,N_9741,N_9554);
or U9894 (N_9894,N_9634,N_9693);
and U9895 (N_9895,N_9542,N_9724);
xor U9896 (N_9896,N_9671,N_9668);
nand U9897 (N_9897,N_9555,N_9735);
or U9898 (N_9898,N_9530,N_9730);
and U9899 (N_9899,N_9529,N_9693);
nand U9900 (N_9900,N_9602,N_9700);
nor U9901 (N_9901,N_9709,N_9647);
xor U9902 (N_9902,N_9691,N_9584);
nand U9903 (N_9903,N_9563,N_9515);
nand U9904 (N_9904,N_9736,N_9679);
or U9905 (N_9905,N_9524,N_9746);
nand U9906 (N_9906,N_9539,N_9672);
nor U9907 (N_9907,N_9575,N_9715);
xnor U9908 (N_9908,N_9694,N_9732);
nor U9909 (N_9909,N_9557,N_9665);
xor U9910 (N_9910,N_9697,N_9583);
nand U9911 (N_9911,N_9644,N_9502);
and U9912 (N_9912,N_9613,N_9501);
xor U9913 (N_9913,N_9626,N_9591);
or U9914 (N_9914,N_9504,N_9723);
or U9915 (N_9915,N_9607,N_9592);
xnor U9916 (N_9916,N_9642,N_9572);
or U9917 (N_9917,N_9521,N_9740);
nand U9918 (N_9918,N_9709,N_9681);
nand U9919 (N_9919,N_9577,N_9649);
or U9920 (N_9920,N_9646,N_9660);
and U9921 (N_9921,N_9568,N_9734);
nor U9922 (N_9922,N_9601,N_9730);
nand U9923 (N_9923,N_9725,N_9545);
and U9924 (N_9924,N_9676,N_9586);
or U9925 (N_9925,N_9714,N_9728);
and U9926 (N_9926,N_9662,N_9509);
nor U9927 (N_9927,N_9512,N_9720);
and U9928 (N_9928,N_9559,N_9739);
nor U9929 (N_9929,N_9633,N_9723);
xnor U9930 (N_9930,N_9626,N_9572);
or U9931 (N_9931,N_9737,N_9569);
xnor U9932 (N_9932,N_9622,N_9636);
nor U9933 (N_9933,N_9719,N_9511);
xor U9934 (N_9934,N_9596,N_9547);
nor U9935 (N_9935,N_9713,N_9551);
and U9936 (N_9936,N_9633,N_9506);
or U9937 (N_9937,N_9691,N_9623);
xnor U9938 (N_9938,N_9629,N_9573);
xor U9939 (N_9939,N_9588,N_9727);
nor U9940 (N_9940,N_9563,N_9714);
and U9941 (N_9941,N_9541,N_9505);
or U9942 (N_9942,N_9645,N_9634);
nor U9943 (N_9943,N_9573,N_9515);
xor U9944 (N_9944,N_9630,N_9552);
xnor U9945 (N_9945,N_9530,N_9577);
nand U9946 (N_9946,N_9615,N_9726);
nand U9947 (N_9947,N_9605,N_9644);
xnor U9948 (N_9948,N_9556,N_9544);
nor U9949 (N_9949,N_9738,N_9631);
nor U9950 (N_9950,N_9636,N_9677);
and U9951 (N_9951,N_9739,N_9539);
and U9952 (N_9952,N_9615,N_9575);
or U9953 (N_9953,N_9502,N_9627);
nand U9954 (N_9954,N_9650,N_9550);
nor U9955 (N_9955,N_9727,N_9673);
and U9956 (N_9956,N_9735,N_9690);
and U9957 (N_9957,N_9576,N_9543);
nor U9958 (N_9958,N_9645,N_9724);
xnor U9959 (N_9959,N_9557,N_9749);
xnor U9960 (N_9960,N_9668,N_9502);
or U9961 (N_9961,N_9507,N_9563);
or U9962 (N_9962,N_9624,N_9563);
nor U9963 (N_9963,N_9574,N_9577);
and U9964 (N_9964,N_9723,N_9508);
and U9965 (N_9965,N_9508,N_9683);
xor U9966 (N_9966,N_9547,N_9742);
and U9967 (N_9967,N_9535,N_9531);
or U9968 (N_9968,N_9571,N_9594);
xor U9969 (N_9969,N_9652,N_9553);
or U9970 (N_9970,N_9508,N_9562);
xor U9971 (N_9971,N_9583,N_9728);
or U9972 (N_9972,N_9548,N_9588);
nand U9973 (N_9973,N_9576,N_9569);
nor U9974 (N_9974,N_9705,N_9538);
nand U9975 (N_9975,N_9501,N_9551);
nand U9976 (N_9976,N_9586,N_9510);
nand U9977 (N_9977,N_9582,N_9559);
and U9978 (N_9978,N_9581,N_9589);
nand U9979 (N_9979,N_9679,N_9697);
or U9980 (N_9980,N_9647,N_9699);
nand U9981 (N_9981,N_9563,N_9686);
xor U9982 (N_9982,N_9696,N_9622);
xnor U9983 (N_9983,N_9699,N_9718);
nor U9984 (N_9984,N_9553,N_9587);
nor U9985 (N_9985,N_9559,N_9629);
nand U9986 (N_9986,N_9561,N_9612);
nor U9987 (N_9987,N_9693,N_9604);
nand U9988 (N_9988,N_9630,N_9573);
xnor U9989 (N_9989,N_9688,N_9548);
nor U9990 (N_9990,N_9695,N_9625);
nand U9991 (N_9991,N_9611,N_9715);
or U9992 (N_9992,N_9617,N_9531);
nand U9993 (N_9993,N_9530,N_9676);
nor U9994 (N_9994,N_9572,N_9558);
xor U9995 (N_9995,N_9612,N_9551);
nand U9996 (N_9996,N_9581,N_9536);
or U9997 (N_9997,N_9705,N_9708);
and U9998 (N_9998,N_9743,N_9525);
xnor U9999 (N_9999,N_9598,N_9690);
nor U10000 (N_10000,N_9945,N_9854);
xnor U10001 (N_10001,N_9757,N_9916);
and U10002 (N_10002,N_9897,N_9834);
xnor U10003 (N_10003,N_9786,N_9882);
and U10004 (N_10004,N_9922,N_9799);
or U10005 (N_10005,N_9852,N_9822);
or U10006 (N_10006,N_9780,N_9766);
and U10007 (N_10007,N_9819,N_9783);
nand U10008 (N_10008,N_9857,N_9840);
nand U10009 (N_10009,N_9870,N_9761);
nand U10010 (N_10010,N_9936,N_9997);
or U10011 (N_10011,N_9896,N_9765);
or U10012 (N_10012,N_9989,N_9774);
nor U10013 (N_10013,N_9807,N_9833);
and U10014 (N_10014,N_9983,N_9888);
and U10015 (N_10015,N_9976,N_9762);
xnor U10016 (N_10016,N_9816,N_9795);
and U10017 (N_10017,N_9917,N_9817);
xor U10018 (N_10018,N_9873,N_9855);
or U10019 (N_10019,N_9994,N_9874);
nor U10020 (N_10020,N_9839,N_9959);
xor U10021 (N_10021,N_9991,N_9810);
nand U10022 (N_10022,N_9778,N_9805);
nand U10023 (N_10023,N_9800,N_9919);
and U10024 (N_10024,N_9825,N_9827);
nor U10025 (N_10025,N_9787,N_9935);
and U10026 (N_10026,N_9954,N_9871);
xnor U10027 (N_10027,N_9963,N_9946);
nor U10028 (N_10028,N_9990,N_9832);
nand U10029 (N_10029,N_9934,N_9821);
or U10030 (N_10030,N_9955,N_9993);
nor U10031 (N_10031,N_9891,N_9909);
xor U10032 (N_10032,N_9998,N_9974);
xor U10033 (N_10033,N_9830,N_9924);
and U10034 (N_10034,N_9932,N_9960);
or U10035 (N_10035,N_9838,N_9767);
xor U10036 (N_10036,N_9950,N_9880);
nand U10037 (N_10037,N_9972,N_9913);
nand U10038 (N_10038,N_9894,N_9753);
nand U10039 (N_10039,N_9881,N_9875);
xnor U10040 (N_10040,N_9943,N_9903);
xor U10041 (N_10041,N_9971,N_9895);
nand U10042 (N_10042,N_9801,N_9904);
and U10043 (N_10043,N_9889,N_9781);
or U10044 (N_10044,N_9771,N_9905);
and U10045 (N_10045,N_9979,N_9802);
nor U10046 (N_10046,N_9804,N_9975);
nor U10047 (N_10047,N_9856,N_9751);
nor U10048 (N_10048,N_9953,N_9829);
xor U10049 (N_10049,N_9847,N_9867);
xnor U10050 (N_10050,N_9773,N_9984);
or U10051 (N_10051,N_9929,N_9844);
and U10052 (N_10052,N_9890,N_9967);
xor U10053 (N_10053,N_9759,N_9811);
nand U10054 (N_10054,N_9938,N_9939);
xor U10055 (N_10055,N_9923,N_9792);
or U10056 (N_10056,N_9865,N_9768);
or U10057 (N_10057,N_9981,N_9914);
and U10058 (N_10058,N_9797,N_9937);
nor U10059 (N_10059,N_9758,N_9784);
xnor U10060 (N_10060,N_9755,N_9898);
nor U10061 (N_10061,N_9878,N_9995);
and U10062 (N_10062,N_9769,N_9837);
nor U10063 (N_10063,N_9956,N_9910);
and U10064 (N_10064,N_9980,N_9925);
nor U10065 (N_10065,N_9970,N_9944);
nor U10066 (N_10066,N_9892,N_9828);
nand U10067 (N_10067,N_9861,N_9920);
nor U10068 (N_10068,N_9899,N_9809);
nand U10069 (N_10069,N_9996,N_9928);
and U10070 (N_10070,N_9763,N_9835);
xor U10071 (N_10071,N_9853,N_9879);
or U10072 (N_10072,N_9777,N_9961);
nand U10073 (N_10073,N_9750,N_9933);
nand U10074 (N_10074,N_9941,N_9788);
nor U10075 (N_10075,N_9864,N_9884);
xnor U10076 (N_10076,N_9973,N_9824);
and U10077 (N_10077,N_9846,N_9947);
or U10078 (N_10078,N_9862,N_9860);
nand U10079 (N_10079,N_9843,N_9812);
and U10080 (N_10080,N_9901,N_9977);
nand U10081 (N_10081,N_9982,N_9915);
xor U10082 (N_10082,N_9776,N_9885);
or U10083 (N_10083,N_9820,N_9948);
and U10084 (N_10084,N_9872,N_9815);
nor U10085 (N_10085,N_9918,N_9887);
xor U10086 (N_10086,N_9876,N_9791);
xor U10087 (N_10087,N_9969,N_9999);
nor U10088 (N_10088,N_9803,N_9931);
or U10089 (N_10089,N_9764,N_9866);
nor U10090 (N_10090,N_9850,N_9851);
and U10091 (N_10091,N_9858,N_9966);
and U10092 (N_10092,N_9782,N_9985);
xor U10093 (N_10093,N_9823,N_9912);
or U10094 (N_10094,N_9779,N_9965);
and U10095 (N_10095,N_9868,N_9806);
xor U10096 (N_10096,N_9798,N_9826);
nand U10097 (N_10097,N_9869,N_9886);
nor U10098 (N_10098,N_9772,N_9789);
nor U10099 (N_10099,N_9849,N_9951);
and U10100 (N_10100,N_9907,N_9814);
or U10101 (N_10101,N_9893,N_9908);
nor U10102 (N_10102,N_9842,N_9785);
nor U10103 (N_10103,N_9877,N_9926);
nor U10104 (N_10104,N_9940,N_9900);
or U10105 (N_10105,N_9911,N_9859);
or U10106 (N_10106,N_9813,N_9831);
xnor U10107 (N_10107,N_9790,N_9770);
and U10108 (N_10108,N_9841,N_9958);
xnor U10109 (N_10109,N_9988,N_9930);
nor U10110 (N_10110,N_9902,N_9756);
nand U10111 (N_10111,N_9754,N_9952);
nor U10112 (N_10112,N_9760,N_9845);
or U10113 (N_10113,N_9962,N_9992);
nand U10114 (N_10114,N_9987,N_9906);
or U10115 (N_10115,N_9752,N_9794);
and U10116 (N_10116,N_9775,N_9808);
and U10117 (N_10117,N_9957,N_9793);
nor U10118 (N_10118,N_9848,N_9949);
nor U10119 (N_10119,N_9796,N_9927);
or U10120 (N_10120,N_9942,N_9921);
and U10121 (N_10121,N_9863,N_9978);
nand U10122 (N_10122,N_9836,N_9968);
nor U10123 (N_10123,N_9986,N_9964);
and U10124 (N_10124,N_9818,N_9883);
nand U10125 (N_10125,N_9822,N_9928);
nor U10126 (N_10126,N_9849,N_9872);
nand U10127 (N_10127,N_9800,N_9810);
or U10128 (N_10128,N_9828,N_9944);
and U10129 (N_10129,N_9958,N_9788);
and U10130 (N_10130,N_9960,N_9956);
and U10131 (N_10131,N_9907,N_9780);
nor U10132 (N_10132,N_9875,N_9869);
nor U10133 (N_10133,N_9957,N_9868);
nand U10134 (N_10134,N_9996,N_9889);
and U10135 (N_10135,N_9888,N_9855);
and U10136 (N_10136,N_9861,N_9976);
nand U10137 (N_10137,N_9813,N_9768);
nor U10138 (N_10138,N_9950,N_9889);
nor U10139 (N_10139,N_9979,N_9935);
or U10140 (N_10140,N_9762,N_9788);
or U10141 (N_10141,N_9939,N_9955);
xor U10142 (N_10142,N_9797,N_9859);
nand U10143 (N_10143,N_9902,N_9842);
nand U10144 (N_10144,N_9907,N_9789);
nand U10145 (N_10145,N_9796,N_9997);
or U10146 (N_10146,N_9906,N_9899);
nor U10147 (N_10147,N_9782,N_9898);
nor U10148 (N_10148,N_9880,N_9963);
and U10149 (N_10149,N_9759,N_9833);
or U10150 (N_10150,N_9804,N_9946);
and U10151 (N_10151,N_9823,N_9948);
nand U10152 (N_10152,N_9906,N_9943);
and U10153 (N_10153,N_9819,N_9969);
nor U10154 (N_10154,N_9874,N_9911);
or U10155 (N_10155,N_9989,N_9779);
nor U10156 (N_10156,N_9927,N_9806);
nand U10157 (N_10157,N_9893,N_9924);
and U10158 (N_10158,N_9948,N_9981);
or U10159 (N_10159,N_9986,N_9911);
or U10160 (N_10160,N_9877,N_9833);
nand U10161 (N_10161,N_9903,N_9923);
or U10162 (N_10162,N_9959,N_9945);
xnor U10163 (N_10163,N_9990,N_9950);
xor U10164 (N_10164,N_9795,N_9893);
nor U10165 (N_10165,N_9826,N_9990);
xnor U10166 (N_10166,N_9852,N_9760);
or U10167 (N_10167,N_9855,N_9933);
or U10168 (N_10168,N_9978,N_9810);
nand U10169 (N_10169,N_9768,N_9947);
nand U10170 (N_10170,N_9757,N_9961);
xor U10171 (N_10171,N_9831,N_9882);
nand U10172 (N_10172,N_9907,N_9764);
nor U10173 (N_10173,N_9883,N_9819);
nand U10174 (N_10174,N_9970,N_9947);
and U10175 (N_10175,N_9953,N_9791);
or U10176 (N_10176,N_9915,N_9991);
nor U10177 (N_10177,N_9937,N_9781);
nand U10178 (N_10178,N_9869,N_9846);
and U10179 (N_10179,N_9838,N_9862);
and U10180 (N_10180,N_9972,N_9816);
or U10181 (N_10181,N_9766,N_9959);
nand U10182 (N_10182,N_9763,N_9866);
nand U10183 (N_10183,N_9939,N_9916);
xnor U10184 (N_10184,N_9841,N_9809);
nand U10185 (N_10185,N_9870,N_9958);
or U10186 (N_10186,N_9831,N_9930);
nor U10187 (N_10187,N_9774,N_9886);
xor U10188 (N_10188,N_9765,N_9834);
xor U10189 (N_10189,N_9790,N_9846);
xnor U10190 (N_10190,N_9987,N_9797);
xor U10191 (N_10191,N_9988,N_9924);
xnor U10192 (N_10192,N_9862,N_9821);
nand U10193 (N_10193,N_9907,N_9852);
nand U10194 (N_10194,N_9801,N_9898);
and U10195 (N_10195,N_9795,N_9994);
nor U10196 (N_10196,N_9876,N_9836);
xor U10197 (N_10197,N_9955,N_9845);
nor U10198 (N_10198,N_9795,N_9982);
xor U10199 (N_10199,N_9856,N_9823);
nor U10200 (N_10200,N_9758,N_9770);
nor U10201 (N_10201,N_9953,N_9900);
and U10202 (N_10202,N_9921,N_9961);
xnor U10203 (N_10203,N_9779,N_9875);
and U10204 (N_10204,N_9938,N_9923);
nand U10205 (N_10205,N_9759,N_9758);
and U10206 (N_10206,N_9895,N_9936);
or U10207 (N_10207,N_9793,N_9969);
or U10208 (N_10208,N_9760,N_9782);
nor U10209 (N_10209,N_9882,N_9901);
xnor U10210 (N_10210,N_9839,N_9982);
nor U10211 (N_10211,N_9973,N_9759);
nand U10212 (N_10212,N_9978,N_9832);
nor U10213 (N_10213,N_9802,N_9881);
xor U10214 (N_10214,N_9778,N_9938);
nand U10215 (N_10215,N_9997,N_9880);
or U10216 (N_10216,N_9933,N_9839);
or U10217 (N_10217,N_9767,N_9819);
nand U10218 (N_10218,N_9979,N_9939);
xor U10219 (N_10219,N_9953,N_9770);
or U10220 (N_10220,N_9782,N_9777);
or U10221 (N_10221,N_9802,N_9767);
or U10222 (N_10222,N_9788,N_9972);
nand U10223 (N_10223,N_9762,N_9799);
xnor U10224 (N_10224,N_9926,N_9845);
xor U10225 (N_10225,N_9960,N_9782);
nor U10226 (N_10226,N_9933,N_9866);
xnor U10227 (N_10227,N_9841,N_9774);
and U10228 (N_10228,N_9961,N_9982);
nand U10229 (N_10229,N_9884,N_9986);
or U10230 (N_10230,N_9974,N_9885);
or U10231 (N_10231,N_9973,N_9829);
nor U10232 (N_10232,N_9756,N_9903);
xor U10233 (N_10233,N_9979,N_9898);
xor U10234 (N_10234,N_9810,N_9852);
nor U10235 (N_10235,N_9890,N_9943);
or U10236 (N_10236,N_9973,N_9863);
and U10237 (N_10237,N_9826,N_9885);
nand U10238 (N_10238,N_9943,N_9783);
xnor U10239 (N_10239,N_9785,N_9958);
and U10240 (N_10240,N_9966,N_9770);
nor U10241 (N_10241,N_9770,N_9793);
nand U10242 (N_10242,N_9839,N_9826);
xnor U10243 (N_10243,N_9833,N_9964);
or U10244 (N_10244,N_9899,N_9938);
and U10245 (N_10245,N_9957,N_9912);
xor U10246 (N_10246,N_9819,N_9908);
nor U10247 (N_10247,N_9752,N_9976);
xnor U10248 (N_10248,N_9985,N_9859);
nand U10249 (N_10249,N_9952,N_9801);
nand U10250 (N_10250,N_10067,N_10191);
and U10251 (N_10251,N_10181,N_10229);
and U10252 (N_10252,N_10010,N_10174);
or U10253 (N_10253,N_10039,N_10060);
nand U10254 (N_10254,N_10127,N_10248);
xor U10255 (N_10255,N_10173,N_10094);
nor U10256 (N_10256,N_10111,N_10091);
nor U10257 (N_10257,N_10080,N_10150);
nor U10258 (N_10258,N_10184,N_10133);
nand U10259 (N_10259,N_10053,N_10047);
nor U10260 (N_10260,N_10114,N_10038);
and U10261 (N_10261,N_10139,N_10102);
nand U10262 (N_10262,N_10126,N_10117);
and U10263 (N_10263,N_10210,N_10044);
nand U10264 (N_10264,N_10175,N_10050);
nand U10265 (N_10265,N_10195,N_10187);
nand U10266 (N_10266,N_10046,N_10239);
or U10267 (N_10267,N_10098,N_10149);
or U10268 (N_10268,N_10221,N_10092);
xnor U10269 (N_10269,N_10024,N_10041);
nand U10270 (N_10270,N_10241,N_10030);
nor U10271 (N_10271,N_10182,N_10160);
nand U10272 (N_10272,N_10021,N_10087);
xnor U10273 (N_10273,N_10151,N_10032);
and U10274 (N_10274,N_10148,N_10162);
nand U10275 (N_10275,N_10085,N_10069);
nor U10276 (N_10276,N_10134,N_10078);
nand U10277 (N_10277,N_10227,N_10016);
nor U10278 (N_10278,N_10129,N_10012);
nor U10279 (N_10279,N_10071,N_10124);
nor U10280 (N_10280,N_10001,N_10142);
and U10281 (N_10281,N_10121,N_10008);
xnor U10282 (N_10282,N_10088,N_10141);
nand U10283 (N_10283,N_10165,N_10109);
and U10284 (N_10284,N_10167,N_10154);
and U10285 (N_10285,N_10140,N_10163);
or U10286 (N_10286,N_10113,N_10058);
and U10287 (N_10287,N_10122,N_10033);
nand U10288 (N_10288,N_10112,N_10236);
nand U10289 (N_10289,N_10043,N_10222);
and U10290 (N_10290,N_10089,N_10093);
xor U10291 (N_10291,N_10152,N_10104);
nand U10292 (N_10292,N_10232,N_10176);
or U10293 (N_10293,N_10011,N_10159);
nor U10294 (N_10294,N_10145,N_10082);
xor U10295 (N_10295,N_10218,N_10027);
nor U10296 (N_10296,N_10100,N_10108);
and U10297 (N_10297,N_10048,N_10237);
and U10298 (N_10298,N_10006,N_10106);
nor U10299 (N_10299,N_10037,N_10065);
nor U10300 (N_10300,N_10186,N_10198);
nor U10301 (N_10301,N_10205,N_10209);
nand U10302 (N_10302,N_10247,N_10005);
and U10303 (N_10303,N_10115,N_10212);
xor U10304 (N_10304,N_10194,N_10119);
nand U10305 (N_10305,N_10243,N_10083);
nor U10306 (N_10306,N_10076,N_10137);
nand U10307 (N_10307,N_10215,N_10015);
nor U10308 (N_10308,N_10063,N_10234);
nor U10309 (N_10309,N_10042,N_10025);
nand U10310 (N_10310,N_10009,N_10073);
or U10311 (N_10311,N_10035,N_10183);
nand U10312 (N_10312,N_10125,N_10128);
and U10313 (N_10313,N_10054,N_10246);
or U10314 (N_10314,N_10017,N_10223);
xor U10315 (N_10315,N_10120,N_10249);
nor U10316 (N_10316,N_10171,N_10014);
and U10317 (N_10317,N_10132,N_10028);
nand U10318 (N_10318,N_10055,N_10007);
nor U10319 (N_10319,N_10095,N_10213);
and U10320 (N_10320,N_10061,N_10189);
or U10321 (N_10321,N_10072,N_10220);
or U10322 (N_10322,N_10177,N_10225);
and U10323 (N_10323,N_10211,N_10003);
nor U10324 (N_10324,N_10203,N_10096);
nand U10325 (N_10325,N_10144,N_10170);
xnor U10326 (N_10326,N_10143,N_10074);
nand U10327 (N_10327,N_10040,N_10034);
nor U10328 (N_10328,N_10097,N_10202);
nor U10329 (N_10329,N_10153,N_10123);
xnor U10330 (N_10330,N_10002,N_10062);
nor U10331 (N_10331,N_10059,N_10192);
xor U10332 (N_10332,N_10118,N_10023);
or U10333 (N_10333,N_10231,N_10190);
or U10334 (N_10334,N_10090,N_10224);
or U10335 (N_10335,N_10110,N_10101);
nor U10336 (N_10336,N_10136,N_10146);
xor U10337 (N_10337,N_10103,N_10138);
or U10338 (N_10338,N_10155,N_10056);
and U10339 (N_10339,N_10193,N_10064);
nor U10340 (N_10340,N_10166,N_10105);
nand U10341 (N_10341,N_10107,N_10199);
or U10342 (N_10342,N_10049,N_10164);
nor U10343 (N_10343,N_10022,N_10244);
xnor U10344 (N_10344,N_10196,N_10219);
nand U10345 (N_10345,N_10045,N_10099);
or U10346 (N_10346,N_10207,N_10131);
and U10347 (N_10347,N_10116,N_10004);
or U10348 (N_10348,N_10086,N_10019);
and U10349 (N_10349,N_10020,N_10057);
xor U10350 (N_10350,N_10208,N_10178);
xor U10351 (N_10351,N_10216,N_10238);
nor U10352 (N_10352,N_10226,N_10235);
nor U10353 (N_10353,N_10180,N_10206);
nand U10354 (N_10354,N_10068,N_10070);
and U10355 (N_10355,N_10135,N_10179);
or U10356 (N_10356,N_10214,N_10233);
nand U10357 (N_10357,N_10051,N_10130);
xor U10358 (N_10358,N_10197,N_10157);
nand U10359 (N_10359,N_10168,N_10169);
nand U10360 (N_10360,N_10156,N_10075);
and U10361 (N_10361,N_10217,N_10204);
or U10362 (N_10362,N_10084,N_10242);
xnor U10363 (N_10363,N_10245,N_10240);
or U10364 (N_10364,N_10200,N_10018);
and U10365 (N_10365,N_10036,N_10228);
and U10366 (N_10366,N_10079,N_10013);
nand U10367 (N_10367,N_10066,N_10000);
nand U10368 (N_10368,N_10029,N_10031);
xnor U10369 (N_10369,N_10230,N_10026);
xnor U10370 (N_10370,N_10188,N_10172);
xor U10371 (N_10371,N_10147,N_10161);
nor U10372 (N_10372,N_10052,N_10158);
nand U10373 (N_10373,N_10077,N_10185);
xor U10374 (N_10374,N_10201,N_10081);
nor U10375 (N_10375,N_10221,N_10184);
nor U10376 (N_10376,N_10201,N_10093);
nand U10377 (N_10377,N_10170,N_10227);
xnor U10378 (N_10378,N_10056,N_10116);
nor U10379 (N_10379,N_10096,N_10099);
or U10380 (N_10380,N_10155,N_10201);
nand U10381 (N_10381,N_10058,N_10021);
nor U10382 (N_10382,N_10085,N_10005);
nor U10383 (N_10383,N_10211,N_10022);
nand U10384 (N_10384,N_10184,N_10127);
nor U10385 (N_10385,N_10173,N_10108);
xor U10386 (N_10386,N_10035,N_10177);
nor U10387 (N_10387,N_10034,N_10190);
xor U10388 (N_10388,N_10129,N_10153);
xor U10389 (N_10389,N_10236,N_10223);
and U10390 (N_10390,N_10180,N_10221);
and U10391 (N_10391,N_10127,N_10200);
or U10392 (N_10392,N_10206,N_10214);
and U10393 (N_10393,N_10193,N_10019);
or U10394 (N_10394,N_10044,N_10127);
nand U10395 (N_10395,N_10218,N_10076);
xor U10396 (N_10396,N_10042,N_10104);
nand U10397 (N_10397,N_10198,N_10022);
nor U10398 (N_10398,N_10207,N_10044);
nor U10399 (N_10399,N_10236,N_10024);
nand U10400 (N_10400,N_10191,N_10212);
xnor U10401 (N_10401,N_10016,N_10085);
xnor U10402 (N_10402,N_10232,N_10079);
nor U10403 (N_10403,N_10056,N_10020);
xnor U10404 (N_10404,N_10190,N_10081);
nand U10405 (N_10405,N_10220,N_10108);
and U10406 (N_10406,N_10129,N_10130);
xnor U10407 (N_10407,N_10142,N_10099);
nand U10408 (N_10408,N_10144,N_10206);
nand U10409 (N_10409,N_10249,N_10169);
xor U10410 (N_10410,N_10191,N_10010);
or U10411 (N_10411,N_10239,N_10202);
nand U10412 (N_10412,N_10185,N_10213);
xor U10413 (N_10413,N_10200,N_10103);
nand U10414 (N_10414,N_10162,N_10223);
nand U10415 (N_10415,N_10242,N_10175);
and U10416 (N_10416,N_10218,N_10010);
or U10417 (N_10417,N_10176,N_10070);
and U10418 (N_10418,N_10223,N_10084);
xor U10419 (N_10419,N_10146,N_10199);
and U10420 (N_10420,N_10072,N_10186);
nor U10421 (N_10421,N_10184,N_10057);
nand U10422 (N_10422,N_10116,N_10071);
nand U10423 (N_10423,N_10105,N_10006);
and U10424 (N_10424,N_10087,N_10224);
or U10425 (N_10425,N_10086,N_10247);
or U10426 (N_10426,N_10017,N_10205);
or U10427 (N_10427,N_10100,N_10204);
xor U10428 (N_10428,N_10159,N_10084);
or U10429 (N_10429,N_10228,N_10026);
nand U10430 (N_10430,N_10228,N_10188);
nand U10431 (N_10431,N_10174,N_10064);
xnor U10432 (N_10432,N_10181,N_10003);
or U10433 (N_10433,N_10127,N_10071);
or U10434 (N_10434,N_10033,N_10057);
xor U10435 (N_10435,N_10005,N_10230);
or U10436 (N_10436,N_10030,N_10155);
xor U10437 (N_10437,N_10057,N_10135);
or U10438 (N_10438,N_10105,N_10174);
or U10439 (N_10439,N_10014,N_10243);
nor U10440 (N_10440,N_10102,N_10042);
and U10441 (N_10441,N_10231,N_10127);
nand U10442 (N_10442,N_10225,N_10148);
nor U10443 (N_10443,N_10123,N_10189);
nand U10444 (N_10444,N_10104,N_10112);
nand U10445 (N_10445,N_10117,N_10185);
and U10446 (N_10446,N_10038,N_10080);
nand U10447 (N_10447,N_10000,N_10062);
nor U10448 (N_10448,N_10147,N_10068);
or U10449 (N_10449,N_10210,N_10066);
or U10450 (N_10450,N_10194,N_10086);
nand U10451 (N_10451,N_10131,N_10220);
and U10452 (N_10452,N_10203,N_10207);
or U10453 (N_10453,N_10201,N_10004);
or U10454 (N_10454,N_10166,N_10081);
or U10455 (N_10455,N_10139,N_10081);
nand U10456 (N_10456,N_10127,N_10169);
nand U10457 (N_10457,N_10050,N_10232);
or U10458 (N_10458,N_10020,N_10132);
or U10459 (N_10459,N_10133,N_10249);
nor U10460 (N_10460,N_10060,N_10175);
or U10461 (N_10461,N_10101,N_10172);
nor U10462 (N_10462,N_10232,N_10170);
or U10463 (N_10463,N_10009,N_10006);
nand U10464 (N_10464,N_10062,N_10149);
nand U10465 (N_10465,N_10033,N_10145);
xor U10466 (N_10466,N_10227,N_10235);
nand U10467 (N_10467,N_10006,N_10088);
nand U10468 (N_10468,N_10137,N_10035);
xor U10469 (N_10469,N_10014,N_10092);
nor U10470 (N_10470,N_10018,N_10031);
and U10471 (N_10471,N_10204,N_10245);
xnor U10472 (N_10472,N_10135,N_10208);
or U10473 (N_10473,N_10188,N_10010);
or U10474 (N_10474,N_10118,N_10235);
nor U10475 (N_10475,N_10142,N_10146);
and U10476 (N_10476,N_10055,N_10165);
nor U10477 (N_10477,N_10106,N_10100);
nand U10478 (N_10478,N_10173,N_10038);
nor U10479 (N_10479,N_10094,N_10039);
and U10480 (N_10480,N_10018,N_10207);
nand U10481 (N_10481,N_10137,N_10079);
and U10482 (N_10482,N_10156,N_10003);
or U10483 (N_10483,N_10123,N_10129);
nand U10484 (N_10484,N_10126,N_10038);
nor U10485 (N_10485,N_10006,N_10024);
and U10486 (N_10486,N_10149,N_10133);
and U10487 (N_10487,N_10075,N_10072);
nor U10488 (N_10488,N_10106,N_10166);
xor U10489 (N_10489,N_10001,N_10226);
or U10490 (N_10490,N_10209,N_10047);
or U10491 (N_10491,N_10059,N_10244);
or U10492 (N_10492,N_10139,N_10137);
or U10493 (N_10493,N_10165,N_10168);
nor U10494 (N_10494,N_10199,N_10036);
nand U10495 (N_10495,N_10139,N_10061);
and U10496 (N_10496,N_10047,N_10232);
xor U10497 (N_10497,N_10040,N_10075);
nor U10498 (N_10498,N_10024,N_10200);
and U10499 (N_10499,N_10187,N_10141);
nand U10500 (N_10500,N_10462,N_10295);
nor U10501 (N_10501,N_10431,N_10325);
or U10502 (N_10502,N_10358,N_10388);
nor U10503 (N_10503,N_10432,N_10287);
and U10504 (N_10504,N_10414,N_10289);
or U10505 (N_10505,N_10298,N_10486);
nand U10506 (N_10506,N_10300,N_10407);
nor U10507 (N_10507,N_10448,N_10277);
nand U10508 (N_10508,N_10267,N_10485);
xnor U10509 (N_10509,N_10250,N_10257);
or U10510 (N_10510,N_10435,N_10284);
xor U10511 (N_10511,N_10335,N_10276);
xnor U10512 (N_10512,N_10425,N_10312);
nor U10513 (N_10513,N_10401,N_10354);
nand U10514 (N_10514,N_10400,N_10308);
xnor U10515 (N_10515,N_10428,N_10282);
nand U10516 (N_10516,N_10447,N_10382);
or U10517 (N_10517,N_10449,N_10331);
or U10518 (N_10518,N_10473,N_10293);
nor U10519 (N_10519,N_10424,N_10412);
nand U10520 (N_10520,N_10367,N_10252);
nand U10521 (N_10521,N_10436,N_10451);
or U10522 (N_10522,N_10415,N_10341);
nor U10523 (N_10523,N_10319,N_10444);
and U10524 (N_10524,N_10480,N_10345);
nor U10525 (N_10525,N_10366,N_10251);
xnor U10526 (N_10526,N_10453,N_10322);
or U10527 (N_10527,N_10303,N_10306);
and U10528 (N_10528,N_10385,N_10361);
or U10529 (N_10529,N_10334,N_10348);
or U10530 (N_10530,N_10314,N_10391);
nor U10531 (N_10531,N_10405,N_10310);
nand U10532 (N_10532,N_10286,N_10418);
or U10533 (N_10533,N_10378,N_10387);
and U10534 (N_10534,N_10454,N_10346);
and U10535 (N_10535,N_10389,N_10355);
or U10536 (N_10536,N_10321,N_10411);
nor U10537 (N_10537,N_10374,N_10307);
xor U10538 (N_10538,N_10259,N_10492);
and U10539 (N_10539,N_10375,N_10445);
nor U10540 (N_10540,N_10403,N_10317);
nand U10541 (N_10541,N_10397,N_10398);
nor U10542 (N_10542,N_10392,N_10404);
xor U10543 (N_10543,N_10281,N_10433);
and U10544 (N_10544,N_10255,N_10406);
nand U10545 (N_10545,N_10477,N_10373);
xor U10546 (N_10546,N_10461,N_10262);
and U10547 (N_10547,N_10470,N_10402);
and U10548 (N_10548,N_10253,N_10323);
nor U10549 (N_10549,N_10288,N_10377);
nor U10550 (N_10550,N_10313,N_10258);
xnor U10551 (N_10551,N_10429,N_10491);
nor U10552 (N_10552,N_10324,N_10296);
or U10553 (N_10553,N_10343,N_10381);
and U10554 (N_10554,N_10439,N_10496);
nand U10555 (N_10555,N_10338,N_10394);
or U10556 (N_10556,N_10364,N_10426);
nand U10557 (N_10557,N_10350,N_10490);
nor U10558 (N_10558,N_10472,N_10476);
xor U10559 (N_10559,N_10292,N_10395);
or U10560 (N_10560,N_10487,N_10427);
xor U10561 (N_10561,N_10318,N_10423);
and U10562 (N_10562,N_10457,N_10383);
nor U10563 (N_10563,N_10356,N_10344);
or U10564 (N_10564,N_10471,N_10488);
or U10565 (N_10565,N_10459,N_10499);
or U10566 (N_10566,N_10489,N_10290);
nand U10567 (N_10567,N_10379,N_10330);
and U10568 (N_10568,N_10393,N_10422);
nor U10569 (N_10569,N_10437,N_10416);
xnor U10570 (N_10570,N_10328,N_10479);
xor U10571 (N_10571,N_10464,N_10305);
nand U10572 (N_10572,N_10481,N_10498);
nor U10573 (N_10573,N_10261,N_10475);
and U10574 (N_10574,N_10274,N_10482);
nand U10575 (N_10575,N_10336,N_10254);
and U10576 (N_10576,N_10376,N_10302);
nor U10577 (N_10577,N_10369,N_10408);
nand U10578 (N_10578,N_10283,N_10465);
or U10579 (N_10579,N_10271,N_10419);
or U10580 (N_10580,N_10359,N_10452);
nand U10581 (N_10581,N_10463,N_10371);
xnor U10582 (N_10582,N_10458,N_10438);
nor U10583 (N_10583,N_10467,N_10370);
or U10584 (N_10584,N_10413,N_10291);
or U10585 (N_10585,N_10396,N_10316);
or U10586 (N_10586,N_10484,N_10493);
nor U10587 (N_10587,N_10269,N_10256);
or U10588 (N_10588,N_10469,N_10311);
and U10589 (N_10589,N_10478,N_10260);
and U10590 (N_10590,N_10363,N_10420);
nand U10591 (N_10591,N_10266,N_10360);
nand U10592 (N_10592,N_10280,N_10326);
and U10593 (N_10593,N_10309,N_10315);
or U10594 (N_10594,N_10333,N_10263);
or U10595 (N_10595,N_10357,N_10299);
nor U10596 (N_10596,N_10434,N_10399);
and U10597 (N_10597,N_10440,N_10327);
xnor U10598 (N_10598,N_10409,N_10332);
nand U10599 (N_10599,N_10304,N_10368);
or U10600 (N_10600,N_10268,N_10297);
and U10601 (N_10601,N_10442,N_10347);
and U10602 (N_10602,N_10329,N_10380);
or U10603 (N_10603,N_10410,N_10272);
and U10604 (N_10604,N_10441,N_10340);
xor U10605 (N_10605,N_10497,N_10468);
nor U10606 (N_10606,N_10372,N_10384);
xor U10607 (N_10607,N_10365,N_10430);
and U10608 (N_10608,N_10349,N_10294);
or U10609 (N_10609,N_10264,N_10450);
xor U10610 (N_10610,N_10320,N_10417);
nand U10611 (N_10611,N_10273,N_10362);
or U10612 (N_10612,N_10421,N_10342);
nor U10613 (N_10613,N_10494,N_10386);
and U10614 (N_10614,N_10446,N_10495);
nor U10615 (N_10615,N_10460,N_10278);
and U10616 (N_10616,N_10353,N_10455);
nor U10617 (N_10617,N_10456,N_10270);
and U10618 (N_10618,N_10351,N_10337);
xnor U10619 (N_10619,N_10301,N_10339);
and U10620 (N_10620,N_10466,N_10474);
nand U10621 (N_10621,N_10275,N_10279);
xor U10622 (N_10622,N_10483,N_10265);
nor U10623 (N_10623,N_10443,N_10352);
nand U10624 (N_10624,N_10390,N_10285);
nor U10625 (N_10625,N_10353,N_10334);
or U10626 (N_10626,N_10267,N_10268);
nor U10627 (N_10627,N_10427,N_10433);
nor U10628 (N_10628,N_10290,N_10341);
xnor U10629 (N_10629,N_10409,N_10410);
nor U10630 (N_10630,N_10265,N_10346);
and U10631 (N_10631,N_10291,N_10295);
xor U10632 (N_10632,N_10263,N_10271);
nor U10633 (N_10633,N_10297,N_10358);
xnor U10634 (N_10634,N_10273,N_10354);
nand U10635 (N_10635,N_10460,N_10366);
and U10636 (N_10636,N_10488,N_10484);
and U10637 (N_10637,N_10414,N_10353);
or U10638 (N_10638,N_10405,N_10460);
nand U10639 (N_10639,N_10462,N_10264);
or U10640 (N_10640,N_10285,N_10434);
xor U10641 (N_10641,N_10444,N_10455);
and U10642 (N_10642,N_10358,N_10255);
nor U10643 (N_10643,N_10477,N_10347);
nand U10644 (N_10644,N_10317,N_10288);
xor U10645 (N_10645,N_10454,N_10288);
or U10646 (N_10646,N_10276,N_10413);
xnor U10647 (N_10647,N_10258,N_10301);
or U10648 (N_10648,N_10327,N_10438);
or U10649 (N_10649,N_10448,N_10461);
and U10650 (N_10650,N_10257,N_10457);
and U10651 (N_10651,N_10349,N_10250);
nor U10652 (N_10652,N_10308,N_10262);
or U10653 (N_10653,N_10474,N_10382);
or U10654 (N_10654,N_10274,N_10336);
and U10655 (N_10655,N_10342,N_10451);
nand U10656 (N_10656,N_10400,N_10352);
or U10657 (N_10657,N_10438,N_10309);
and U10658 (N_10658,N_10409,N_10362);
or U10659 (N_10659,N_10371,N_10342);
nand U10660 (N_10660,N_10394,N_10474);
or U10661 (N_10661,N_10430,N_10450);
xor U10662 (N_10662,N_10496,N_10443);
nor U10663 (N_10663,N_10449,N_10315);
and U10664 (N_10664,N_10485,N_10269);
or U10665 (N_10665,N_10263,N_10491);
and U10666 (N_10666,N_10301,N_10400);
xnor U10667 (N_10667,N_10429,N_10485);
and U10668 (N_10668,N_10464,N_10477);
and U10669 (N_10669,N_10422,N_10401);
nor U10670 (N_10670,N_10292,N_10447);
and U10671 (N_10671,N_10479,N_10281);
nor U10672 (N_10672,N_10464,N_10279);
nand U10673 (N_10673,N_10444,N_10313);
and U10674 (N_10674,N_10423,N_10478);
or U10675 (N_10675,N_10424,N_10487);
xnor U10676 (N_10676,N_10404,N_10432);
or U10677 (N_10677,N_10422,N_10445);
xnor U10678 (N_10678,N_10476,N_10345);
and U10679 (N_10679,N_10363,N_10285);
and U10680 (N_10680,N_10308,N_10493);
nand U10681 (N_10681,N_10392,N_10332);
and U10682 (N_10682,N_10273,N_10499);
nand U10683 (N_10683,N_10460,N_10395);
nor U10684 (N_10684,N_10275,N_10299);
nor U10685 (N_10685,N_10283,N_10432);
and U10686 (N_10686,N_10454,N_10360);
or U10687 (N_10687,N_10378,N_10328);
nand U10688 (N_10688,N_10384,N_10485);
nand U10689 (N_10689,N_10333,N_10471);
nor U10690 (N_10690,N_10265,N_10287);
nor U10691 (N_10691,N_10402,N_10393);
and U10692 (N_10692,N_10390,N_10397);
xnor U10693 (N_10693,N_10276,N_10362);
and U10694 (N_10694,N_10489,N_10389);
and U10695 (N_10695,N_10395,N_10302);
nand U10696 (N_10696,N_10316,N_10416);
xnor U10697 (N_10697,N_10258,N_10260);
or U10698 (N_10698,N_10482,N_10464);
nand U10699 (N_10699,N_10432,N_10477);
nor U10700 (N_10700,N_10323,N_10465);
or U10701 (N_10701,N_10361,N_10353);
or U10702 (N_10702,N_10450,N_10370);
nand U10703 (N_10703,N_10433,N_10316);
xnor U10704 (N_10704,N_10386,N_10419);
and U10705 (N_10705,N_10450,N_10445);
nor U10706 (N_10706,N_10485,N_10441);
or U10707 (N_10707,N_10467,N_10395);
xor U10708 (N_10708,N_10298,N_10279);
and U10709 (N_10709,N_10301,N_10465);
or U10710 (N_10710,N_10407,N_10484);
or U10711 (N_10711,N_10266,N_10476);
nand U10712 (N_10712,N_10264,N_10312);
nor U10713 (N_10713,N_10293,N_10263);
nor U10714 (N_10714,N_10359,N_10342);
or U10715 (N_10715,N_10434,N_10352);
xor U10716 (N_10716,N_10485,N_10338);
or U10717 (N_10717,N_10416,N_10490);
nand U10718 (N_10718,N_10364,N_10322);
xnor U10719 (N_10719,N_10347,N_10344);
or U10720 (N_10720,N_10294,N_10311);
nor U10721 (N_10721,N_10284,N_10462);
nand U10722 (N_10722,N_10258,N_10366);
xor U10723 (N_10723,N_10446,N_10317);
nand U10724 (N_10724,N_10251,N_10309);
or U10725 (N_10725,N_10269,N_10460);
xor U10726 (N_10726,N_10484,N_10363);
nor U10727 (N_10727,N_10437,N_10380);
and U10728 (N_10728,N_10446,N_10337);
nor U10729 (N_10729,N_10347,N_10260);
and U10730 (N_10730,N_10479,N_10310);
nand U10731 (N_10731,N_10289,N_10360);
nor U10732 (N_10732,N_10349,N_10350);
and U10733 (N_10733,N_10413,N_10345);
xor U10734 (N_10734,N_10301,N_10375);
nand U10735 (N_10735,N_10322,N_10398);
xor U10736 (N_10736,N_10299,N_10398);
or U10737 (N_10737,N_10464,N_10334);
or U10738 (N_10738,N_10465,N_10483);
or U10739 (N_10739,N_10329,N_10356);
or U10740 (N_10740,N_10335,N_10413);
nor U10741 (N_10741,N_10439,N_10411);
nand U10742 (N_10742,N_10441,N_10368);
or U10743 (N_10743,N_10359,N_10472);
nor U10744 (N_10744,N_10377,N_10391);
nor U10745 (N_10745,N_10273,N_10295);
xor U10746 (N_10746,N_10314,N_10485);
and U10747 (N_10747,N_10322,N_10301);
xnor U10748 (N_10748,N_10463,N_10384);
nor U10749 (N_10749,N_10490,N_10420);
nor U10750 (N_10750,N_10638,N_10581);
xor U10751 (N_10751,N_10680,N_10624);
xor U10752 (N_10752,N_10658,N_10704);
and U10753 (N_10753,N_10571,N_10747);
nand U10754 (N_10754,N_10739,N_10625);
or U10755 (N_10755,N_10531,N_10661);
nand U10756 (N_10756,N_10708,N_10699);
nor U10757 (N_10757,N_10645,N_10698);
and U10758 (N_10758,N_10582,N_10735);
xnor U10759 (N_10759,N_10605,N_10722);
xor U10760 (N_10760,N_10578,N_10682);
or U10761 (N_10761,N_10541,N_10547);
or U10762 (N_10762,N_10600,N_10542);
xor U10763 (N_10763,N_10595,N_10672);
xor U10764 (N_10764,N_10715,N_10709);
xor U10765 (N_10765,N_10586,N_10726);
xnor U10766 (N_10766,N_10730,N_10617);
or U10767 (N_10767,N_10639,N_10630);
nand U10768 (N_10768,N_10740,N_10669);
and U10769 (N_10769,N_10681,N_10685);
xnor U10770 (N_10770,N_10666,N_10599);
nor U10771 (N_10771,N_10532,N_10543);
nand U10772 (N_10772,N_10559,N_10626);
and U10773 (N_10773,N_10741,N_10511);
or U10774 (N_10774,N_10662,N_10513);
nand U10775 (N_10775,N_10644,N_10696);
nor U10776 (N_10776,N_10728,N_10727);
and U10777 (N_10777,N_10703,N_10505);
nor U10778 (N_10778,N_10620,N_10663);
nor U10779 (N_10779,N_10636,N_10604);
and U10780 (N_10780,N_10554,N_10563);
and U10781 (N_10781,N_10594,N_10634);
nand U10782 (N_10782,N_10652,N_10635);
xnor U10783 (N_10783,N_10549,N_10508);
nor U10784 (N_10784,N_10688,N_10621);
nor U10785 (N_10785,N_10514,N_10623);
or U10786 (N_10786,N_10517,N_10567);
and U10787 (N_10787,N_10614,N_10520);
nand U10788 (N_10788,N_10647,N_10646);
or U10789 (N_10789,N_10712,N_10710);
nand U10790 (N_10790,N_10526,N_10673);
nor U10791 (N_10791,N_10684,N_10707);
and U10792 (N_10792,N_10743,N_10602);
and U10793 (N_10793,N_10558,N_10568);
xnor U10794 (N_10794,N_10535,N_10603);
nand U10795 (N_10795,N_10628,N_10540);
or U10796 (N_10796,N_10742,N_10748);
nand U10797 (N_10797,N_10731,N_10653);
and U10798 (N_10798,N_10702,N_10587);
and U10799 (N_10799,N_10598,N_10637);
nand U10800 (N_10800,N_10577,N_10544);
xnor U10801 (N_10801,N_10711,N_10575);
xnor U10802 (N_10802,N_10631,N_10590);
or U10803 (N_10803,N_10525,N_10537);
nor U10804 (N_10804,N_10700,N_10725);
nor U10805 (N_10805,N_10523,N_10665);
nor U10806 (N_10806,N_10601,N_10713);
nor U10807 (N_10807,N_10534,N_10503);
nor U10808 (N_10808,N_10643,N_10689);
xor U10809 (N_10809,N_10649,N_10611);
nand U10810 (N_10810,N_10576,N_10619);
or U10811 (N_10811,N_10719,N_10548);
or U10812 (N_10812,N_10519,N_10550);
nand U10813 (N_10813,N_10717,N_10580);
and U10814 (N_10814,N_10648,N_10524);
nand U10815 (N_10815,N_10610,N_10509);
or U10816 (N_10816,N_10512,N_10705);
nand U10817 (N_10817,N_10687,N_10676);
nor U10818 (N_10818,N_10612,N_10627);
nor U10819 (N_10819,N_10695,N_10588);
xor U10820 (N_10820,N_10527,N_10596);
or U10821 (N_10821,N_10608,N_10690);
and U10822 (N_10822,N_10570,N_10655);
nand U10823 (N_10823,N_10716,N_10516);
or U10824 (N_10824,N_10553,N_10555);
xor U10825 (N_10825,N_10538,N_10664);
nor U10826 (N_10826,N_10723,N_10574);
or U10827 (N_10827,N_10675,N_10736);
nand U10828 (N_10828,N_10515,N_10733);
and U10829 (N_10829,N_10502,N_10691);
or U10830 (N_10830,N_10651,N_10592);
and U10831 (N_10831,N_10654,N_10714);
nand U10832 (N_10832,N_10668,N_10724);
nand U10833 (N_10833,N_10583,N_10607);
nand U10834 (N_10834,N_10706,N_10674);
or U10835 (N_10835,N_10679,N_10545);
or U10836 (N_10836,N_10530,N_10718);
or U10837 (N_10837,N_10616,N_10501);
or U10838 (N_10838,N_10734,N_10609);
nor U10839 (N_10839,N_10539,N_10678);
nor U10840 (N_10840,N_10642,N_10506);
xnor U10841 (N_10841,N_10591,N_10650);
xnor U10842 (N_10842,N_10572,N_10660);
and U10843 (N_10843,N_10677,N_10618);
or U10844 (N_10844,N_10615,N_10640);
and U10845 (N_10845,N_10613,N_10552);
or U10846 (N_10846,N_10504,N_10507);
and U10847 (N_10847,N_10671,N_10729);
nor U10848 (N_10848,N_10584,N_10686);
xnor U10849 (N_10849,N_10749,N_10697);
and U10850 (N_10850,N_10683,N_10597);
or U10851 (N_10851,N_10629,N_10529);
xor U10852 (N_10852,N_10657,N_10561);
xnor U10853 (N_10853,N_10641,N_10556);
or U10854 (N_10854,N_10565,N_10573);
and U10855 (N_10855,N_10633,N_10500);
nand U10856 (N_10856,N_10528,N_10701);
nor U10857 (N_10857,N_10737,N_10546);
and U10858 (N_10858,N_10694,N_10557);
and U10859 (N_10859,N_10510,N_10522);
xor U10860 (N_10860,N_10656,N_10670);
xor U10861 (N_10861,N_10585,N_10518);
and U10862 (N_10862,N_10745,N_10593);
or U10863 (N_10863,N_10521,N_10744);
nor U10864 (N_10864,N_10566,N_10569);
and U10865 (N_10865,N_10746,N_10693);
xor U10866 (N_10866,N_10721,N_10533);
and U10867 (N_10867,N_10632,N_10667);
or U10868 (N_10868,N_10589,N_10564);
xor U10869 (N_10869,N_10659,N_10551);
nand U10870 (N_10870,N_10606,N_10562);
nor U10871 (N_10871,N_10536,N_10732);
nand U10872 (N_10872,N_10560,N_10579);
nor U10873 (N_10873,N_10622,N_10692);
and U10874 (N_10874,N_10720,N_10738);
xnor U10875 (N_10875,N_10516,N_10724);
nand U10876 (N_10876,N_10639,N_10567);
and U10877 (N_10877,N_10653,N_10522);
or U10878 (N_10878,N_10560,N_10710);
nand U10879 (N_10879,N_10609,N_10616);
xor U10880 (N_10880,N_10662,N_10718);
nor U10881 (N_10881,N_10525,N_10545);
nand U10882 (N_10882,N_10656,N_10619);
or U10883 (N_10883,N_10643,N_10626);
nor U10884 (N_10884,N_10576,N_10675);
and U10885 (N_10885,N_10692,N_10600);
and U10886 (N_10886,N_10560,N_10561);
nor U10887 (N_10887,N_10546,N_10703);
nor U10888 (N_10888,N_10737,N_10568);
and U10889 (N_10889,N_10569,N_10542);
and U10890 (N_10890,N_10629,N_10617);
nand U10891 (N_10891,N_10557,N_10567);
and U10892 (N_10892,N_10690,N_10549);
nand U10893 (N_10893,N_10559,N_10608);
and U10894 (N_10894,N_10511,N_10502);
nor U10895 (N_10895,N_10652,N_10738);
and U10896 (N_10896,N_10545,N_10701);
or U10897 (N_10897,N_10669,N_10569);
nor U10898 (N_10898,N_10676,N_10642);
xnor U10899 (N_10899,N_10610,N_10573);
xor U10900 (N_10900,N_10644,N_10532);
xor U10901 (N_10901,N_10548,N_10522);
or U10902 (N_10902,N_10711,N_10678);
nor U10903 (N_10903,N_10725,N_10741);
and U10904 (N_10904,N_10550,N_10746);
xnor U10905 (N_10905,N_10551,N_10708);
nand U10906 (N_10906,N_10724,N_10635);
xor U10907 (N_10907,N_10580,N_10543);
or U10908 (N_10908,N_10698,N_10614);
nor U10909 (N_10909,N_10705,N_10523);
xor U10910 (N_10910,N_10541,N_10539);
xnor U10911 (N_10911,N_10618,N_10746);
or U10912 (N_10912,N_10645,N_10676);
nand U10913 (N_10913,N_10511,N_10668);
or U10914 (N_10914,N_10691,N_10571);
nor U10915 (N_10915,N_10514,N_10630);
and U10916 (N_10916,N_10743,N_10616);
and U10917 (N_10917,N_10591,N_10680);
and U10918 (N_10918,N_10644,N_10702);
nand U10919 (N_10919,N_10500,N_10648);
nor U10920 (N_10920,N_10712,N_10552);
and U10921 (N_10921,N_10615,N_10516);
and U10922 (N_10922,N_10566,N_10645);
nor U10923 (N_10923,N_10606,N_10726);
and U10924 (N_10924,N_10610,N_10639);
or U10925 (N_10925,N_10555,N_10695);
or U10926 (N_10926,N_10608,N_10745);
nand U10927 (N_10927,N_10531,N_10712);
xor U10928 (N_10928,N_10500,N_10697);
or U10929 (N_10929,N_10546,N_10600);
nand U10930 (N_10930,N_10542,N_10583);
and U10931 (N_10931,N_10696,N_10619);
and U10932 (N_10932,N_10620,N_10695);
nor U10933 (N_10933,N_10510,N_10537);
nand U10934 (N_10934,N_10737,N_10506);
nand U10935 (N_10935,N_10616,N_10515);
or U10936 (N_10936,N_10561,N_10619);
nor U10937 (N_10937,N_10537,N_10711);
and U10938 (N_10938,N_10684,N_10625);
nand U10939 (N_10939,N_10736,N_10686);
xnor U10940 (N_10940,N_10584,N_10579);
or U10941 (N_10941,N_10525,N_10665);
nor U10942 (N_10942,N_10575,N_10739);
xor U10943 (N_10943,N_10603,N_10542);
xor U10944 (N_10944,N_10615,N_10581);
or U10945 (N_10945,N_10500,N_10649);
nor U10946 (N_10946,N_10685,N_10712);
xor U10947 (N_10947,N_10739,N_10543);
or U10948 (N_10948,N_10624,N_10746);
nor U10949 (N_10949,N_10697,N_10650);
nor U10950 (N_10950,N_10703,N_10711);
nor U10951 (N_10951,N_10555,N_10581);
nor U10952 (N_10952,N_10568,N_10684);
nor U10953 (N_10953,N_10576,N_10643);
and U10954 (N_10954,N_10641,N_10609);
nor U10955 (N_10955,N_10550,N_10620);
or U10956 (N_10956,N_10501,N_10592);
nor U10957 (N_10957,N_10721,N_10527);
nor U10958 (N_10958,N_10579,N_10660);
nand U10959 (N_10959,N_10688,N_10568);
nand U10960 (N_10960,N_10655,N_10639);
and U10961 (N_10961,N_10546,N_10542);
xnor U10962 (N_10962,N_10509,N_10660);
and U10963 (N_10963,N_10607,N_10501);
nand U10964 (N_10964,N_10692,N_10519);
and U10965 (N_10965,N_10739,N_10694);
nand U10966 (N_10966,N_10681,N_10743);
and U10967 (N_10967,N_10519,N_10564);
nor U10968 (N_10968,N_10531,N_10555);
xnor U10969 (N_10969,N_10718,N_10697);
nor U10970 (N_10970,N_10715,N_10727);
nor U10971 (N_10971,N_10598,N_10587);
nand U10972 (N_10972,N_10641,N_10722);
nand U10973 (N_10973,N_10624,N_10721);
nor U10974 (N_10974,N_10697,N_10603);
nor U10975 (N_10975,N_10537,N_10542);
and U10976 (N_10976,N_10699,N_10531);
xor U10977 (N_10977,N_10659,N_10680);
nand U10978 (N_10978,N_10663,N_10527);
nand U10979 (N_10979,N_10549,N_10717);
nor U10980 (N_10980,N_10588,N_10500);
nand U10981 (N_10981,N_10746,N_10716);
or U10982 (N_10982,N_10649,N_10505);
nor U10983 (N_10983,N_10734,N_10667);
or U10984 (N_10984,N_10654,N_10692);
and U10985 (N_10985,N_10553,N_10559);
xnor U10986 (N_10986,N_10630,N_10554);
xor U10987 (N_10987,N_10711,N_10521);
and U10988 (N_10988,N_10749,N_10698);
nor U10989 (N_10989,N_10617,N_10561);
nor U10990 (N_10990,N_10526,N_10729);
nor U10991 (N_10991,N_10516,N_10672);
nand U10992 (N_10992,N_10687,N_10721);
nor U10993 (N_10993,N_10504,N_10599);
or U10994 (N_10994,N_10665,N_10609);
nand U10995 (N_10995,N_10612,N_10537);
or U10996 (N_10996,N_10738,N_10677);
nor U10997 (N_10997,N_10711,N_10524);
xor U10998 (N_10998,N_10660,N_10523);
nor U10999 (N_10999,N_10507,N_10563);
and U11000 (N_11000,N_10794,N_10990);
xnor U11001 (N_11001,N_10804,N_10833);
xor U11002 (N_11002,N_10974,N_10819);
nand U11003 (N_11003,N_10936,N_10762);
or U11004 (N_11004,N_10820,N_10981);
xor U11005 (N_11005,N_10834,N_10816);
or U11006 (N_11006,N_10867,N_10785);
nor U11007 (N_11007,N_10971,N_10943);
and U11008 (N_11008,N_10826,N_10975);
and U11009 (N_11009,N_10821,N_10907);
xnor U11010 (N_11010,N_10814,N_10933);
or U11011 (N_11011,N_10817,N_10830);
nor U11012 (N_11012,N_10846,N_10925);
nor U11013 (N_11013,N_10866,N_10876);
nand U11014 (N_11014,N_10859,N_10945);
or U11015 (N_11015,N_10844,N_10827);
nand U11016 (N_11016,N_10849,N_10960);
nand U11017 (N_11017,N_10966,N_10767);
xor U11018 (N_11018,N_10803,N_10951);
nand U11019 (N_11019,N_10777,N_10993);
nand U11020 (N_11020,N_10940,N_10939);
and U11021 (N_11021,N_10902,N_10929);
nor U11022 (N_11022,N_10901,N_10930);
or U11023 (N_11023,N_10841,N_10786);
nor U11024 (N_11024,N_10835,N_10875);
or U11025 (N_11025,N_10838,N_10905);
nand U11026 (N_11026,N_10997,N_10904);
nand U11027 (N_11027,N_10917,N_10825);
or U11028 (N_11028,N_10967,N_10832);
xor U11029 (N_11029,N_10949,N_10758);
or U11030 (N_11030,N_10801,N_10999);
and U11031 (N_11031,N_10870,N_10822);
nand U11032 (N_11032,N_10934,N_10815);
nand U11033 (N_11033,N_10800,N_10784);
or U11034 (N_11034,N_10911,N_10855);
nand U11035 (N_11035,N_10884,N_10813);
xnor U11036 (N_11036,N_10985,N_10980);
or U11037 (N_11037,N_10845,N_10941);
xnor U11038 (N_11038,N_10984,N_10898);
nor U11039 (N_11039,N_10989,N_10824);
xnor U11040 (N_11040,N_10788,N_10897);
xnor U11041 (N_11041,N_10969,N_10783);
nand U11042 (N_11042,N_10995,N_10873);
or U11043 (N_11043,N_10903,N_10948);
or U11044 (N_11044,N_10922,N_10836);
xor U11045 (N_11045,N_10955,N_10893);
and U11046 (N_11046,N_10802,N_10991);
nor U11047 (N_11047,N_10896,N_10750);
and U11048 (N_11048,N_10760,N_10938);
or U11049 (N_11049,N_10973,N_10850);
xnor U11050 (N_11050,N_10775,N_10842);
nand U11051 (N_11051,N_10914,N_10753);
nand U11052 (N_11052,N_10912,N_10976);
nand U11053 (N_11053,N_10840,N_10772);
nor U11054 (N_11054,N_10810,N_10755);
nor U11055 (N_11055,N_10769,N_10751);
xor U11056 (N_11056,N_10868,N_10871);
nand U11057 (N_11057,N_10890,N_10956);
and U11058 (N_11058,N_10831,N_10878);
or U11059 (N_11059,N_10752,N_10920);
nand U11060 (N_11060,N_10950,N_10952);
and U11061 (N_11061,N_10795,N_10858);
and U11062 (N_11062,N_10906,N_10774);
or U11063 (N_11063,N_10926,N_10857);
nor U11064 (N_11064,N_10910,N_10860);
or U11065 (N_11065,N_10882,N_10970);
nor U11066 (N_11066,N_10927,N_10759);
nand U11067 (N_11067,N_10895,N_10765);
nand U11068 (N_11068,N_10796,N_10894);
nand U11069 (N_11069,N_10880,N_10961);
or U11070 (N_11070,N_10754,N_10812);
and U11071 (N_11071,N_10965,N_10928);
and U11072 (N_11072,N_10761,N_10983);
or U11073 (N_11073,N_10996,N_10916);
nor U11074 (N_11074,N_10944,N_10856);
nand U11075 (N_11075,N_10918,N_10942);
nand U11076 (N_11076,N_10828,N_10768);
xnor U11077 (N_11077,N_10978,N_10865);
and U11078 (N_11078,N_10988,N_10776);
nor U11079 (N_11079,N_10771,N_10964);
and U11080 (N_11080,N_10924,N_10848);
xnor U11081 (N_11081,N_10839,N_10998);
and U11082 (N_11082,N_10992,N_10883);
nand U11083 (N_11083,N_10770,N_10935);
nand U11084 (N_11084,N_10915,N_10958);
xnor U11085 (N_11085,N_10852,N_10874);
nor U11086 (N_11086,N_10766,N_10888);
or U11087 (N_11087,N_10863,N_10909);
xor U11088 (N_11088,N_10847,N_10864);
or U11089 (N_11089,N_10778,N_10986);
and U11090 (N_11090,N_10879,N_10877);
or U11091 (N_11091,N_10982,N_10932);
nor U11092 (N_11092,N_10799,N_10843);
nand U11093 (N_11093,N_10931,N_10886);
and U11094 (N_11094,N_10963,N_10946);
or U11095 (N_11095,N_10793,N_10881);
and U11096 (N_11096,N_10962,N_10891);
xnor U11097 (N_11097,N_10790,N_10862);
xnor U11098 (N_11098,N_10829,N_10763);
nand U11099 (N_11099,N_10807,N_10947);
or U11100 (N_11100,N_10954,N_10957);
nand U11101 (N_11101,N_10837,N_10764);
or U11102 (N_11102,N_10851,N_10809);
nor U11103 (N_11103,N_10811,N_10861);
nand U11104 (N_11104,N_10923,N_10805);
nor U11105 (N_11105,N_10853,N_10780);
nand U11106 (N_11106,N_10885,N_10977);
and U11107 (N_11107,N_10937,N_10968);
or U11108 (N_11108,N_10869,N_10791);
and U11109 (N_11109,N_10921,N_10773);
or U11110 (N_11110,N_10757,N_10913);
or U11111 (N_11111,N_10854,N_10782);
or U11112 (N_11112,N_10779,N_10756);
nand U11113 (N_11113,N_10919,N_10889);
and U11114 (N_11114,N_10787,N_10887);
xor U11115 (N_11115,N_10892,N_10953);
and U11116 (N_11116,N_10908,N_10900);
and U11117 (N_11117,N_10899,N_10808);
and U11118 (N_11118,N_10872,N_10798);
and U11119 (N_11119,N_10987,N_10797);
or U11120 (N_11120,N_10823,N_10959);
nand U11121 (N_11121,N_10972,N_10806);
and U11122 (N_11122,N_10979,N_10789);
nor U11123 (N_11123,N_10792,N_10818);
nand U11124 (N_11124,N_10994,N_10781);
nand U11125 (N_11125,N_10830,N_10865);
nand U11126 (N_11126,N_10762,N_10799);
nand U11127 (N_11127,N_10772,N_10997);
and U11128 (N_11128,N_10907,N_10884);
xnor U11129 (N_11129,N_10815,N_10975);
or U11130 (N_11130,N_10917,N_10971);
nor U11131 (N_11131,N_10855,N_10983);
nor U11132 (N_11132,N_10908,N_10994);
xor U11133 (N_11133,N_10929,N_10982);
and U11134 (N_11134,N_10993,N_10753);
or U11135 (N_11135,N_10756,N_10864);
or U11136 (N_11136,N_10975,N_10978);
or U11137 (N_11137,N_10990,N_10889);
nor U11138 (N_11138,N_10834,N_10798);
xor U11139 (N_11139,N_10809,N_10885);
nor U11140 (N_11140,N_10871,N_10794);
or U11141 (N_11141,N_10858,N_10903);
and U11142 (N_11142,N_10940,N_10985);
nor U11143 (N_11143,N_10859,N_10772);
xor U11144 (N_11144,N_10817,N_10994);
and U11145 (N_11145,N_10879,N_10970);
or U11146 (N_11146,N_10896,N_10946);
and U11147 (N_11147,N_10921,N_10809);
nor U11148 (N_11148,N_10751,N_10966);
and U11149 (N_11149,N_10922,N_10832);
and U11150 (N_11150,N_10814,N_10982);
nand U11151 (N_11151,N_10761,N_10847);
or U11152 (N_11152,N_10955,N_10843);
nor U11153 (N_11153,N_10891,N_10902);
or U11154 (N_11154,N_10820,N_10750);
and U11155 (N_11155,N_10821,N_10916);
nor U11156 (N_11156,N_10762,N_10848);
and U11157 (N_11157,N_10808,N_10809);
or U11158 (N_11158,N_10954,N_10979);
nand U11159 (N_11159,N_10942,N_10970);
xor U11160 (N_11160,N_10774,N_10898);
nand U11161 (N_11161,N_10792,N_10864);
and U11162 (N_11162,N_10894,N_10965);
nand U11163 (N_11163,N_10955,N_10979);
and U11164 (N_11164,N_10972,N_10915);
xor U11165 (N_11165,N_10938,N_10849);
nand U11166 (N_11166,N_10913,N_10841);
nand U11167 (N_11167,N_10825,N_10822);
nand U11168 (N_11168,N_10771,N_10873);
nor U11169 (N_11169,N_10989,N_10785);
nor U11170 (N_11170,N_10894,N_10832);
and U11171 (N_11171,N_10922,N_10888);
and U11172 (N_11172,N_10774,N_10961);
xor U11173 (N_11173,N_10905,N_10971);
nand U11174 (N_11174,N_10920,N_10895);
xnor U11175 (N_11175,N_10874,N_10903);
or U11176 (N_11176,N_10827,N_10892);
or U11177 (N_11177,N_10765,N_10976);
or U11178 (N_11178,N_10816,N_10893);
nand U11179 (N_11179,N_10898,N_10750);
xor U11180 (N_11180,N_10782,N_10967);
xor U11181 (N_11181,N_10992,N_10813);
xor U11182 (N_11182,N_10963,N_10926);
xor U11183 (N_11183,N_10757,N_10788);
and U11184 (N_11184,N_10840,N_10962);
or U11185 (N_11185,N_10868,N_10759);
and U11186 (N_11186,N_10839,N_10965);
and U11187 (N_11187,N_10853,N_10916);
or U11188 (N_11188,N_10759,N_10804);
nand U11189 (N_11189,N_10905,N_10963);
and U11190 (N_11190,N_10922,N_10840);
nor U11191 (N_11191,N_10843,N_10860);
nand U11192 (N_11192,N_10871,N_10770);
xnor U11193 (N_11193,N_10873,N_10918);
nor U11194 (N_11194,N_10812,N_10941);
or U11195 (N_11195,N_10894,N_10798);
xnor U11196 (N_11196,N_10798,N_10881);
nor U11197 (N_11197,N_10969,N_10914);
or U11198 (N_11198,N_10802,N_10941);
and U11199 (N_11199,N_10885,N_10926);
or U11200 (N_11200,N_10862,N_10821);
or U11201 (N_11201,N_10938,N_10895);
nand U11202 (N_11202,N_10870,N_10821);
and U11203 (N_11203,N_10861,N_10840);
nor U11204 (N_11204,N_10791,N_10996);
nor U11205 (N_11205,N_10809,N_10811);
and U11206 (N_11206,N_10824,N_10872);
and U11207 (N_11207,N_10998,N_10901);
or U11208 (N_11208,N_10884,N_10810);
nor U11209 (N_11209,N_10769,N_10772);
xor U11210 (N_11210,N_10754,N_10976);
and U11211 (N_11211,N_10900,N_10782);
and U11212 (N_11212,N_10928,N_10890);
nand U11213 (N_11213,N_10883,N_10983);
nand U11214 (N_11214,N_10980,N_10956);
nand U11215 (N_11215,N_10767,N_10773);
or U11216 (N_11216,N_10762,N_10885);
or U11217 (N_11217,N_10853,N_10859);
xnor U11218 (N_11218,N_10868,N_10977);
nand U11219 (N_11219,N_10854,N_10861);
nand U11220 (N_11220,N_10777,N_10959);
or U11221 (N_11221,N_10932,N_10971);
nand U11222 (N_11222,N_10867,N_10830);
and U11223 (N_11223,N_10815,N_10907);
or U11224 (N_11224,N_10809,N_10821);
and U11225 (N_11225,N_10827,N_10889);
nor U11226 (N_11226,N_10814,N_10987);
xnor U11227 (N_11227,N_10965,N_10837);
nor U11228 (N_11228,N_10834,N_10810);
nor U11229 (N_11229,N_10900,N_10935);
nor U11230 (N_11230,N_10839,N_10877);
and U11231 (N_11231,N_10968,N_10876);
nor U11232 (N_11232,N_10908,N_10791);
and U11233 (N_11233,N_10778,N_10926);
xnor U11234 (N_11234,N_10991,N_10926);
nor U11235 (N_11235,N_10751,N_10789);
and U11236 (N_11236,N_10898,N_10965);
nand U11237 (N_11237,N_10890,N_10907);
or U11238 (N_11238,N_10765,N_10910);
or U11239 (N_11239,N_10866,N_10764);
nor U11240 (N_11240,N_10978,N_10863);
nor U11241 (N_11241,N_10795,N_10879);
nor U11242 (N_11242,N_10765,N_10939);
nand U11243 (N_11243,N_10756,N_10871);
xnor U11244 (N_11244,N_10875,N_10978);
nand U11245 (N_11245,N_10936,N_10979);
or U11246 (N_11246,N_10875,N_10916);
or U11247 (N_11247,N_10927,N_10857);
or U11248 (N_11248,N_10894,N_10999);
and U11249 (N_11249,N_10760,N_10848);
xnor U11250 (N_11250,N_11128,N_11088);
xnor U11251 (N_11251,N_11188,N_11075);
and U11252 (N_11252,N_11074,N_11096);
or U11253 (N_11253,N_11005,N_11195);
nand U11254 (N_11254,N_11127,N_11191);
xnor U11255 (N_11255,N_11172,N_11139);
and U11256 (N_11256,N_11019,N_11123);
nor U11257 (N_11257,N_11197,N_11061);
and U11258 (N_11258,N_11109,N_11176);
nand U11259 (N_11259,N_11163,N_11017);
xnor U11260 (N_11260,N_11065,N_11168);
xor U11261 (N_11261,N_11084,N_11090);
xnor U11262 (N_11262,N_11186,N_11080);
xor U11263 (N_11263,N_11102,N_11018);
nand U11264 (N_11264,N_11151,N_11104);
and U11265 (N_11265,N_11094,N_11210);
nand U11266 (N_11266,N_11231,N_11027);
and U11267 (N_11267,N_11241,N_11125);
nor U11268 (N_11268,N_11122,N_11066);
or U11269 (N_11269,N_11047,N_11246);
nor U11270 (N_11270,N_11048,N_11242);
nand U11271 (N_11271,N_11154,N_11085);
and U11272 (N_11272,N_11067,N_11112);
nand U11273 (N_11273,N_11240,N_11069);
and U11274 (N_11274,N_11129,N_11220);
xor U11275 (N_11275,N_11082,N_11032);
and U11276 (N_11276,N_11148,N_11175);
xor U11277 (N_11277,N_11086,N_11223);
nand U11278 (N_11278,N_11189,N_11010);
nor U11279 (N_11279,N_11143,N_11155);
and U11280 (N_11280,N_11092,N_11198);
xor U11281 (N_11281,N_11238,N_11161);
and U11282 (N_11282,N_11239,N_11033);
nor U11283 (N_11283,N_11101,N_11152);
xor U11284 (N_11284,N_11037,N_11056);
and U11285 (N_11285,N_11059,N_11167);
nand U11286 (N_11286,N_11212,N_11170);
xnor U11287 (N_11287,N_11180,N_11157);
nand U11288 (N_11288,N_11034,N_11205);
and U11289 (N_11289,N_11146,N_11221);
nand U11290 (N_11290,N_11029,N_11124);
nor U11291 (N_11291,N_11153,N_11110);
nor U11292 (N_11292,N_11014,N_11055);
and U11293 (N_11293,N_11068,N_11016);
or U11294 (N_11294,N_11095,N_11135);
nor U11295 (N_11295,N_11007,N_11041);
and U11296 (N_11296,N_11162,N_11229);
and U11297 (N_11297,N_11166,N_11036);
xnor U11298 (N_11298,N_11165,N_11156);
xor U11299 (N_11299,N_11012,N_11169);
nand U11300 (N_11300,N_11024,N_11142);
nand U11301 (N_11301,N_11177,N_11228);
or U11302 (N_11302,N_11057,N_11118);
nand U11303 (N_11303,N_11171,N_11051);
and U11304 (N_11304,N_11028,N_11040);
or U11305 (N_11305,N_11131,N_11247);
nand U11306 (N_11306,N_11207,N_11022);
xnor U11307 (N_11307,N_11062,N_11236);
and U11308 (N_11308,N_11244,N_11081);
or U11309 (N_11309,N_11203,N_11216);
nand U11310 (N_11310,N_11204,N_11064);
nor U11311 (N_11311,N_11008,N_11174);
and U11312 (N_11312,N_11181,N_11200);
and U11313 (N_11313,N_11230,N_11083);
xor U11314 (N_11314,N_11179,N_11234);
xnor U11315 (N_11315,N_11249,N_11093);
and U11316 (N_11316,N_11073,N_11183);
or U11317 (N_11317,N_11126,N_11144);
nand U11318 (N_11318,N_11076,N_11091);
and U11319 (N_11319,N_11114,N_11025);
or U11320 (N_11320,N_11020,N_11209);
and U11321 (N_11321,N_11026,N_11190);
and U11322 (N_11322,N_11050,N_11199);
and U11323 (N_11323,N_11023,N_11078);
or U11324 (N_11324,N_11134,N_11053);
and U11325 (N_11325,N_11201,N_11219);
nand U11326 (N_11326,N_11087,N_11117);
nand U11327 (N_11327,N_11098,N_11141);
and U11328 (N_11328,N_11235,N_11009);
or U11329 (N_11329,N_11149,N_11206);
and U11330 (N_11330,N_11079,N_11248);
nor U11331 (N_11331,N_11196,N_11213);
and U11332 (N_11332,N_11077,N_11097);
nand U11333 (N_11333,N_11105,N_11035);
nand U11334 (N_11334,N_11136,N_11211);
nand U11335 (N_11335,N_11138,N_11044);
nand U11336 (N_11336,N_11237,N_11232);
nand U11337 (N_11337,N_11130,N_11021);
nand U11338 (N_11338,N_11039,N_11063);
and U11339 (N_11339,N_11115,N_11045);
xnor U11340 (N_11340,N_11222,N_11160);
or U11341 (N_11341,N_11011,N_11107);
nand U11342 (N_11342,N_11015,N_11215);
nand U11343 (N_11343,N_11178,N_11046);
nor U11344 (N_11344,N_11106,N_11187);
nor U11345 (N_11345,N_11225,N_11003);
or U11346 (N_11346,N_11054,N_11070);
nand U11347 (N_11347,N_11182,N_11132);
nand U11348 (N_11348,N_11071,N_11089);
xor U11349 (N_11349,N_11173,N_11208);
nand U11350 (N_11350,N_11030,N_11243);
xnor U11351 (N_11351,N_11214,N_11145);
nor U11352 (N_11352,N_11159,N_11194);
xnor U11353 (N_11353,N_11052,N_11158);
and U11354 (N_11354,N_11072,N_11164);
xor U11355 (N_11355,N_11113,N_11137);
nand U11356 (N_11356,N_11224,N_11111);
or U11357 (N_11357,N_11147,N_11049);
or U11358 (N_11358,N_11100,N_11193);
and U11359 (N_11359,N_11116,N_11004);
nand U11360 (N_11360,N_11002,N_11031);
or U11361 (N_11361,N_11013,N_11043);
nand U11362 (N_11362,N_11038,N_11006);
or U11363 (N_11363,N_11103,N_11184);
and U11364 (N_11364,N_11001,N_11108);
and U11365 (N_11365,N_11119,N_11227);
and U11366 (N_11366,N_11042,N_11202);
nand U11367 (N_11367,N_11000,N_11192);
and U11368 (N_11368,N_11058,N_11150);
xor U11369 (N_11369,N_11226,N_11060);
and U11370 (N_11370,N_11245,N_11133);
and U11371 (N_11371,N_11185,N_11217);
or U11372 (N_11372,N_11233,N_11121);
nand U11373 (N_11373,N_11140,N_11218);
or U11374 (N_11374,N_11120,N_11099);
nand U11375 (N_11375,N_11182,N_11243);
or U11376 (N_11376,N_11044,N_11160);
xnor U11377 (N_11377,N_11159,N_11013);
nor U11378 (N_11378,N_11232,N_11205);
or U11379 (N_11379,N_11234,N_11243);
and U11380 (N_11380,N_11238,N_11147);
nand U11381 (N_11381,N_11158,N_11165);
nor U11382 (N_11382,N_11194,N_11210);
xor U11383 (N_11383,N_11030,N_11191);
nor U11384 (N_11384,N_11126,N_11106);
and U11385 (N_11385,N_11169,N_11087);
nor U11386 (N_11386,N_11214,N_11170);
nor U11387 (N_11387,N_11113,N_11246);
xnor U11388 (N_11388,N_11049,N_11212);
or U11389 (N_11389,N_11238,N_11129);
nand U11390 (N_11390,N_11043,N_11032);
nand U11391 (N_11391,N_11022,N_11027);
and U11392 (N_11392,N_11002,N_11249);
xnor U11393 (N_11393,N_11225,N_11046);
and U11394 (N_11394,N_11059,N_11055);
nand U11395 (N_11395,N_11199,N_11098);
nor U11396 (N_11396,N_11181,N_11216);
nand U11397 (N_11397,N_11098,N_11140);
nand U11398 (N_11398,N_11081,N_11024);
nand U11399 (N_11399,N_11181,N_11012);
xor U11400 (N_11400,N_11076,N_11088);
and U11401 (N_11401,N_11179,N_11090);
nor U11402 (N_11402,N_11001,N_11086);
nand U11403 (N_11403,N_11164,N_11005);
nor U11404 (N_11404,N_11092,N_11144);
or U11405 (N_11405,N_11062,N_11123);
nand U11406 (N_11406,N_11199,N_11039);
or U11407 (N_11407,N_11070,N_11126);
and U11408 (N_11408,N_11074,N_11173);
and U11409 (N_11409,N_11092,N_11017);
xor U11410 (N_11410,N_11231,N_11149);
xor U11411 (N_11411,N_11069,N_11222);
nand U11412 (N_11412,N_11182,N_11157);
or U11413 (N_11413,N_11105,N_11116);
or U11414 (N_11414,N_11013,N_11038);
and U11415 (N_11415,N_11239,N_11062);
and U11416 (N_11416,N_11014,N_11041);
or U11417 (N_11417,N_11164,N_11006);
or U11418 (N_11418,N_11050,N_11122);
nor U11419 (N_11419,N_11232,N_11024);
nor U11420 (N_11420,N_11151,N_11144);
and U11421 (N_11421,N_11212,N_11025);
and U11422 (N_11422,N_11147,N_11235);
xnor U11423 (N_11423,N_11081,N_11235);
nand U11424 (N_11424,N_11157,N_11101);
xnor U11425 (N_11425,N_11241,N_11025);
or U11426 (N_11426,N_11121,N_11231);
and U11427 (N_11427,N_11054,N_11006);
xnor U11428 (N_11428,N_11038,N_11231);
xnor U11429 (N_11429,N_11233,N_11189);
nand U11430 (N_11430,N_11007,N_11244);
and U11431 (N_11431,N_11093,N_11219);
or U11432 (N_11432,N_11062,N_11089);
xnor U11433 (N_11433,N_11126,N_11215);
and U11434 (N_11434,N_11212,N_11021);
and U11435 (N_11435,N_11155,N_11010);
xor U11436 (N_11436,N_11046,N_11051);
xnor U11437 (N_11437,N_11248,N_11204);
or U11438 (N_11438,N_11176,N_11002);
nand U11439 (N_11439,N_11113,N_11034);
xnor U11440 (N_11440,N_11034,N_11004);
and U11441 (N_11441,N_11065,N_11200);
nand U11442 (N_11442,N_11032,N_11141);
nand U11443 (N_11443,N_11066,N_11054);
and U11444 (N_11444,N_11038,N_11094);
nor U11445 (N_11445,N_11175,N_11180);
nand U11446 (N_11446,N_11178,N_11216);
nand U11447 (N_11447,N_11013,N_11120);
or U11448 (N_11448,N_11080,N_11012);
nor U11449 (N_11449,N_11111,N_11021);
and U11450 (N_11450,N_11165,N_11132);
xnor U11451 (N_11451,N_11188,N_11059);
nor U11452 (N_11452,N_11225,N_11086);
or U11453 (N_11453,N_11096,N_11068);
nor U11454 (N_11454,N_11074,N_11178);
and U11455 (N_11455,N_11028,N_11123);
and U11456 (N_11456,N_11014,N_11095);
nand U11457 (N_11457,N_11065,N_11194);
xor U11458 (N_11458,N_11181,N_11233);
xnor U11459 (N_11459,N_11148,N_11022);
xnor U11460 (N_11460,N_11020,N_11149);
and U11461 (N_11461,N_11054,N_11199);
nor U11462 (N_11462,N_11181,N_11051);
or U11463 (N_11463,N_11142,N_11188);
nor U11464 (N_11464,N_11152,N_11015);
nor U11465 (N_11465,N_11248,N_11005);
and U11466 (N_11466,N_11242,N_11206);
and U11467 (N_11467,N_11204,N_11043);
and U11468 (N_11468,N_11090,N_11186);
xor U11469 (N_11469,N_11103,N_11115);
nor U11470 (N_11470,N_11065,N_11222);
and U11471 (N_11471,N_11065,N_11009);
and U11472 (N_11472,N_11131,N_11092);
nand U11473 (N_11473,N_11123,N_11217);
and U11474 (N_11474,N_11171,N_11234);
or U11475 (N_11475,N_11165,N_11028);
and U11476 (N_11476,N_11148,N_11222);
nor U11477 (N_11477,N_11140,N_11086);
nor U11478 (N_11478,N_11150,N_11156);
xnor U11479 (N_11479,N_11030,N_11212);
nor U11480 (N_11480,N_11129,N_11244);
or U11481 (N_11481,N_11207,N_11163);
nand U11482 (N_11482,N_11084,N_11201);
nor U11483 (N_11483,N_11205,N_11249);
nand U11484 (N_11484,N_11184,N_11051);
xnor U11485 (N_11485,N_11192,N_11126);
xnor U11486 (N_11486,N_11045,N_11044);
xor U11487 (N_11487,N_11238,N_11044);
or U11488 (N_11488,N_11112,N_11178);
and U11489 (N_11489,N_11074,N_11042);
or U11490 (N_11490,N_11160,N_11141);
nand U11491 (N_11491,N_11115,N_11226);
or U11492 (N_11492,N_11240,N_11116);
nand U11493 (N_11493,N_11161,N_11075);
xnor U11494 (N_11494,N_11009,N_11152);
nor U11495 (N_11495,N_11162,N_11042);
nand U11496 (N_11496,N_11036,N_11233);
nand U11497 (N_11497,N_11102,N_11155);
nor U11498 (N_11498,N_11184,N_11046);
nand U11499 (N_11499,N_11050,N_11225);
nand U11500 (N_11500,N_11294,N_11449);
and U11501 (N_11501,N_11495,N_11253);
nand U11502 (N_11502,N_11380,N_11435);
or U11503 (N_11503,N_11350,N_11298);
nor U11504 (N_11504,N_11358,N_11252);
or U11505 (N_11505,N_11328,N_11457);
nor U11506 (N_11506,N_11333,N_11446);
or U11507 (N_11507,N_11254,N_11475);
xnor U11508 (N_11508,N_11264,N_11351);
or U11509 (N_11509,N_11400,N_11444);
or U11510 (N_11510,N_11267,N_11386);
xnor U11511 (N_11511,N_11291,N_11327);
and U11512 (N_11512,N_11472,N_11462);
xor U11513 (N_11513,N_11366,N_11322);
nand U11514 (N_11514,N_11332,N_11293);
nor U11515 (N_11515,N_11408,N_11371);
nor U11516 (N_11516,N_11301,N_11389);
or U11517 (N_11517,N_11492,N_11278);
and U11518 (N_11518,N_11348,N_11474);
or U11519 (N_11519,N_11312,N_11274);
xnor U11520 (N_11520,N_11478,N_11349);
and U11521 (N_11521,N_11467,N_11407);
nor U11522 (N_11522,N_11316,N_11279);
or U11523 (N_11523,N_11439,N_11260);
nand U11524 (N_11524,N_11423,N_11417);
and U11525 (N_11525,N_11497,N_11481);
nor U11526 (N_11526,N_11356,N_11255);
nor U11527 (N_11527,N_11344,N_11436);
nand U11528 (N_11528,N_11412,N_11454);
xor U11529 (N_11529,N_11392,N_11415);
and U11530 (N_11530,N_11266,N_11460);
or U11531 (N_11531,N_11370,N_11448);
nor U11532 (N_11532,N_11490,N_11486);
nand U11533 (N_11533,N_11487,N_11288);
nand U11534 (N_11534,N_11307,N_11355);
xnor U11535 (N_11535,N_11480,N_11450);
and U11536 (N_11536,N_11336,N_11281);
and U11537 (N_11537,N_11270,N_11447);
or U11538 (N_11538,N_11424,N_11445);
nor U11539 (N_11539,N_11429,N_11305);
and U11540 (N_11540,N_11277,N_11455);
nor U11541 (N_11541,N_11364,N_11414);
or U11542 (N_11542,N_11477,N_11426);
and U11543 (N_11543,N_11363,N_11499);
nor U11544 (N_11544,N_11297,N_11342);
nand U11545 (N_11545,N_11384,N_11304);
and U11546 (N_11546,N_11362,N_11319);
nand U11547 (N_11547,N_11416,N_11265);
nor U11548 (N_11548,N_11498,N_11465);
or U11549 (N_11549,N_11313,N_11388);
and U11550 (N_11550,N_11359,N_11276);
nor U11551 (N_11551,N_11343,N_11334);
xor U11552 (N_11552,N_11339,N_11357);
nand U11553 (N_11553,N_11483,N_11300);
or U11554 (N_11554,N_11311,N_11482);
and U11555 (N_11555,N_11451,N_11420);
or U11556 (N_11556,N_11430,N_11250);
or U11557 (N_11557,N_11489,N_11393);
and U11558 (N_11558,N_11368,N_11296);
xnor U11559 (N_11559,N_11317,N_11282);
xor U11560 (N_11560,N_11273,N_11418);
or U11561 (N_11561,N_11361,N_11367);
or U11562 (N_11562,N_11470,N_11346);
nand U11563 (N_11563,N_11256,N_11268);
and U11564 (N_11564,N_11369,N_11459);
or U11565 (N_11565,N_11461,N_11428);
xor U11566 (N_11566,N_11394,N_11320);
nand U11567 (N_11567,N_11354,N_11377);
and U11568 (N_11568,N_11272,N_11330);
nand U11569 (N_11569,N_11390,N_11405);
or U11570 (N_11570,N_11262,N_11374);
nor U11571 (N_11571,N_11401,N_11329);
nor U11572 (N_11572,N_11431,N_11473);
xor U11573 (N_11573,N_11468,N_11458);
nand U11574 (N_11574,N_11299,N_11494);
xnor U11575 (N_11575,N_11463,N_11290);
or U11576 (N_11576,N_11289,N_11421);
nor U11577 (N_11577,N_11440,N_11442);
or U11578 (N_11578,N_11466,N_11432);
nor U11579 (N_11579,N_11464,N_11485);
or U11580 (N_11580,N_11365,N_11353);
xnor U11581 (N_11581,N_11258,N_11391);
nor U11582 (N_11582,N_11402,N_11425);
nor U11583 (N_11583,N_11360,N_11398);
and U11584 (N_11584,N_11437,N_11271);
xnor U11585 (N_11585,N_11285,N_11341);
nor U11586 (N_11586,N_11441,N_11403);
xnor U11587 (N_11587,N_11345,N_11337);
and U11588 (N_11588,N_11324,N_11280);
and U11589 (N_11589,N_11385,N_11269);
nand U11590 (N_11590,N_11406,N_11292);
xnor U11591 (N_11591,N_11382,N_11409);
and U11592 (N_11592,N_11335,N_11443);
nand U11593 (N_11593,N_11383,N_11493);
nor U11594 (N_11594,N_11308,N_11326);
or U11595 (N_11595,N_11438,N_11373);
or U11596 (N_11596,N_11427,N_11309);
or U11597 (N_11597,N_11379,N_11479);
nor U11598 (N_11598,N_11314,N_11331);
nor U11599 (N_11599,N_11395,N_11275);
xor U11600 (N_11600,N_11413,N_11376);
nor U11601 (N_11601,N_11310,N_11315);
or U11602 (N_11602,N_11484,N_11257);
or U11603 (N_11603,N_11488,N_11338);
nor U11604 (N_11604,N_11419,N_11302);
nand U11605 (N_11605,N_11306,N_11404);
and U11606 (N_11606,N_11286,N_11387);
or U11607 (N_11607,N_11287,N_11347);
and U11608 (N_11608,N_11375,N_11452);
nor U11609 (N_11609,N_11456,N_11471);
and U11610 (N_11610,N_11340,N_11476);
and U11611 (N_11611,N_11378,N_11453);
xnor U11612 (N_11612,N_11323,N_11251);
xnor U11613 (N_11613,N_11410,N_11422);
or U11614 (N_11614,N_11433,N_11352);
and U11615 (N_11615,N_11469,N_11325);
nor U11616 (N_11616,N_11284,N_11397);
and U11617 (N_11617,N_11321,N_11396);
xnor U11618 (N_11618,N_11261,N_11263);
or U11619 (N_11619,N_11399,N_11411);
and U11620 (N_11620,N_11372,N_11496);
nand U11621 (N_11621,N_11318,N_11381);
nor U11622 (N_11622,N_11303,N_11283);
or U11623 (N_11623,N_11259,N_11491);
xnor U11624 (N_11624,N_11434,N_11295);
or U11625 (N_11625,N_11443,N_11373);
nand U11626 (N_11626,N_11400,N_11304);
nand U11627 (N_11627,N_11417,N_11315);
and U11628 (N_11628,N_11373,N_11485);
and U11629 (N_11629,N_11263,N_11313);
or U11630 (N_11630,N_11277,N_11379);
nor U11631 (N_11631,N_11258,N_11289);
or U11632 (N_11632,N_11320,N_11408);
and U11633 (N_11633,N_11281,N_11415);
xor U11634 (N_11634,N_11472,N_11382);
nand U11635 (N_11635,N_11362,N_11361);
nand U11636 (N_11636,N_11390,N_11414);
xor U11637 (N_11637,N_11341,N_11310);
nand U11638 (N_11638,N_11443,N_11294);
and U11639 (N_11639,N_11469,N_11455);
nor U11640 (N_11640,N_11346,N_11380);
or U11641 (N_11641,N_11288,N_11277);
and U11642 (N_11642,N_11316,N_11444);
nand U11643 (N_11643,N_11425,N_11440);
nand U11644 (N_11644,N_11381,N_11321);
or U11645 (N_11645,N_11427,N_11315);
or U11646 (N_11646,N_11364,N_11466);
and U11647 (N_11647,N_11329,N_11270);
xor U11648 (N_11648,N_11257,N_11362);
xor U11649 (N_11649,N_11460,N_11258);
nand U11650 (N_11650,N_11341,N_11449);
or U11651 (N_11651,N_11274,N_11323);
and U11652 (N_11652,N_11269,N_11441);
xnor U11653 (N_11653,N_11387,N_11405);
or U11654 (N_11654,N_11310,N_11388);
nand U11655 (N_11655,N_11366,N_11421);
and U11656 (N_11656,N_11471,N_11499);
and U11657 (N_11657,N_11460,N_11288);
or U11658 (N_11658,N_11386,N_11431);
nand U11659 (N_11659,N_11400,N_11435);
nand U11660 (N_11660,N_11283,N_11473);
nand U11661 (N_11661,N_11352,N_11262);
nand U11662 (N_11662,N_11320,N_11481);
nor U11663 (N_11663,N_11272,N_11432);
nor U11664 (N_11664,N_11354,N_11452);
nor U11665 (N_11665,N_11343,N_11421);
nand U11666 (N_11666,N_11309,N_11454);
and U11667 (N_11667,N_11408,N_11321);
nor U11668 (N_11668,N_11385,N_11488);
nor U11669 (N_11669,N_11333,N_11318);
and U11670 (N_11670,N_11270,N_11393);
and U11671 (N_11671,N_11321,N_11460);
nor U11672 (N_11672,N_11342,N_11363);
or U11673 (N_11673,N_11309,N_11490);
or U11674 (N_11674,N_11440,N_11256);
or U11675 (N_11675,N_11324,N_11476);
or U11676 (N_11676,N_11430,N_11429);
and U11677 (N_11677,N_11474,N_11420);
and U11678 (N_11678,N_11453,N_11283);
xnor U11679 (N_11679,N_11405,N_11479);
nor U11680 (N_11680,N_11429,N_11287);
and U11681 (N_11681,N_11310,N_11486);
nand U11682 (N_11682,N_11325,N_11448);
and U11683 (N_11683,N_11316,N_11424);
nor U11684 (N_11684,N_11497,N_11276);
nand U11685 (N_11685,N_11311,N_11275);
and U11686 (N_11686,N_11272,N_11388);
and U11687 (N_11687,N_11424,N_11456);
nor U11688 (N_11688,N_11369,N_11415);
or U11689 (N_11689,N_11294,N_11347);
or U11690 (N_11690,N_11416,N_11380);
or U11691 (N_11691,N_11416,N_11366);
nand U11692 (N_11692,N_11275,N_11279);
nand U11693 (N_11693,N_11277,N_11297);
nor U11694 (N_11694,N_11373,N_11400);
nor U11695 (N_11695,N_11487,N_11492);
and U11696 (N_11696,N_11376,N_11441);
or U11697 (N_11697,N_11284,N_11371);
nand U11698 (N_11698,N_11459,N_11324);
and U11699 (N_11699,N_11425,N_11347);
nor U11700 (N_11700,N_11486,N_11404);
xnor U11701 (N_11701,N_11429,N_11351);
and U11702 (N_11702,N_11425,N_11269);
and U11703 (N_11703,N_11390,N_11458);
xor U11704 (N_11704,N_11398,N_11349);
xor U11705 (N_11705,N_11283,N_11485);
xor U11706 (N_11706,N_11468,N_11318);
and U11707 (N_11707,N_11374,N_11290);
xnor U11708 (N_11708,N_11493,N_11491);
or U11709 (N_11709,N_11451,N_11387);
nand U11710 (N_11710,N_11306,N_11485);
and U11711 (N_11711,N_11497,N_11357);
or U11712 (N_11712,N_11251,N_11253);
nor U11713 (N_11713,N_11344,N_11425);
or U11714 (N_11714,N_11471,N_11288);
or U11715 (N_11715,N_11490,N_11400);
and U11716 (N_11716,N_11357,N_11391);
xnor U11717 (N_11717,N_11338,N_11394);
xor U11718 (N_11718,N_11424,N_11433);
nor U11719 (N_11719,N_11269,N_11413);
nor U11720 (N_11720,N_11360,N_11344);
xor U11721 (N_11721,N_11383,N_11300);
nor U11722 (N_11722,N_11385,N_11402);
xor U11723 (N_11723,N_11291,N_11322);
nand U11724 (N_11724,N_11438,N_11290);
nor U11725 (N_11725,N_11490,N_11396);
xor U11726 (N_11726,N_11447,N_11255);
nand U11727 (N_11727,N_11471,N_11427);
nand U11728 (N_11728,N_11301,N_11491);
xor U11729 (N_11729,N_11473,N_11297);
nand U11730 (N_11730,N_11338,N_11392);
nand U11731 (N_11731,N_11256,N_11291);
and U11732 (N_11732,N_11377,N_11300);
and U11733 (N_11733,N_11446,N_11356);
and U11734 (N_11734,N_11359,N_11356);
xnor U11735 (N_11735,N_11304,N_11380);
xnor U11736 (N_11736,N_11278,N_11390);
nor U11737 (N_11737,N_11356,N_11312);
and U11738 (N_11738,N_11467,N_11359);
nand U11739 (N_11739,N_11261,N_11275);
or U11740 (N_11740,N_11416,N_11250);
nand U11741 (N_11741,N_11318,N_11408);
nor U11742 (N_11742,N_11482,N_11432);
nand U11743 (N_11743,N_11285,N_11495);
nor U11744 (N_11744,N_11279,N_11456);
or U11745 (N_11745,N_11374,N_11334);
nor U11746 (N_11746,N_11261,N_11304);
and U11747 (N_11747,N_11367,N_11363);
nand U11748 (N_11748,N_11286,N_11252);
or U11749 (N_11749,N_11497,N_11485);
nor U11750 (N_11750,N_11640,N_11736);
and U11751 (N_11751,N_11688,N_11698);
or U11752 (N_11752,N_11522,N_11566);
and U11753 (N_11753,N_11587,N_11631);
xor U11754 (N_11754,N_11741,N_11641);
or U11755 (N_11755,N_11711,N_11635);
xor U11756 (N_11756,N_11662,N_11732);
nor U11757 (N_11757,N_11636,N_11626);
nor U11758 (N_11758,N_11530,N_11694);
xnor U11759 (N_11759,N_11632,N_11514);
xor U11760 (N_11760,N_11511,N_11739);
xnor U11761 (N_11761,N_11619,N_11655);
xor U11762 (N_11762,N_11745,N_11706);
nand U11763 (N_11763,N_11531,N_11661);
xnor U11764 (N_11764,N_11502,N_11695);
xor U11765 (N_11765,N_11679,N_11692);
xor U11766 (N_11766,N_11669,N_11513);
nor U11767 (N_11767,N_11535,N_11659);
xnor U11768 (N_11768,N_11547,N_11570);
xnor U11769 (N_11769,N_11515,N_11568);
or U11770 (N_11770,N_11521,N_11671);
or U11771 (N_11771,N_11528,N_11508);
xor U11772 (N_11772,N_11561,N_11576);
nor U11773 (N_11773,N_11684,N_11562);
xor U11774 (N_11774,N_11586,N_11743);
nor U11775 (N_11775,N_11554,N_11581);
nand U11776 (N_11776,N_11746,N_11606);
or U11777 (N_11777,N_11733,N_11708);
xor U11778 (N_11778,N_11505,N_11724);
nor U11779 (N_11779,N_11593,N_11716);
nor U11780 (N_11780,N_11569,N_11689);
and U11781 (N_11781,N_11742,N_11678);
xnor U11782 (N_11782,N_11548,N_11611);
nor U11783 (N_11783,N_11633,N_11721);
or U11784 (N_11784,N_11627,N_11500);
nor U11785 (N_11785,N_11556,N_11507);
nand U11786 (N_11786,N_11539,N_11729);
nand U11787 (N_11787,N_11592,N_11697);
xor U11788 (N_11788,N_11524,N_11674);
and U11789 (N_11789,N_11610,N_11728);
nand U11790 (N_11790,N_11552,N_11579);
and U11791 (N_11791,N_11544,N_11532);
nand U11792 (N_11792,N_11555,N_11625);
and U11793 (N_11793,N_11677,N_11558);
nor U11794 (N_11794,N_11720,N_11649);
and U11795 (N_11795,N_11598,N_11596);
nand U11796 (N_11796,N_11506,N_11526);
xor U11797 (N_11797,N_11654,N_11693);
nor U11798 (N_11798,N_11701,N_11509);
or U11799 (N_11799,N_11747,N_11685);
xor U11800 (N_11800,N_11503,N_11668);
xor U11801 (N_11801,N_11715,N_11714);
and U11802 (N_11802,N_11559,N_11622);
and U11803 (N_11803,N_11608,N_11696);
xnor U11804 (N_11804,N_11510,N_11638);
nand U11805 (N_11805,N_11525,N_11546);
and U11806 (N_11806,N_11718,N_11577);
nand U11807 (N_11807,N_11597,N_11734);
or U11808 (N_11808,N_11660,N_11519);
nor U11809 (N_11809,N_11523,N_11700);
or U11810 (N_11810,N_11717,N_11571);
and U11811 (N_11811,N_11628,N_11712);
xnor U11812 (N_11812,N_11642,N_11595);
or U11813 (N_11813,N_11735,N_11545);
and U11814 (N_11814,N_11675,N_11629);
nor U11815 (N_11815,N_11560,N_11719);
nor U11816 (N_11816,N_11614,N_11713);
xnor U11817 (N_11817,N_11603,N_11550);
or U11818 (N_11818,N_11630,N_11551);
nor U11819 (N_11819,N_11578,N_11590);
nor U11820 (N_11820,N_11637,N_11541);
xnor U11821 (N_11821,N_11722,N_11613);
nand U11822 (N_11822,N_11563,N_11617);
nand U11823 (N_11823,N_11599,N_11725);
nor U11824 (N_11824,N_11749,N_11501);
xnor U11825 (N_11825,N_11537,N_11594);
nand U11826 (N_11826,N_11564,N_11740);
xor U11827 (N_11827,N_11676,N_11691);
and U11828 (N_11828,N_11527,N_11621);
nor U11829 (N_11829,N_11601,N_11602);
and U11830 (N_11830,N_11686,N_11699);
or U11831 (N_11831,N_11682,N_11647);
nor U11832 (N_11832,N_11543,N_11517);
xnor U11833 (N_11833,N_11656,N_11644);
nor U11834 (N_11834,N_11585,N_11520);
nand U11835 (N_11835,N_11573,N_11643);
and U11836 (N_11836,N_11582,N_11604);
or U11837 (N_11837,N_11567,N_11710);
nor U11838 (N_11838,N_11723,N_11575);
or U11839 (N_11839,N_11727,N_11646);
xnor U11840 (N_11840,N_11534,N_11565);
and U11841 (N_11841,N_11516,N_11730);
xor U11842 (N_11842,N_11624,N_11650);
nand U11843 (N_11843,N_11738,N_11683);
nor U11844 (N_11844,N_11652,N_11612);
nor U11845 (N_11845,N_11690,N_11672);
or U11846 (N_11846,N_11648,N_11623);
nor U11847 (N_11847,N_11580,N_11687);
xnor U11848 (N_11848,N_11744,N_11673);
nand U11849 (N_11849,N_11572,N_11707);
and U11850 (N_11850,N_11615,N_11518);
xnor U11851 (N_11851,N_11704,N_11589);
nor U11852 (N_11852,N_11663,N_11726);
nor U11853 (N_11853,N_11666,N_11645);
nand U11854 (N_11854,N_11607,N_11731);
or U11855 (N_11855,N_11538,N_11653);
xor U11856 (N_11856,N_11591,N_11600);
nor U11857 (N_11857,N_11557,N_11609);
xor U11858 (N_11858,N_11605,N_11574);
nand U11859 (N_11859,N_11620,N_11705);
nor U11860 (N_11860,N_11639,N_11504);
nand U11861 (N_11861,N_11512,N_11542);
nor U11862 (N_11862,N_11681,N_11709);
nor U11863 (N_11863,N_11549,N_11703);
and U11864 (N_11864,N_11651,N_11553);
nand U11865 (N_11865,N_11583,N_11737);
nand U11866 (N_11866,N_11667,N_11657);
xnor U11867 (N_11867,N_11584,N_11616);
or U11868 (N_11868,N_11670,N_11540);
and U11869 (N_11869,N_11748,N_11588);
nand U11870 (N_11870,N_11680,N_11634);
xor U11871 (N_11871,N_11665,N_11702);
and U11872 (N_11872,N_11658,N_11533);
or U11873 (N_11873,N_11664,N_11536);
xor U11874 (N_11874,N_11618,N_11529);
xnor U11875 (N_11875,N_11564,N_11608);
xnor U11876 (N_11876,N_11653,N_11596);
xnor U11877 (N_11877,N_11743,N_11642);
xor U11878 (N_11878,N_11700,N_11652);
and U11879 (N_11879,N_11510,N_11564);
xnor U11880 (N_11880,N_11749,N_11724);
nor U11881 (N_11881,N_11699,N_11689);
nor U11882 (N_11882,N_11588,N_11520);
nand U11883 (N_11883,N_11626,N_11501);
nand U11884 (N_11884,N_11532,N_11568);
xor U11885 (N_11885,N_11696,N_11543);
nor U11886 (N_11886,N_11596,N_11548);
and U11887 (N_11887,N_11711,N_11648);
nand U11888 (N_11888,N_11733,N_11589);
and U11889 (N_11889,N_11677,N_11685);
xnor U11890 (N_11890,N_11570,N_11709);
nor U11891 (N_11891,N_11572,N_11616);
nand U11892 (N_11892,N_11677,N_11571);
or U11893 (N_11893,N_11586,N_11506);
nand U11894 (N_11894,N_11609,N_11550);
and U11895 (N_11895,N_11583,N_11668);
and U11896 (N_11896,N_11694,N_11710);
or U11897 (N_11897,N_11642,N_11608);
or U11898 (N_11898,N_11590,N_11640);
xor U11899 (N_11899,N_11705,N_11582);
and U11900 (N_11900,N_11523,N_11512);
nand U11901 (N_11901,N_11552,N_11622);
xor U11902 (N_11902,N_11680,N_11701);
and U11903 (N_11903,N_11658,N_11653);
nand U11904 (N_11904,N_11550,N_11644);
or U11905 (N_11905,N_11727,N_11682);
nor U11906 (N_11906,N_11695,N_11545);
or U11907 (N_11907,N_11569,N_11648);
nand U11908 (N_11908,N_11587,N_11543);
nor U11909 (N_11909,N_11663,N_11504);
or U11910 (N_11910,N_11527,N_11544);
nand U11911 (N_11911,N_11726,N_11701);
or U11912 (N_11912,N_11717,N_11700);
xnor U11913 (N_11913,N_11516,N_11589);
xor U11914 (N_11914,N_11709,N_11697);
nand U11915 (N_11915,N_11568,N_11578);
or U11916 (N_11916,N_11740,N_11519);
nor U11917 (N_11917,N_11647,N_11584);
xnor U11918 (N_11918,N_11533,N_11692);
nor U11919 (N_11919,N_11546,N_11693);
xor U11920 (N_11920,N_11689,N_11545);
and U11921 (N_11921,N_11718,N_11543);
xor U11922 (N_11922,N_11566,N_11592);
nand U11923 (N_11923,N_11635,N_11556);
or U11924 (N_11924,N_11661,N_11611);
and U11925 (N_11925,N_11617,N_11635);
nand U11926 (N_11926,N_11588,N_11547);
xnor U11927 (N_11927,N_11700,N_11531);
xor U11928 (N_11928,N_11619,N_11515);
nor U11929 (N_11929,N_11731,N_11506);
nor U11930 (N_11930,N_11656,N_11725);
xor U11931 (N_11931,N_11667,N_11647);
nand U11932 (N_11932,N_11650,N_11513);
nand U11933 (N_11933,N_11720,N_11583);
xor U11934 (N_11934,N_11743,N_11505);
nand U11935 (N_11935,N_11679,N_11739);
or U11936 (N_11936,N_11669,N_11745);
xnor U11937 (N_11937,N_11747,N_11588);
nand U11938 (N_11938,N_11576,N_11555);
and U11939 (N_11939,N_11591,N_11686);
nand U11940 (N_11940,N_11614,N_11604);
nand U11941 (N_11941,N_11648,N_11566);
or U11942 (N_11942,N_11519,N_11518);
or U11943 (N_11943,N_11598,N_11619);
nand U11944 (N_11944,N_11674,N_11647);
or U11945 (N_11945,N_11518,N_11749);
and U11946 (N_11946,N_11644,N_11620);
and U11947 (N_11947,N_11719,N_11604);
nand U11948 (N_11948,N_11682,N_11532);
nor U11949 (N_11949,N_11551,N_11508);
xnor U11950 (N_11950,N_11723,N_11618);
xor U11951 (N_11951,N_11683,N_11536);
or U11952 (N_11952,N_11738,N_11720);
nor U11953 (N_11953,N_11662,N_11717);
nor U11954 (N_11954,N_11653,N_11670);
nor U11955 (N_11955,N_11689,N_11530);
nand U11956 (N_11956,N_11617,N_11551);
or U11957 (N_11957,N_11713,N_11745);
nor U11958 (N_11958,N_11611,N_11594);
or U11959 (N_11959,N_11746,N_11607);
and U11960 (N_11960,N_11691,N_11711);
or U11961 (N_11961,N_11506,N_11705);
and U11962 (N_11962,N_11717,N_11593);
nand U11963 (N_11963,N_11705,N_11551);
or U11964 (N_11964,N_11536,N_11706);
and U11965 (N_11965,N_11680,N_11686);
xnor U11966 (N_11966,N_11616,N_11652);
or U11967 (N_11967,N_11705,N_11621);
nand U11968 (N_11968,N_11657,N_11545);
nand U11969 (N_11969,N_11676,N_11744);
nand U11970 (N_11970,N_11506,N_11682);
nor U11971 (N_11971,N_11697,N_11530);
and U11972 (N_11972,N_11668,N_11522);
or U11973 (N_11973,N_11735,N_11581);
nand U11974 (N_11974,N_11654,N_11722);
or U11975 (N_11975,N_11569,N_11662);
or U11976 (N_11976,N_11617,N_11604);
nor U11977 (N_11977,N_11522,N_11635);
and U11978 (N_11978,N_11659,N_11500);
and U11979 (N_11979,N_11548,N_11568);
xor U11980 (N_11980,N_11548,N_11575);
nand U11981 (N_11981,N_11601,N_11576);
or U11982 (N_11982,N_11503,N_11650);
and U11983 (N_11983,N_11678,N_11548);
or U11984 (N_11984,N_11606,N_11737);
or U11985 (N_11985,N_11726,N_11691);
xnor U11986 (N_11986,N_11518,N_11740);
nand U11987 (N_11987,N_11748,N_11735);
and U11988 (N_11988,N_11519,N_11527);
or U11989 (N_11989,N_11540,N_11632);
or U11990 (N_11990,N_11519,N_11551);
and U11991 (N_11991,N_11702,N_11740);
xnor U11992 (N_11992,N_11579,N_11569);
nor U11993 (N_11993,N_11635,N_11721);
or U11994 (N_11994,N_11652,N_11735);
or U11995 (N_11995,N_11595,N_11698);
nor U11996 (N_11996,N_11701,N_11544);
nor U11997 (N_11997,N_11747,N_11501);
nor U11998 (N_11998,N_11564,N_11540);
nor U11999 (N_11999,N_11570,N_11699);
xnor U12000 (N_12000,N_11829,N_11819);
or U12001 (N_12001,N_11772,N_11934);
and U12002 (N_12002,N_11959,N_11806);
and U12003 (N_12003,N_11856,N_11902);
and U12004 (N_12004,N_11993,N_11897);
nor U12005 (N_12005,N_11820,N_11945);
nor U12006 (N_12006,N_11999,N_11953);
xor U12007 (N_12007,N_11997,N_11796);
and U12008 (N_12008,N_11888,N_11940);
and U12009 (N_12009,N_11903,N_11781);
and U12010 (N_12010,N_11987,N_11963);
nor U12011 (N_12011,N_11865,N_11957);
xor U12012 (N_12012,N_11962,N_11761);
and U12013 (N_12013,N_11803,N_11815);
or U12014 (N_12014,N_11822,N_11810);
and U12015 (N_12015,N_11935,N_11768);
nor U12016 (N_12016,N_11956,N_11925);
xnor U12017 (N_12017,N_11920,N_11871);
and U12018 (N_12018,N_11978,N_11980);
nor U12019 (N_12019,N_11771,N_11840);
and U12020 (N_12020,N_11793,N_11916);
nor U12021 (N_12021,N_11949,N_11757);
or U12022 (N_12022,N_11944,N_11850);
and U12023 (N_12023,N_11992,N_11870);
xor U12024 (N_12024,N_11782,N_11910);
nor U12025 (N_12025,N_11911,N_11839);
or U12026 (N_12026,N_11842,N_11816);
xor U12027 (N_12027,N_11784,N_11979);
nor U12028 (N_12028,N_11844,N_11891);
nand U12029 (N_12029,N_11947,N_11926);
or U12030 (N_12030,N_11809,N_11893);
nand U12031 (N_12031,N_11973,N_11798);
or U12032 (N_12032,N_11831,N_11795);
xnor U12033 (N_12033,N_11833,N_11814);
and U12034 (N_12034,N_11885,N_11900);
and U12035 (N_12035,N_11960,N_11834);
or U12036 (N_12036,N_11951,N_11948);
and U12037 (N_12037,N_11882,N_11994);
nand U12038 (N_12038,N_11848,N_11984);
and U12039 (N_12039,N_11936,N_11824);
xor U12040 (N_12040,N_11847,N_11790);
xnor U12041 (N_12041,N_11913,N_11879);
nand U12042 (N_12042,N_11912,N_11905);
xnor U12043 (N_12043,N_11867,N_11752);
nand U12044 (N_12044,N_11895,N_11812);
or U12045 (N_12045,N_11939,N_11838);
or U12046 (N_12046,N_11898,N_11989);
and U12047 (N_12047,N_11883,N_11769);
nor U12048 (N_12048,N_11933,N_11862);
or U12049 (N_12049,N_11818,N_11884);
nor U12050 (N_12050,N_11914,N_11841);
xor U12051 (N_12051,N_11909,N_11968);
or U12052 (N_12052,N_11958,N_11899);
nor U12053 (N_12053,N_11828,N_11876);
and U12054 (N_12054,N_11808,N_11779);
nor U12055 (N_12055,N_11765,N_11763);
or U12056 (N_12056,N_11794,N_11890);
nand U12057 (N_12057,N_11878,N_11907);
and U12058 (N_12058,N_11915,N_11858);
nor U12059 (N_12059,N_11930,N_11860);
nor U12060 (N_12060,N_11777,N_11754);
nand U12061 (N_12061,N_11800,N_11990);
xor U12062 (N_12062,N_11826,N_11985);
or U12063 (N_12063,N_11955,N_11801);
nor U12064 (N_12064,N_11863,N_11766);
nor U12065 (N_12065,N_11886,N_11887);
nor U12066 (N_12066,N_11889,N_11918);
nand U12067 (N_12067,N_11943,N_11773);
xnor U12068 (N_12068,N_11789,N_11965);
nand U12069 (N_12069,N_11908,N_11821);
nand U12070 (N_12070,N_11869,N_11767);
nor U12071 (N_12071,N_11775,N_11976);
xnor U12072 (N_12072,N_11921,N_11830);
nor U12073 (N_12073,N_11866,N_11991);
nand U12074 (N_12074,N_11881,N_11966);
and U12075 (N_12075,N_11785,N_11995);
nand U12076 (N_12076,N_11832,N_11974);
or U12077 (N_12077,N_11807,N_11857);
nand U12078 (N_12078,N_11927,N_11788);
and U12079 (N_12079,N_11792,N_11837);
and U12080 (N_12080,N_11791,N_11846);
or U12081 (N_12081,N_11952,N_11859);
or U12082 (N_12082,N_11864,N_11758);
or U12083 (N_12083,N_11932,N_11937);
and U12084 (N_12084,N_11854,N_11946);
and U12085 (N_12085,N_11780,N_11760);
nor U12086 (N_12086,N_11970,N_11770);
and U12087 (N_12087,N_11917,N_11880);
nor U12088 (N_12088,N_11983,N_11762);
nand U12089 (N_12089,N_11804,N_11924);
or U12090 (N_12090,N_11877,N_11988);
nor U12091 (N_12091,N_11892,N_11929);
nand U12092 (N_12092,N_11904,N_11823);
or U12093 (N_12093,N_11753,N_11755);
and U12094 (N_12094,N_11817,N_11906);
nand U12095 (N_12095,N_11996,N_11799);
or U12096 (N_12096,N_11855,N_11835);
nand U12097 (N_12097,N_11853,N_11836);
and U12098 (N_12098,N_11813,N_11825);
and U12099 (N_12099,N_11961,N_11827);
xor U12100 (N_12100,N_11778,N_11802);
or U12101 (N_12101,N_11969,N_11861);
and U12102 (N_12102,N_11851,N_11972);
xor U12103 (N_12103,N_11922,N_11923);
nor U12104 (N_12104,N_11986,N_11931);
nor U12105 (N_12105,N_11852,N_11805);
nand U12106 (N_12106,N_11894,N_11942);
xor U12107 (N_12107,N_11750,N_11783);
nand U12108 (N_12108,N_11971,N_11843);
or U12109 (N_12109,N_11845,N_11975);
xnor U12110 (N_12110,N_11849,N_11982);
nor U12111 (N_12111,N_11797,N_11811);
xor U12112 (N_12112,N_11774,N_11872);
or U12113 (N_12113,N_11787,N_11751);
xor U12114 (N_12114,N_11873,N_11764);
or U12115 (N_12115,N_11950,N_11977);
or U12116 (N_12116,N_11759,N_11868);
or U12117 (N_12117,N_11938,N_11998);
nand U12118 (N_12118,N_11928,N_11776);
xor U12119 (N_12119,N_11964,N_11919);
nand U12120 (N_12120,N_11875,N_11896);
and U12121 (N_12121,N_11901,N_11981);
nand U12122 (N_12122,N_11786,N_11941);
nor U12123 (N_12123,N_11874,N_11756);
and U12124 (N_12124,N_11954,N_11967);
nor U12125 (N_12125,N_11834,N_11911);
nand U12126 (N_12126,N_11819,N_11876);
nor U12127 (N_12127,N_11882,N_11918);
or U12128 (N_12128,N_11991,N_11921);
or U12129 (N_12129,N_11783,N_11755);
or U12130 (N_12130,N_11854,N_11759);
nand U12131 (N_12131,N_11828,N_11965);
nor U12132 (N_12132,N_11946,N_11954);
and U12133 (N_12133,N_11841,N_11797);
nand U12134 (N_12134,N_11980,N_11897);
or U12135 (N_12135,N_11915,N_11816);
or U12136 (N_12136,N_11982,N_11752);
xor U12137 (N_12137,N_11989,N_11867);
nand U12138 (N_12138,N_11996,N_11848);
nor U12139 (N_12139,N_11787,N_11833);
nor U12140 (N_12140,N_11951,N_11878);
and U12141 (N_12141,N_11922,N_11821);
xnor U12142 (N_12142,N_11921,N_11833);
xnor U12143 (N_12143,N_11944,N_11815);
nor U12144 (N_12144,N_11753,N_11902);
and U12145 (N_12145,N_11757,N_11766);
xnor U12146 (N_12146,N_11805,N_11894);
or U12147 (N_12147,N_11873,N_11891);
nor U12148 (N_12148,N_11975,N_11756);
nor U12149 (N_12149,N_11773,N_11909);
or U12150 (N_12150,N_11750,N_11975);
xnor U12151 (N_12151,N_11913,N_11780);
nor U12152 (N_12152,N_11811,N_11899);
or U12153 (N_12153,N_11891,N_11989);
or U12154 (N_12154,N_11769,N_11953);
nand U12155 (N_12155,N_11999,N_11978);
nand U12156 (N_12156,N_11976,N_11904);
nand U12157 (N_12157,N_11873,N_11770);
nor U12158 (N_12158,N_11818,N_11969);
nor U12159 (N_12159,N_11991,N_11886);
or U12160 (N_12160,N_11816,N_11956);
nor U12161 (N_12161,N_11789,N_11782);
nor U12162 (N_12162,N_11805,N_11893);
or U12163 (N_12163,N_11876,N_11903);
and U12164 (N_12164,N_11839,N_11919);
nor U12165 (N_12165,N_11992,N_11942);
nand U12166 (N_12166,N_11814,N_11934);
nand U12167 (N_12167,N_11780,N_11909);
nor U12168 (N_12168,N_11761,N_11912);
or U12169 (N_12169,N_11958,N_11967);
nor U12170 (N_12170,N_11919,N_11760);
and U12171 (N_12171,N_11975,N_11868);
nand U12172 (N_12172,N_11925,N_11959);
xnor U12173 (N_12173,N_11996,N_11885);
and U12174 (N_12174,N_11776,N_11864);
nor U12175 (N_12175,N_11840,N_11891);
xor U12176 (N_12176,N_11984,N_11943);
xnor U12177 (N_12177,N_11889,N_11869);
and U12178 (N_12178,N_11841,N_11784);
and U12179 (N_12179,N_11886,N_11817);
xor U12180 (N_12180,N_11869,N_11989);
nor U12181 (N_12181,N_11973,N_11921);
xnor U12182 (N_12182,N_11755,N_11955);
nand U12183 (N_12183,N_11872,N_11933);
and U12184 (N_12184,N_11798,N_11935);
nand U12185 (N_12185,N_11762,N_11772);
and U12186 (N_12186,N_11848,N_11853);
nand U12187 (N_12187,N_11983,N_11797);
nand U12188 (N_12188,N_11790,N_11902);
or U12189 (N_12189,N_11952,N_11982);
nand U12190 (N_12190,N_11962,N_11785);
xnor U12191 (N_12191,N_11876,N_11825);
nor U12192 (N_12192,N_11894,N_11964);
xor U12193 (N_12193,N_11809,N_11938);
and U12194 (N_12194,N_11961,N_11893);
nor U12195 (N_12195,N_11755,N_11808);
or U12196 (N_12196,N_11783,N_11925);
xnor U12197 (N_12197,N_11934,N_11897);
and U12198 (N_12198,N_11806,N_11909);
nand U12199 (N_12199,N_11994,N_11791);
or U12200 (N_12200,N_11800,N_11840);
or U12201 (N_12201,N_11949,N_11762);
xor U12202 (N_12202,N_11998,N_11971);
and U12203 (N_12203,N_11814,N_11898);
xor U12204 (N_12204,N_11924,N_11766);
and U12205 (N_12205,N_11999,N_11926);
nor U12206 (N_12206,N_11807,N_11975);
xor U12207 (N_12207,N_11967,N_11831);
or U12208 (N_12208,N_11785,N_11964);
and U12209 (N_12209,N_11853,N_11999);
or U12210 (N_12210,N_11868,N_11883);
or U12211 (N_12211,N_11954,N_11950);
and U12212 (N_12212,N_11802,N_11955);
or U12213 (N_12213,N_11933,N_11984);
and U12214 (N_12214,N_11830,N_11932);
or U12215 (N_12215,N_11983,N_11798);
and U12216 (N_12216,N_11798,N_11916);
or U12217 (N_12217,N_11866,N_11788);
and U12218 (N_12218,N_11810,N_11971);
and U12219 (N_12219,N_11817,N_11909);
xnor U12220 (N_12220,N_11763,N_11959);
nor U12221 (N_12221,N_11845,N_11758);
nand U12222 (N_12222,N_11815,N_11752);
nand U12223 (N_12223,N_11778,N_11849);
nor U12224 (N_12224,N_11764,N_11991);
or U12225 (N_12225,N_11916,N_11915);
xnor U12226 (N_12226,N_11792,N_11820);
nand U12227 (N_12227,N_11933,N_11759);
xnor U12228 (N_12228,N_11869,N_11926);
and U12229 (N_12229,N_11760,N_11946);
and U12230 (N_12230,N_11855,N_11916);
and U12231 (N_12231,N_11801,N_11923);
nand U12232 (N_12232,N_11886,N_11762);
or U12233 (N_12233,N_11933,N_11845);
nand U12234 (N_12234,N_11769,N_11817);
nand U12235 (N_12235,N_11809,N_11773);
or U12236 (N_12236,N_11842,N_11921);
or U12237 (N_12237,N_11886,N_11910);
xor U12238 (N_12238,N_11781,N_11954);
xnor U12239 (N_12239,N_11884,N_11994);
or U12240 (N_12240,N_11781,N_11784);
or U12241 (N_12241,N_11867,N_11852);
or U12242 (N_12242,N_11947,N_11804);
or U12243 (N_12243,N_11983,N_11984);
xor U12244 (N_12244,N_11856,N_11952);
and U12245 (N_12245,N_11953,N_11975);
nor U12246 (N_12246,N_11794,N_11858);
and U12247 (N_12247,N_11813,N_11788);
xor U12248 (N_12248,N_11824,N_11881);
nand U12249 (N_12249,N_11773,N_11874);
and U12250 (N_12250,N_12197,N_12121);
xnor U12251 (N_12251,N_12224,N_12072);
or U12252 (N_12252,N_12071,N_12226);
and U12253 (N_12253,N_12150,N_12138);
and U12254 (N_12254,N_12187,N_12149);
nor U12255 (N_12255,N_12122,N_12008);
and U12256 (N_12256,N_12109,N_12044);
nor U12257 (N_12257,N_12087,N_12170);
and U12258 (N_12258,N_12006,N_12098);
and U12259 (N_12259,N_12180,N_12240);
or U12260 (N_12260,N_12235,N_12068);
xnor U12261 (N_12261,N_12141,N_12178);
nor U12262 (N_12262,N_12196,N_12153);
and U12263 (N_12263,N_12175,N_12214);
or U12264 (N_12264,N_12229,N_12011);
nand U12265 (N_12265,N_12022,N_12212);
or U12266 (N_12266,N_12085,N_12078);
and U12267 (N_12267,N_12115,N_12216);
nand U12268 (N_12268,N_12119,N_12094);
xnor U12269 (N_12269,N_12101,N_12038);
or U12270 (N_12270,N_12207,N_12206);
nor U12271 (N_12271,N_12057,N_12051);
nand U12272 (N_12272,N_12107,N_12102);
or U12273 (N_12273,N_12120,N_12043);
and U12274 (N_12274,N_12129,N_12190);
and U12275 (N_12275,N_12118,N_12185);
nand U12276 (N_12276,N_12053,N_12001);
nor U12277 (N_12277,N_12033,N_12025);
xnor U12278 (N_12278,N_12227,N_12135);
and U12279 (N_12279,N_12169,N_12213);
and U12280 (N_12280,N_12160,N_12188);
nand U12281 (N_12281,N_12082,N_12243);
nor U12282 (N_12282,N_12161,N_12158);
nand U12283 (N_12283,N_12090,N_12154);
nand U12284 (N_12284,N_12238,N_12172);
nand U12285 (N_12285,N_12209,N_12124);
xnor U12286 (N_12286,N_12177,N_12027);
xor U12287 (N_12287,N_12063,N_12110);
nor U12288 (N_12288,N_12249,N_12097);
nand U12289 (N_12289,N_12136,N_12152);
nor U12290 (N_12290,N_12123,N_12201);
and U12291 (N_12291,N_12205,N_12099);
and U12292 (N_12292,N_12009,N_12003);
xnor U12293 (N_12293,N_12058,N_12193);
or U12294 (N_12294,N_12244,N_12017);
nor U12295 (N_12295,N_12225,N_12164);
nand U12296 (N_12296,N_12145,N_12080);
or U12297 (N_12297,N_12245,N_12093);
nand U12298 (N_12298,N_12112,N_12042);
and U12299 (N_12299,N_12079,N_12041);
xor U12300 (N_12300,N_12050,N_12039);
nand U12301 (N_12301,N_12073,N_12021);
nand U12302 (N_12302,N_12151,N_12202);
and U12303 (N_12303,N_12204,N_12139);
and U12304 (N_12304,N_12155,N_12059);
nand U12305 (N_12305,N_12174,N_12234);
nor U12306 (N_12306,N_12131,N_12052);
nand U12307 (N_12307,N_12246,N_12007);
and U12308 (N_12308,N_12159,N_12211);
nand U12309 (N_12309,N_12130,N_12166);
nand U12310 (N_12310,N_12069,N_12032);
or U12311 (N_12311,N_12132,N_12077);
nand U12312 (N_12312,N_12182,N_12076);
nand U12313 (N_12313,N_12013,N_12140);
and U12314 (N_12314,N_12000,N_12142);
xor U12315 (N_12315,N_12221,N_12127);
nor U12316 (N_12316,N_12026,N_12031);
nor U12317 (N_12317,N_12030,N_12239);
and U12318 (N_12318,N_12198,N_12200);
and U12319 (N_12319,N_12012,N_12126);
nor U12320 (N_12320,N_12179,N_12067);
nand U12321 (N_12321,N_12125,N_12148);
xor U12322 (N_12322,N_12208,N_12064);
xor U12323 (N_12323,N_12114,N_12228);
xor U12324 (N_12324,N_12014,N_12055);
nand U12325 (N_12325,N_12091,N_12035);
xor U12326 (N_12326,N_12181,N_12070);
xnor U12327 (N_12327,N_12222,N_12242);
or U12328 (N_12328,N_12019,N_12168);
nand U12329 (N_12329,N_12100,N_12117);
and U12330 (N_12330,N_12106,N_12113);
or U12331 (N_12331,N_12195,N_12066);
nand U12332 (N_12332,N_12074,N_12247);
nor U12333 (N_12333,N_12005,N_12194);
and U12334 (N_12334,N_12049,N_12108);
or U12335 (N_12335,N_12144,N_12040);
or U12336 (N_12336,N_12086,N_12056);
and U12337 (N_12337,N_12111,N_12215);
and U12338 (N_12338,N_12105,N_12116);
xor U12339 (N_12339,N_12023,N_12037);
nand U12340 (N_12340,N_12219,N_12223);
xor U12341 (N_12341,N_12015,N_12048);
xnor U12342 (N_12342,N_12203,N_12165);
or U12343 (N_12343,N_12248,N_12232);
nand U12344 (N_12344,N_12104,N_12157);
or U12345 (N_12345,N_12220,N_12137);
or U12346 (N_12346,N_12083,N_12065);
or U12347 (N_12347,N_12103,N_12089);
or U12348 (N_12348,N_12075,N_12147);
xnor U12349 (N_12349,N_12231,N_12241);
or U12350 (N_12350,N_12191,N_12028);
xor U12351 (N_12351,N_12081,N_12210);
and U12352 (N_12352,N_12237,N_12236);
nor U12353 (N_12353,N_12199,N_12146);
and U12354 (N_12354,N_12002,N_12016);
nand U12355 (N_12355,N_12045,N_12060);
xnor U12356 (N_12356,N_12133,N_12128);
and U12357 (N_12357,N_12171,N_12096);
xnor U12358 (N_12358,N_12143,N_12029);
nand U12359 (N_12359,N_12046,N_12134);
nor U12360 (N_12360,N_12062,N_12189);
nand U12361 (N_12361,N_12186,N_12218);
nand U12362 (N_12362,N_12176,N_12047);
nor U12363 (N_12363,N_12054,N_12061);
or U12364 (N_12364,N_12010,N_12163);
xnor U12365 (N_12365,N_12217,N_12084);
or U12366 (N_12366,N_12156,N_12230);
xor U12367 (N_12367,N_12183,N_12034);
or U12368 (N_12368,N_12167,N_12162);
nand U12369 (N_12369,N_12036,N_12095);
and U12370 (N_12370,N_12018,N_12192);
and U12371 (N_12371,N_12024,N_12088);
and U12372 (N_12372,N_12233,N_12004);
xor U12373 (N_12373,N_12184,N_12092);
nor U12374 (N_12374,N_12020,N_12173);
xor U12375 (N_12375,N_12076,N_12194);
nor U12376 (N_12376,N_12166,N_12202);
and U12377 (N_12377,N_12051,N_12193);
xnor U12378 (N_12378,N_12146,N_12027);
nand U12379 (N_12379,N_12031,N_12231);
or U12380 (N_12380,N_12087,N_12196);
nand U12381 (N_12381,N_12200,N_12073);
or U12382 (N_12382,N_12058,N_12039);
or U12383 (N_12383,N_12146,N_12246);
nor U12384 (N_12384,N_12244,N_12139);
or U12385 (N_12385,N_12240,N_12161);
or U12386 (N_12386,N_12157,N_12231);
and U12387 (N_12387,N_12009,N_12091);
nand U12388 (N_12388,N_12248,N_12106);
and U12389 (N_12389,N_12138,N_12189);
xnor U12390 (N_12390,N_12231,N_12189);
or U12391 (N_12391,N_12079,N_12056);
and U12392 (N_12392,N_12068,N_12240);
nor U12393 (N_12393,N_12169,N_12080);
or U12394 (N_12394,N_12194,N_12044);
nand U12395 (N_12395,N_12093,N_12166);
xnor U12396 (N_12396,N_12154,N_12035);
xor U12397 (N_12397,N_12083,N_12137);
xnor U12398 (N_12398,N_12176,N_12223);
xnor U12399 (N_12399,N_12011,N_12121);
nor U12400 (N_12400,N_12014,N_12009);
nand U12401 (N_12401,N_12094,N_12176);
nand U12402 (N_12402,N_12193,N_12021);
nor U12403 (N_12403,N_12028,N_12144);
xor U12404 (N_12404,N_12141,N_12174);
nand U12405 (N_12405,N_12164,N_12238);
nand U12406 (N_12406,N_12181,N_12229);
and U12407 (N_12407,N_12115,N_12003);
nand U12408 (N_12408,N_12105,N_12159);
and U12409 (N_12409,N_12140,N_12016);
or U12410 (N_12410,N_12147,N_12122);
or U12411 (N_12411,N_12124,N_12032);
or U12412 (N_12412,N_12168,N_12055);
xnor U12413 (N_12413,N_12183,N_12142);
xor U12414 (N_12414,N_12161,N_12218);
or U12415 (N_12415,N_12032,N_12165);
or U12416 (N_12416,N_12247,N_12134);
xnor U12417 (N_12417,N_12238,N_12182);
nor U12418 (N_12418,N_12204,N_12056);
nand U12419 (N_12419,N_12031,N_12123);
nor U12420 (N_12420,N_12228,N_12125);
nand U12421 (N_12421,N_12244,N_12041);
and U12422 (N_12422,N_12214,N_12168);
and U12423 (N_12423,N_12078,N_12126);
xnor U12424 (N_12424,N_12048,N_12041);
xnor U12425 (N_12425,N_12148,N_12034);
and U12426 (N_12426,N_12115,N_12220);
nor U12427 (N_12427,N_12157,N_12216);
and U12428 (N_12428,N_12056,N_12116);
nand U12429 (N_12429,N_12151,N_12130);
or U12430 (N_12430,N_12160,N_12018);
nand U12431 (N_12431,N_12231,N_12137);
and U12432 (N_12432,N_12015,N_12237);
and U12433 (N_12433,N_12040,N_12142);
and U12434 (N_12434,N_12046,N_12186);
xor U12435 (N_12435,N_12095,N_12141);
xnor U12436 (N_12436,N_12098,N_12166);
nor U12437 (N_12437,N_12240,N_12182);
or U12438 (N_12438,N_12238,N_12121);
nand U12439 (N_12439,N_12189,N_12181);
or U12440 (N_12440,N_12211,N_12016);
xnor U12441 (N_12441,N_12047,N_12100);
and U12442 (N_12442,N_12038,N_12037);
nor U12443 (N_12443,N_12081,N_12105);
nor U12444 (N_12444,N_12215,N_12034);
nand U12445 (N_12445,N_12018,N_12197);
nor U12446 (N_12446,N_12116,N_12224);
or U12447 (N_12447,N_12241,N_12056);
xnor U12448 (N_12448,N_12225,N_12126);
or U12449 (N_12449,N_12024,N_12240);
or U12450 (N_12450,N_12233,N_12121);
and U12451 (N_12451,N_12055,N_12237);
nor U12452 (N_12452,N_12192,N_12217);
nand U12453 (N_12453,N_12207,N_12112);
nor U12454 (N_12454,N_12206,N_12071);
and U12455 (N_12455,N_12137,N_12049);
nor U12456 (N_12456,N_12130,N_12110);
and U12457 (N_12457,N_12019,N_12124);
or U12458 (N_12458,N_12008,N_12082);
nand U12459 (N_12459,N_12014,N_12245);
nand U12460 (N_12460,N_12051,N_12174);
or U12461 (N_12461,N_12241,N_12018);
nand U12462 (N_12462,N_12132,N_12141);
nand U12463 (N_12463,N_12180,N_12060);
nor U12464 (N_12464,N_12229,N_12108);
nor U12465 (N_12465,N_12236,N_12086);
xor U12466 (N_12466,N_12145,N_12171);
or U12467 (N_12467,N_12128,N_12191);
or U12468 (N_12468,N_12005,N_12131);
xnor U12469 (N_12469,N_12129,N_12220);
nor U12470 (N_12470,N_12222,N_12076);
xor U12471 (N_12471,N_12122,N_12074);
or U12472 (N_12472,N_12070,N_12051);
nand U12473 (N_12473,N_12108,N_12183);
or U12474 (N_12474,N_12035,N_12066);
and U12475 (N_12475,N_12002,N_12200);
or U12476 (N_12476,N_12101,N_12010);
nand U12477 (N_12477,N_12238,N_12073);
nand U12478 (N_12478,N_12221,N_12107);
xnor U12479 (N_12479,N_12043,N_12226);
xor U12480 (N_12480,N_12245,N_12195);
or U12481 (N_12481,N_12176,N_12038);
nand U12482 (N_12482,N_12103,N_12229);
xnor U12483 (N_12483,N_12125,N_12176);
xnor U12484 (N_12484,N_12231,N_12024);
xor U12485 (N_12485,N_12082,N_12025);
and U12486 (N_12486,N_12095,N_12072);
and U12487 (N_12487,N_12183,N_12044);
nand U12488 (N_12488,N_12043,N_12246);
or U12489 (N_12489,N_12076,N_12191);
nor U12490 (N_12490,N_12182,N_12111);
or U12491 (N_12491,N_12053,N_12119);
nand U12492 (N_12492,N_12223,N_12207);
nor U12493 (N_12493,N_12187,N_12010);
and U12494 (N_12494,N_12096,N_12140);
nand U12495 (N_12495,N_12193,N_12075);
xor U12496 (N_12496,N_12025,N_12161);
and U12497 (N_12497,N_12127,N_12059);
xnor U12498 (N_12498,N_12108,N_12238);
xnor U12499 (N_12499,N_12066,N_12215);
and U12500 (N_12500,N_12470,N_12356);
nand U12501 (N_12501,N_12403,N_12329);
xnor U12502 (N_12502,N_12434,N_12266);
nor U12503 (N_12503,N_12400,N_12259);
or U12504 (N_12504,N_12467,N_12254);
or U12505 (N_12505,N_12280,N_12339);
xnor U12506 (N_12506,N_12278,N_12317);
xnor U12507 (N_12507,N_12458,N_12461);
nand U12508 (N_12508,N_12355,N_12474);
nor U12509 (N_12509,N_12493,N_12426);
xor U12510 (N_12510,N_12386,N_12272);
nor U12511 (N_12511,N_12437,N_12391);
and U12512 (N_12512,N_12387,N_12480);
nor U12513 (N_12513,N_12430,N_12463);
xor U12514 (N_12514,N_12489,N_12442);
and U12515 (N_12515,N_12353,N_12452);
and U12516 (N_12516,N_12364,N_12395);
and U12517 (N_12517,N_12378,N_12481);
xor U12518 (N_12518,N_12326,N_12441);
or U12519 (N_12519,N_12252,N_12439);
and U12520 (N_12520,N_12340,N_12308);
nand U12521 (N_12521,N_12371,N_12344);
and U12522 (N_12522,N_12392,N_12389);
and U12523 (N_12523,N_12343,N_12492);
and U12524 (N_12524,N_12438,N_12388);
nand U12525 (N_12525,N_12327,N_12465);
xor U12526 (N_12526,N_12486,N_12269);
nand U12527 (N_12527,N_12490,N_12302);
or U12528 (N_12528,N_12296,N_12449);
nor U12529 (N_12529,N_12484,N_12423);
nand U12530 (N_12530,N_12276,N_12447);
nor U12531 (N_12531,N_12348,N_12306);
or U12532 (N_12532,N_12363,N_12337);
xnor U12533 (N_12533,N_12401,N_12390);
xnor U12534 (N_12534,N_12301,N_12381);
xnor U12535 (N_12535,N_12373,N_12468);
and U12536 (N_12536,N_12498,N_12315);
and U12537 (N_12537,N_12271,N_12451);
and U12538 (N_12538,N_12385,N_12455);
and U12539 (N_12539,N_12435,N_12411);
and U12540 (N_12540,N_12314,N_12405);
or U12541 (N_12541,N_12375,N_12478);
nand U12542 (N_12542,N_12473,N_12257);
nor U12543 (N_12543,N_12349,N_12475);
nand U12544 (N_12544,N_12454,N_12347);
nand U12545 (N_12545,N_12305,N_12270);
and U12546 (N_12546,N_12338,N_12415);
nand U12547 (N_12547,N_12304,N_12361);
xnor U12548 (N_12548,N_12383,N_12459);
and U12549 (N_12549,N_12487,N_12393);
nor U12550 (N_12550,N_12333,N_12497);
or U12551 (N_12551,N_12288,N_12346);
and U12552 (N_12552,N_12477,N_12352);
or U12553 (N_12553,N_12402,N_12299);
or U12554 (N_12554,N_12289,N_12494);
nand U12555 (N_12555,N_12376,N_12444);
and U12556 (N_12556,N_12313,N_12495);
xnor U12557 (N_12557,N_12491,N_12482);
and U12558 (N_12558,N_12483,N_12418);
nor U12559 (N_12559,N_12425,N_12287);
nand U12560 (N_12560,N_12292,N_12342);
xnor U12561 (N_12561,N_12443,N_12382);
nor U12562 (N_12562,N_12283,N_12377);
or U12563 (N_12563,N_12414,N_12307);
nand U12564 (N_12564,N_12290,N_12407);
nand U12565 (N_12565,N_12496,N_12319);
nand U12566 (N_12566,N_12499,N_12294);
or U12567 (N_12567,N_12323,N_12331);
nand U12568 (N_12568,N_12253,N_12408);
nor U12569 (N_12569,N_12255,N_12433);
nor U12570 (N_12570,N_12469,N_12429);
xnor U12571 (N_12571,N_12309,N_12396);
nor U12572 (N_12572,N_12261,N_12281);
nor U12573 (N_12573,N_12398,N_12300);
or U12574 (N_12574,N_12360,N_12421);
xnor U12575 (N_12575,N_12431,N_12419);
nor U12576 (N_12576,N_12357,N_12291);
or U12577 (N_12577,N_12420,N_12324);
and U12578 (N_12578,N_12298,N_12359);
xor U12579 (N_12579,N_12273,N_12256);
nand U12580 (N_12580,N_12303,N_12264);
nand U12581 (N_12581,N_12422,N_12328);
or U12582 (N_12582,N_12410,N_12274);
nor U12583 (N_12583,N_12354,N_12251);
or U12584 (N_12584,N_12413,N_12404);
nor U12585 (N_12585,N_12464,N_12368);
xnor U12586 (N_12586,N_12310,N_12440);
or U12587 (N_12587,N_12267,N_12262);
nor U12588 (N_12588,N_12330,N_12379);
nand U12589 (N_12589,N_12286,N_12406);
and U12590 (N_12590,N_12295,N_12318);
or U12591 (N_12591,N_12427,N_12312);
nor U12592 (N_12592,N_12350,N_12372);
and U12593 (N_12593,N_12268,N_12263);
and U12594 (N_12594,N_12471,N_12394);
or U12595 (N_12595,N_12453,N_12334);
nand U12596 (N_12596,N_12336,N_12428);
xnor U12597 (N_12597,N_12397,N_12358);
and U12598 (N_12598,N_12448,N_12279);
nand U12599 (N_12599,N_12409,N_12335);
xor U12600 (N_12600,N_12366,N_12457);
or U12601 (N_12601,N_12436,N_12380);
and U12602 (N_12602,N_12369,N_12265);
nor U12603 (N_12603,N_12450,N_12362);
or U12604 (N_12604,N_12432,N_12332);
or U12605 (N_12605,N_12285,N_12462);
nor U12606 (N_12606,N_12250,N_12424);
nand U12607 (N_12607,N_12320,N_12311);
nand U12608 (N_12608,N_12399,N_12446);
nand U12609 (N_12609,N_12260,N_12345);
or U12610 (N_12610,N_12485,N_12472);
nand U12611 (N_12611,N_12325,N_12258);
nor U12612 (N_12612,N_12316,N_12284);
nor U12613 (N_12613,N_12417,N_12416);
xnor U12614 (N_12614,N_12322,N_12277);
xnor U12615 (N_12615,N_12321,N_12466);
nor U12616 (N_12616,N_12367,N_12365);
nor U12617 (N_12617,N_12293,N_12460);
and U12618 (N_12618,N_12488,N_12412);
or U12619 (N_12619,N_12445,N_12282);
nand U12620 (N_12620,N_12456,N_12351);
nor U12621 (N_12621,N_12341,N_12479);
and U12622 (N_12622,N_12297,N_12370);
or U12623 (N_12623,N_12476,N_12384);
or U12624 (N_12624,N_12374,N_12275);
xor U12625 (N_12625,N_12394,N_12365);
nor U12626 (N_12626,N_12291,N_12295);
nor U12627 (N_12627,N_12488,N_12328);
xnor U12628 (N_12628,N_12380,N_12258);
xor U12629 (N_12629,N_12326,N_12345);
and U12630 (N_12630,N_12417,N_12309);
and U12631 (N_12631,N_12401,N_12314);
or U12632 (N_12632,N_12378,N_12321);
xor U12633 (N_12633,N_12402,N_12420);
nand U12634 (N_12634,N_12424,N_12354);
and U12635 (N_12635,N_12269,N_12308);
nor U12636 (N_12636,N_12408,N_12364);
nor U12637 (N_12637,N_12322,N_12386);
nor U12638 (N_12638,N_12282,N_12471);
or U12639 (N_12639,N_12270,N_12489);
xnor U12640 (N_12640,N_12410,N_12435);
or U12641 (N_12641,N_12459,N_12333);
and U12642 (N_12642,N_12422,N_12401);
xnor U12643 (N_12643,N_12307,N_12383);
nand U12644 (N_12644,N_12288,N_12321);
xor U12645 (N_12645,N_12319,N_12310);
and U12646 (N_12646,N_12287,N_12410);
nor U12647 (N_12647,N_12346,N_12432);
or U12648 (N_12648,N_12372,N_12453);
nor U12649 (N_12649,N_12309,N_12329);
xnor U12650 (N_12650,N_12465,N_12355);
and U12651 (N_12651,N_12384,N_12348);
or U12652 (N_12652,N_12363,N_12394);
or U12653 (N_12653,N_12347,N_12398);
or U12654 (N_12654,N_12446,N_12349);
nor U12655 (N_12655,N_12374,N_12368);
nor U12656 (N_12656,N_12374,N_12391);
nand U12657 (N_12657,N_12492,N_12270);
xnor U12658 (N_12658,N_12414,N_12402);
nand U12659 (N_12659,N_12330,N_12328);
nand U12660 (N_12660,N_12292,N_12275);
xor U12661 (N_12661,N_12459,N_12435);
or U12662 (N_12662,N_12299,N_12391);
nor U12663 (N_12663,N_12266,N_12351);
xnor U12664 (N_12664,N_12461,N_12415);
and U12665 (N_12665,N_12466,N_12265);
nand U12666 (N_12666,N_12329,N_12460);
nand U12667 (N_12667,N_12486,N_12359);
nand U12668 (N_12668,N_12466,N_12250);
and U12669 (N_12669,N_12284,N_12389);
and U12670 (N_12670,N_12491,N_12464);
nor U12671 (N_12671,N_12470,N_12337);
nand U12672 (N_12672,N_12475,N_12452);
nand U12673 (N_12673,N_12487,N_12294);
and U12674 (N_12674,N_12419,N_12360);
nand U12675 (N_12675,N_12471,N_12312);
nor U12676 (N_12676,N_12437,N_12362);
nand U12677 (N_12677,N_12491,N_12432);
or U12678 (N_12678,N_12385,N_12472);
nand U12679 (N_12679,N_12296,N_12465);
nand U12680 (N_12680,N_12259,N_12358);
and U12681 (N_12681,N_12296,N_12354);
nor U12682 (N_12682,N_12263,N_12397);
nor U12683 (N_12683,N_12391,N_12420);
nor U12684 (N_12684,N_12320,N_12345);
nand U12685 (N_12685,N_12277,N_12372);
or U12686 (N_12686,N_12367,N_12320);
nor U12687 (N_12687,N_12386,N_12292);
and U12688 (N_12688,N_12455,N_12490);
xnor U12689 (N_12689,N_12277,N_12483);
xor U12690 (N_12690,N_12472,N_12409);
or U12691 (N_12691,N_12357,N_12411);
or U12692 (N_12692,N_12340,N_12349);
nand U12693 (N_12693,N_12287,N_12400);
and U12694 (N_12694,N_12325,N_12339);
or U12695 (N_12695,N_12366,N_12454);
and U12696 (N_12696,N_12339,N_12330);
xor U12697 (N_12697,N_12267,N_12295);
and U12698 (N_12698,N_12384,N_12372);
nor U12699 (N_12699,N_12408,N_12464);
and U12700 (N_12700,N_12412,N_12417);
or U12701 (N_12701,N_12387,N_12445);
xor U12702 (N_12702,N_12321,N_12315);
and U12703 (N_12703,N_12413,N_12256);
nand U12704 (N_12704,N_12469,N_12470);
or U12705 (N_12705,N_12498,N_12324);
xor U12706 (N_12706,N_12454,N_12374);
and U12707 (N_12707,N_12339,N_12260);
nand U12708 (N_12708,N_12271,N_12390);
xnor U12709 (N_12709,N_12424,N_12359);
or U12710 (N_12710,N_12262,N_12261);
nand U12711 (N_12711,N_12439,N_12265);
nor U12712 (N_12712,N_12325,N_12318);
or U12713 (N_12713,N_12424,N_12448);
and U12714 (N_12714,N_12482,N_12463);
or U12715 (N_12715,N_12384,N_12256);
nor U12716 (N_12716,N_12250,N_12494);
xnor U12717 (N_12717,N_12440,N_12353);
nand U12718 (N_12718,N_12387,N_12355);
xnor U12719 (N_12719,N_12350,N_12344);
nand U12720 (N_12720,N_12480,N_12341);
and U12721 (N_12721,N_12298,N_12416);
nor U12722 (N_12722,N_12344,N_12340);
and U12723 (N_12723,N_12317,N_12435);
xnor U12724 (N_12724,N_12353,N_12468);
and U12725 (N_12725,N_12463,N_12488);
nor U12726 (N_12726,N_12280,N_12389);
and U12727 (N_12727,N_12485,N_12319);
and U12728 (N_12728,N_12386,N_12336);
nand U12729 (N_12729,N_12252,N_12275);
or U12730 (N_12730,N_12345,N_12378);
nand U12731 (N_12731,N_12469,N_12440);
xor U12732 (N_12732,N_12259,N_12361);
or U12733 (N_12733,N_12432,N_12327);
or U12734 (N_12734,N_12274,N_12279);
nor U12735 (N_12735,N_12355,N_12316);
and U12736 (N_12736,N_12279,N_12414);
xor U12737 (N_12737,N_12332,N_12435);
or U12738 (N_12738,N_12445,N_12490);
or U12739 (N_12739,N_12491,N_12316);
xnor U12740 (N_12740,N_12262,N_12426);
nor U12741 (N_12741,N_12390,N_12306);
nand U12742 (N_12742,N_12358,N_12409);
nand U12743 (N_12743,N_12340,N_12342);
nand U12744 (N_12744,N_12271,N_12256);
nand U12745 (N_12745,N_12419,N_12441);
or U12746 (N_12746,N_12492,N_12341);
and U12747 (N_12747,N_12497,N_12299);
nor U12748 (N_12748,N_12285,N_12379);
nor U12749 (N_12749,N_12266,N_12325);
nand U12750 (N_12750,N_12694,N_12638);
and U12751 (N_12751,N_12551,N_12583);
and U12752 (N_12752,N_12637,N_12507);
or U12753 (N_12753,N_12514,N_12639);
xor U12754 (N_12754,N_12568,N_12600);
nand U12755 (N_12755,N_12605,N_12730);
xor U12756 (N_12756,N_12528,N_12555);
xor U12757 (N_12757,N_12698,N_12721);
or U12758 (N_12758,N_12575,N_12641);
nand U12759 (N_12759,N_12517,N_12561);
or U12760 (N_12760,N_12526,N_12500);
xnor U12761 (N_12761,N_12562,N_12736);
or U12762 (N_12762,N_12683,N_12520);
or U12763 (N_12763,N_12717,N_12589);
or U12764 (N_12764,N_12640,N_12682);
and U12765 (N_12765,N_12739,N_12665);
nand U12766 (N_12766,N_12627,N_12588);
or U12767 (N_12767,N_12710,N_12548);
or U12768 (N_12768,N_12731,N_12614);
and U12769 (N_12769,N_12655,N_12693);
or U12770 (N_12770,N_12625,N_12644);
or U12771 (N_12771,N_12673,N_12632);
nor U12772 (N_12772,N_12530,N_12704);
nor U12773 (N_12773,N_12656,N_12580);
xnor U12774 (N_12774,N_12607,N_12697);
nand U12775 (N_12775,N_12572,N_12689);
and U12776 (N_12776,N_12746,N_12578);
and U12777 (N_12777,N_12635,N_12552);
or U12778 (N_12778,N_12601,N_12684);
xor U12779 (N_12779,N_12504,N_12599);
or U12780 (N_12780,N_12603,N_12587);
xor U12781 (N_12781,N_12700,N_12690);
and U12782 (N_12782,N_12557,N_12711);
xnor U12783 (N_12783,N_12544,N_12716);
or U12784 (N_12784,N_12612,N_12604);
xor U12785 (N_12785,N_12705,N_12509);
xor U12786 (N_12786,N_12707,N_12747);
xnor U12787 (N_12787,N_12525,N_12606);
nand U12788 (N_12788,N_12592,N_12608);
nand U12789 (N_12789,N_12681,N_12680);
and U12790 (N_12790,N_12687,N_12560);
nor U12791 (N_12791,N_12633,N_12718);
nand U12792 (N_12792,N_12506,N_12543);
and U12793 (N_12793,N_12631,N_12537);
and U12794 (N_12794,N_12740,N_12676);
and U12795 (N_12795,N_12685,N_12737);
or U12796 (N_12796,N_12724,N_12674);
and U12797 (N_12797,N_12553,N_12550);
xor U12798 (N_12798,N_12518,N_12649);
nor U12799 (N_12799,N_12563,N_12692);
or U12800 (N_12800,N_12725,N_12558);
xor U12801 (N_12801,N_12715,N_12738);
nor U12802 (N_12802,N_12667,N_12547);
nor U12803 (N_12803,N_12659,N_12722);
xor U12804 (N_12804,N_12577,N_12733);
and U12805 (N_12805,N_12597,N_12559);
nand U12806 (N_12806,N_12732,N_12523);
and U12807 (N_12807,N_12686,N_12611);
xor U12808 (N_12808,N_12616,N_12519);
nor U12809 (N_12809,N_12657,N_12566);
or U12810 (N_12810,N_12708,N_12505);
or U12811 (N_12811,N_12675,N_12648);
nand U12812 (N_12812,N_12510,N_12695);
nand U12813 (N_12813,N_12565,N_12669);
xnor U12814 (N_12814,N_12654,N_12629);
and U12815 (N_12815,N_12582,N_12713);
or U12816 (N_12816,N_12748,N_12642);
nand U12817 (N_12817,N_12653,N_12501);
nor U12818 (N_12818,N_12743,N_12539);
nor U12819 (N_12819,N_12726,N_12742);
nor U12820 (N_12820,N_12609,N_12630);
and U12821 (N_12821,N_12508,N_12613);
and U12822 (N_12822,N_12643,N_12661);
xnor U12823 (N_12823,N_12541,N_12679);
nor U12824 (N_12824,N_12594,N_12668);
or U12825 (N_12825,N_12720,N_12513);
or U12826 (N_12826,N_12650,N_12749);
xor U12827 (N_12827,N_12574,N_12729);
nor U12828 (N_12828,N_12696,N_12586);
xor U12829 (N_12829,N_12556,N_12634);
xnor U12830 (N_12830,N_12735,N_12590);
or U12831 (N_12831,N_12615,N_12670);
nor U12832 (N_12832,N_12533,N_12534);
nor U12833 (N_12833,N_12521,N_12663);
or U12834 (N_12834,N_12502,N_12529);
or U12835 (N_12835,N_12744,N_12598);
nand U12836 (N_12836,N_12712,N_12527);
xnor U12837 (N_12837,N_12546,N_12522);
xor U12838 (N_12838,N_12677,N_12573);
nand U12839 (N_12839,N_12628,N_12734);
and U12840 (N_12840,N_12535,N_12512);
nor U12841 (N_12841,N_12549,N_12503);
xnor U12842 (N_12842,N_12623,N_12678);
xor U12843 (N_12843,N_12564,N_12727);
xor U12844 (N_12844,N_12542,N_12621);
nand U12845 (N_12845,N_12531,N_12741);
xor U12846 (N_12846,N_12540,N_12524);
nand U12847 (N_12847,N_12709,N_12719);
or U12848 (N_12848,N_12622,N_12723);
nor U12849 (N_12849,N_12536,N_12602);
xnor U12850 (N_12850,N_12596,N_12591);
nand U12851 (N_12851,N_12701,N_12664);
and U12852 (N_12852,N_12620,N_12579);
xnor U12853 (N_12853,N_12645,N_12728);
nor U12854 (N_12854,N_12745,N_12666);
nor U12855 (N_12855,N_12545,N_12617);
or U12856 (N_12856,N_12570,N_12511);
and U12857 (N_12857,N_12658,N_12532);
or U12858 (N_12858,N_12515,N_12569);
nor U12859 (N_12859,N_12699,N_12702);
xnor U12860 (N_12860,N_12538,N_12567);
and U12861 (N_12861,N_12652,N_12626);
and U12862 (N_12862,N_12624,N_12593);
xor U12863 (N_12863,N_12581,N_12595);
nor U12864 (N_12864,N_12554,N_12619);
and U12865 (N_12865,N_12576,N_12703);
or U12866 (N_12866,N_12671,N_12516);
xor U12867 (N_12867,N_12660,N_12585);
nor U12868 (N_12868,N_12610,N_12647);
or U12869 (N_12869,N_12584,N_12571);
and U12870 (N_12870,N_12662,N_12688);
nor U12871 (N_12871,N_12651,N_12646);
or U12872 (N_12872,N_12691,N_12636);
or U12873 (N_12873,N_12714,N_12672);
nand U12874 (N_12874,N_12706,N_12618);
nand U12875 (N_12875,N_12696,N_12550);
xor U12876 (N_12876,N_12553,N_12668);
and U12877 (N_12877,N_12524,N_12657);
or U12878 (N_12878,N_12621,N_12676);
xnor U12879 (N_12879,N_12732,N_12660);
xor U12880 (N_12880,N_12540,N_12642);
or U12881 (N_12881,N_12519,N_12649);
or U12882 (N_12882,N_12630,N_12573);
nor U12883 (N_12883,N_12714,N_12645);
nor U12884 (N_12884,N_12514,N_12569);
and U12885 (N_12885,N_12571,N_12680);
nand U12886 (N_12886,N_12613,N_12532);
and U12887 (N_12887,N_12694,N_12716);
nor U12888 (N_12888,N_12592,N_12654);
nand U12889 (N_12889,N_12594,N_12628);
or U12890 (N_12890,N_12577,N_12582);
xnor U12891 (N_12891,N_12643,N_12570);
nand U12892 (N_12892,N_12613,N_12641);
xnor U12893 (N_12893,N_12521,N_12515);
and U12894 (N_12894,N_12653,N_12576);
nand U12895 (N_12895,N_12699,N_12738);
or U12896 (N_12896,N_12743,N_12543);
xnor U12897 (N_12897,N_12595,N_12733);
or U12898 (N_12898,N_12624,N_12576);
nand U12899 (N_12899,N_12585,N_12627);
or U12900 (N_12900,N_12620,N_12530);
nand U12901 (N_12901,N_12723,N_12704);
or U12902 (N_12902,N_12657,N_12526);
and U12903 (N_12903,N_12714,N_12737);
xor U12904 (N_12904,N_12627,N_12660);
and U12905 (N_12905,N_12580,N_12735);
and U12906 (N_12906,N_12700,N_12516);
xor U12907 (N_12907,N_12737,N_12604);
or U12908 (N_12908,N_12534,N_12577);
nor U12909 (N_12909,N_12738,N_12735);
or U12910 (N_12910,N_12591,N_12605);
xor U12911 (N_12911,N_12619,N_12715);
xnor U12912 (N_12912,N_12688,N_12709);
nor U12913 (N_12913,N_12640,N_12637);
or U12914 (N_12914,N_12676,N_12567);
and U12915 (N_12915,N_12696,N_12661);
and U12916 (N_12916,N_12614,N_12635);
xor U12917 (N_12917,N_12553,N_12744);
xnor U12918 (N_12918,N_12739,N_12534);
nor U12919 (N_12919,N_12530,N_12714);
or U12920 (N_12920,N_12511,N_12671);
or U12921 (N_12921,N_12744,N_12603);
nor U12922 (N_12922,N_12663,N_12718);
nand U12923 (N_12923,N_12541,N_12689);
xnor U12924 (N_12924,N_12540,N_12595);
xnor U12925 (N_12925,N_12548,N_12515);
and U12926 (N_12926,N_12508,N_12728);
xor U12927 (N_12927,N_12613,N_12553);
or U12928 (N_12928,N_12525,N_12692);
nand U12929 (N_12929,N_12627,N_12744);
or U12930 (N_12930,N_12523,N_12664);
or U12931 (N_12931,N_12669,N_12590);
or U12932 (N_12932,N_12621,N_12689);
nand U12933 (N_12933,N_12729,N_12630);
or U12934 (N_12934,N_12588,N_12696);
xnor U12935 (N_12935,N_12667,N_12626);
and U12936 (N_12936,N_12533,N_12554);
nor U12937 (N_12937,N_12533,N_12504);
nor U12938 (N_12938,N_12502,N_12538);
nand U12939 (N_12939,N_12654,N_12605);
nand U12940 (N_12940,N_12713,N_12561);
nor U12941 (N_12941,N_12678,N_12685);
nor U12942 (N_12942,N_12652,N_12675);
and U12943 (N_12943,N_12556,N_12543);
xnor U12944 (N_12944,N_12736,N_12522);
nor U12945 (N_12945,N_12704,N_12616);
nand U12946 (N_12946,N_12609,N_12703);
and U12947 (N_12947,N_12704,N_12747);
and U12948 (N_12948,N_12730,N_12685);
nand U12949 (N_12949,N_12696,N_12736);
nand U12950 (N_12950,N_12551,N_12600);
and U12951 (N_12951,N_12659,N_12706);
nand U12952 (N_12952,N_12519,N_12521);
nor U12953 (N_12953,N_12705,N_12563);
nand U12954 (N_12954,N_12730,N_12644);
xnor U12955 (N_12955,N_12699,N_12613);
or U12956 (N_12956,N_12670,N_12563);
xor U12957 (N_12957,N_12543,N_12586);
and U12958 (N_12958,N_12720,N_12527);
or U12959 (N_12959,N_12707,N_12574);
and U12960 (N_12960,N_12606,N_12595);
nand U12961 (N_12961,N_12579,N_12674);
or U12962 (N_12962,N_12579,N_12626);
and U12963 (N_12963,N_12652,N_12539);
nand U12964 (N_12964,N_12722,N_12634);
nor U12965 (N_12965,N_12677,N_12740);
and U12966 (N_12966,N_12670,N_12526);
or U12967 (N_12967,N_12611,N_12582);
nand U12968 (N_12968,N_12551,N_12604);
nand U12969 (N_12969,N_12627,N_12529);
or U12970 (N_12970,N_12565,N_12724);
and U12971 (N_12971,N_12664,N_12736);
or U12972 (N_12972,N_12625,N_12693);
nand U12973 (N_12973,N_12540,N_12526);
or U12974 (N_12974,N_12518,N_12654);
or U12975 (N_12975,N_12640,N_12716);
and U12976 (N_12976,N_12561,N_12533);
nor U12977 (N_12977,N_12517,N_12534);
xnor U12978 (N_12978,N_12654,N_12628);
nor U12979 (N_12979,N_12523,N_12722);
nand U12980 (N_12980,N_12628,N_12721);
nor U12981 (N_12981,N_12585,N_12564);
or U12982 (N_12982,N_12737,N_12744);
or U12983 (N_12983,N_12659,N_12600);
nor U12984 (N_12984,N_12569,N_12617);
xnor U12985 (N_12985,N_12677,N_12643);
or U12986 (N_12986,N_12571,N_12518);
xnor U12987 (N_12987,N_12560,N_12505);
nor U12988 (N_12988,N_12636,N_12578);
xor U12989 (N_12989,N_12733,N_12534);
nor U12990 (N_12990,N_12529,N_12679);
nor U12991 (N_12991,N_12706,N_12504);
xor U12992 (N_12992,N_12648,N_12510);
and U12993 (N_12993,N_12551,N_12743);
nand U12994 (N_12994,N_12577,N_12670);
nand U12995 (N_12995,N_12521,N_12512);
xor U12996 (N_12996,N_12543,N_12618);
xnor U12997 (N_12997,N_12558,N_12712);
or U12998 (N_12998,N_12500,N_12611);
or U12999 (N_12999,N_12685,N_12502);
nor U13000 (N_13000,N_12861,N_12977);
nand U13001 (N_13001,N_12800,N_12950);
or U13002 (N_13002,N_12821,N_12920);
nor U13003 (N_13003,N_12995,N_12960);
or U13004 (N_13004,N_12796,N_12825);
xor U13005 (N_13005,N_12917,N_12873);
and U13006 (N_13006,N_12828,N_12914);
or U13007 (N_13007,N_12848,N_12923);
and U13008 (N_13008,N_12753,N_12774);
and U13009 (N_13009,N_12801,N_12813);
or U13010 (N_13010,N_12795,N_12954);
xnor U13011 (N_13011,N_12969,N_12755);
or U13012 (N_13012,N_12927,N_12953);
xor U13013 (N_13013,N_12872,N_12929);
or U13014 (N_13014,N_12834,N_12829);
xor U13015 (N_13015,N_12901,N_12967);
and U13016 (N_13016,N_12990,N_12905);
or U13017 (N_13017,N_12868,N_12996);
and U13018 (N_13018,N_12896,N_12810);
nand U13019 (N_13019,N_12997,N_12938);
and U13020 (N_13020,N_12856,N_12999);
or U13021 (N_13021,N_12935,N_12855);
xor U13022 (N_13022,N_12945,N_12946);
or U13023 (N_13023,N_12915,N_12936);
or U13024 (N_13024,N_12754,N_12817);
nand U13025 (N_13025,N_12980,N_12998);
or U13026 (N_13026,N_12773,N_12879);
and U13027 (N_13027,N_12762,N_12830);
or U13028 (N_13028,N_12832,N_12906);
and U13029 (N_13029,N_12952,N_12798);
or U13030 (N_13030,N_12932,N_12888);
or U13031 (N_13031,N_12892,N_12765);
nand U13032 (N_13032,N_12948,N_12860);
nand U13033 (N_13033,N_12957,N_12891);
or U13034 (N_13034,N_12840,N_12910);
xnor U13035 (N_13035,N_12956,N_12781);
nor U13036 (N_13036,N_12939,N_12852);
xor U13037 (N_13037,N_12993,N_12972);
nor U13038 (N_13038,N_12907,N_12772);
nor U13039 (N_13039,N_12770,N_12783);
nor U13040 (N_13040,N_12898,N_12925);
or U13041 (N_13041,N_12794,N_12839);
and U13042 (N_13042,N_12989,N_12858);
nand U13043 (N_13043,N_12761,N_12809);
xor U13044 (N_13044,N_12822,N_12846);
and U13045 (N_13045,N_12869,N_12862);
or U13046 (N_13046,N_12885,N_12787);
nand U13047 (N_13047,N_12756,N_12978);
nor U13048 (N_13048,N_12790,N_12806);
xor U13049 (N_13049,N_12912,N_12877);
or U13050 (N_13050,N_12926,N_12937);
or U13051 (N_13051,N_12897,N_12820);
nor U13052 (N_13052,N_12786,N_12833);
nand U13053 (N_13053,N_12766,N_12962);
nand U13054 (N_13054,N_12951,N_12853);
xor U13055 (N_13055,N_12793,N_12902);
or U13056 (N_13056,N_12802,N_12850);
nor U13057 (N_13057,N_12865,N_12991);
nand U13058 (N_13058,N_12924,N_12921);
xor U13059 (N_13059,N_12780,N_12771);
or U13060 (N_13060,N_12894,N_12941);
nor U13061 (N_13061,N_12768,N_12875);
or U13062 (N_13062,N_12911,N_12985);
or U13063 (N_13063,N_12874,N_12867);
nor U13064 (N_13064,N_12982,N_12788);
or U13065 (N_13065,N_12988,N_12965);
and U13066 (N_13066,N_12889,N_12931);
nand U13067 (N_13067,N_12994,N_12973);
and U13068 (N_13068,N_12750,N_12971);
xor U13069 (N_13069,N_12797,N_12958);
and U13070 (N_13070,N_12949,N_12792);
or U13071 (N_13071,N_12984,N_12823);
xnor U13072 (N_13072,N_12849,N_12784);
nand U13073 (N_13073,N_12827,N_12818);
xnor U13074 (N_13074,N_12777,N_12887);
nand U13075 (N_13075,N_12871,N_12838);
nand U13076 (N_13076,N_12987,N_12979);
or U13077 (N_13077,N_12763,N_12816);
xor U13078 (N_13078,N_12808,N_12961);
nor U13079 (N_13079,N_12942,N_12864);
nand U13080 (N_13080,N_12963,N_12851);
nor U13081 (N_13081,N_12970,N_12815);
nor U13082 (N_13082,N_12769,N_12758);
nor U13083 (N_13083,N_12841,N_12854);
nand U13084 (N_13084,N_12890,N_12908);
nand U13085 (N_13085,N_12992,N_12779);
xor U13086 (N_13086,N_12981,N_12955);
xor U13087 (N_13087,N_12842,N_12976);
or U13088 (N_13088,N_12799,N_12884);
nor U13089 (N_13089,N_12947,N_12843);
nand U13090 (N_13090,N_12857,N_12778);
or U13091 (N_13091,N_12803,N_12876);
nor U13092 (N_13092,N_12928,N_12882);
or U13093 (N_13093,N_12986,N_12776);
xnor U13094 (N_13094,N_12764,N_12807);
and U13095 (N_13095,N_12811,N_12805);
and U13096 (N_13096,N_12863,N_12943);
or U13097 (N_13097,N_12964,N_12944);
and U13098 (N_13098,N_12909,N_12752);
and U13099 (N_13099,N_12878,N_12886);
xor U13100 (N_13100,N_12785,N_12918);
nand U13101 (N_13101,N_12968,N_12893);
xnor U13102 (N_13102,N_12959,N_12767);
and U13103 (N_13103,N_12916,N_12966);
and U13104 (N_13104,N_12844,N_12775);
nand U13105 (N_13105,N_12975,N_12934);
nor U13106 (N_13106,N_12940,N_12826);
and U13107 (N_13107,N_12757,N_12847);
nand U13108 (N_13108,N_12751,N_12759);
and U13109 (N_13109,N_12974,N_12819);
and U13110 (N_13110,N_12804,N_12899);
nand U13111 (N_13111,N_12866,N_12895);
and U13112 (N_13112,N_12760,N_12837);
nand U13113 (N_13113,N_12883,N_12933);
nand U13114 (N_13114,N_12983,N_12904);
nor U13115 (N_13115,N_12831,N_12913);
nand U13116 (N_13116,N_12859,N_12791);
nor U13117 (N_13117,N_12814,N_12824);
and U13118 (N_13118,N_12845,N_12836);
xnor U13119 (N_13119,N_12922,N_12919);
nor U13120 (N_13120,N_12870,N_12930);
xnor U13121 (N_13121,N_12881,N_12782);
nand U13122 (N_13122,N_12835,N_12880);
nor U13123 (N_13123,N_12900,N_12789);
nor U13124 (N_13124,N_12903,N_12812);
xnor U13125 (N_13125,N_12971,N_12884);
and U13126 (N_13126,N_12861,N_12797);
and U13127 (N_13127,N_12990,N_12957);
and U13128 (N_13128,N_12816,N_12754);
nand U13129 (N_13129,N_12840,N_12837);
or U13130 (N_13130,N_12893,N_12766);
xor U13131 (N_13131,N_12862,N_12839);
or U13132 (N_13132,N_12753,N_12914);
xor U13133 (N_13133,N_12941,N_12779);
nand U13134 (N_13134,N_12819,N_12827);
and U13135 (N_13135,N_12800,N_12921);
and U13136 (N_13136,N_12940,N_12851);
nor U13137 (N_13137,N_12985,N_12854);
and U13138 (N_13138,N_12957,N_12857);
xor U13139 (N_13139,N_12941,N_12892);
nand U13140 (N_13140,N_12880,N_12962);
and U13141 (N_13141,N_12918,N_12831);
nor U13142 (N_13142,N_12768,N_12880);
or U13143 (N_13143,N_12996,N_12903);
nor U13144 (N_13144,N_12772,N_12921);
or U13145 (N_13145,N_12836,N_12877);
or U13146 (N_13146,N_12792,N_12846);
or U13147 (N_13147,N_12974,N_12867);
nor U13148 (N_13148,N_12841,N_12787);
and U13149 (N_13149,N_12924,N_12937);
or U13150 (N_13150,N_12890,N_12783);
or U13151 (N_13151,N_12938,N_12759);
nor U13152 (N_13152,N_12992,N_12960);
xor U13153 (N_13153,N_12859,N_12752);
and U13154 (N_13154,N_12910,N_12900);
xnor U13155 (N_13155,N_12922,N_12829);
nor U13156 (N_13156,N_12854,N_12865);
nor U13157 (N_13157,N_12950,N_12806);
and U13158 (N_13158,N_12861,N_12857);
and U13159 (N_13159,N_12754,N_12792);
nor U13160 (N_13160,N_12922,N_12979);
nand U13161 (N_13161,N_12804,N_12836);
and U13162 (N_13162,N_12982,N_12861);
and U13163 (N_13163,N_12933,N_12980);
xor U13164 (N_13164,N_12963,N_12959);
xor U13165 (N_13165,N_12916,N_12908);
nand U13166 (N_13166,N_12803,N_12879);
or U13167 (N_13167,N_12956,N_12837);
nand U13168 (N_13168,N_12939,N_12922);
xnor U13169 (N_13169,N_12965,N_12898);
xnor U13170 (N_13170,N_12856,N_12967);
nor U13171 (N_13171,N_12789,N_12880);
nand U13172 (N_13172,N_12800,N_12979);
xor U13173 (N_13173,N_12852,N_12780);
nor U13174 (N_13174,N_12877,N_12800);
or U13175 (N_13175,N_12974,N_12832);
nor U13176 (N_13176,N_12784,N_12946);
xor U13177 (N_13177,N_12971,N_12866);
nand U13178 (N_13178,N_12987,N_12950);
and U13179 (N_13179,N_12948,N_12866);
xor U13180 (N_13180,N_12771,N_12941);
xnor U13181 (N_13181,N_12982,N_12814);
xor U13182 (N_13182,N_12977,N_12894);
nand U13183 (N_13183,N_12818,N_12985);
or U13184 (N_13184,N_12999,N_12783);
xor U13185 (N_13185,N_12846,N_12776);
xnor U13186 (N_13186,N_12933,N_12920);
nand U13187 (N_13187,N_12791,N_12750);
or U13188 (N_13188,N_12881,N_12808);
nand U13189 (N_13189,N_12923,N_12872);
and U13190 (N_13190,N_12971,N_12967);
nand U13191 (N_13191,N_12791,N_12850);
or U13192 (N_13192,N_12838,N_12842);
and U13193 (N_13193,N_12920,N_12796);
xor U13194 (N_13194,N_12915,N_12916);
or U13195 (N_13195,N_12778,N_12913);
or U13196 (N_13196,N_12863,N_12811);
nand U13197 (N_13197,N_12816,N_12819);
or U13198 (N_13198,N_12980,N_12976);
nor U13199 (N_13199,N_12763,N_12753);
and U13200 (N_13200,N_12860,N_12751);
xor U13201 (N_13201,N_12859,N_12972);
nor U13202 (N_13202,N_12971,N_12832);
xnor U13203 (N_13203,N_12990,N_12863);
or U13204 (N_13204,N_12903,N_12859);
and U13205 (N_13205,N_12892,N_12948);
or U13206 (N_13206,N_12896,N_12794);
nand U13207 (N_13207,N_12823,N_12955);
nand U13208 (N_13208,N_12778,N_12898);
or U13209 (N_13209,N_12951,N_12986);
and U13210 (N_13210,N_12968,N_12972);
nor U13211 (N_13211,N_12777,N_12927);
xnor U13212 (N_13212,N_12777,N_12978);
or U13213 (N_13213,N_12760,N_12770);
or U13214 (N_13214,N_12964,N_12982);
nor U13215 (N_13215,N_12919,N_12949);
and U13216 (N_13216,N_12809,N_12864);
nand U13217 (N_13217,N_12873,N_12786);
and U13218 (N_13218,N_12856,N_12986);
xor U13219 (N_13219,N_12906,N_12843);
or U13220 (N_13220,N_12807,N_12930);
and U13221 (N_13221,N_12952,N_12904);
nor U13222 (N_13222,N_12932,N_12919);
xnor U13223 (N_13223,N_12965,N_12918);
or U13224 (N_13224,N_12943,N_12906);
nand U13225 (N_13225,N_12961,N_12952);
and U13226 (N_13226,N_12818,N_12822);
xor U13227 (N_13227,N_12980,N_12769);
xnor U13228 (N_13228,N_12968,N_12824);
or U13229 (N_13229,N_12948,N_12979);
xor U13230 (N_13230,N_12920,N_12761);
or U13231 (N_13231,N_12918,N_12875);
or U13232 (N_13232,N_12821,N_12991);
and U13233 (N_13233,N_12813,N_12948);
nor U13234 (N_13234,N_12924,N_12802);
nand U13235 (N_13235,N_12755,N_12784);
xnor U13236 (N_13236,N_12877,N_12934);
or U13237 (N_13237,N_12806,N_12980);
or U13238 (N_13238,N_12890,N_12856);
and U13239 (N_13239,N_12846,N_12910);
xor U13240 (N_13240,N_12976,N_12870);
xor U13241 (N_13241,N_12976,N_12844);
or U13242 (N_13242,N_12989,N_12996);
xor U13243 (N_13243,N_12893,N_12863);
nor U13244 (N_13244,N_12900,N_12851);
or U13245 (N_13245,N_12783,N_12896);
or U13246 (N_13246,N_12903,N_12800);
nand U13247 (N_13247,N_12863,N_12796);
nor U13248 (N_13248,N_12944,N_12994);
nor U13249 (N_13249,N_12764,N_12956);
xnor U13250 (N_13250,N_13149,N_13184);
nand U13251 (N_13251,N_13081,N_13224);
and U13252 (N_13252,N_13174,N_13194);
nand U13253 (N_13253,N_13239,N_13100);
xor U13254 (N_13254,N_13124,N_13021);
nor U13255 (N_13255,N_13136,N_13034);
or U13256 (N_13256,N_13162,N_13178);
xnor U13257 (N_13257,N_13023,N_13175);
nand U13258 (N_13258,N_13070,N_13120);
xor U13259 (N_13259,N_13092,N_13153);
xor U13260 (N_13260,N_13051,N_13222);
xor U13261 (N_13261,N_13139,N_13106);
or U13262 (N_13262,N_13059,N_13074);
or U13263 (N_13263,N_13009,N_13128);
nor U13264 (N_13264,N_13165,N_13007);
xnor U13265 (N_13265,N_13216,N_13179);
and U13266 (N_13266,N_13082,N_13014);
nor U13267 (N_13267,N_13122,N_13160);
nor U13268 (N_13268,N_13039,N_13111);
nand U13269 (N_13269,N_13025,N_13248);
nand U13270 (N_13270,N_13126,N_13215);
xnor U13271 (N_13271,N_13036,N_13033);
nor U13272 (N_13272,N_13119,N_13209);
or U13273 (N_13273,N_13037,N_13094);
and U13274 (N_13274,N_13105,N_13097);
xor U13275 (N_13275,N_13156,N_13202);
xnor U13276 (N_13276,N_13107,N_13029);
and U13277 (N_13277,N_13217,N_13137);
or U13278 (N_13278,N_13205,N_13158);
xor U13279 (N_13279,N_13032,N_13008);
and U13280 (N_13280,N_13109,N_13071);
xor U13281 (N_13281,N_13161,N_13212);
xnor U13282 (N_13282,N_13242,N_13044);
or U13283 (N_13283,N_13190,N_13129);
and U13284 (N_13284,N_13235,N_13241);
xor U13285 (N_13285,N_13141,N_13134);
nand U13286 (N_13286,N_13026,N_13056);
nand U13287 (N_13287,N_13176,N_13062);
nor U13288 (N_13288,N_13063,N_13113);
xor U13289 (N_13289,N_13168,N_13200);
or U13290 (N_13290,N_13110,N_13146);
xnor U13291 (N_13291,N_13166,N_13022);
or U13292 (N_13292,N_13041,N_13127);
xnor U13293 (N_13293,N_13079,N_13091);
or U13294 (N_13294,N_13047,N_13028);
and U13295 (N_13295,N_13229,N_13171);
and U13296 (N_13296,N_13104,N_13201);
or U13297 (N_13297,N_13228,N_13077);
and U13298 (N_13298,N_13154,N_13024);
nor U13299 (N_13299,N_13230,N_13005);
and U13300 (N_13300,N_13157,N_13232);
nor U13301 (N_13301,N_13078,N_13196);
nand U13302 (N_13302,N_13043,N_13214);
nand U13303 (N_13303,N_13225,N_13131);
nor U13304 (N_13304,N_13012,N_13083);
nand U13305 (N_13305,N_13031,N_13116);
nand U13306 (N_13306,N_13052,N_13017);
nand U13307 (N_13307,N_13140,N_13173);
and U13308 (N_13308,N_13006,N_13181);
or U13309 (N_13309,N_13151,N_13125);
and U13310 (N_13310,N_13203,N_13084);
xor U13311 (N_13311,N_13223,N_13233);
or U13312 (N_13312,N_13088,N_13069);
or U13313 (N_13313,N_13053,N_13093);
or U13314 (N_13314,N_13170,N_13226);
nand U13315 (N_13315,N_13045,N_13066);
nand U13316 (N_13316,N_13090,N_13213);
nand U13317 (N_13317,N_13159,N_13011);
xor U13318 (N_13318,N_13003,N_13210);
and U13319 (N_13319,N_13085,N_13048);
nand U13320 (N_13320,N_13187,N_13193);
nand U13321 (N_13321,N_13087,N_13246);
xor U13322 (N_13322,N_13015,N_13204);
or U13323 (N_13323,N_13143,N_13095);
nor U13324 (N_13324,N_13046,N_13080);
or U13325 (N_13325,N_13133,N_13211);
nor U13326 (N_13326,N_13183,N_13010);
or U13327 (N_13327,N_13065,N_13114);
xnor U13328 (N_13328,N_13054,N_13221);
nor U13329 (N_13329,N_13227,N_13050);
nand U13330 (N_13330,N_13000,N_13020);
nand U13331 (N_13331,N_13167,N_13138);
and U13332 (N_13332,N_13002,N_13188);
xnor U13333 (N_13333,N_13199,N_13099);
nor U13334 (N_13334,N_13150,N_13042);
or U13335 (N_13335,N_13013,N_13058);
and U13336 (N_13336,N_13185,N_13240);
nor U13337 (N_13337,N_13191,N_13061);
nand U13338 (N_13338,N_13049,N_13089);
or U13339 (N_13339,N_13019,N_13067);
xor U13340 (N_13340,N_13231,N_13247);
and U13341 (N_13341,N_13234,N_13206);
nor U13342 (N_13342,N_13197,N_13064);
and U13343 (N_13343,N_13198,N_13102);
and U13344 (N_13344,N_13072,N_13177);
nand U13345 (N_13345,N_13238,N_13182);
nand U13346 (N_13346,N_13144,N_13180);
and U13347 (N_13347,N_13004,N_13245);
or U13348 (N_13348,N_13218,N_13244);
xor U13349 (N_13349,N_13121,N_13132);
nor U13350 (N_13350,N_13172,N_13016);
nand U13351 (N_13351,N_13055,N_13207);
xor U13352 (N_13352,N_13117,N_13057);
and U13353 (N_13353,N_13068,N_13220);
nor U13354 (N_13354,N_13147,N_13195);
nand U13355 (N_13355,N_13018,N_13236);
and U13356 (N_13356,N_13115,N_13145);
nand U13357 (N_13357,N_13076,N_13249);
nor U13358 (N_13358,N_13038,N_13130);
or U13359 (N_13359,N_13243,N_13030);
xnor U13360 (N_13360,N_13075,N_13192);
or U13361 (N_13361,N_13101,N_13096);
xor U13362 (N_13362,N_13103,N_13123);
and U13363 (N_13363,N_13148,N_13164);
or U13364 (N_13364,N_13237,N_13001);
or U13365 (N_13365,N_13040,N_13155);
and U13366 (N_13366,N_13112,N_13152);
and U13367 (N_13367,N_13098,N_13118);
xnor U13368 (N_13368,N_13086,N_13142);
nor U13369 (N_13369,N_13027,N_13208);
nand U13370 (N_13370,N_13219,N_13169);
nor U13371 (N_13371,N_13189,N_13135);
and U13372 (N_13372,N_13163,N_13060);
or U13373 (N_13373,N_13035,N_13108);
xor U13374 (N_13374,N_13073,N_13186);
xnor U13375 (N_13375,N_13075,N_13058);
xor U13376 (N_13376,N_13098,N_13201);
xnor U13377 (N_13377,N_13136,N_13072);
and U13378 (N_13378,N_13042,N_13218);
nand U13379 (N_13379,N_13119,N_13110);
xor U13380 (N_13380,N_13215,N_13191);
or U13381 (N_13381,N_13144,N_13095);
or U13382 (N_13382,N_13107,N_13044);
nor U13383 (N_13383,N_13188,N_13214);
nand U13384 (N_13384,N_13138,N_13085);
and U13385 (N_13385,N_13087,N_13232);
nor U13386 (N_13386,N_13077,N_13172);
xnor U13387 (N_13387,N_13193,N_13071);
nand U13388 (N_13388,N_13245,N_13002);
xnor U13389 (N_13389,N_13139,N_13186);
and U13390 (N_13390,N_13172,N_13165);
or U13391 (N_13391,N_13050,N_13040);
and U13392 (N_13392,N_13189,N_13210);
xnor U13393 (N_13393,N_13158,N_13193);
xor U13394 (N_13394,N_13122,N_13133);
nand U13395 (N_13395,N_13011,N_13208);
xor U13396 (N_13396,N_13221,N_13072);
and U13397 (N_13397,N_13078,N_13173);
xor U13398 (N_13398,N_13192,N_13200);
xor U13399 (N_13399,N_13225,N_13007);
xnor U13400 (N_13400,N_13073,N_13149);
or U13401 (N_13401,N_13135,N_13200);
and U13402 (N_13402,N_13052,N_13149);
nand U13403 (N_13403,N_13131,N_13191);
and U13404 (N_13404,N_13229,N_13015);
xnor U13405 (N_13405,N_13046,N_13035);
and U13406 (N_13406,N_13012,N_13106);
or U13407 (N_13407,N_13097,N_13030);
nand U13408 (N_13408,N_13136,N_13198);
and U13409 (N_13409,N_13045,N_13180);
nor U13410 (N_13410,N_13200,N_13117);
or U13411 (N_13411,N_13102,N_13071);
nand U13412 (N_13412,N_13116,N_13062);
nor U13413 (N_13413,N_13161,N_13200);
or U13414 (N_13414,N_13188,N_13128);
nor U13415 (N_13415,N_13192,N_13063);
and U13416 (N_13416,N_13004,N_13081);
xnor U13417 (N_13417,N_13210,N_13196);
xnor U13418 (N_13418,N_13227,N_13232);
nor U13419 (N_13419,N_13229,N_13110);
nor U13420 (N_13420,N_13135,N_13142);
nand U13421 (N_13421,N_13110,N_13061);
and U13422 (N_13422,N_13099,N_13161);
or U13423 (N_13423,N_13213,N_13001);
nand U13424 (N_13424,N_13110,N_13149);
nand U13425 (N_13425,N_13154,N_13173);
nor U13426 (N_13426,N_13119,N_13084);
nand U13427 (N_13427,N_13202,N_13195);
and U13428 (N_13428,N_13117,N_13086);
or U13429 (N_13429,N_13054,N_13151);
nand U13430 (N_13430,N_13173,N_13218);
and U13431 (N_13431,N_13100,N_13174);
nand U13432 (N_13432,N_13220,N_13096);
and U13433 (N_13433,N_13230,N_13071);
nand U13434 (N_13434,N_13087,N_13108);
nor U13435 (N_13435,N_13068,N_13150);
or U13436 (N_13436,N_13155,N_13182);
nor U13437 (N_13437,N_13010,N_13199);
xnor U13438 (N_13438,N_13033,N_13008);
and U13439 (N_13439,N_13165,N_13014);
or U13440 (N_13440,N_13032,N_13069);
or U13441 (N_13441,N_13179,N_13030);
or U13442 (N_13442,N_13082,N_13176);
xnor U13443 (N_13443,N_13053,N_13150);
nand U13444 (N_13444,N_13209,N_13227);
xnor U13445 (N_13445,N_13054,N_13018);
nor U13446 (N_13446,N_13031,N_13199);
nor U13447 (N_13447,N_13002,N_13217);
nor U13448 (N_13448,N_13047,N_13129);
nand U13449 (N_13449,N_13102,N_13002);
xor U13450 (N_13450,N_13142,N_13046);
or U13451 (N_13451,N_13143,N_13249);
and U13452 (N_13452,N_13117,N_13008);
nand U13453 (N_13453,N_13088,N_13200);
or U13454 (N_13454,N_13211,N_13146);
nand U13455 (N_13455,N_13024,N_13057);
and U13456 (N_13456,N_13118,N_13237);
xnor U13457 (N_13457,N_13177,N_13235);
nand U13458 (N_13458,N_13006,N_13037);
and U13459 (N_13459,N_13098,N_13167);
nor U13460 (N_13460,N_13177,N_13200);
nor U13461 (N_13461,N_13093,N_13097);
nand U13462 (N_13462,N_13019,N_13088);
or U13463 (N_13463,N_13100,N_13193);
nand U13464 (N_13464,N_13150,N_13015);
nor U13465 (N_13465,N_13155,N_13195);
nor U13466 (N_13466,N_13249,N_13219);
nor U13467 (N_13467,N_13115,N_13243);
nand U13468 (N_13468,N_13114,N_13139);
nor U13469 (N_13469,N_13065,N_13223);
and U13470 (N_13470,N_13208,N_13173);
xor U13471 (N_13471,N_13097,N_13130);
nand U13472 (N_13472,N_13241,N_13216);
nor U13473 (N_13473,N_13108,N_13117);
and U13474 (N_13474,N_13144,N_13207);
xnor U13475 (N_13475,N_13087,N_13220);
nand U13476 (N_13476,N_13032,N_13108);
nor U13477 (N_13477,N_13002,N_13171);
xnor U13478 (N_13478,N_13114,N_13222);
nor U13479 (N_13479,N_13116,N_13177);
or U13480 (N_13480,N_13228,N_13204);
nand U13481 (N_13481,N_13152,N_13208);
nor U13482 (N_13482,N_13031,N_13242);
nor U13483 (N_13483,N_13116,N_13003);
or U13484 (N_13484,N_13134,N_13101);
nor U13485 (N_13485,N_13070,N_13065);
nand U13486 (N_13486,N_13139,N_13023);
xor U13487 (N_13487,N_13221,N_13227);
and U13488 (N_13488,N_13150,N_13006);
or U13489 (N_13489,N_13100,N_13112);
and U13490 (N_13490,N_13149,N_13071);
nand U13491 (N_13491,N_13164,N_13143);
or U13492 (N_13492,N_13011,N_13249);
xor U13493 (N_13493,N_13007,N_13082);
nand U13494 (N_13494,N_13143,N_13151);
or U13495 (N_13495,N_13227,N_13138);
or U13496 (N_13496,N_13218,N_13003);
nand U13497 (N_13497,N_13106,N_13095);
nor U13498 (N_13498,N_13078,N_13209);
xor U13499 (N_13499,N_13241,N_13208);
or U13500 (N_13500,N_13254,N_13328);
nor U13501 (N_13501,N_13450,N_13326);
xor U13502 (N_13502,N_13394,N_13415);
and U13503 (N_13503,N_13344,N_13346);
nand U13504 (N_13504,N_13358,N_13263);
nand U13505 (N_13505,N_13362,N_13476);
nor U13506 (N_13506,N_13436,N_13386);
and U13507 (N_13507,N_13469,N_13342);
nor U13508 (N_13508,N_13286,N_13492);
and U13509 (N_13509,N_13434,N_13266);
xor U13510 (N_13510,N_13473,N_13491);
and U13511 (N_13511,N_13417,N_13451);
or U13512 (N_13512,N_13317,N_13462);
nor U13513 (N_13513,N_13308,N_13453);
nor U13514 (N_13514,N_13290,N_13371);
or U13515 (N_13515,N_13384,N_13423);
or U13516 (N_13516,N_13457,N_13425);
nand U13517 (N_13517,N_13259,N_13400);
or U13518 (N_13518,N_13255,N_13474);
nor U13519 (N_13519,N_13332,N_13442);
nand U13520 (N_13520,N_13305,N_13275);
and U13521 (N_13521,N_13370,N_13419);
and U13522 (N_13522,N_13281,N_13452);
xnor U13523 (N_13523,N_13265,N_13416);
xor U13524 (N_13524,N_13282,N_13293);
or U13525 (N_13525,N_13338,N_13264);
xnor U13526 (N_13526,N_13253,N_13294);
xor U13527 (N_13527,N_13279,N_13257);
or U13528 (N_13528,N_13349,N_13427);
nor U13529 (N_13529,N_13373,N_13289);
and U13530 (N_13530,N_13356,N_13463);
and U13531 (N_13531,N_13260,N_13341);
nor U13532 (N_13532,N_13420,N_13331);
xnor U13533 (N_13533,N_13385,N_13489);
xnor U13534 (N_13534,N_13418,N_13430);
nor U13535 (N_13535,N_13399,N_13404);
xnor U13536 (N_13536,N_13449,N_13359);
and U13537 (N_13537,N_13318,N_13475);
or U13538 (N_13538,N_13488,N_13322);
xnor U13539 (N_13539,N_13313,N_13296);
xnor U13540 (N_13540,N_13273,N_13262);
xor U13541 (N_13541,N_13319,N_13292);
and U13542 (N_13542,N_13377,N_13479);
and U13543 (N_13543,N_13432,N_13464);
xnor U13544 (N_13544,N_13276,N_13390);
and U13545 (N_13545,N_13304,N_13440);
nand U13546 (N_13546,N_13334,N_13340);
or U13547 (N_13547,N_13306,N_13354);
or U13548 (N_13548,N_13446,N_13287);
nand U13549 (N_13549,N_13407,N_13443);
and U13550 (N_13550,N_13277,N_13361);
or U13551 (N_13551,N_13398,N_13363);
nand U13552 (N_13552,N_13393,N_13312);
or U13553 (N_13553,N_13366,N_13378);
xnor U13554 (N_13554,N_13498,N_13261);
and U13555 (N_13555,N_13278,N_13499);
xor U13556 (N_13556,N_13320,N_13483);
nor U13557 (N_13557,N_13468,N_13480);
xnor U13558 (N_13558,N_13395,N_13329);
and U13559 (N_13559,N_13347,N_13481);
nor U13560 (N_13560,N_13337,N_13327);
xor U13561 (N_13561,N_13323,N_13343);
or U13562 (N_13562,N_13402,N_13309);
and U13563 (N_13563,N_13381,N_13274);
or U13564 (N_13564,N_13497,N_13321);
xnor U13565 (N_13565,N_13369,N_13471);
or U13566 (N_13566,N_13314,N_13297);
and U13567 (N_13567,N_13397,N_13339);
nor U13568 (N_13568,N_13350,N_13303);
nand U13569 (N_13569,N_13403,N_13269);
nand U13570 (N_13570,N_13439,N_13258);
nor U13571 (N_13571,N_13298,N_13285);
nand U13572 (N_13572,N_13335,N_13428);
and U13573 (N_13573,N_13267,N_13360);
xnor U13574 (N_13574,N_13250,N_13272);
nor U13575 (N_13575,N_13352,N_13355);
xor U13576 (N_13576,N_13301,N_13494);
nand U13577 (N_13577,N_13429,N_13367);
or U13578 (N_13578,N_13484,N_13421);
nand U13579 (N_13579,N_13495,N_13299);
or U13580 (N_13580,N_13380,N_13316);
xnor U13581 (N_13581,N_13383,N_13412);
xor U13582 (N_13582,N_13409,N_13372);
nor U13583 (N_13583,N_13368,N_13477);
and U13584 (N_13584,N_13283,N_13379);
and U13585 (N_13585,N_13365,N_13325);
nand U13586 (N_13586,N_13351,N_13447);
or U13587 (N_13587,N_13490,N_13467);
and U13588 (N_13588,N_13410,N_13461);
nor U13589 (N_13589,N_13311,N_13315);
nand U13590 (N_13590,N_13396,N_13268);
nor U13591 (N_13591,N_13310,N_13435);
nor U13592 (N_13592,N_13433,N_13458);
and U13593 (N_13593,N_13405,N_13441);
or U13594 (N_13594,N_13413,N_13391);
and U13595 (N_13595,N_13460,N_13376);
nor U13596 (N_13596,N_13389,N_13382);
xnor U13597 (N_13597,N_13375,N_13401);
nand U13598 (N_13598,N_13388,N_13353);
and U13599 (N_13599,N_13387,N_13493);
or U13600 (N_13600,N_13459,N_13324);
and U13601 (N_13601,N_13348,N_13445);
or U13602 (N_13602,N_13431,N_13496);
nor U13603 (N_13603,N_13288,N_13426);
and U13604 (N_13604,N_13437,N_13252);
xor U13605 (N_13605,N_13251,N_13465);
or U13606 (N_13606,N_13336,N_13411);
xnor U13607 (N_13607,N_13454,N_13295);
nor U13608 (N_13608,N_13270,N_13374);
and U13609 (N_13609,N_13364,N_13448);
nor U13610 (N_13610,N_13470,N_13422);
or U13611 (N_13611,N_13300,N_13456);
xnor U13612 (N_13612,N_13291,N_13438);
nor U13613 (N_13613,N_13414,N_13408);
and U13614 (N_13614,N_13485,N_13486);
and U13615 (N_13615,N_13280,N_13284);
or U13616 (N_13616,N_13307,N_13271);
nand U13617 (N_13617,N_13256,N_13444);
and U13618 (N_13618,N_13330,N_13472);
and U13619 (N_13619,N_13466,N_13487);
xor U13620 (N_13620,N_13406,N_13392);
xor U13621 (N_13621,N_13302,N_13478);
or U13622 (N_13622,N_13357,N_13482);
or U13623 (N_13623,N_13333,N_13455);
and U13624 (N_13624,N_13345,N_13424);
nor U13625 (N_13625,N_13456,N_13469);
and U13626 (N_13626,N_13345,N_13489);
and U13627 (N_13627,N_13271,N_13464);
nand U13628 (N_13628,N_13484,N_13276);
xor U13629 (N_13629,N_13493,N_13279);
xnor U13630 (N_13630,N_13253,N_13382);
or U13631 (N_13631,N_13312,N_13418);
nand U13632 (N_13632,N_13400,N_13288);
nor U13633 (N_13633,N_13299,N_13430);
nor U13634 (N_13634,N_13346,N_13461);
or U13635 (N_13635,N_13405,N_13418);
nand U13636 (N_13636,N_13437,N_13447);
nor U13637 (N_13637,N_13259,N_13380);
or U13638 (N_13638,N_13412,N_13262);
xnor U13639 (N_13639,N_13358,N_13435);
and U13640 (N_13640,N_13473,N_13356);
or U13641 (N_13641,N_13286,N_13370);
nand U13642 (N_13642,N_13364,N_13345);
xor U13643 (N_13643,N_13434,N_13351);
and U13644 (N_13644,N_13274,N_13408);
xnor U13645 (N_13645,N_13387,N_13473);
xnor U13646 (N_13646,N_13268,N_13258);
and U13647 (N_13647,N_13268,N_13483);
and U13648 (N_13648,N_13456,N_13312);
xor U13649 (N_13649,N_13323,N_13340);
and U13650 (N_13650,N_13286,N_13410);
nor U13651 (N_13651,N_13268,N_13308);
and U13652 (N_13652,N_13355,N_13381);
nand U13653 (N_13653,N_13329,N_13257);
and U13654 (N_13654,N_13330,N_13310);
and U13655 (N_13655,N_13314,N_13474);
and U13656 (N_13656,N_13289,N_13277);
and U13657 (N_13657,N_13466,N_13355);
nor U13658 (N_13658,N_13497,N_13251);
and U13659 (N_13659,N_13492,N_13260);
nand U13660 (N_13660,N_13386,N_13375);
or U13661 (N_13661,N_13341,N_13455);
or U13662 (N_13662,N_13375,N_13461);
or U13663 (N_13663,N_13473,N_13345);
xnor U13664 (N_13664,N_13342,N_13353);
and U13665 (N_13665,N_13347,N_13275);
or U13666 (N_13666,N_13375,N_13422);
nor U13667 (N_13667,N_13323,N_13413);
and U13668 (N_13668,N_13403,N_13450);
or U13669 (N_13669,N_13311,N_13254);
nor U13670 (N_13670,N_13474,N_13389);
nor U13671 (N_13671,N_13295,N_13379);
nand U13672 (N_13672,N_13464,N_13474);
nor U13673 (N_13673,N_13322,N_13262);
nor U13674 (N_13674,N_13479,N_13350);
nand U13675 (N_13675,N_13290,N_13326);
xor U13676 (N_13676,N_13455,N_13330);
xnor U13677 (N_13677,N_13419,N_13393);
nand U13678 (N_13678,N_13332,N_13303);
nor U13679 (N_13679,N_13432,N_13405);
xor U13680 (N_13680,N_13321,N_13401);
xnor U13681 (N_13681,N_13275,N_13494);
xor U13682 (N_13682,N_13426,N_13311);
nor U13683 (N_13683,N_13250,N_13447);
nor U13684 (N_13684,N_13378,N_13364);
or U13685 (N_13685,N_13453,N_13426);
and U13686 (N_13686,N_13274,N_13393);
nor U13687 (N_13687,N_13287,N_13451);
nand U13688 (N_13688,N_13355,N_13443);
or U13689 (N_13689,N_13481,N_13352);
or U13690 (N_13690,N_13426,N_13433);
nand U13691 (N_13691,N_13287,N_13488);
xnor U13692 (N_13692,N_13312,N_13304);
and U13693 (N_13693,N_13451,N_13335);
or U13694 (N_13694,N_13386,N_13443);
nor U13695 (N_13695,N_13406,N_13404);
nor U13696 (N_13696,N_13309,N_13412);
xor U13697 (N_13697,N_13415,N_13455);
or U13698 (N_13698,N_13474,N_13258);
nand U13699 (N_13699,N_13265,N_13272);
nor U13700 (N_13700,N_13363,N_13318);
xor U13701 (N_13701,N_13340,N_13352);
xnor U13702 (N_13702,N_13282,N_13317);
or U13703 (N_13703,N_13322,N_13388);
nor U13704 (N_13704,N_13443,N_13321);
xor U13705 (N_13705,N_13356,N_13313);
or U13706 (N_13706,N_13288,N_13313);
nand U13707 (N_13707,N_13303,N_13299);
nor U13708 (N_13708,N_13487,N_13410);
nand U13709 (N_13709,N_13451,N_13462);
nand U13710 (N_13710,N_13464,N_13379);
and U13711 (N_13711,N_13394,N_13275);
nor U13712 (N_13712,N_13294,N_13252);
nor U13713 (N_13713,N_13260,N_13257);
nor U13714 (N_13714,N_13291,N_13382);
or U13715 (N_13715,N_13295,N_13394);
and U13716 (N_13716,N_13314,N_13380);
xnor U13717 (N_13717,N_13373,N_13383);
nand U13718 (N_13718,N_13364,N_13401);
or U13719 (N_13719,N_13427,N_13336);
nor U13720 (N_13720,N_13341,N_13321);
nor U13721 (N_13721,N_13278,N_13401);
or U13722 (N_13722,N_13381,N_13431);
nor U13723 (N_13723,N_13265,N_13299);
or U13724 (N_13724,N_13423,N_13491);
xor U13725 (N_13725,N_13472,N_13465);
xor U13726 (N_13726,N_13278,N_13435);
nor U13727 (N_13727,N_13385,N_13297);
nand U13728 (N_13728,N_13499,N_13272);
and U13729 (N_13729,N_13272,N_13407);
nand U13730 (N_13730,N_13298,N_13453);
or U13731 (N_13731,N_13466,N_13400);
nand U13732 (N_13732,N_13284,N_13270);
nor U13733 (N_13733,N_13307,N_13343);
xnor U13734 (N_13734,N_13318,N_13497);
xnor U13735 (N_13735,N_13426,N_13484);
xor U13736 (N_13736,N_13458,N_13475);
and U13737 (N_13737,N_13453,N_13285);
or U13738 (N_13738,N_13469,N_13454);
nand U13739 (N_13739,N_13449,N_13437);
nor U13740 (N_13740,N_13334,N_13251);
nand U13741 (N_13741,N_13353,N_13487);
and U13742 (N_13742,N_13269,N_13368);
nor U13743 (N_13743,N_13440,N_13467);
nor U13744 (N_13744,N_13360,N_13384);
and U13745 (N_13745,N_13283,N_13260);
and U13746 (N_13746,N_13436,N_13362);
and U13747 (N_13747,N_13471,N_13495);
nand U13748 (N_13748,N_13302,N_13378);
xor U13749 (N_13749,N_13299,N_13312);
xnor U13750 (N_13750,N_13715,N_13576);
or U13751 (N_13751,N_13607,N_13537);
and U13752 (N_13752,N_13746,N_13684);
or U13753 (N_13753,N_13631,N_13596);
nand U13754 (N_13754,N_13729,N_13527);
nor U13755 (N_13755,N_13720,N_13690);
or U13756 (N_13756,N_13740,N_13653);
and U13757 (N_13757,N_13515,N_13736);
nor U13758 (N_13758,N_13745,N_13541);
and U13759 (N_13759,N_13591,N_13513);
xor U13760 (N_13760,N_13711,N_13521);
and U13761 (N_13761,N_13622,N_13669);
and U13762 (N_13762,N_13635,N_13639);
xor U13763 (N_13763,N_13712,N_13553);
xnor U13764 (N_13764,N_13749,N_13662);
nand U13765 (N_13765,N_13713,N_13504);
nor U13766 (N_13766,N_13636,N_13608);
or U13767 (N_13767,N_13678,N_13721);
or U13768 (N_13768,N_13701,N_13546);
nand U13769 (N_13769,N_13612,N_13585);
or U13770 (N_13770,N_13747,N_13681);
nand U13771 (N_13771,N_13718,N_13531);
nor U13772 (N_13772,N_13675,N_13544);
or U13773 (N_13773,N_13558,N_13547);
or U13774 (N_13774,N_13658,N_13647);
nand U13775 (N_13775,N_13672,N_13642);
and U13776 (N_13776,N_13543,N_13510);
and U13777 (N_13777,N_13560,N_13624);
xnor U13778 (N_13778,N_13522,N_13698);
nand U13779 (N_13779,N_13643,N_13732);
nand U13780 (N_13780,N_13676,N_13691);
xnor U13781 (N_13781,N_13630,N_13735);
and U13782 (N_13782,N_13739,N_13589);
xnor U13783 (N_13783,N_13707,N_13696);
and U13784 (N_13784,N_13501,N_13551);
and U13785 (N_13785,N_13562,N_13697);
xor U13786 (N_13786,N_13660,N_13529);
and U13787 (N_13787,N_13533,N_13657);
and U13788 (N_13788,N_13604,N_13619);
nor U13789 (N_13789,N_13623,N_13683);
xor U13790 (N_13790,N_13561,N_13569);
xor U13791 (N_13791,N_13679,N_13530);
and U13792 (N_13792,N_13606,N_13629);
nor U13793 (N_13793,N_13526,N_13656);
and U13794 (N_13794,N_13689,N_13685);
or U13795 (N_13795,N_13620,N_13525);
or U13796 (N_13796,N_13725,N_13563);
or U13797 (N_13797,N_13613,N_13556);
and U13798 (N_13798,N_13542,N_13634);
and U13799 (N_13799,N_13644,N_13733);
nor U13800 (N_13800,N_13555,N_13540);
nor U13801 (N_13801,N_13700,N_13570);
xnor U13802 (N_13802,N_13580,N_13655);
xnor U13803 (N_13803,N_13605,N_13584);
and U13804 (N_13804,N_13706,N_13695);
xor U13805 (N_13805,N_13516,N_13566);
nor U13806 (N_13806,N_13550,N_13661);
or U13807 (N_13807,N_13595,N_13677);
xnor U13808 (N_13808,N_13523,N_13659);
xnor U13809 (N_13809,N_13668,N_13500);
nand U13810 (N_13810,N_13719,N_13680);
nor U13811 (N_13811,N_13709,N_13552);
nand U13812 (N_13812,N_13667,N_13625);
and U13813 (N_13813,N_13666,N_13694);
xnor U13814 (N_13814,N_13723,N_13615);
nor U13815 (N_13815,N_13532,N_13524);
nor U13816 (N_13816,N_13617,N_13693);
or U13817 (N_13817,N_13512,N_13616);
or U13818 (N_13818,N_13650,N_13599);
xnor U13819 (N_13819,N_13534,N_13559);
and U13820 (N_13820,N_13600,N_13572);
or U13821 (N_13821,N_13536,N_13614);
nand U13822 (N_13822,N_13633,N_13673);
nand U13823 (N_13823,N_13727,N_13734);
nor U13824 (N_13824,N_13628,N_13593);
nor U13825 (N_13825,N_13507,N_13519);
xor U13826 (N_13826,N_13538,N_13575);
and U13827 (N_13827,N_13654,N_13603);
or U13828 (N_13828,N_13621,N_13671);
and U13829 (N_13829,N_13687,N_13705);
and U13830 (N_13830,N_13743,N_13646);
or U13831 (N_13831,N_13598,N_13640);
nand U13832 (N_13832,N_13539,N_13511);
and U13833 (N_13833,N_13557,N_13688);
nor U13834 (N_13834,N_13549,N_13641);
nor U13835 (N_13835,N_13602,N_13577);
xnor U13836 (N_13836,N_13514,N_13737);
nor U13837 (N_13837,N_13545,N_13573);
and U13838 (N_13838,N_13583,N_13742);
and U13839 (N_13839,N_13748,N_13590);
nand U13840 (N_13840,N_13651,N_13611);
xnor U13841 (N_13841,N_13638,N_13565);
nor U13842 (N_13842,N_13664,N_13518);
or U13843 (N_13843,N_13509,N_13674);
or U13844 (N_13844,N_13665,N_13503);
and U13845 (N_13845,N_13564,N_13710);
xor U13846 (N_13846,N_13682,N_13609);
nand U13847 (N_13847,N_13726,N_13571);
or U13848 (N_13848,N_13722,N_13738);
nand U13849 (N_13849,N_13692,N_13535);
xnor U13850 (N_13850,N_13730,N_13744);
xor U13851 (N_13851,N_13508,N_13601);
nor U13852 (N_13852,N_13502,N_13567);
and U13853 (N_13853,N_13582,N_13649);
or U13854 (N_13854,N_13717,N_13704);
or U13855 (N_13855,N_13626,N_13716);
xor U13856 (N_13856,N_13592,N_13548);
or U13857 (N_13857,N_13632,N_13618);
and U13858 (N_13858,N_13702,N_13506);
and U13859 (N_13859,N_13741,N_13554);
or U13860 (N_13860,N_13597,N_13581);
nand U13861 (N_13861,N_13594,N_13587);
or U13862 (N_13862,N_13588,N_13728);
nand U13863 (N_13863,N_13708,N_13648);
xor U13864 (N_13864,N_13578,N_13610);
xnor U13865 (N_13865,N_13505,N_13670);
nand U13866 (N_13866,N_13703,N_13637);
nor U13867 (N_13867,N_13568,N_13579);
and U13868 (N_13868,N_13699,N_13652);
nand U13869 (N_13869,N_13686,N_13724);
nor U13870 (N_13870,N_13663,N_13517);
and U13871 (N_13871,N_13520,N_13574);
and U13872 (N_13872,N_13645,N_13586);
nor U13873 (N_13873,N_13627,N_13528);
nand U13874 (N_13874,N_13714,N_13731);
xnor U13875 (N_13875,N_13583,N_13685);
xor U13876 (N_13876,N_13691,N_13662);
xor U13877 (N_13877,N_13691,N_13703);
xnor U13878 (N_13878,N_13749,N_13573);
xnor U13879 (N_13879,N_13647,N_13619);
nand U13880 (N_13880,N_13584,N_13650);
or U13881 (N_13881,N_13666,N_13710);
nor U13882 (N_13882,N_13562,N_13727);
nand U13883 (N_13883,N_13678,N_13523);
nor U13884 (N_13884,N_13596,N_13594);
and U13885 (N_13885,N_13575,N_13580);
and U13886 (N_13886,N_13525,N_13505);
and U13887 (N_13887,N_13666,N_13733);
or U13888 (N_13888,N_13731,N_13710);
xnor U13889 (N_13889,N_13540,N_13678);
xor U13890 (N_13890,N_13521,N_13610);
and U13891 (N_13891,N_13722,N_13683);
xnor U13892 (N_13892,N_13564,N_13673);
and U13893 (N_13893,N_13594,N_13644);
and U13894 (N_13894,N_13691,N_13693);
xnor U13895 (N_13895,N_13736,N_13501);
or U13896 (N_13896,N_13608,N_13576);
nor U13897 (N_13897,N_13613,N_13650);
xor U13898 (N_13898,N_13692,N_13613);
and U13899 (N_13899,N_13599,N_13543);
or U13900 (N_13900,N_13633,N_13655);
nand U13901 (N_13901,N_13635,N_13512);
and U13902 (N_13902,N_13658,N_13709);
xnor U13903 (N_13903,N_13674,N_13569);
nand U13904 (N_13904,N_13610,N_13736);
or U13905 (N_13905,N_13618,N_13527);
or U13906 (N_13906,N_13506,N_13598);
nor U13907 (N_13907,N_13656,N_13516);
and U13908 (N_13908,N_13613,N_13684);
nand U13909 (N_13909,N_13716,N_13674);
and U13910 (N_13910,N_13602,N_13654);
nand U13911 (N_13911,N_13591,N_13741);
nand U13912 (N_13912,N_13710,N_13741);
xor U13913 (N_13913,N_13602,N_13671);
and U13914 (N_13914,N_13547,N_13549);
xor U13915 (N_13915,N_13552,N_13723);
and U13916 (N_13916,N_13627,N_13742);
nor U13917 (N_13917,N_13626,N_13574);
xnor U13918 (N_13918,N_13518,N_13520);
nand U13919 (N_13919,N_13714,N_13555);
xor U13920 (N_13920,N_13733,N_13561);
xnor U13921 (N_13921,N_13661,N_13620);
and U13922 (N_13922,N_13683,N_13594);
nand U13923 (N_13923,N_13525,N_13533);
nand U13924 (N_13924,N_13582,N_13516);
and U13925 (N_13925,N_13544,N_13512);
xor U13926 (N_13926,N_13685,N_13517);
and U13927 (N_13927,N_13601,N_13649);
nor U13928 (N_13928,N_13621,N_13609);
and U13929 (N_13929,N_13640,N_13588);
nor U13930 (N_13930,N_13678,N_13711);
and U13931 (N_13931,N_13682,N_13549);
and U13932 (N_13932,N_13545,N_13630);
and U13933 (N_13933,N_13541,N_13577);
nor U13934 (N_13934,N_13730,N_13567);
xnor U13935 (N_13935,N_13511,N_13640);
xor U13936 (N_13936,N_13688,N_13693);
or U13937 (N_13937,N_13550,N_13633);
nand U13938 (N_13938,N_13688,N_13682);
and U13939 (N_13939,N_13560,N_13519);
or U13940 (N_13940,N_13616,N_13717);
nor U13941 (N_13941,N_13512,N_13682);
or U13942 (N_13942,N_13629,N_13687);
or U13943 (N_13943,N_13636,N_13583);
or U13944 (N_13944,N_13541,N_13678);
and U13945 (N_13945,N_13512,N_13547);
nand U13946 (N_13946,N_13598,N_13714);
xnor U13947 (N_13947,N_13740,N_13552);
nor U13948 (N_13948,N_13581,N_13637);
or U13949 (N_13949,N_13558,N_13664);
or U13950 (N_13950,N_13627,N_13746);
or U13951 (N_13951,N_13623,N_13741);
nand U13952 (N_13952,N_13523,N_13506);
nor U13953 (N_13953,N_13623,N_13554);
nor U13954 (N_13954,N_13721,N_13647);
xor U13955 (N_13955,N_13625,N_13564);
nor U13956 (N_13956,N_13506,N_13705);
or U13957 (N_13957,N_13528,N_13552);
or U13958 (N_13958,N_13630,N_13687);
nor U13959 (N_13959,N_13524,N_13566);
and U13960 (N_13960,N_13515,N_13620);
nor U13961 (N_13961,N_13514,N_13713);
or U13962 (N_13962,N_13533,N_13703);
xor U13963 (N_13963,N_13512,N_13625);
nand U13964 (N_13964,N_13621,N_13557);
xnor U13965 (N_13965,N_13636,N_13682);
xor U13966 (N_13966,N_13737,N_13662);
or U13967 (N_13967,N_13749,N_13541);
nor U13968 (N_13968,N_13736,N_13657);
nor U13969 (N_13969,N_13523,N_13603);
nand U13970 (N_13970,N_13502,N_13548);
nand U13971 (N_13971,N_13674,N_13659);
and U13972 (N_13972,N_13727,N_13534);
xnor U13973 (N_13973,N_13656,N_13569);
nand U13974 (N_13974,N_13540,N_13562);
xor U13975 (N_13975,N_13545,N_13613);
nand U13976 (N_13976,N_13660,N_13566);
or U13977 (N_13977,N_13506,N_13557);
xor U13978 (N_13978,N_13574,N_13592);
nand U13979 (N_13979,N_13688,N_13712);
nor U13980 (N_13980,N_13671,N_13529);
xor U13981 (N_13981,N_13684,N_13537);
xor U13982 (N_13982,N_13509,N_13554);
nor U13983 (N_13983,N_13558,N_13673);
xor U13984 (N_13984,N_13693,N_13653);
or U13985 (N_13985,N_13569,N_13578);
and U13986 (N_13986,N_13634,N_13577);
nor U13987 (N_13987,N_13578,N_13563);
and U13988 (N_13988,N_13636,N_13689);
nor U13989 (N_13989,N_13722,N_13633);
nor U13990 (N_13990,N_13684,N_13650);
nor U13991 (N_13991,N_13614,N_13608);
nor U13992 (N_13992,N_13735,N_13596);
nand U13993 (N_13993,N_13510,N_13686);
xnor U13994 (N_13994,N_13677,N_13747);
nor U13995 (N_13995,N_13505,N_13673);
or U13996 (N_13996,N_13627,N_13573);
or U13997 (N_13997,N_13513,N_13716);
and U13998 (N_13998,N_13604,N_13557);
nand U13999 (N_13999,N_13613,N_13539);
xnor U14000 (N_14000,N_13845,N_13815);
nor U14001 (N_14001,N_13956,N_13888);
or U14002 (N_14002,N_13876,N_13880);
nor U14003 (N_14003,N_13847,N_13823);
nand U14004 (N_14004,N_13899,N_13891);
or U14005 (N_14005,N_13821,N_13933);
nand U14006 (N_14006,N_13841,N_13837);
nand U14007 (N_14007,N_13895,N_13762);
nor U14008 (N_14008,N_13921,N_13819);
or U14009 (N_14009,N_13926,N_13976);
nor U14010 (N_14010,N_13767,N_13804);
and U14011 (N_14011,N_13958,N_13860);
nand U14012 (N_14012,N_13853,N_13934);
or U14013 (N_14013,N_13817,N_13828);
xnor U14014 (N_14014,N_13941,N_13961);
and U14015 (N_14015,N_13945,N_13893);
or U14016 (N_14016,N_13826,N_13839);
and U14017 (N_14017,N_13766,N_13808);
nor U14018 (N_14018,N_13981,N_13750);
nor U14019 (N_14019,N_13781,N_13843);
nand U14020 (N_14020,N_13756,N_13970);
nor U14021 (N_14021,N_13792,N_13890);
or U14022 (N_14022,N_13922,N_13832);
or U14023 (N_14023,N_13835,N_13783);
nand U14024 (N_14024,N_13807,N_13829);
or U14025 (N_14025,N_13963,N_13882);
or U14026 (N_14026,N_13915,N_13789);
nor U14027 (N_14027,N_13866,N_13753);
and U14028 (N_14028,N_13889,N_13858);
nand U14029 (N_14029,N_13770,N_13869);
or U14030 (N_14030,N_13814,N_13831);
or U14031 (N_14031,N_13992,N_13914);
or U14032 (N_14032,N_13944,N_13947);
nand U14033 (N_14033,N_13959,N_13946);
xor U14034 (N_14034,N_13928,N_13885);
and U14035 (N_14035,N_13952,N_13902);
nand U14036 (N_14036,N_13898,N_13862);
xor U14037 (N_14037,N_13769,N_13780);
or U14038 (N_14038,N_13938,N_13875);
nor U14039 (N_14039,N_13951,N_13972);
nor U14040 (N_14040,N_13910,N_13818);
or U14041 (N_14041,N_13751,N_13916);
or U14042 (N_14042,N_13846,N_13986);
and U14043 (N_14043,N_13903,N_13897);
and U14044 (N_14044,N_13840,N_13948);
and U14045 (N_14045,N_13881,N_13811);
xnor U14046 (N_14046,N_13854,N_13791);
xor U14047 (N_14047,N_13975,N_13793);
xnor U14048 (N_14048,N_13803,N_13939);
nor U14049 (N_14049,N_13787,N_13870);
or U14050 (N_14050,N_13852,N_13937);
nor U14051 (N_14051,N_13964,N_13772);
nor U14052 (N_14052,N_13824,N_13873);
or U14053 (N_14053,N_13782,N_13918);
xor U14054 (N_14054,N_13949,N_13901);
nand U14055 (N_14055,N_13844,N_13812);
xor U14056 (N_14056,N_13872,N_13940);
xor U14057 (N_14057,N_13834,N_13987);
or U14058 (N_14058,N_13919,N_13871);
xnor U14059 (N_14059,N_13950,N_13813);
nand U14060 (N_14060,N_13884,N_13966);
and U14061 (N_14061,N_13758,N_13773);
nand U14062 (N_14062,N_13996,N_13927);
and U14063 (N_14063,N_13822,N_13864);
xnor U14064 (N_14064,N_13760,N_13931);
and U14065 (N_14065,N_13763,N_13994);
nand U14066 (N_14066,N_13920,N_13932);
nand U14067 (N_14067,N_13974,N_13816);
nor U14068 (N_14068,N_13968,N_13833);
xnor U14069 (N_14069,N_13776,N_13985);
nand U14070 (N_14070,N_13953,N_13957);
nor U14071 (N_14071,N_13930,N_13993);
xor U14072 (N_14072,N_13861,N_13809);
nand U14073 (N_14073,N_13923,N_13806);
nand U14074 (N_14074,N_13863,N_13757);
and U14075 (N_14075,N_13983,N_13779);
and U14076 (N_14076,N_13942,N_13797);
nand U14077 (N_14077,N_13984,N_13795);
or U14078 (N_14078,N_13790,N_13905);
xor U14079 (N_14079,N_13786,N_13755);
or U14080 (N_14080,N_13973,N_13785);
xor U14081 (N_14081,N_13764,N_13925);
and U14082 (N_14082,N_13851,N_13857);
nand U14083 (N_14083,N_13802,N_13894);
xor U14084 (N_14084,N_13887,N_13859);
nor U14085 (N_14085,N_13917,N_13825);
or U14086 (N_14086,N_13849,N_13874);
xnor U14087 (N_14087,N_13877,N_13886);
nor U14088 (N_14088,N_13868,N_13896);
and U14089 (N_14089,N_13913,N_13954);
or U14090 (N_14090,N_13867,N_13892);
xnor U14091 (N_14091,N_13778,N_13759);
xor U14092 (N_14092,N_13788,N_13799);
or U14093 (N_14093,N_13924,N_13798);
nand U14094 (N_14094,N_13969,N_13962);
or U14095 (N_14095,N_13908,N_13912);
xor U14096 (N_14096,N_13906,N_13754);
nand U14097 (N_14097,N_13988,N_13827);
xor U14098 (N_14098,N_13929,N_13768);
nor U14099 (N_14099,N_13999,N_13907);
xor U14100 (N_14100,N_13982,N_13800);
or U14101 (N_14101,N_13796,N_13960);
and U14102 (N_14102,N_13943,N_13794);
or U14103 (N_14103,N_13878,N_13911);
nor U14104 (N_14104,N_13842,N_13855);
nand U14105 (N_14105,N_13991,N_13900);
and U14106 (N_14106,N_13967,N_13904);
or U14107 (N_14107,N_13850,N_13980);
nor U14108 (N_14108,N_13978,N_13801);
nand U14109 (N_14109,N_13830,N_13998);
nor U14110 (N_14110,N_13836,N_13761);
nor U14111 (N_14111,N_13971,N_13856);
nor U14112 (N_14112,N_13883,N_13965);
xnor U14113 (N_14113,N_13990,N_13997);
nand U14114 (N_14114,N_13936,N_13820);
nor U14115 (N_14115,N_13935,N_13909);
nand U14116 (N_14116,N_13805,N_13784);
xor U14117 (N_14117,N_13955,N_13810);
or U14118 (N_14118,N_13979,N_13879);
nor U14119 (N_14119,N_13995,N_13775);
nand U14120 (N_14120,N_13777,N_13989);
and U14121 (N_14121,N_13838,N_13848);
or U14122 (N_14122,N_13774,N_13771);
xnor U14123 (N_14123,N_13752,N_13977);
nor U14124 (N_14124,N_13865,N_13765);
nor U14125 (N_14125,N_13873,N_13915);
nor U14126 (N_14126,N_13923,N_13965);
nor U14127 (N_14127,N_13876,N_13940);
xnor U14128 (N_14128,N_13969,N_13839);
nor U14129 (N_14129,N_13854,N_13852);
and U14130 (N_14130,N_13870,N_13761);
nand U14131 (N_14131,N_13782,N_13910);
nor U14132 (N_14132,N_13772,N_13884);
nor U14133 (N_14133,N_13853,N_13960);
nand U14134 (N_14134,N_13844,N_13777);
nor U14135 (N_14135,N_13984,N_13893);
nand U14136 (N_14136,N_13922,N_13770);
and U14137 (N_14137,N_13836,N_13989);
and U14138 (N_14138,N_13972,N_13944);
nor U14139 (N_14139,N_13842,N_13813);
or U14140 (N_14140,N_13975,N_13884);
or U14141 (N_14141,N_13901,N_13792);
xnor U14142 (N_14142,N_13850,N_13810);
nor U14143 (N_14143,N_13848,N_13956);
nand U14144 (N_14144,N_13987,N_13938);
xor U14145 (N_14145,N_13774,N_13872);
and U14146 (N_14146,N_13894,N_13785);
xnor U14147 (N_14147,N_13879,N_13892);
or U14148 (N_14148,N_13960,N_13862);
xor U14149 (N_14149,N_13842,N_13983);
or U14150 (N_14150,N_13954,N_13925);
or U14151 (N_14151,N_13790,N_13841);
and U14152 (N_14152,N_13922,N_13957);
and U14153 (N_14153,N_13958,N_13781);
or U14154 (N_14154,N_13917,N_13868);
and U14155 (N_14155,N_13776,N_13934);
nor U14156 (N_14156,N_13993,N_13800);
or U14157 (N_14157,N_13803,N_13804);
or U14158 (N_14158,N_13832,N_13753);
and U14159 (N_14159,N_13813,N_13796);
xnor U14160 (N_14160,N_13925,N_13886);
nor U14161 (N_14161,N_13929,N_13859);
and U14162 (N_14162,N_13853,N_13756);
xor U14163 (N_14163,N_13760,N_13802);
nand U14164 (N_14164,N_13806,N_13794);
or U14165 (N_14165,N_13995,N_13820);
and U14166 (N_14166,N_13815,N_13990);
nand U14167 (N_14167,N_13836,N_13763);
xnor U14168 (N_14168,N_13953,N_13803);
and U14169 (N_14169,N_13995,N_13885);
xor U14170 (N_14170,N_13931,N_13833);
and U14171 (N_14171,N_13847,N_13879);
nand U14172 (N_14172,N_13983,N_13900);
xor U14173 (N_14173,N_13833,N_13995);
xnor U14174 (N_14174,N_13905,N_13805);
xnor U14175 (N_14175,N_13910,N_13895);
xor U14176 (N_14176,N_13877,N_13897);
or U14177 (N_14177,N_13925,N_13867);
xor U14178 (N_14178,N_13983,N_13889);
nand U14179 (N_14179,N_13960,N_13859);
xor U14180 (N_14180,N_13947,N_13892);
nor U14181 (N_14181,N_13890,N_13974);
and U14182 (N_14182,N_13886,N_13809);
xor U14183 (N_14183,N_13886,N_13799);
or U14184 (N_14184,N_13775,N_13803);
nand U14185 (N_14185,N_13799,N_13884);
nand U14186 (N_14186,N_13960,N_13974);
nand U14187 (N_14187,N_13884,N_13854);
or U14188 (N_14188,N_13840,N_13803);
and U14189 (N_14189,N_13853,N_13812);
xor U14190 (N_14190,N_13938,N_13796);
xor U14191 (N_14191,N_13779,N_13896);
or U14192 (N_14192,N_13936,N_13864);
nand U14193 (N_14193,N_13913,N_13794);
nor U14194 (N_14194,N_13814,N_13868);
or U14195 (N_14195,N_13843,N_13750);
xor U14196 (N_14196,N_13772,N_13798);
nor U14197 (N_14197,N_13939,N_13774);
nor U14198 (N_14198,N_13909,N_13769);
nor U14199 (N_14199,N_13973,N_13968);
nand U14200 (N_14200,N_13907,N_13911);
and U14201 (N_14201,N_13956,N_13828);
xor U14202 (N_14202,N_13806,N_13770);
nor U14203 (N_14203,N_13835,N_13999);
nor U14204 (N_14204,N_13842,N_13893);
nand U14205 (N_14205,N_13969,N_13764);
nand U14206 (N_14206,N_13970,N_13822);
xnor U14207 (N_14207,N_13841,N_13856);
and U14208 (N_14208,N_13814,N_13946);
nor U14209 (N_14209,N_13983,N_13851);
or U14210 (N_14210,N_13957,N_13764);
nor U14211 (N_14211,N_13993,N_13994);
xor U14212 (N_14212,N_13983,N_13866);
nand U14213 (N_14213,N_13833,N_13792);
xnor U14214 (N_14214,N_13941,N_13766);
xnor U14215 (N_14215,N_13845,N_13999);
or U14216 (N_14216,N_13940,N_13965);
xor U14217 (N_14217,N_13789,N_13754);
nor U14218 (N_14218,N_13861,N_13800);
nand U14219 (N_14219,N_13838,N_13925);
and U14220 (N_14220,N_13803,N_13856);
or U14221 (N_14221,N_13972,N_13874);
xor U14222 (N_14222,N_13805,N_13950);
nor U14223 (N_14223,N_13811,N_13943);
xnor U14224 (N_14224,N_13790,N_13913);
nand U14225 (N_14225,N_13825,N_13863);
nor U14226 (N_14226,N_13902,N_13802);
nand U14227 (N_14227,N_13892,N_13838);
nor U14228 (N_14228,N_13782,N_13905);
nand U14229 (N_14229,N_13958,N_13914);
and U14230 (N_14230,N_13778,N_13874);
or U14231 (N_14231,N_13768,N_13932);
nand U14232 (N_14232,N_13902,N_13795);
nor U14233 (N_14233,N_13866,N_13763);
nor U14234 (N_14234,N_13791,N_13910);
nand U14235 (N_14235,N_13883,N_13926);
and U14236 (N_14236,N_13937,N_13794);
and U14237 (N_14237,N_13936,N_13999);
nand U14238 (N_14238,N_13979,N_13922);
nor U14239 (N_14239,N_13891,N_13992);
nor U14240 (N_14240,N_13806,N_13801);
and U14241 (N_14241,N_13772,N_13922);
and U14242 (N_14242,N_13810,N_13919);
nor U14243 (N_14243,N_13863,N_13993);
and U14244 (N_14244,N_13805,N_13948);
nor U14245 (N_14245,N_13879,N_13920);
nor U14246 (N_14246,N_13888,N_13958);
and U14247 (N_14247,N_13868,N_13807);
and U14248 (N_14248,N_13803,N_13870);
xor U14249 (N_14249,N_13827,N_13896);
nand U14250 (N_14250,N_14142,N_14134);
nand U14251 (N_14251,N_14021,N_14120);
or U14252 (N_14252,N_14136,N_14248);
or U14253 (N_14253,N_14217,N_14143);
nand U14254 (N_14254,N_14177,N_14215);
nor U14255 (N_14255,N_14137,N_14161);
nand U14256 (N_14256,N_14247,N_14230);
nor U14257 (N_14257,N_14125,N_14099);
and U14258 (N_14258,N_14117,N_14153);
nor U14259 (N_14259,N_14184,N_14123);
nand U14260 (N_14260,N_14237,N_14246);
nand U14261 (N_14261,N_14218,N_14027);
xnor U14262 (N_14262,N_14231,N_14007);
nor U14263 (N_14263,N_14204,N_14176);
nor U14264 (N_14264,N_14210,N_14188);
or U14265 (N_14265,N_14243,N_14050);
nor U14266 (N_14266,N_14135,N_14108);
or U14267 (N_14267,N_14180,N_14014);
nand U14268 (N_14268,N_14070,N_14115);
or U14269 (N_14269,N_14226,N_14138);
or U14270 (N_14270,N_14025,N_14061);
or U14271 (N_14271,N_14057,N_14082);
nand U14272 (N_14272,N_14102,N_14018);
and U14273 (N_14273,N_14078,N_14097);
nor U14274 (N_14274,N_14095,N_14200);
nand U14275 (N_14275,N_14132,N_14091);
xor U14276 (N_14276,N_14076,N_14022);
or U14277 (N_14277,N_14089,N_14009);
or U14278 (N_14278,N_14221,N_14029);
or U14279 (N_14279,N_14058,N_14175);
xor U14280 (N_14280,N_14150,N_14185);
nor U14281 (N_14281,N_14077,N_14220);
nand U14282 (N_14282,N_14186,N_14166);
xor U14283 (N_14283,N_14028,N_14212);
or U14284 (N_14284,N_14206,N_14229);
or U14285 (N_14285,N_14208,N_14074);
and U14286 (N_14286,N_14244,N_14182);
nor U14287 (N_14287,N_14201,N_14242);
xor U14288 (N_14288,N_14171,N_14181);
or U14289 (N_14289,N_14065,N_14158);
or U14290 (N_14290,N_14066,N_14084);
nor U14291 (N_14291,N_14227,N_14017);
and U14292 (N_14292,N_14056,N_14020);
or U14293 (N_14293,N_14036,N_14189);
nand U14294 (N_14294,N_14047,N_14122);
nand U14295 (N_14295,N_14163,N_14000);
xor U14296 (N_14296,N_14059,N_14178);
xnor U14297 (N_14297,N_14039,N_14087);
or U14298 (N_14298,N_14053,N_14196);
or U14299 (N_14299,N_14052,N_14241);
nand U14300 (N_14300,N_14010,N_14041);
or U14301 (N_14301,N_14006,N_14033);
and U14302 (N_14302,N_14239,N_14155);
or U14303 (N_14303,N_14249,N_14160);
or U14304 (N_14304,N_14035,N_14207);
nor U14305 (N_14305,N_14026,N_14044);
xor U14306 (N_14306,N_14075,N_14159);
nor U14307 (N_14307,N_14124,N_14148);
xnor U14308 (N_14308,N_14126,N_14034);
or U14309 (N_14309,N_14019,N_14024);
or U14310 (N_14310,N_14232,N_14104);
and U14311 (N_14311,N_14110,N_14173);
xor U14312 (N_14312,N_14112,N_14149);
and U14313 (N_14313,N_14079,N_14068);
and U14314 (N_14314,N_14168,N_14111);
nor U14315 (N_14315,N_14013,N_14245);
and U14316 (N_14316,N_14202,N_14015);
or U14317 (N_14317,N_14005,N_14129);
nand U14318 (N_14318,N_14085,N_14045);
or U14319 (N_14319,N_14170,N_14098);
xor U14320 (N_14320,N_14187,N_14071);
nand U14321 (N_14321,N_14154,N_14001);
nand U14322 (N_14322,N_14234,N_14139);
nor U14323 (N_14323,N_14004,N_14109);
and U14324 (N_14324,N_14203,N_14011);
and U14325 (N_14325,N_14198,N_14191);
or U14326 (N_14326,N_14146,N_14116);
xor U14327 (N_14327,N_14038,N_14127);
nor U14328 (N_14328,N_14179,N_14069);
or U14329 (N_14329,N_14133,N_14023);
nor U14330 (N_14330,N_14096,N_14048);
and U14331 (N_14331,N_14209,N_14062);
and U14332 (N_14332,N_14157,N_14063);
nand U14333 (N_14333,N_14167,N_14031);
nor U14334 (N_14334,N_14222,N_14238);
nand U14335 (N_14335,N_14080,N_14114);
nand U14336 (N_14336,N_14092,N_14088);
nand U14337 (N_14337,N_14030,N_14172);
and U14338 (N_14338,N_14037,N_14216);
xnor U14339 (N_14339,N_14223,N_14140);
nor U14340 (N_14340,N_14086,N_14032);
nor U14341 (N_14341,N_14118,N_14093);
xnor U14342 (N_14342,N_14016,N_14156);
and U14343 (N_14343,N_14240,N_14072);
nor U14344 (N_14344,N_14003,N_14054);
nand U14345 (N_14345,N_14183,N_14219);
or U14346 (N_14346,N_14169,N_14121);
nand U14347 (N_14347,N_14081,N_14049);
xnor U14348 (N_14348,N_14197,N_14012);
nand U14349 (N_14349,N_14214,N_14233);
nor U14350 (N_14350,N_14194,N_14046);
xnor U14351 (N_14351,N_14107,N_14235);
nand U14352 (N_14352,N_14147,N_14100);
and U14353 (N_14353,N_14103,N_14141);
and U14354 (N_14354,N_14174,N_14040);
or U14355 (N_14355,N_14060,N_14211);
or U14356 (N_14356,N_14144,N_14131);
nand U14357 (N_14357,N_14193,N_14083);
and U14358 (N_14358,N_14199,N_14090);
xnor U14359 (N_14359,N_14094,N_14165);
xnor U14360 (N_14360,N_14119,N_14067);
nor U14361 (N_14361,N_14073,N_14051);
xor U14362 (N_14362,N_14236,N_14225);
xnor U14363 (N_14363,N_14205,N_14130);
nand U14364 (N_14364,N_14113,N_14162);
nor U14365 (N_14365,N_14055,N_14164);
nor U14366 (N_14366,N_14002,N_14043);
nand U14367 (N_14367,N_14152,N_14101);
nand U14368 (N_14368,N_14195,N_14105);
or U14369 (N_14369,N_14228,N_14106);
xor U14370 (N_14370,N_14145,N_14042);
nand U14371 (N_14371,N_14151,N_14008);
xor U14372 (N_14372,N_14224,N_14064);
nor U14373 (N_14373,N_14213,N_14190);
xnor U14374 (N_14374,N_14128,N_14192);
or U14375 (N_14375,N_14024,N_14159);
nor U14376 (N_14376,N_14210,N_14043);
nor U14377 (N_14377,N_14190,N_14223);
and U14378 (N_14378,N_14030,N_14077);
and U14379 (N_14379,N_14084,N_14101);
nand U14380 (N_14380,N_14150,N_14146);
nand U14381 (N_14381,N_14059,N_14104);
or U14382 (N_14382,N_14134,N_14032);
nand U14383 (N_14383,N_14182,N_14170);
xor U14384 (N_14384,N_14202,N_14167);
and U14385 (N_14385,N_14181,N_14037);
nor U14386 (N_14386,N_14171,N_14108);
and U14387 (N_14387,N_14114,N_14125);
or U14388 (N_14388,N_14116,N_14063);
and U14389 (N_14389,N_14009,N_14095);
xnor U14390 (N_14390,N_14089,N_14149);
nand U14391 (N_14391,N_14034,N_14217);
or U14392 (N_14392,N_14036,N_14133);
nor U14393 (N_14393,N_14242,N_14175);
and U14394 (N_14394,N_14179,N_14158);
xor U14395 (N_14395,N_14247,N_14004);
nand U14396 (N_14396,N_14106,N_14184);
or U14397 (N_14397,N_14183,N_14064);
or U14398 (N_14398,N_14065,N_14095);
nor U14399 (N_14399,N_14136,N_14221);
nor U14400 (N_14400,N_14069,N_14229);
or U14401 (N_14401,N_14094,N_14174);
nand U14402 (N_14402,N_14007,N_14245);
nand U14403 (N_14403,N_14060,N_14202);
xor U14404 (N_14404,N_14217,N_14130);
nand U14405 (N_14405,N_14031,N_14137);
or U14406 (N_14406,N_14099,N_14102);
or U14407 (N_14407,N_14007,N_14111);
nand U14408 (N_14408,N_14214,N_14004);
and U14409 (N_14409,N_14074,N_14104);
xor U14410 (N_14410,N_14220,N_14119);
nand U14411 (N_14411,N_14017,N_14069);
nor U14412 (N_14412,N_14033,N_14119);
nor U14413 (N_14413,N_14186,N_14081);
nand U14414 (N_14414,N_14230,N_14154);
and U14415 (N_14415,N_14034,N_14101);
nand U14416 (N_14416,N_14117,N_14185);
nand U14417 (N_14417,N_14229,N_14160);
and U14418 (N_14418,N_14180,N_14187);
and U14419 (N_14419,N_14006,N_14241);
nor U14420 (N_14420,N_14128,N_14147);
xor U14421 (N_14421,N_14074,N_14112);
and U14422 (N_14422,N_14048,N_14132);
xor U14423 (N_14423,N_14248,N_14201);
nor U14424 (N_14424,N_14160,N_14094);
nand U14425 (N_14425,N_14041,N_14113);
nand U14426 (N_14426,N_14105,N_14247);
or U14427 (N_14427,N_14015,N_14100);
nor U14428 (N_14428,N_14158,N_14208);
xnor U14429 (N_14429,N_14119,N_14166);
nand U14430 (N_14430,N_14130,N_14166);
nand U14431 (N_14431,N_14103,N_14144);
xor U14432 (N_14432,N_14040,N_14034);
nor U14433 (N_14433,N_14129,N_14124);
or U14434 (N_14434,N_14017,N_14115);
nor U14435 (N_14435,N_14137,N_14111);
xor U14436 (N_14436,N_14200,N_14140);
nand U14437 (N_14437,N_14164,N_14231);
or U14438 (N_14438,N_14034,N_14182);
nor U14439 (N_14439,N_14062,N_14036);
xor U14440 (N_14440,N_14093,N_14059);
or U14441 (N_14441,N_14204,N_14227);
or U14442 (N_14442,N_14053,N_14037);
nor U14443 (N_14443,N_14213,N_14102);
nand U14444 (N_14444,N_14118,N_14182);
and U14445 (N_14445,N_14195,N_14217);
nor U14446 (N_14446,N_14082,N_14204);
xor U14447 (N_14447,N_14074,N_14099);
or U14448 (N_14448,N_14099,N_14088);
nor U14449 (N_14449,N_14018,N_14121);
or U14450 (N_14450,N_14046,N_14205);
nand U14451 (N_14451,N_14194,N_14215);
nor U14452 (N_14452,N_14232,N_14187);
nand U14453 (N_14453,N_14122,N_14173);
nand U14454 (N_14454,N_14050,N_14211);
nand U14455 (N_14455,N_14167,N_14044);
nand U14456 (N_14456,N_14114,N_14073);
nand U14457 (N_14457,N_14119,N_14233);
or U14458 (N_14458,N_14207,N_14160);
xnor U14459 (N_14459,N_14108,N_14207);
and U14460 (N_14460,N_14006,N_14169);
nand U14461 (N_14461,N_14028,N_14247);
nor U14462 (N_14462,N_14225,N_14071);
xnor U14463 (N_14463,N_14107,N_14110);
or U14464 (N_14464,N_14164,N_14026);
or U14465 (N_14465,N_14030,N_14188);
or U14466 (N_14466,N_14141,N_14152);
nand U14467 (N_14467,N_14013,N_14150);
or U14468 (N_14468,N_14236,N_14113);
or U14469 (N_14469,N_14004,N_14001);
or U14470 (N_14470,N_14194,N_14055);
or U14471 (N_14471,N_14240,N_14063);
nor U14472 (N_14472,N_14170,N_14152);
and U14473 (N_14473,N_14163,N_14135);
nor U14474 (N_14474,N_14079,N_14003);
or U14475 (N_14475,N_14044,N_14095);
nor U14476 (N_14476,N_14014,N_14091);
nor U14477 (N_14477,N_14043,N_14006);
nand U14478 (N_14478,N_14188,N_14234);
xnor U14479 (N_14479,N_14024,N_14028);
nor U14480 (N_14480,N_14171,N_14236);
nand U14481 (N_14481,N_14108,N_14018);
nor U14482 (N_14482,N_14144,N_14002);
and U14483 (N_14483,N_14135,N_14242);
and U14484 (N_14484,N_14246,N_14124);
nand U14485 (N_14485,N_14192,N_14111);
or U14486 (N_14486,N_14163,N_14073);
nand U14487 (N_14487,N_14245,N_14021);
nand U14488 (N_14488,N_14132,N_14078);
and U14489 (N_14489,N_14172,N_14234);
or U14490 (N_14490,N_14176,N_14149);
nand U14491 (N_14491,N_14100,N_14029);
xnor U14492 (N_14492,N_14204,N_14123);
and U14493 (N_14493,N_14247,N_14033);
or U14494 (N_14494,N_14153,N_14047);
nor U14495 (N_14495,N_14035,N_14149);
or U14496 (N_14496,N_14022,N_14105);
xor U14497 (N_14497,N_14063,N_14096);
nor U14498 (N_14498,N_14016,N_14087);
and U14499 (N_14499,N_14043,N_14172);
xnor U14500 (N_14500,N_14327,N_14424);
nand U14501 (N_14501,N_14454,N_14464);
and U14502 (N_14502,N_14340,N_14477);
xnor U14503 (N_14503,N_14484,N_14402);
nand U14504 (N_14504,N_14453,N_14400);
or U14505 (N_14505,N_14342,N_14421);
nand U14506 (N_14506,N_14428,N_14472);
nand U14507 (N_14507,N_14352,N_14299);
nand U14508 (N_14508,N_14333,N_14292);
or U14509 (N_14509,N_14480,N_14481);
and U14510 (N_14510,N_14398,N_14304);
and U14511 (N_14511,N_14335,N_14356);
nand U14512 (N_14512,N_14431,N_14281);
xnor U14513 (N_14513,N_14300,N_14377);
or U14514 (N_14514,N_14358,N_14283);
and U14515 (N_14515,N_14364,N_14257);
nand U14516 (N_14516,N_14478,N_14267);
nand U14517 (N_14517,N_14379,N_14265);
or U14518 (N_14518,N_14380,N_14361);
nand U14519 (N_14519,N_14291,N_14282);
xor U14520 (N_14520,N_14371,N_14355);
and U14521 (N_14521,N_14451,N_14486);
or U14522 (N_14522,N_14445,N_14331);
xnor U14523 (N_14523,N_14313,N_14404);
and U14524 (N_14524,N_14423,N_14301);
and U14525 (N_14525,N_14479,N_14251);
or U14526 (N_14526,N_14418,N_14348);
xor U14527 (N_14527,N_14397,N_14288);
nor U14528 (N_14528,N_14466,N_14334);
and U14529 (N_14529,N_14269,N_14250);
nor U14530 (N_14530,N_14337,N_14420);
nor U14531 (N_14531,N_14272,N_14280);
nand U14532 (N_14532,N_14483,N_14277);
nor U14533 (N_14533,N_14318,N_14261);
xor U14534 (N_14534,N_14349,N_14383);
nor U14535 (N_14535,N_14344,N_14363);
and U14536 (N_14536,N_14490,N_14390);
xor U14537 (N_14537,N_14471,N_14290);
nor U14538 (N_14538,N_14434,N_14307);
nand U14539 (N_14539,N_14436,N_14403);
xnor U14540 (N_14540,N_14416,N_14297);
nor U14541 (N_14541,N_14323,N_14298);
and U14542 (N_14542,N_14316,N_14387);
and U14543 (N_14543,N_14394,N_14305);
nand U14544 (N_14544,N_14378,N_14275);
or U14545 (N_14545,N_14346,N_14467);
or U14546 (N_14546,N_14293,N_14422);
xnor U14547 (N_14547,N_14351,N_14432);
xnor U14548 (N_14548,N_14336,N_14311);
nor U14549 (N_14549,N_14399,N_14449);
nor U14550 (N_14550,N_14463,N_14494);
nor U14551 (N_14551,N_14252,N_14369);
or U14552 (N_14552,N_14274,N_14462);
nand U14553 (N_14553,N_14469,N_14262);
xnor U14554 (N_14554,N_14286,N_14381);
xnor U14555 (N_14555,N_14401,N_14429);
or U14556 (N_14556,N_14408,N_14295);
or U14557 (N_14557,N_14446,N_14360);
nand U14558 (N_14558,N_14433,N_14461);
nor U14559 (N_14559,N_14350,N_14465);
nor U14560 (N_14560,N_14302,N_14441);
nor U14561 (N_14561,N_14343,N_14444);
nor U14562 (N_14562,N_14310,N_14296);
or U14563 (N_14563,N_14263,N_14285);
nor U14564 (N_14564,N_14289,N_14317);
and U14565 (N_14565,N_14332,N_14443);
nor U14566 (N_14566,N_14357,N_14492);
or U14567 (N_14567,N_14457,N_14417);
nor U14568 (N_14568,N_14468,N_14459);
nor U14569 (N_14569,N_14324,N_14495);
or U14570 (N_14570,N_14329,N_14393);
or U14571 (N_14571,N_14406,N_14448);
xor U14572 (N_14572,N_14386,N_14435);
nor U14573 (N_14573,N_14496,N_14359);
or U14574 (N_14574,N_14354,N_14419);
nor U14575 (N_14575,N_14396,N_14376);
nand U14576 (N_14576,N_14470,N_14312);
or U14577 (N_14577,N_14372,N_14455);
nor U14578 (N_14578,N_14430,N_14279);
nand U14579 (N_14579,N_14266,N_14338);
nand U14580 (N_14580,N_14414,N_14411);
xnor U14581 (N_14581,N_14440,N_14498);
and U14582 (N_14582,N_14270,N_14384);
or U14583 (N_14583,N_14388,N_14491);
nor U14584 (N_14584,N_14320,N_14341);
nor U14585 (N_14585,N_14438,N_14370);
or U14586 (N_14586,N_14409,N_14294);
nand U14587 (N_14587,N_14273,N_14450);
xnor U14588 (N_14588,N_14322,N_14460);
and U14589 (N_14589,N_14405,N_14258);
nand U14590 (N_14590,N_14278,N_14452);
xnor U14591 (N_14591,N_14382,N_14412);
xor U14592 (N_14592,N_14328,N_14407);
or U14593 (N_14593,N_14447,N_14395);
xnor U14594 (N_14594,N_14489,N_14306);
and U14595 (N_14595,N_14437,N_14315);
nand U14596 (N_14596,N_14497,N_14392);
or U14597 (N_14597,N_14439,N_14391);
or U14598 (N_14598,N_14389,N_14345);
nand U14599 (N_14599,N_14314,N_14365);
and U14600 (N_14600,N_14259,N_14385);
xnor U14601 (N_14601,N_14366,N_14326);
xor U14602 (N_14602,N_14442,N_14271);
nor U14603 (N_14603,N_14264,N_14260);
nor U14604 (N_14604,N_14287,N_14488);
nand U14605 (N_14605,N_14308,N_14373);
and U14606 (N_14606,N_14493,N_14415);
nor U14607 (N_14607,N_14368,N_14476);
or U14608 (N_14608,N_14253,N_14319);
or U14609 (N_14609,N_14276,N_14475);
nand U14610 (N_14610,N_14303,N_14410);
and U14611 (N_14611,N_14413,N_14309);
and U14612 (N_14612,N_14367,N_14485);
nand U14613 (N_14613,N_14330,N_14321);
nor U14614 (N_14614,N_14254,N_14482);
nor U14615 (N_14615,N_14347,N_14375);
or U14616 (N_14616,N_14458,N_14474);
or U14617 (N_14617,N_14325,N_14284);
nand U14618 (N_14618,N_14256,N_14255);
nand U14619 (N_14619,N_14426,N_14353);
or U14620 (N_14620,N_14456,N_14374);
or U14621 (N_14621,N_14487,N_14425);
nand U14622 (N_14622,N_14339,N_14499);
or U14623 (N_14623,N_14268,N_14362);
and U14624 (N_14624,N_14473,N_14427);
nor U14625 (N_14625,N_14484,N_14426);
and U14626 (N_14626,N_14432,N_14423);
and U14627 (N_14627,N_14376,N_14489);
or U14628 (N_14628,N_14464,N_14266);
xor U14629 (N_14629,N_14391,N_14462);
and U14630 (N_14630,N_14415,N_14405);
xor U14631 (N_14631,N_14323,N_14358);
xor U14632 (N_14632,N_14495,N_14419);
nor U14633 (N_14633,N_14255,N_14449);
xor U14634 (N_14634,N_14293,N_14297);
nor U14635 (N_14635,N_14450,N_14417);
or U14636 (N_14636,N_14304,N_14477);
xor U14637 (N_14637,N_14337,N_14489);
nor U14638 (N_14638,N_14321,N_14267);
or U14639 (N_14639,N_14311,N_14260);
xnor U14640 (N_14640,N_14442,N_14417);
or U14641 (N_14641,N_14322,N_14339);
or U14642 (N_14642,N_14485,N_14495);
or U14643 (N_14643,N_14459,N_14414);
or U14644 (N_14644,N_14439,N_14456);
or U14645 (N_14645,N_14277,N_14359);
and U14646 (N_14646,N_14335,N_14334);
xnor U14647 (N_14647,N_14416,N_14360);
xnor U14648 (N_14648,N_14426,N_14436);
xnor U14649 (N_14649,N_14372,N_14382);
nand U14650 (N_14650,N_14260,N_14288);
or U14651 (N_14651,N_14412,N_14361);
nor U14652 (N_14652,N_14399,N_14287);
nor U14653 (N_14653,N_14492,N_14317);
xor U14654 (N_14654,N_14278,N_14294);
xor U14655 (N_14655,N_14286,N_14434);
xnor U14656 (N_14656,N_14411,N_14383);
and U14657 (N_14657,N_14408,N_14327);
and U14658 (N_14658,N_14438,N_14442);
or U14659 (N_14659,N_14251,N_14345);
nand U14660 (N_14660,N_14265,N_14366);
or U14661 (N_14661,N_14347,N_14443);
xor U14662 (N_14662,N_14274,N_14498);
xor U14663 (N_14663,N_14498,N_14305);
or U14664 (N_14664,N_14255,N_14335);
nand U14665 (N_14665,N_14357,N_14298);
xnor U14666 (N_14666,N_14354,N_14379);
nor U14667 (N_14667,N_14306,N_14421);
xor U14668 (N_14668,N_14442,N_14327);
nand U14669 (N_14669,N_14347,N_14447);
or U14670 (N_14670,N_14287,N_14483);
or U14671 (N_14671,N_14322,N_14408);
and U14672 (N_14672,N_14259,N_14265);
or U14673 (N_14673,N_14365,N_14384);
nand U14674 (N_14674,N_14411,N_14300);
nand U14675 (N_14675,N_14343,N_14488);
xor U14676 (N_14676,N_14453,N_14473);
or U14677 (N_14677,N_14472,N_14315);
xor U14678 (N_14678,N_14466,N_14450);
nand U14679 (N_14679,N_14289,N_14381);
xor U14680 (N_14680,N_14317,N_14462);
nand U14681 (N_14681,N_14433,N_14281);
nand U14682 (N_14682,N_14453,N_14299);
and U14683 (N_14683,N_14475,N_14414);
nor U14684 (N_14684,N_14482,N_14285);
and U14685 (N_14685,N_14263,N_14409);
xnor U14686 (N_14686,N_14414,N_14336);
xnor U14687 (N_14687,N_14455,N_14486);
xor U14688 (N_14688,N_14269,N_14437);
xnor U14689 (N_14689,N_14389,N_14316);
or U14690 (N_14690,N_14451,N_14417);
and U14691 (N_14691,N_14315,N_14390);
xnor U14692 (N_14692,N_14314,N_14418);
nand U14693 (N_14693,N_14429,N_14442);
nor U14694 (N_14694,N_14485,N_14274);
and U14695 (N_14695,N_14251,N_14419);
nand U14696 (N_14696,N_14471,N_14278);
and U14697 (N_14697,N_14387,N_14334);
xnor U14698 (N_14698,N_14323,N_14338);
and U14699 (N_14699,N_14292,N_14400);
or U14700 (N_14700,N_14465,N_14361);
nand U14701 (N_14701,N_14462,N_14461);
nand U14702 (N_14702,N_14291,N_14439);
xnor U14703 (N_14703,N_14403,N_14405);
xnor U14704 (N_14704,N_14361,N_14331);
xnor U14705 (N_14705,N_14369,N_14452);
nor U14706 (N_14706,N_14379,N_14374);
or U14707 (N_14707,N_14256,N_14405);
nand U14708 (N_14708,N_14378,N_14293);
or U14709 (N_14709,N_14488,N_14336);
nor U14710 (N_14710,N_14298,N_14480);
or U14711 (N_14711,N_14390,N_14368);
xor U14712 (N_14712,N_14436,N_14369);
nor U14713 (N_14713,N_14298,N_14327);
nand U14714 (N_14714,N_14295,N_14470);
nand U14715 (N_14715,N_14413,N_14486);
or U14716 (N_14716,N_14416,N_14400);
nor U14717 (N_14717,N_14274,N_14469);
and U14718 (N_14718,N_14467,N_14446);
nor U14719 (N_14719,N_14359,N_14442);
xnor U14720 (N_14720,N_14304,N_14469);
or U14721 (N_14721,N_14445,N_14473);
and U14722 (N_14722,N_14413,N_14333);
and U14723 (N_14723,N_14315,N_14319);
and U14724 (N_14724,N_14263,N_14326);
or U14725 (N_14725,N_14355,N_14360);
nor U14726 (N_14726,N_14277,N_14347);
or U14727 (N_14727,N_14265,N_14457);
nor U14728 (N_14728,N_14299,N_14260);
or U14729 (N_14729,N_14320,N_14359);
or U14730 (N_14730,N_14499,N_14304);
xor U14731 (N_14731,N_14316,N_14325);
and U14732 (N_14732,N_14477,N_14486);
and U14733 (N_14733,N_14421,N_14388);
nor U14734 (N_14734,N_14473,N_14483);
or U14735 (N_14735,N_14418,N_14440);
xnor U14736 (N_14736,N_14361,N_14492);
nor U14737 (N_14737,N_14276,N_14479);
and U14738 (N_14738,N_14381,N_14299);
nor U14739 (N_14739,N_14385,N_14340);
nand U14740 (N_14740,N_14390,N_14310);
nand U14741 (N_14741,N_14471,N_14266);
xnor U14742 (N_14742,N_14455,N_14271);
xor U14743 (N_14743,N_14490,N_14275);
or U14744 (N_14744,N_14381,N_14482);
or U14745 (N_14745,N_14316,N_14408);
nor U14746 (N_14746,N_14339,N_14389);
nand U14747 (N_14747,N_14493,N_14251);
or U14748 (N_14748,N_14261,N_14298);
nor U14749 (N_14749,N_14269,N_14468);
nand U14750 (N_14750,N_14621,N_14636);
and U14751 (N_14751,N_14554,N_14715);
and U14752 (N_14752,N_14524,N_14687);
and U14753 (N_14753,N_14637,N_14586);
or U14754 (N_14754,N_14702,N_14571);
xnor U14755 (N_14755,N_14657,N_14596);
xor U14756 (N_14756,N_14622,N_14726);
or U14757 (N_14757,N_14503,N_14609);
xnor U14758 (N_14758,N_14602,N_14658);
or U14759 (N_14759,N_14717,N_14635);
and U14760 (N_14760,N_14588,N_14545);
or U14761 (N_14761,N_14612,N_14703);
and U14762 (N_14762,N_14732,N_14599);
xnor U14763 (N_14763,N_14564,N_14600);
nor U14764 (N_14764,N_14616,N_14679);
and U14765 (N_14765,N_14525,N_14744);
and U14766 (N_14766,N_14513,N_14649);
xnor U14767 (N_14767,N_14573,N_14695);
and U14768 (N_14768,N_14688,N_14631);
nor U14769 (N_14769,N_14537,N_14562);
or U14770 (N_14770,N_14730,N_14652);
nand U14771 (N_14771,N_14686,N_14561);
xor U14772 (N_14772,N_14729,N_14711);
nor U14773 (N_14773,N_14639,N_14601);
nand U14774 (N_14774,N_14510,N_14713);
and U14775 (N_14775,N_14748,N_14556);
nand U14776 (N_14776,N_14705,N_14589);
nand U14777 (N_14777,N_14745,N_14535);
or U14778 (N_14778,N_14625,N_14617);
nor U14779 (N_14779,N_14663,N_14646);
and U14780 (N_14780,N_14552,N_14570);
or U14781 (N_14781,N_14704,N_14664);
and U14782 (N_14782,N_14644,N_14615);
or U14783 (N_14783,N_14712,N_14611);
nor U14784 (N_14784,N_14632,N_14605);
and U14785 (N_14785,N_14551,N_14707);
or U14786 (N_14786,N_14590,N_14643);
xor U14787 (N_14787,N_14743,N_14576);
or U14788 (N_14788,N_14579,N_14574);
nand U14789 (N_14789,N_14697,N_14529);
xnor U14790 (N_14790,N_14553,N_14502);
and U14791 (N_14791,N_14698,N_14547);
nand U14792 (N_14792,N_14647,N_14549);
and U14793 (N_14793,N_14534,N_14683);
nand U14794 (N_14794,N_14651,N_14634);
xnor U14795 (N_14795,N_14685,N_14624);
xnor U14796 (N_14796,N_14681,N_14735);
nand U14797 (N_14797,N_14608,N_14520);
nor U14798 (N_14798,N_14515,N_14559);
or U14799 (N_14799,N_14580,N_14640);
xnor U14800 (N_14800,N_14566,N_14665);
xor U14801 (N_14801,N_14655,N_14747);
xor U14802 (N_14802,N_14613,N_14544);
xor U14803 (N_14803,N_14509,N_14699);
nand U14804 (N_14804,N_14741,N_14678);
xnor U14805 (N_14805,N_14514,N_14528);
nand U14806 (N_14806,N_14505,N_14530);
nor U14807 (N_14807,N_14680,N_14533);
nand U14808 (N_14808,N_14626,N_14749);
nor U14809 (N_14809,N_14565,N_14746);
nor U14810 (N_14810,N_14662,N_14583);
and U14811 (N_14811,N_14512,N_14569);
nor U14812 (N_14812,N_14708,N_14740);
nor U14813 (N_14813,N_14661,N_14560);
nor U14814 (N_14814,N_14592,N_14610);
xor U14815 (N_14815,N_14674,N_14511);
and U14816 (N_14816,N_14519,N_14557);
or U14817 (N_14817,N_14618,N_14669);
nor U14818 (N_14818,N_14736,N_14696);
or U14819 (N_14819,N_14721,N_14693);
nor U14820 (N_14820,N_14656,N_14734);
nor U14821 (N_14821,N_14603,N_14676);
or U14822 (N_14822,N_14720,N_14706);
or U14823 (N_14823,N_14714,N_14595);
nand U14824 (N_14824,N_14710,N_14733);
nand U14825 (N_14825,N_14543,N_14725);
nand U14826 (N_14826,N_14587,N_14585);
or U14827 (N_14827,N_14629,N_14539);
nor U14828 (N_14828,N_14682,N_14538);
xor U14829 (N_14829,N_14563,N_14568);
or U14830 (N_14830,N_14653,N_14659);
nor U14831 (N_14831,N_14517,N_14728);
xor U14832 (N_14832,N_14521,N_14722);
nor U14833 (N_14833,N_14550,N_14555);
and U14834 (N_14834,N_14623,N_14516);
or U14835 (N_14835,N_14532,N_14670);
nor U14836 (N_14836,N_14597,N_14719);
and U14837 (N_14837,N_14591,N_14723);
xor U14838 (N_14838,N_14654,N_14642);
and U14839 (N_14839,N_14598,N_14526);
nor U14840 (N_14840,N_14593,N_14645);
nand U14841 (N_14841,N_14508,N_14718);
and U14842 (N_14842,N_14667,N_14518);
nand U14843 (N_14843,N_14506,N_14541);
nor U14844 (N_14844,N_14650,N_14738);
nand U14845 (N_14845,N_14501,N_14572);
nor U14846 (N_14846,N_14523,N_14677);
and U14847 (N_14847,N_14700,N_14507);
or U14848 (N_14848,N_14727,N_14668);
nand U14849 (N_14849,N_14522,N_14641);
nand U14850 (N_14850,N_14716,N_14731);
nor U14851 (N_14851,N_14673,N_14578);
nand U14852 (N_14852,N_14604,N_14607);
and U14853 (N_14853,N_14504,N_14739);
and U14854 (N_14854,N_14582,N_14584);
xnor U14855 (N_14855,N_14575,N_14660);
nand U14856 (N_14856,N_14689,N_14527);
and U14857 (N_14857,N_14633,N_14724);
and U14858 (N_14858,N_14671,N_14531);
and U14859 (N_14859,N_14675,N_14548);
xor U14860 (N_14860,N_14691,N_14536);
xor U14861 (N_14861,N_14648,N_14694);
xor U14862 (N_14862,N_14692,N_14684);
or U14863 (N_14863,N_14619,N_14709);
or U14864 (N_14864,N_14594,N_14628);
xnor U14865 (N_14865,N_14558,N_14742);
nand U14866 (N_14866,N_14638,N_14606);
and U14867 (N_14867,N_14567,N_14500);
and U14868 (N_14868,N_14690,N_14627);
nor U14869 (N_14869,N_14546,N_14614);
or U14870 (N_14870,N_14672,N_14581);
and U14871 (N_14871,N_14620,N_14701);
or U14872 (N_14872,N_14737,N_14542);
nand U14873 (N_14873,N_14666,N_14577);
and U14874 (N_14874,N_14540,N_14630);
and U14875 (N_14875,N_14707,N_14676);
and U14876 (N_14876,N_14685,N_14692);
or U14877 (N_14877,N_14686,N_14535);
nor U14878 (N_14878,N_14705,N_14577);
nand U14879 (N_14879,N_14562,N_14524);
or U14880 (N_14880,N_14563,N_14516);
xnor U14881 (N_14881,N_14660,N_14730);
xor U14882 (N_14882,N_14661,N_14558);
or U14883 (N_14883,N_14653,N_14540);
or U14884 (N_14884,N_14693,N_14618);
and U14885 (N_14885,N_14645,N_14554);
xnor U14886 (N_14886,N_14616,N_14654);
or U14887 (N_14887,N_14718,N_14523);
and U14888 (N_14888,N_14516,N_14698);
xnor U14889 (N_14889,N_14541,N_14720);
xor U14890 (N_14890,N_14507,N_14560);
nor U14891 (N_14891,N_14675,N_14608);
nand U14892 (N_14892,N_14617,N_14686);
and U14893 (N_14893,N_14702,N_14585);
or U14894 (N_14894,N_14562,N_14744);
nand U14895 (N_14895,N_14646,N_14657);
nor U14896 (N_14896,N_14736,N_14744);
and U14897 (N_14897,N_14610,N_14736);
and U14898 (N_14898,N_14662,N_14746);
nand U14899 (N_14899,N_14550,N_14586);
or U14900 (N_14900,N_14516,N_14699);
or U14901 (N_14901,N_14598,N_14694);
xor U14902 (N_14902,N_14500,N_14635);
xor U14903 (N_14903,N_14742,N_14633);
nand U14904 (N_14904,N_14548,N_14732);
and U14905 (N_14905,N_14606,N_14727);
nand U14906 (N_14906,N_14615,N_14613);
nand U14907 (N_14907,N_14639,N_14544);
nor U14908 (N_14908,N_14593,N_14710);
or U14909 (N_14909,N_14693,N_14565);
nand U14910 (N_14910,N_14698,N_14651);
or U14911 (N_14911,N_14727,N_14725);
and U14912 (N_14912,N_14565,N_14712);
nor U14913 (N_14913,N_14552,N_14636);
xnor U14914 (N_14914,N_14644,N_14633);
xnor U14915 (N_14915,N_14629,N_14531);
nor U14916 (N_14916,N_14664,N_14502);
or U14917 (N_14917,N_14715,N_14743);
or U14918 (N_14918,N_14566,N_14524);
xor U14919 (N_14919,N_14669,N_14580);
nor U14920 (N_14920,N_14577,N_14560);
nand U14921 (N_14921,N_14695,N_14729);
xnor U14922 (N_14922,N_14674,N_14551);
or U14923 (N_14923,N_14639,N_14736);
or U14924 (N_14924,N_14597,N_14734);
nor U14925 (N_14925,N_14677,N_14747);
nor U14926 (N_14926,N_14506,N_14522);
nor U14927 (N_14927,N_14700,N_14734);
and U14928 (N_14928,N_14688,N_14712);
and U14929 (N_14929,N_14596,N_14665);
nand U14930 (N_14930,N_14698,N_14505);
and U14931 (N_14931,N_14704,N_14500);
or U14932 (N_14932,N_14546,N_14740);
xnor U14933 (N_14933,N_14527,N_14575);
and U14934 (N_14934,N_14503,N_14533);
nand U14935 (N_14935,N_14634,N_14509);
and U14936 (N_14936,N_14578,N_14614);
xnor U14937 (N_14937,N_14652,N_14604);
nor U14938 (N_14938,N_14502,N_14717);
and U14939 (N_14939,N_14653,N_14647);
nand U14940 (N_14940,N_14532,N_14538);
xor U14941 (N_14941,N_14623,N_14645);
nor U14942 (N_14942,N_14597,N_14569);
or U14943 (N_14943,N_14696,N_14612);
and U14944 (N_14944,N_14677,N_14695);
nor U14945 (N_14945,N_14729,N_14657);
nand U14946 (N_14946,N_14638,N_14619);
nand U14947 (N_14947,N_14704,N_14734);
xnor U14948 (N_14948,N_14694,N_14640);
and U14949 (N_14949,N_14645,N_14565);
xnor U14950 (N_14950,N_14668,N_14580);
nand U14951 (N_14951,N_14675,N_14727);
xnor U14952 (N_14952,N_14627,N_14726);
xor U14953 (N_14953,N_14522,N_14532);
nor U14954 (N_14954,N_14715,N_14623);
xor U14955 (N_14955,N_14661,N_14656);
and U14956 (N_14956,N_14556,N_14600);
nor U14957 (N_14957,N_14544,N_14568);
and U14958 (N_14958,N_14714,N_14597);
xnor U14959 (N_14959,N_14632,N_14637);
xnor U14960 (N_14960,N_14581,N_14619);
nor U14961 (N_14961,N_14525,N_14725);
xnor U14962 (N_14962,N_14504,N_14590);
nand U14963 (N_14963,N_14520,N_14721);
and U14964 (N_14964,N_14527,N_14520);
or U14965 (N_14965,N_14612,N_14583);
nand U14966 (N_14966,N_14508,N_14529);
xnor U14967 (N_14967,N_14716,N_14650);
xnor U14968 (N_14968,N_14696,N_14627);
and U14969 (N_14969,N_14720,N_14546);
or U14970 (N_14970,N_14528,N_14705);
and U14971 (N_14971,N_14697,N_14634);
xnor U14972 (N_14972,N_14603,N_14543);
and U14973 (N_14973,N_14558,N_14543);
and U14974 (N_14974,N_14714,N_14600);
or U14975 (N_14975,N_14646,N_14572);
nor U14976 (N_14976,N_14587,N_14543);
nand U14977 (N_14977,N_14684,N_14677);
and U14978 (N_14978,N_14524,N_14676);
and U14979 (N_14979,N_14572,N_14689);
nand U14980 (N_14980,N_14703,N_14724);
or U14981 (N_14981,N_14547,N_14588);
nor U14982 (N_14982,N_14570,N_14624);
nor U14983 (N_14983,N_14736,N_14508);
and U14984 (N_14984,N_14742,N_14578);
and U14985 (N_14985,N_14730,N_14654);
and U14986 (N_14986,N_14613,N_14744);
or U14987 (N_14987,N_14685,N_14706);
and U14988 (N_14988,N_14594,N_14688);
xor U14989 (N_14989,N_14562,N_14543);
xor U14990 (N_14990,N_14664,N_14535);
and U14991 (N_14991,N_14549,N_14528);
xnor U14992 (N_14992,N_14534,N_14738);
nand U14993 (N_14993,N_14694,N_14602);
nand U14994 (N_14994,N_14705,N_14616);
nor U14995 (N_14995,N_14606,N_14683);
nor U14996 (N_14996,N_14584,N_14699);
nand U14997 (N_14997,N_14616,N_14661);
and U14998 (N_14998,N_14543,N_14685);
and U14999 (N_14999,N_14572,N_14567);
nand U15000 (N_15000,N_14934,N_14916);
nor U15001 (N_15001,N_14824,N_14911);
or U15002 (N_15002,N_14986,N_14878);
nor U15003 (N_15003,N_14872,N_14964);
nand U15004 (N_15004,N_14929,N_14790);
xor U15005 (N_15005,N_14910,N_14975);
nor U15006 (N_15006,N_14927,N_14861);
or U15007 (N_15007,N_14832,N_14945);
nor U15008 (N_15008,N_14864,N_14999);
nand U15009 (N_15009,N_14923,N_14865);
and U15010 (N_15010,N_14845,N_14785);
nand U15011 (N_15011,N_14781,N_14802);
nor U15012 (N_15012,N_14848,N_14826);
or U15013 (N_15013,N_14919,N_14853);
or U15014 (N_15014,N_14901,N_14813);
or U15015 (N_15015,N_14834,N_14961);
nand U15016 (N_15016,N_14993,N_14833);
or U15017 (N_15017,N_14760,N_14970);
nor U15018 (N_15018,N_14963,N_14799);
and U15019 (N_15019,N_14909,N_14974);
xor U15020 (N_15020,N_14792,N_14873);
nor U15021 (N_15021,N_14756,N_14943);
nand U15022 (N_15022,N_14948,N_14795);
nor U15023 (N_15023,N_14844,N_14763);
and U15024 (N_15024,N_14958,N_14817);
nand U15025 (N_15025,N_14761,N_14820);
xor U15026 (N_15026,N_14891,N_14973);
nor U15027 (N_15027,N_14828,N_14941);
or U15028 (N_15028,N_14764,N_14808);
nand U15029 (N_15029,N_14827,N_14972);
nor U15030 (N_15030,N_14996,N_14947);
and U15031 (N_15031,N_14871,N_14825);
nor U15032 (N_15032,N_14855,N_14841);
nand U15033 (N_15033,N_14881,N_14937);
or U15034 (N_15034,N_14750,N_14954);
nor U15035 (N_15035,N_14959,N_14866);
and U15036 (N_15036,N_14857,N_14976);
nand U15037 (N_15037,N_14752,N_14770);
and U15038 (N_15038,N_14779,N_14774);
xnor U15039 (N_15039,N_14821,N_14899);
xnor U15040 (N_15040,N_14846,N_14907);
or U15041 (N_15041,N_14940,N_14896);
or U15042 (N_15042,N_14843,N_14982);
and U15043 (N_15043,N_14854,N_14860);
or U15044 (N_15044,N_14862,N_14997);
and U15045 (N_15045,N_14879,N_14884);
nand U15046 (N_15046,N_14776,N_14762);
and U15047 (N_15047,N_14890,N_14849);
and U15048 (N_15048,N_14998,N_14882);
nand U15049 (N_15049,N_14992,N_14912);
or U15050 (N_15050,N_14939,N_14793);
nand U15051 (N_15051,N_14930,N_14874);
xnor U15052 (N_15052,N_14782,N_14960);
or U15053 (N_15053,N_14903,N_14822);
or U15054 (N_15054,N_14801,N_14967);
xnor U15055 (N_15055,N_14783,N_14755);
and U15056 (N_15056,N_14900,N_14758);
nand U15057 (N_15057,N_14778,N_14754);
nand U15058 (N_15058,N_14794,N_14914);
xnor U15059 (N_15059,N_14966,N_14991);
nor U15060 (N_15060,N_14815,N_14938);
or U15061 (N_15061,N_14810,N_14892);
and U15062 (N_15062,N_14955,N_14788);
xor U15063 (N_15063,N_14906,N_14765);
nor U15064 (N_15064,N_14935,N_14859);
and U15065 (N_15065,N_14831,N_14789);
and U15066 (N_15066,N_14842,N_14894);
nor U15067 (N_15067,N_14918,N_14889);
nand U15068 (N_15068,N_14771,N_14800);
nor U15069 (N_15069,N_14951,N_14987);
nand U15070 (N_15070,N_14913,N_14944);
or U15071 (N_15071,N_14766,N_14805);
or U15072 (N_15072,N_14759,N_14753);
nor U15073 (N_15073,N_14921,N_14971);
nand U15074 (N_15074,N_14988,N_14983);
nor U15075 (N_15075,N_14990,N_14953);
nor U15076 (N_15076,N_14751,N_14819);
xnor U15077 (N_15077,N_14870,N_14980);
nor U15078 (N_15078,N_14984,N_14995);
xnor U15079 (N_15079,N_14769,N_14847);
xnor U15080 (N_15080,N_14979,N_14804);
nand U15081 (N_15081,N_14823,N_14933);
or U15082 (N_15082,N_14829,N_14768);
and U15083 (N_15083,N_14787,N_14786);
and U15084 (N_15084,N_14887,N_14968);
nand U15085 (N_15085,N_14920,N_14888);
and U15086 (N_15086,N_14868,N_14839);
and U15087 (N_15087,N_14856,N_14956);
nand U15088 (N_15088,N_14917,N_14893);
nor U15089 (N_15089,N_14780,N_14798);
nand U15090 (N_15090,N_14994,N_14812);
nor U15091 (N_15091,N_14978,N_14818);
or U15092 (N_15092,N_14942,N_14952);
xor U15093 (N_15093,N_14876,N_14809);
or U15094 (N_15094,N_14925,N_14869);
xnor U15095 (N_15095,N_14965,N_14904);
and U15096 (N_15096,N_14877,N_14924);
nor U15097 (N_15097,N_14796,N_14928);
nand U15098 (N_15098,N_14836,N_14757);
xnor U15099 (N_15099,N_14977,N_14807);
nor U15100 (N_15100,N_14905,N_14867);
or U15101 (N_15101,N_14897,N_14806);
or U15102 (N_15102,N_14858,N_14772);
and U15103 (N_15103,N_14915,N_14931);
nand U15104 (N_15104,N_14773,N_14850);
nand U15105 (N_15105,N_14830,N_14803);
nor U15106 (N_15106,N_14814,N_14898);
nand U15107 (N_15107,N_14949,N_14885);
or U15108 (N_15108,N_14775,N_14946);
nand U15109 (N_15109,N_14835,N_14989);
nand U15110 (N_15110,N_14784,N_14852);
and U15111 (N_15111,N_14886,N_14895);
and U15112 (N_15112,N_14875,N_14863);
or U15113 (N_15113,N_14902,N_14981);
or U15114 (N_15114,N_14791,N_14926);
nand U15115 (N_15115,N_14932,N_14811);
xnor U15116 (N_15116,N_14908,N_14851);
xor U15117 (N_15117,N_14883,N_14816);
xor U15118 (N_15118,N_14840,N_14962);
and U15119 (N_15119,N_14936,N_14922);
xnor U15120 (N_15120,N_14797,N_14880);
or U15121 (N_15121,N_14969,N_14767);
nor U15122 (N_15122,N_14777,N_14838);
xnor U15123 (N_15123,N_14950,N_14985);
xor U15124 (N_15124,N_14837,N_14957);
nand U15125 (N_15125,N_14789,N_14784);
and U15126 (N_15126,N_14893,N_14846);
and U15127 (N_15127,N_14756,N_14841);
nand U15128 (N_15128,N_14827,N_14830);
nand U15129 (N_15129,N_14843,N_14895);
and U15130 (N_15130,N_14892,N_14814);
and U15131 (N_15131,N_14755,N_14962);
nand U15132 (N_15132,N_14793,N_14969);
or U15133 (N_15133,N_14883,N_14970);
or U15134 (N_15134,N_14886,N_14935);
and U15135 (N_15135,N_14902,N_14883);
nand U15136 (N_15136,N_14966,N_14788);
nand U15137 (N_15137,N_14898,N_14987);
xor U15138 (N_15138,N_14835,N_14882);
xor U15139 (N_15139,N_14950,N_14751);
xnor U15140 (N_15140,N_14913,N_14775);
nor U15141 (N_15141,N_14919,N_14864);
xor U15142 (N_15142,N_14824,N_14916);
nand U15143 (N_15143,N_14892,N_14797);
nor U15144 (N_15144,N_14791,N_14796);
or U15145 (N_15145,N_14962,N_14765);
nand U15146 (N_15146,N_14859,N_14845);
and U15147 (N_15147,N_14916,N_14757);
nor U15148 (N_15148,N_14852,N_14947);
nor U15149 (N_15149,N_14927,N_14779);
xnor U15150 (N_15150,N_14965,N_14866);
nand U15151 (N_15151,N_14952,N_14853);
and U15152 (N_15152,N_14752,N_14786);
xnor U15153 (N_15153,N_14858,N_14871);
or U15154 (N_15154,N_14826,N_14852);
xnor U15155 (N_15155,N_14780,N_14943);
and U15156 (N_15156,N_14890,N_14841);
nand U15157 (N_15157,N_14841,N_14919);
or U15158 (N_15158,N_14926,N_14987);
or U15159 (N_15159,N_14926,N_14883);
nand U15160 (N_15160,N_14800,N_14783);
nor U15161 (N_15161,N_14989,N_14873);
and U15162 (N_15162,N_14803,N_14891);
nor U15163 (N_15163,N_14984,N_14999);
or U15164 (N_15164,N_14855,N_14870);
and U15165 (N_15165,N_14767,N_14816);
xor U15166 (N_15166,N_14889,N_14970);
and U15167 (N_15167,N_14811,N_14761);
and U15168 (N_15168,N_14951,N_14904);
and U15169 (N_15169,N_14899,N_14878);
nand U15170 (N_15170,N_14984,N_14775);
and U15171 (N_15171,N_14819,N_14818);
nand U15172 (N_15172,N_14797,N_14757);
or U15173 (N_15173,N_14751,N_14993);
xnor U15174 (N_15174,N_14790,N_14902);
or U15175 (N_15175,N_14964,N_14841);
nand U15176 (N_15176,N_14853,N_14956);
and U15177 (N_15177,N_14783,N_14940);
or U15178 (N_15178,N_14894,N_14853);
or U15179 (N_15179,N_14968,N_14869);
xnor U15180 (N_15180,N_14917,N_14877);
xor U15181 (N_15181,N_14944,N_14959);
and U15182 (N_15182,N_14847,N_14887);
nand U15183 (N_15183,N_14991,N_14850);
nand U15184 (N_15184,N_14985,N_14887);
xnor U15185 (N_15185,N_14762,N_14936);
nor U15186 (N_15186,N_14797,N_14918);
and U15187 (N_15187,N_14875,N_14785);
or U15188 (N_15188,N_14772,N_14750);
and U15189 (N_15189,N_14955,N_14841);
nand U15190 (N_15190,N_14968,N_14801);
and U15191 (N_15191,N_14971,N_14770);
nor U15192 (N_15192,N_14910,N_14786);
nand U15193 (N_15193,N_14848,N_14806);
xor U15194 (N_15194,N_14988,N_14897);
or U15195 (N_15195,N_14927,N_14964);
nand U15196 (N_15196,N_14870,N_14784);
xor U15197 (N_15197,N_14781,N_14972);
xor U15198 (N_15198,N_14857,N_14818);
nand U15199 (N_15199,N_14751,N_14793);
and U15200 (N_15200,N_14771,N_14998);
nand U15201 (N_15201,N_14867,N_14913);
nor U15202 (N_15202,N_14801,N_14848);
or U15203 (N_15203,N_14955,N_14753);
nand U15204 (N_15204,N_14987,N_14762);
nand U15205 (N_15205,N_14921,N_14853);
xnor U15206 (N_15206,N_14949,N_14864);
nand U15207 (N_15207,N_14955,N_14783);
and U15208 (N_15208,N_14830,N_14911);
or U15209 (N_15209,N_14888,N_14750);
nor U15210 (N_15210,N_14996,N_14828);
xor U15211 (N_15211,N_14760,N_14974);
or U15212 (N_15212,N_14831,N_14970);
or U15213 (N_15213,N_14967,N_14894);
xnor U15214 (N_15214,N_14978,N_14952);
nand U15215 (N_15215,N_14827,N_14941);
nor U15216 (N_15216,N_14821,N_14965);
or U15217 (N_15217,N_14923,N_14931);
and U15218 (N_15218,N_14992,N_14847);
nor U15219 (N_15219,N_14859,N_14799);
xor U15220 (N_15220,N_14929,N_14809);
nor U15221 (N_15221,N_14905,N_14904);
or U15222 (N_15222,N_14799,N_14830);
nor U15223 (N_15223,N_14789,N_14764);
or U15224 (N_15224,N_14912,N_14920);
and U15225 (N_15225,N_14992,N_14928);
xnor U15226 (N_15226,N_14845,N_14773);
nand U15227 (N_15227,N_14799,N_14803);
xnor U15228 (N_15228,N_14995,N_14785);
or U15229 (N_15229,N_14854,N_14823);
or U15230 (N_15230,N_14987,N_14828);
nor U15231 (N_15231,N_14897,N_14917);
nand U15232 (N_15232,N_14827,N_14894);
nand U15233 (N_15233,N_14864,N_14905);
or U15234 (N_15234,N_14750,N_14845);
xnor U15235 (N_15235,N_14876,N_14995);
nor U15236 (N_15236,N_14841,N_14940);
nor U15237 (N_15237,N_14855,N_14930);
and U15238 (N_15238,N_14915,N_14800);
nand U15239 (N_15239,N_14923,N_14908);
and U15240 (N_15240,N_14893,N_14963);
nor U15241 (N_15241,N_14934,N_14834);
xor U15242 (N_15242,N_14983,N_14772);
xnor U15243 (N_15243,N_14914,N_14917);
nor U15244 (N_15244,N_14894,N_14794);
nor U15245 (N_15245,N_14824,N_14907);
and U15246 (N_15246,N_14910,N_14846);
nand U15247 (N_15247,N_14849,N_14938);
nor U15248 (N_15248,N_14775,N_14925);
or U15249 (N_15249,N_14929,N_14956);
and U15250 (N_15250,N_15195,N_15150);
and U15251 (N_15251,N_15073,N_15038);
nor U15252 (N_15252,N_15063,N_15170);
nand U15253 (N_15253,N_15103,N_15010);
nand U15254 (N_15254,N_15119,N_15231);
or U15255 (N_15255,N_15031,N_15015);
nand U15256 (N_15256,N_15002,N_15186);
or U15257 (N_15257,N_15076,N_15071);
or U15258 (N_15258,N_15207,N_15190);
nor U15259 (N_15259,N_15023,N_15104);
nor U15260 (N_15260,N_15155,N_15222);
nor U15261 (N_15261,N_15235,N_15118);
nand U15262 (N_15262,N_15134,N_15246);
or U15263 (N_15263,N_15078,N_15029);
xor U15264 (N_15264,N_15218,N_15021);
nand U15265 (N_15265,N_15234,N_15097);
or U15266 (N_15266,N_15072,N_15171);
xnor U15267 (N_15267,N_15042,N_15243);
nor U15268 (N_15268,N_15056,N_15146);
nand U15269 (N_15269,N_15004,N_15140);
and U15270 (N_15270,N_15033,N_15001);
and U15271 (N_15271,N_15201,N_15233);
nor U15272 (N_15272,N_15088,N_15249);
xnor U15273 (N_15273,N_15153,N_15161);
nand U15274 (N_15274,N_15123,N_15093);
or U15275 (N_15275,N_15035,N_15247);
nor U15276 (N_15276,N_15084,N_15160);
or U15277 (N_15277,N_15232,N_15107);
xor U15278 (N_15278,N_15239,N_15180);
nand U15279 (N_15279,N_15205,N_15040);
nand U15280 (N_15280,N_15053,N_15047);
xor U15281 (N_15281,N_15112,N_15227);
or U15282 (N_15282,N_15157,N_15037);
nor U15283 (N_15283,N_15085,N_15086);
xnor U15284 (N_15284,N_15109,N_15177);
nand U15285 (N_15285,N_15049,N_15028);
xnor U15286 (N_15286,N_15100,N_15238);
nor U15287 (N_15287,N_15012,N_15151);
or U15288 (N_15288,N_15025,N_15237);
xor U15289 (N_15289,N_15051,N_15189);
or U15290 (N_15290,N_15115,N_15041);
nor U15291 (N_15291,N_15193,N_15198);
nor U15292 (N_15292,N_15060,N_15122);
and U15293 (N_15293,N_15216,N_15054);
xor U15294 (N_15294,N_15163,N_15217);
nand U15295 (N_15295,N_15050,N_15081);
xnor U15296 (N_15296,N_15080,N_15143);
nor U15297 (N_15297,N_15066,N_15101);
nand U15298 (N_15298,N_15077,N_15057);
or U15299 (N_15299,N_15075,N_15202);
xor U15300 (N_15300,N_15114,N_15067);
and U15301 (N_15301,N_15181,N_15007);
and U15302 (N_15302,N_15108,N_15148);
nor U15303 (N_15303,N_15131,N_15182);
nor U15304 (N_15304,N_15110,N_15124);
and U15305 (N_15305,N_15069,N_15090);
nor U15306 (N_15306,N_15045,N_15221);
xor U15307 (N_15307,N_15199,N_15185);
or U15308 (N_15308,N_15164,N_15242);
or U15309 (N_15309,N_15011,N_15194);
nor U15310 (N_15310,N_15070,N_15200);
nor U15311 (N_15311,N_15089,N_15154);
xor U15312 (N_15312,N_15027,N_15026);
nor U15313 (N_15313,N_15174,N_15228);
nor U15314 (N_15314,N_15208,N_15014);
and U15315 (N_15315,N_15064,N_15149);
and U15316 (N_15316,N_15229,N_15017);
or U15317 (N_15317,N_15020,N_15032);
xor U15318 (N_15318,N_15166,N_15136);
nor U15319 (N_15319,N_15046,N_15209);
xnor U15320 (N_15320,N_15219,N_15137);
xor U15321 (N_15321,N_15102,N_15224);
nor U15322 (N_15322,N_15203,N_15039);
xnor U15323 (N_15323,N_15223,N_15142);
nand U15324 (N_15324,N_15248,N_15175);
and U15325 (N_15325,N_15133,N_15183);
or U15326 (N_15326,N_15152,N_15048);
nand U15327 (N_15327,N_15132,N_15003);
and U15328 (N_15328,N_15236,N_15144);
nand U15329 (N_15329,N_15240,N_15068);
xor U15330 (N_15330,N_15117,N_15120);
and U15331 (N_15331,N_15214,N_15024);
xnor U15332 (N_15332,N_15168,N_15096);
nand U15333 (N_15333,N_15135,N_15098);
xor U15334 (N_15334,N_15055,N_15074);
xnor U15335 (N_15335,N_15082,N_15094);
xor U15336 (N_15336,N_15187,N_15044);
xnor U15337 (N_15337,N_15092,N_15197);
or U15338 (N_15338,N_15206,N_15006);
xnor U15339 (N_15339,N_15139,N_15178);
xor U15340 (N_15340,N_15127,N_15106);
xor U15341 (N_15341,N_15022,N_15169);
and U15342 (N_15342,N_15125,N_15220);
nor U15343 (N_15343,N_15113,N_15213);
and U15344 (N_15344,N_15147,N_15167);
nor U15345 (N_15345,N_15244,N_15009);
nand U15346 (N_15346,N_15034,N_15138);
or U15347 (N_15347,N_15212,N_15000);
nor U15348 (N_15348,N_15019,N_15173);
and U15349 (N_15349,N_15005,N_15105);
nand U15350 (N_15350,N_15016,N_15162);
xnor U15351 (N_15351,N_15192,N_15059);
or U15352 (N_15352,N_15145,N_15065);
nor U15353 (N_15353,N_15188,N_15018);
and U15354 (N_15354,N_15156,N_15083);
xnor U15355 (N_15355,N_15211,N_15062);
and U15356 (N_15356,N_15095,N_15129);
or U15357 (N_15357,N_15241,N_15191);
xnor U15358 (N_15358,N_15225,N_15226);
and U15359 (N_15359,N_15245,N_15091);
xor U15360 (N_15360,N_15141,N_15043);
nor U15361 (N_15361,N_15058,N_15196);
nand U15362 (N_15362,N_15204,N_15052);
or U15363 (N_15363,N_15215,N_15165);
or U15364 (N_15364,N_15210,N_15116);
nor U15365 (N_15365,N_15121,N_15111);
nand U15366 (N_15366,N_15230,N_15130);
and U15367 (N_15367,N_15013,N_15008);
nor U15368 (N_15368,N_15158,N_15079);
nor U15369 (N_15369,N_15172,N_15126);
or U15370 (N_15370,N_15176,N_15184);
xnor U15371 (N_15371,N_15128,N_15087);
xor U15372 (N_15372,N_15030,N_15159);
nor U15373 (N_15373,N_15099,N_15036);
xnor U15374 (N_15374,N_15061,N_15179);
nor U15375 (N_15375,N_15180,N_15144);
and U15376 (N_15376,N_15141,N_15106);
and U15377 (N_15377,N_15162,N_15197);
or U15378 (N_15378,N_15008,N_15036);
or U15379 (N_15379,N_15204,N_15110);
or U15380 (N_15380,N_15053,N_15021);
or U15381 (N_15381,N_15129,N_15056);
xnor U15382 (N_15382,N_15228,N_15020);
nand U15383 (N_15383,N_15044,N_15048);
and U15384 (N_15384,N_15033,N_15165);
xnor U15385 (N_15385,N_15013,N_15087);
or U15386 (N_15386,N_15053,N_15037);
or U15387 (N_15387,N_15142,N_15119);
nor U15388 (N_15388,N_15118,N_15115);
xor U15389 (N_15389,N_15218,N_15009);
and U15390 (N_15390,N_15165,N_15016);
xor U15391 (N_15391,N_15003,N_15072);
and U15392 (N_15392,N_15011,N_15067);
and U15393 (N_15393,N_15216,N_15058);
nand U15394 (N_15394,N_15042,N_15207);
nor U15395 (N_15395,N_15066,N_15106);
nand U15396 (N_15396,N_15013,N_15125);
and U15397 (N_15397,N_15248,N_15150);
and U15398 (N_15398,N_15240,N_15141);
nand U15399 (N_15399,N_15173,N_15221);
or U15400 (N_15400,N_15114,N_15214);
nand U15401 (N_15401,N_15167,N_15001);
nand U15402 (N_15402,N_15120,N_15037);
nand U15403 (N_15403,N_15200,N_15210);
nand U15404 (N_15404,N_15060,N_15010);
xor U15405 (N_15405,N_15249,N_15147);
nor U15406 (N_15406,N_15059,N_15097);
or U15407 (N_15407,N_15216,N_15116);
or U15408 (N_15408,N_15051,N_15242);
nor U15409 (N_15409,N_15026,N_15239);
nor U15410 (N_15410,N_15145,N_15158);
or U15411 (N_15411,N_15022,N_15200);
nor U15412 (N_15412,N_15234,N_15007);
xor U15413 (N_15413,N_15025,N_15062);
nor U15414 (N_15414,N_15046,N_15077);
xor U15415 (N_15415,N_15222,N_15142);
or U15416 (N_15416,N_15065,N_15113);
nand U15417 (N_15417,N_15036,N_15112);
and U15418 (N_15418,N_15004,N_15189);
or U15419 (N_15419,N_15027,N_15182);
and U15420 (N_15420,N_15083,N_15087);
and U15421 (N_15421,N_15032,N_15061);
nor U15422 (N_15422,N_15094,N_15225);
and U15423 (N_15423,N_15146,N_15132);
xor U15424 (N_15424,N_15216,N_15076);
nor U15425 (N_15425,N_15104,N_15214);
or U15426 (N_15426,N_15107,N_15196);
or U15427 (N_15427,N_15101,N_15226);
and U15428 (N_15428,N_15069,N_15058);
or U15429 (N_15429,N_15242,N_15152);
nand U15430 (N_15430,N_15078,N_15224);
xor U15431 (N_15431,N_15151,N_15219);
xor U15432 (N_15432,N_15118,N_15045);
nor U15433 (N_15433,N_15120,N_15013);
xor U15434 (N_15434,N_15052,N_15149);
or U15435 (N_15435,N_15015,N_15098);
xnor U15436 (N_15436,N_15098,N_15222);
or U15437 (N_15437,N_15223,N_15195);
xor U15438 (N_15438,N_15100,N_15227);
and U15439 (N_15439,N_15167,N_15115);
nor U15440 (N_15440,N_15045,N_15173);
or U15441 (N_15441,N_15196,N_15096);
xor U15442 (N_15442,N_15007,N_15232);
or U15443 (N_15443,N_15164,N_15146);
xnor U15444 (N_15444,N_15077,N_15082);
or U15445 (N_15445,N_15070,N_15016);
xor U15446 (N_15446,N_15143,N_15200);
nand U15447 (N_15447,N_15016,N_15231);
or U15448 (N_15448,N_15042,N_15083);
nor U15449 (N_15449,N_15125,N_15207);
xor U15450 (N_15450,N_15066,N_15175);
and U15451 (N_15451,N_15229,N_15170);
nor U15452 (N_15452,N_15084,N_15149);
or U15453 (N_15453,N_15075,N_15208);
xnor U15454 (N_15454,N_15133,N_15171);
xor U15455 (N_15455,N_15089,N_15178);
or U15456 (N_15456,N_15076,N_15080);
nand U15457 (N_15457,N_15162,N_15056);
and U15458 (N_15458,N_15219,N_15193);
or U15459 (N_15459,N_15090,N_15112);
nor U15460 (N_15460,N_15220,N_15029);
xnor U15461 (N_15461,N_15010,N_15069);
or U15462 (N_15462,N_15208,N_15151);
nor U15463 (N_15463,N_15040,N_15182);
xnor U15464 (N_15464,N_15034,N_15122);
xor U15465 (N_15465,N_15034,N_15091);
nand U15466 (N_15466,N_15099,N_15149);
and U15467 (N_15467,N_15066,N_15232);
xnor U15468 (N_15468,N_15048,N_15204);
or U15469 (N_15469,N_15154,N_15190);
nand U15470 (N_15470,N_15053,N_15138);
or U15471 (N_15471,N_15170,N_15143);
or U15472 (N_15472,N_15062,N_15181);
or U15473 (N_15473,N_15163,N_15186);
and U15474 (N_15474,N_15138,N_15098);
and U15475 (N_15475,N_15213,N_15012);
nand U15476 (N_15476,N_15216,N_15214);
xnor U15477 (N_15477,N_15148,N_15228);
xor U15478 (N_15478,N_15129,N_15236);
nand U15479 (N_15479,N_15125,N_15172);
nand U15480 (N_15480,N_15157,N_15005);
and U15481 (N_15481,N_15054,N_15238);
xor U15482 (N_15482,N_15140,N_15057);
xor U15483 (N_15483,N_15219,N_15119);
or U15484 (N_15484,N_15046,N_15145);
and U15485 (N_15485,N_15092,N_15078);
nand U15486 (N_15486,N_15109,N_15128);
nor U15487 (N_15487,N_15146,N_15028);
or U15488 (N_15488,N_15213,N_15150);
xor U15489 (N_15489,N_15241,N_15023);
nor U15490 (N_15490,N_15130,N_15163);
nand U15491 (N_15491,N_15025,N_15029);
or U15492 (N_15492,N_15021,N_15132);
and U15493 (N_15493,N_15220,N_15111);
or U15494 (N_15494,N_15014,N_15202);
or U15495 (N_15495,N_15156,N_15199);
xnor U15496 (N_15496,N_15080,N_15040);
and U15497 (N_15497,N_15181,N_15060);
xnor U15498 (N_15498,N_15063,N_15142);
and U15499 (N_15499,N_15224,N_15046);
and U15500 (N_15500,N_15350,N_15392);
xor U15501 (N_15501,N_15287,N_15343);
xnor U15502 (N_15502,N_15474,N_15494);
or U15503 (N_15503,N_15446,N_15498);
and U15504 (N_15504,N_15303,N_15420);
and U15505 (N_15505,N_15449,N_15497);
and U15506 (N_15506,N_15486,N_15275);
and U15507 (N_15507,N_15262,N_15280);
and U15508 (N_15508,N_15269,N_15396);
nor U15509 (N_15509,N_15376,N_15489);
xnor U15510 (N_15510,N_15456,N_15306);
and U15511 (N_15511,N_15296,N_15441);
or U15512 (N_15512,N_15437,N_15381);
xnor U15513 (N_15513,N_15468,N_15423);
and U15514 (N_15514,N_15373,N_15279);
or U15515 (N_15515,N_15499,N_15254);
xnor U15516 (N_15516,N_15355,N_15271);
nor U15517 (N_15517,N_15490,N_15365);
and U15518 (N_15518,N_15375,N_15337);
nor U15519 (N_15519,N_15487,N_15290);
nand U15520 (N_15520,N_15266,N_15388);
nor U15521 (N_15521,N_15444,N_15384);
nand U15522 (N_15522,N_15305,N_15410);
and U15523 (N_15523,N_15327,N_15276);
nor U15524 (N_15524,N_15480,N_15263);
nand U15525 (N_15525,N_15292,N_15430);
nand U15526 (N_15526,N_15323,N_15251);
nor U15527 (N_15527,N_15493,N_15464);
xor U15528 (N_15528,N_15418,N_15301);
nand U15529 (N_15529,N_15378,N_15286);
nand U15530 (N_15530,N_15492,N_15409);
nand U15531 (N_15531,N_15435,N_15316);
or U15532 (N_15532,N_15330,N_15436);
xnor U15533 (N_15533,N_15288,N_15377);
nand U15534 (N_15534,N_15320,N_15479);
nand U15535 (N_15535,N_15427,N_15344);
xor U15536 (N_15536,N_15260,N_15340);
xnor U15537 (N_15537,N_15358,N_15372);
and U15538 (N_15538,N_15360,N_15397);
xor U15539 (N_15539,N_15349,N_15447);
nor U15540 (N_15540,N_15407,N_15453);
or U15541 (N_15541,N_15440,N_15332);
nor U15542 (N_15542,N_15465,N_15382);
nor U15543 (N_15543,N_15282,N_15258);
and U15544 (N_15544,N_15411,N_15253);
and U15545 (N_15545,N_15272,N_15293);
nor U15546 (N_15546,N_15270,N_15485);
nand U15547 (N_15547,N_15257,N_15277);
nor U15548 (N_15548,N_15267,N_15475);
or U15549 (N_15549,N_15256,N_15307);
and U15550 (N_15550,N_15426,N_15273);
nor U15551 (N_15551,N_15317,N_15419);
and U15552 (N_15552,N_15405,N_15471);
nand U15553 (N_15553,N_15359,N_15429);
or U15554 (N_15554,N_15398,N_15477);
or U15555 (N_15555,N_15297,N_15434);
or U15556 (N_15556,N_15342,N_15472);
xor U15557 (N_15557,N_15274,N_15348);
nand U15558 (N_15558,N_15466,N_15404);
or U15559 (N_15559,N_15285,N_15473);
or U15560 (N_15560,N_15321,N_15283);
nor U15561 (N_15561,N_15463,N_15338);
xnor U15562 (N_15562,N_15354,N_15457);
or U15563 (N_15563,N_15281,N_15268);
nand U15564 (N_15564,N_15425,N_15302);
nor U15565 (N_15565,N_15361,N_15461);
nor U15566 (N_15566,N_15390,N_15328);
and U15567 (N_15567,N_15408,N_15250);
and U15568 (N_15568,N_15364,N_15326);
nor U15569 (N_15569,N_15433,N_15439);
and U15570 (N_15570,N_15368,N_15482);
nand U15571 (N_15571,N_15393,N_15413);
nand U15572 (N_15572,N_15289,N_15476);
xnor U15573 (N_15573,N_15265,N_15451);
nor U15574 (N_15574,N_15367,N_15389);
nor U15575 (N_15575,N_15469,N_15278);
nor U15576 (N_15576,N_15385,N_15394);
and U15577 (N_15577,N_15264,N_15450);
xor U15578 (N_15578,N_15333,N_15255);
nor U15579 (N_15579,N_15379,N_15324);
or U15580 (N_15580,N_15318,N_15334);
nor U15581 (N_15581,N_15417,N_15462);
or U15582 (N_15582,N_15366,N_15496);
and U15583 (N_15583,N_15402,N_15294);
and U15584 (N_15584,N_15415,N_15403);
or U15585 (N_15585,N_15319,N_15495);
nand U15586 (N_15586,N_15443,N_15458);
or U15587 (N_15587,N_15484,N_15295);
nand U15588 (N_15588,N_15298,N_15353);
nor U15589 (N_15589,N_15454,N_15261);
and U15590 (N_15590,N_15470,N_15357);
xnor U15591 (N_15591,N_15452,N_15478);
nor U15592 (N_15592,N_15406,N_15336);
or U15593 (N_15593,N_15455,N_15335);
nor U15594 (N_15594,N_15339,N_15481);
nor U15595 (N_15595,N_15414,N_15346);
nand U15596 (N_15596,N_15448,N_15421);
nand U15597 (N_15597,N_15284,N_15445);
and U15598 (N_15598,N_15299,N_15308);
and U15599 (N_15599,N_15362,N_15309);
nor U15600 (N_15600,N_15325,N_15467);
and U15601 (N_15601,N_15363,N_15431);
and U15602 (N_15602,N_15345,N_15459);
and U15603 (N_15603,N_15347,N_15311);
nor U15604 (N_15604,N_15483,N_15300);
nor U15605 (N_15605,N_15386,N_15329);
xor U15606 (N_15606,N_15424,N_15387);
and U15607 (N_15607,N_15442,N_15304);
nand U15608 (N_15608,N_15374,N_15460);
nand U15609 (N_15609,N_15356,N_15400);
or U15610 (N_15610,N_15438,N_15313);
nor U15611 (N_15611,N_15351,N_15401);
and U15612 (N_15612,N_15341,N_15395);
xor U15613 (N_15613,N_15371,N_15369);
xnor U15614 (N_15614,N_15491,N_15312);
and U15615 (N_15615,N_15416,N_15380);
and U15616 (N_15616,N_15488,N_15428);
nor U15617 (N_15617,N_15291,N_15412);
and U15618 (N_15618,N_15422,N_15310);
nand U15619 (N_15619,N_15315,N_15314);
xor U15620 (N_15620,N_15399,N_15331);
and U15621 (N_15621,N_15383,N_15370);
or U15622 (N_15622,N_15322,N_15352);
and U15623 (N_15623,N_15391,N_15432);
xnor U15624 (N_15624,N_15252,N_15259);
nor U15625 (N_15625,N_15289,N_15458);
or U15626 (N_15626,N_15402,N_15368);
and U15627 (N_15627,N_15277,N_15372);
nor U15628 (N_15628,N_15433,N_15267);
nor U15629 (N_15629,N_15434,N_15294);
nor U15630 (N_15630,N_15327,N_15361);
xor U15631 (N_15631,N_15317,N_15420);
nor U15632 (N_15632,N_15258,N_15435);
nor U15633 (N_15633,N_15373,N_15466);
nand U15634 (N_15634,N_15373,N_15348);
xnor U15635 (N_15635,N_15403,N_15452);
nor U15636 (N_15636,N_15481,N_15454);
or U15637 (N_15637,N_15461,N_15256);
and U15638 (N_15638,N_15438,N_15461);
nand U15639 (N_15639,N_15370,N_15314);
xnor U15640 (N_15640,N_15356,N_15427);
or U15641 (N_15641,N_15271,N_15278);
and U15642 (N_15642,N_15407,N_15290);
nand U15643 (N_15643,N_15303,N_15381);
nand U15644 (N_15644,N_15351,N_15426);
xnor U15645 (N_15645,N_15337,N_15489);
xor U15646 (N_15646,N_15421,N_15308);
or U15647 (N_15647,N_15460,N_15439);
and U15648 (N_15648,N_15366,N_15371);
nand U15649 (N_15649,N_15256,N_15261);
and U15650 (N_15650,N_15470,N_15378);
xnor U15651 (N_15651,N_15320,N_15335);
and U15652 (N_15652,N_15376,N_15325);
nor U15653 (N_15653,N_15469,N_15263);
xnor U15654 (N_15654,N_15492,N_15260);
xnor U15655 (N_15655,N_15457,N_15426);
or U15656 (N_15656,N_15439,N_15459);
xor U15657 (N_15657,N_15332,N_15460);
or U15658 (N_15658,N_15341,N_15491);
xor U15659 (N_15659,N_15325,N_15433);
xor U15660 (N_15660,N_15297,N_15253);
or U15661 (N_15661,N_15334,N_15315);
nor U15662 (N_15662,N_15268,N_15296);
xnor U15663 (N_15663,N_15391,N_15309);
and U15664 (N_15664,N_15456,N_15285);
and U15665 (N_15665,N_15485,N_15456);
or U15666 (N_15666,N_15359,N_15375);
or U15667 (N_15667,N_15261,N_15413);
and U15668 (N_15668,N_15251,N_15300);
and U15669 (N_15669,N_15423,N_15467);
nor U15670 (N_15670,N_15451,N_15303);
xor U15671 (N_15671,N_15361,N_15311);
nand U15672 (N_15672,N_15357,N_15404);
or U15673 (N_15673,N_15432,N_15497);
and U15674 (N_15674,N_15275,N_15436);
and U15675 (N_15675,N_15277,N_15394);
xnor U15676 (N_15676,N_15467,N_15309);
xor U15677 (N_15677,N_15285,N_15454);
or U15678 (N_15678,N_15289,N_15251);
nand U15679 (N_15679,N_15354,N_15361);
or U15680 (N_15680,N_15261,N_15303);
nand U15681 (N_15681,N_15310,N_15338);
xor U15682 (N_15682,N_15347,N_15459);
nand U15683 (N_15683,N_15422,N_15278);
nor U15684 (N_15684,N_15256,N_15303);
nor U15685 (N_15685,N_15295,N_15314);
nor U15686 (N_15686,N_15484,N_15453);
nand U15687 (N_15687,N_15454,N_15359);
xor U15688 (N_15688,N_15385,N_15316);
nand U15689 (N_15689,N_15342,N_15273);
or U15690 (N_15690,N_15274,N_15347);
nor U15691 (N_15691,N_15377,N_15482);
nand U15692 (N_15692,N_15497,N_15334);
nand U15693 (N_15693,N_15377,N_15398);
nand U15694 (N_15694,N_15369,N_15277);
and U15695 (N_15695,N_15331,N_15318);
and U15696 (N_15696,N_15388,N_15339);
and U15697 (N_15697,N_15458,N_15269);
or U15698 (N_15698,N_15270,N_15315);
xnor U15699 (N_15699,N_15481,N_15384);
and U15700 (N_15700,N_15342,N_15265);
nand U15701 (N_15701,N_15313,N_15408);
and U15702 (N_15702,N_15472,N_15395);
nor U15703 (N_15703,N_15376,N_15294);
or U15704 (N_15704,N_15331,N_15465);
or U15705 (N_15705,N_15407,N_15472);
and U15706 (N_15706,N_15272,N_15376);
and U15707 (N_15707,N_15299,N_15446);
nand U15708 (N_15708,N_15384,N_15292);
and U15709 (N_15709,N_15291,N_15475);
nor U15710 (N_15710,N_15303,N_15346);
nand U15711 (N_15711,N_15276,N_15459);
nor U15712 (N_15712,N_15480,N_15371);
or U15713 (N_15713,N_15494,N_15377);
xnor U15714 (N_15714,N_15399,N_15383);
nand U15715 (N_15715,N_15448,N_15400);
xor U15716 (N_15716,N_15256,N_15335);
or U15717 (N_15717,N_15492,N_15277);
xnor U15718 (N_15718,N_15345,N_15463);
and U15719 (N_15719,N_15443,N_15317);
xor U15720 (N_15720,N_15457,N_15326);
xor U15721 (N_15721,N_15476,N_15281);
nand U15722 (N_15722,N_15420,N_15490);
nor U15723 (N_15723,N_15333,N_15360);
xnor U15724 (N_15724,N_15256,N_15419);
and U15725 (N_15725,N_15322,N_15257);
nor U15726 (N_15726,N_15315,N_15358);
xnor U15727 (N_15727,N_15254,N_15359);
or U15728 (N_15728,N_15351,N_15342);
nand U15729 (N_15729,N_15257,N_15392);
nand U15730 (N_15730,N_15384,N_15472);
nand U15731 (N_15731,N_15404,N_15471);
nor U15732 (N_15732,N_15457,N_15299);
nor U15733 (N_15733,N_15487,N_15494);
and U15734 (N_15734,N_15351,N_15455);
xor U15735 (N_15735,N_15479,N_15321);
or U15736 (N_15736,N_15309,N_15320);
xor U15737 (N_15737,N_15483,N_15384);
or U15738 (N_15738,N_15479,N_15365);
xnor U15739 (N_15739,N_15255,N_15251);
or U15740 (N_15740,N_15446,N_15494);
xnor U15741 (N_15741,N_15279,N_15499);
nor U15742 (N_15742,N_15409,N_15436);
nand U15743 (N_15743,N_15395,N_15270);
nor U15744 (N_15744,N_15418,N_15315);
or U15745 (N_15745,N_15454,N_15414);
or U15746 (N_15746,N_15420,N_15295);
nor U15747 (N_15747,N_15475,N_15353);
nand U15748 (N_15748,N_15299,N_15355);
nor U15749 (N_15749,N_15387,N_15320);
nand U15750 (N_15750,N_15619,N_15602);
or U15751 (N_15751,N_15631,N_15668);
xnor U15752 (N_15752,N_15712,N_15688);
xor U15753 (N_15753,N_15696,N_15669);
xor U15754 (N_15754,N_15566,N_15747);
xor U15755 (N_15755,N_15636,N_15689);
nand U15756 (N_15756,N_15629,N_15730);
nand U15757 (N_15757,N_15722,N_15522);
nand U15758 (N_15758,N_15561,N_15701);
nor U15759 (N_15759,N_15560,N_15516);
xnor U15760 (N_15760,N_15505,N_15657);
xnor U15761 (N_15761,N_15533,N_15732);
nor U15762 (N_15762,N_15726,N_15659);
and U15763 (N_15763,N_15695,N_15616);
nand U15764 (N_15764,N_15655,N_15585);
nor U15765 (N_15765,N_15690,N_15511);
nand U15766 (N_15766,N_15582,N_15581);
and U15767 (N_15767,N_15627,N_15645);
or U15768 (N_15768,N_15683,N_15502);
nand U15769 (N_15769,N_15596,N_15628);
or U15770 (N_15770,N_15654,N_15548);
or U15771 (N_15771,N_15698,N_15664);
and U15772 (N_15772,N_15643,N_15575);
and U15773 (N_15773,N_15630,N_15592);
nor U15774 (N_15774,N_15598,N_15684);
nor U15775 (N_15775,N_15620,N_15617);
xor U15776 (N_15776,N_15538,N_15546);
nor U15777 (N_15777,N_15715,N_15680);
nand U15778 (N_15778,N_15625,N_15723);
nand U15779 (N_15779,N_15749,N_15651);
or U15780 (N_15780,N_15624,N_15681);
nand U15781 (N_15781,N_15674,N_15536);
nor U15782 (N_15782,N_15742,N_15648);
or U15783 (N_15783,N_15621,N_15554);
nor U15784 (N_15784,N_15593,N_15504);
nor U15785 (N_15785,N_15608,N_15559);
xnor U15786 (N_15786,N_15740,N_15633);
xnor U15787 (N_15787,N_15594,N_15580);
or U15788 (N_15788,N_15507,N_15512);
and U15789 (N_15789,N_15686,N_15545);
or U15790 (N_15790,N_15589,N_15597);
xor U15791 (N_15791,N_15720,N_15708);
and U15792 (N_15792,N_15642,N_15524);
and U15793 (N_15793,N_15635,N_15532);
nand U15794 (N_15794,N_15662,N_15705);
xor U15795 (N_15795,N_15703,N_15601);
nand U15796 (N_15796,N_15550,N_15738);
xnor U15797 (N_15797,N_15564,N_15676);
or U15798 (N_15798,N_15724,N_15562);
nor U15799 (N_15799,N_15711,N_15661);
nand U15800 (N_15800,N_15650,N_15685);
and U15801 (N_15801,N_15614,N_15634);
nor U15802 (N_15802,N_15599,N_15671);
or U15803 (N_15803,N_15518,N_15539);
nor U15804 (N_15804,N_15544,N_15748);
or U15805 (N_15805,N_15509,N_15534);
nand U15806 (N_15806,N_15541,N_15741);
nor U15807 (N_15807,N_15666,N_15728);
xor U15808 (N_15808,N_15658,N_15530);
and U15809 (N_15809,N_15605,N_15653);
or U15810 (N_15810,N_15535,N_15514);
nand U15811 (N_15811,N_15610,N_15637);
or U15812 (N_15812,N_15571,N_15691);
nor U15813 (N_15813,N_15604,N_15727);
and U15814 (N_15814,N_15672,N_15743);
and U15815 (N_15815,N_15503,N_15660);
xor U15816 (N_15816,N_15713,N_15697);
nand U15817 (N_15817,N_15734,N_15579);
and U15818 (N_15818,N_15557,N_15739);
nor U15819 (N_15819,N_15542,N_15649);
nor U15820 (N_15820,N_15652,N_15641);
and U15821 (N_15821,N_15521,N_15547);
nor U15822 (N_15822,N_15632,N_15717);
nor U15823 (N_15823,N_15626,N_15744);
xor U15824 (N_15824,N_15588,N_15563);
xnor U15825 (N_15825,N_15549,N_15615);
or U15826 (N_15826,N_15706,N_15577);
nand U15827 (N_15827,N_15737,N_15687);
nand U15828 (N_15828,N_15667,N_15607);
and U15829 (N_15829,N_15523,N_15520);
nor U15830 (N_15830,N_15731,N_15693);
nand U15831 (N_15831,N_15515,N_15510);
nand U15832 (N_15832,N_15600,N_15553);
and U15833 (N_15833,N_15555,N_15551);
nor U15834 (N_15834,N_15573,N_15568);
xor U15835 (N_15835,N_15500,N_15736);
xor U15836 (N_15836,N_15718,N_15572);
nor U15837 (N_15837,N_15525,N_15665);
nand U15838 (N_15838,N_15584,N_15663);
xnor U15839 (N_15839,N_15513,N_15576);
xor U15840 (N_15840,N_15638,N_15714);
and U15841 (N_15841,N_15506,N_15611);
or U15842 (N_15842,N_15517,N_15565);
nor U15843 (N_15843,N_15746,N_15719);
and U15844 (N_15844,N_15699,N_15733);
nor U15845 (N_15845,N_15745,N_15639);
xor U15846 (N_15846,N_15528,N_15569);
nor U15847 (N_15847,N_15692,N_15640);
nor U15848 (N_15848,N_15526,N_15670);
nor U15849 (N_15849,N_15537,N_15735);
and U15850 (N_15850,N_15729,N_15501);
or U15851 (N_15851,N_15700,N_15587);
nor U15852 (N_15852,N_15519,N_15583);
nor U15853 (N_15853,N_15647,N_15702);
nor U15854 (N_15854,N_15558,N_15578);
nand U15855 (N_15855,N_15531,N_15552);
nor U15856 (N_15856,N_15567,N_15622);
and U15857 (N_15857,N_15694,N_15704);
nand U15858 (N_15858,N_15603,N_15710);
nand U15859 (N_15859,N_15623,N_15716);
and U15860 (N_15860,N_15679,N_15707);
nor U15861 (N_15861,N_15606,N_15543);
nor U15862 (N_15862,N_15556,N_15590);
nor U15863 (N_15863,N_15612,N_15709);
or U15864 (N_15864,N_15595,N_15678);
and U15865 (N_15865,N_15656,N_15591);
nand U15866 (N_15866,N_15618,N_15508);
nor U15867 (N_15867,N_15677,N_15586);
nor U15868 (N_15868,N_15675,N_15725);
and U15869 (N_15869,N_15540,N_15682);
nand U15870 (N_15870,N_15527,N_15613);
nor U15871 (N_15871,N_15574,N_15721);
nor U15872 (N_15872,N_15529,N_15673);
nor U15873 (N_15873,N_15570,N_15646);
and U15874 (N_15874,N_15644,N_15609);
and U15875 (N_15875,N_15716,N_15638);
nor U15876 (N_15876,N_15511,N_15633);
xor U15877 (N_15877,N_15543,N_15643);
nand U15878 (N_15878,N_15567,N_15549);
nand U15879 (N_15879,N_15504,N_15717);
and U15880 (N_15880,N_15607,N_15554);
or U15881 (N_15881,N_15623,N_15727);
nand U15882 (N_15882,N_15639,N_15720);
nand U15883 (N_15883,N_15704,N_15563);
or U15884 (N_15884,N_15689,N_15592);
and U15885 (N_15885,N_15515,N_15633);
or U15886 (N_15886,N_15744,N_15701);
or U15887 (N_15887,N_15539,N_15725);
or U15888 (N_15888,N_15743,N_15641);
nand U15889 (N_15889,N_15651,N_15672);
xnor U15890 (N_15890,N_15658,N_15705);
xnor U15891 (N_15891,N_15565,N_15669);
xor U15892 (N_15892,N_15503,N_15555);
nand U15893 (N_15893,N_15642,N_15721);
nor U15894 (N_15894,N_15500,N_15559);
xor U15895 (N_15895,N_15732,N_15694);
or U15896 (N_15896,N_15641,N_15538);
nand U15897 (N_15897,N_15734,N_15626);
or U15898 (N_15898,N_15521,N_15681);
xnor U15899 (N_15899,N_15550,N_15630);
and U15900 (N_15900,N_15618,N_15654);
nand U15901 (N_15901,N_15714,N_15721);
and U15902 (N_15902,N_15726,N_15531);
or U15903 (N_15903,N_15537,N_15714);
nand U15904 (N_15904,N_15735,N_15699);
xnor U15905 (N_15905,N_15567,N_15668);
or U15906 (N_15906,N_15673,N_15654);
nand U15907 (N_15907,N_15560,N_15692);
and U15908 (N_15908,N_15708,N_15573);
or U15909 (N_15909,N_15656,N_15541);
nor U15910 (N_15910,N_15678,N_15746);
or U15911 (N_15911,N_15672,N_15614);
or U15912 (N_15912,N_15634,N_15731);
and U15913 (N_15913,N_15588,N_15670);
and U15914 (N_15914,N_15581,N_15556);
xnor U15915 (N_15915,N_15559,N_15539);
xnor U15916 (N_15916,N_15556,N_15739);
nor U15917 (N_15917,N_15703,N_15687);
nor U15918 (N_15918,N_15523,N_15502);
nor U15919 (N_15919,N_15730,N_15671);
nand U15920 (N_15920,N_15529,N_15699);
or U15921 (N_15921,N_15571,N_15700);
or U15922 (N_15922,N_15690,N_15596);
xor U15923 (N_15923,N_15581,N_15680);
nor U15924 (N_15924,N_15691,N_15578);
nor U15925 (N_15925,N_15690,N_15641);
or U15926 (N_15926,N_15671,N_15578);
nand U15927 (N_15927,N_15598,N_15667);
nor U15928 (N_15928,N_15681,N_15625);
xnor U15929 (N_15929,N_15530,N_15726);
nor U15930 (N_15930,N_15612,N_15710);
nor U15931 (N_15931,N_15507,N_15718);
or U15932 (N_15932,N_15655,N_15513);
nand U15933 (N_15933,N_15555,N_15697);
and U15934 (N_15934,N_15621,N_15598);
and U15935 (N_15935,N_15670,N_15507);
xor U15936 (N_15936,N_15630,N_15627);
or U15937 (N_15937,N_15650,N_15638);
xnor U15938 (N_15938,N_15596,N_15602);
xor U15939 (N_15939,N_15628,N_15568);
or U15940 (N_15940,N_15508,N_15706);
nand U15941 (N_15941,N_15530,N_15534);
or U15942 (N_15942,N_15504,N_15656);
nor U15943 (N_15943,N_15722,N_15689);
xor U15944 (N_15944,N_15581,N_15726);
and U15945 (N_15945,N_15630,N_15738);
xnor U15946 (N_15946,N_15510,N_15561);
or U15947 (N_15947,N_15513,N_15582);
nor U15948 (N_15948,N_15599,N_15675);
or U15949 (N_15949,N_15658,N_15594);
and U15950 (N_15950,N_15723,N_15694);
and U15951 (N_15951,N_15572,N_15744);
or U15952 (N_15952,N_15684,N_15735);
and U15953 (N_15953,N_15589,N_15743);
nor U15954 (N_15954,N_15577,N_15683);
nor U15955 (N_15955,N_15642,N_15545);
or U15956 (N_15956,N_15588,N_15575);
or U15957 (N_15957,N_15652,N_15604);
xnor U15958 (N_15958,N_15516,N_15670);
and U15959 (N_15959,N_15548,N_15612);
and U15960 (N_15960,N_15614,N_15536);
and U15961 (N_15961,N_15650,N_15677);
xnor U15962 (N_15962,N_15719,N_15685);
nor U15963 (N_15963,N_15670,N_15613);
or U15964 (N_15964,N_15623,N_15502);
or U15965 (N_15965,N_15507,N_15553);
nand U15966 (N_15966,N_15554,N_15644);
nor U15967 (N_15967,N_15747,N_15741);
nand U15968 (N_15968,N_15502,N_15576);
and U15969 (N_15969,N_15665,N_15748);
nor U15970 (N_15970,N_15607,N_15600);
or U15971 (N_15971,N_15666,N_15648);
nor U15972 (N_15972,N_15632,N_15707);
nor U15973 (N_15973,N_15552,N_15682);
and U15974 (N_15974,N_15510,N_15575);
nand U15975 (N_15975,N_15537,N_15672);
or U15976 (N_15976,N_15558,N_15510);
nor U15977 (N_15977,N_15676,N_15728);
xor U15978 (N_15978,N_15735,N_15742);
or U15979 (N_15979,N_15580,N_15597);
and U15980 (N_15980,N_15697,N_15602);
and U15981 (N_15981,N_15606,N_15558);
nor U15982 (N_15982,N_15570,N_15633);
and U15983 (N_15983,N_15729,N_15682);
or U15984 (N_15984,N_15545,N_15633);
and U15985 (N_15985,N_15630,N_15604);
and U15986 (N_15986,N_15541,N_15748);
nand U15987 (N_15987,N_15654,N_15634);
nand U15988 (N_15988,N_15727,N_15617);
xor U15989 (N_15989,N_15736,N_15734);
xor U15990 (N_15990,N_15656,N_15604);
and U15991 (N_15991,N_15633,N_15548);
or U15992 (N_15992,N_15661,N_15646);
xor U15993 (N_15993,N_15512,N_15622);
nand U15994 (N_15994,N_15659,N_15601);
nor U15995 (N_15995,N_15679,N_15518);
nand U15996 (N_15996,N_15690,N_15739);
nand U15997 (N_15997,N_15699,N_15533);
nand U15998 (N_15998,N_15553,N_15721);
or U15999 (N_15999,N_15626,N_15572);
xnor U16000 (N_16000,N_15795,N_15962);
nand U16001 (N_16001,N_15882,N_15838);
nor U16002 (N_16002,N_15863,N_15868);
and U16003 (N_16003,N_15827,N_15821);
nand U16004 (N_16004,N_15818,N_15981);
and U16005 (N_16005,N_15770,N_15820);
and U16006 (N_16006,N_15757,N_15831);
nor U16007 (N_16007,N_15855,N_15991);
xor U16008 (N_16008,N_15799,N_15925);
and U16009 (N_16009,N_15853,N_15811);
or U16010 (N_16010,N_15850,N_15994);
xnor U16011 (N_16011,N_15780,N_15928);
or U16012 (N_16012,N_15946,N_15963);
nand U16013 (N_16013,N_15935,N_15776);
and U16014 (N_16014,N_15901,N_15913);
and U16015 (N_16015,N_15889,N_15950);
and U16016 (N_16016,N_15974,N_15986);
nor U16017 (N_16017,N_15971,N_15816);
or U16018 (N_16018,N_15980,N_15947);
nand U16019 (N_16019,N_15989,N_15835);
nand U16020 (N_16020,N_15752,N_15807);
xor U16021 (N_16021,N_15937,N_15839);
or U16022 (N_16022,N_15871,N_15824);
or U16023 (N_16023,N_15990,N_15765);
and U16024 (N_16024,N_15886,N_15829);
and U16025 (N_16025,N_15786,N_15953);
or U16026 (N_16026,N_15851,N_15885);
and U16027 (N_16027,N_15764,N_15781);
or U16028 (N_16028,N_15905,N_15970);
and U16029 (N_16029,N_15858,N_15761);
nand U16030 (N_16030,N_15856,N_15783);
and U16031 (N_16031,N_15862,N_15973);
nor U16032 (N_16032,N_15967,N_15857);
and U16033 (N_16033,N_15959,N_15791);
xnor U16034 (N_16034,N_15903,N_15992);
nor U16035 (N_16035,N_15792,N_15773);
nand U16036 (N_16036,N_15812,N_15993);
or U16037 (N_16037,N_15750,N_15978);
nand U16038 (N_16038,N_15859,N_15785);
and U16039 (N_16039,N_15880,N_15830);
nor U16040 (N_16040,N_15846,N_15890);
xnor U16041 (N_16041,N_15883,N_15975);
nor U16042 (N_16042,N_15922,N_15768);
nand U16043 (N_16043,N_15904,N_15976);
xnor U16044 (N_16044,N_15865,N_15819);
nor U16045 (N_16045,N_15805,N_15794);
and U16046 (N_16046,N_15837,N_15879);
nor U16047 (N_16047,N_15930,N_15876);
nor U16048 (N_16048,N_15877,N_15775);
nand U16049 (N_16049,N_15808,N_15849);
nor U16050 (N_16050,N_15996,N_15875);
xnor U16051 (N_16051,N_15893,N_15860);
xor U16052 (N_16052,N_15809,N_15919);
xnor U16053 (N_16053,N_15822,N_15940);
and U16054 (N_16054,N_15798,N_15836);
or U16055 (N_16055,N_15949,N_15756);
nand U16056 (N_16056,N_15987,N_15977);
nor U16057 (N_16057,N_15834,N_15958);
nor U16058 (N_16058,N_15934,N_15972);
and U16059 (N_16059,N_15910,N_15844);
or U16060 (N_16060,N_15870,N_15897);
nor U16061 (N_16061,N_15938,N_15810);
nand U16062 (N_16062,N_15888,N_15823);
or U16063 (N_16063,N_15840,N_15793);
nand U16064 (N_16064,N_15833,N_15997);
nand U16065 (N_16065,N_15847,N_15891);
nor U16066 (N_16066,N_15814,N_15941);
or U16067 (N_16067,N_15927,N_15983);
and U16068 (N_16068,N_15912,N_15936);
and U16069 (N_16069,N_15804,N_15926);
nand U16070 (N_16070,N_15777,N_15796);
xnor U16071 (N_16071,N_15920,N_15769);
nor U16072 (N_16072,N_15921,N_15852);
and U16073 (N_16073,N_15828,N_15755);
nand U16074 (N_16074,N_15861,N_15762);
or U16075 (N_16075,N_15969,N_15841);
and U16076 (N_16076,N_15968,N_15939);
or U16077 (N_16077,N_15867,N_15918);
nor U16078 (N_16078,N_15767,N_15894);
xor U16079 (N_16079,N_15874,N_15848);
xnor U16080 (N_16080,N_15909,N_15943);
nand U16081 (N_16081,N_15806,N_15944);
or U16082 (N_16082,N_15782,N_15933);
nor U16083 (N_16083,N_15758,N_15982);
nand U16084 (N_16084,N_15759,N_15908);
xor U16085 (N_16085,N_15900,N_15952);
or U16086 (N_16086,N_15789,N_15898);
nand U16087 (N_16087,N_15787,N_15788);
xnor U16088 (N_16088,N_15988,N_15774);
nand U16089 (N_16089,N_15881,N_15896);
nor U16090 (N_16090,N_15966,N_15832);
or U16091 (N_16091,N_15801,N_15914);
nor U16092 (N_16092,N_15948,N_15955);
or U16093 (N_16093,N_15779,N_15778);
xnor U16094 (N_16094,N_15895,N_15817);
and U16095 (N_16095,N_15979,N_15751);
nand U16096 (N_16096,N_15924,N_15771);
nand U16097 (N_16097,N_15956,N_15866);
nor U16098 (N_16098,N_15999,N_15873);
nand U16099 (N_16099,N_15864,N_15916);
xor U16100 (N_16100,N_15984,N_15842);
nor U16101 (N_16101,N_15887,N_15878);
nand U16102 (N_16102,N_15872,N_15964);
and U16103 (N_16103,N_15854,N_15985);
nand U16104 (N_16104,N_15825,N_15826);
and U16105 (N_16105,N_15954,N_15965);
or U16106 (N_16106,N_15957,N_15766);
or U16107 (N_16107,N_15803,N_15760);
xor U16108 (N_16108,N_15763,N_15754);
nor U16109 (N_16109,N_15784,N_15869);
and U16110 (N_16110,N_15800,N_15961);
or U16111 (N_16111,N_15945,N_15911);
nand U16112 (N_16112,N_15995,N_15892);
or U16113 (N_16113,N_15998,N_15931);
nor U16114 (N_16114,N_15902,N_15884);
or U16115 (N_16115,N_15917,N_15797);
nand U16116 (N_16116,N_15815,N_15951);
or U16117 (N_16117,N_15960,N_15942);
xor U16118 (N_16118,N_15906,N_15843);
or U16119 (N_16119,N_15772,N_15929);
nor U16120 (N_16120,N_15915,N_15932);
and U16121 (N_16121,N_15899,N_15802);
xnor U16122 (N_16122,N_15790,N_15907);
and U16123 (N_16123,N_15923,N_15753);
nand U16124 (N_16124,N_15845,N_15813);
or U16125 (N_16125,N_15970,N_15878);
or U16126 (N_16126,N_15842,N_15772);
or U16127 (N_16127,N_15878,N_15830);
and U16128 (N_16128,N_15792,N_15979);
xnor U16129 (N_16129,N_15840,N_15826);
nor U16130 (N_16130,N_15754,N_15978);
nand U16131 (N_16131,N_15810,N_15906);
or U16132 (N_16132,N_15752,N_15876);
nand U16133 (N_16133,N_15859,N_15793);
xnor U16134 (N_16134,N_15931,N_15934);
xor U16135 (N_16135,N_15875,N_15978);
and U16136 (N_16136,N_15978,N_15973);
nor U16137 (N_16137,N_15821,N_15937);
xor U16138 (N_16138,N_15928,N_15950);
and U16139 (N_16139,N_15866,N_15926);
and U16140 (N_16140,N_15861,N_15885);
and U16141 (N_16141,N_15896,N_15939);
or U16142 (N_16142,N_15910,N_15761);
nor U16143 (N_16143,N_15837,N_15934);
and U16144 (N_16144,N_15928,N_15776);
nor U16145 (N_16145,N_15802,N_15904);
xnor U16146 (N_16146,N_15931,N_15762);
and U16147 (N_16147,N_15924,N_15896);
xor U16148 (N_16148,N_15970,N_15898);
xnor U16149 (N_16149,N_15997,N_15879);
nand U16150 (N_16150,N_15817,N_15981);
and U16151 (N_16151,N_15811,N_15918);
or U16152 (N_16152,N_15869,N_15863);
nand U16153 (N_16153,N_15983,N_15765);
and U16154 (N_16154,N_15918,N_15885);
and U16155 (N_16155,N_15919,N_15948);
nand U16156 (N_16156,N_15807,N_15909);
nor U16157 (N_16157,N_15942,N_15948);
xor U16158 (N_16158,N_15877,N_15807);
xnor U16159 (N_16159,N_15836,N_15940);
nor U16160 (N_16160,N_15861,N_15803);
nand U16161 (N_16161,N_15772,N_15830);
and U16162 (N_16162,N_15831,N_15948);
nand U16163 (N_16163,N_15821,N_15976);
xor U16164 (N_16164,N_15785,N_15820);
nand U16165 (N_16165,N_15937,N_15771);
nor U16166 (N_16166,N_15974,N_15998);
xnor U16167 (N_16167,N_15878,N_15966);
nand U16168 (N_16168,N_15848,N_15937);
nor U16169 (N_16169,N_15982,N_15766);
and U16170 (N_16170,N_15885,N_15984);
or U16171 (N_16171,N_15928,N_15953);
or U16172 (N_16172,N_15780,N_15952);
xor U16173 (N_16173,N_15920,N_15869);
and U16174 (N_16174,N_15927,N_15820);
and U16175 (N_16175,N_15827,N_15842);
or U16176 (N_16176,N_15885,N_15824);
or U16177 (N_16177,N_15969,N_15979);
nor U16178 (N_16178,N_15765,N_15836);
nor U16179 (N_16179,N_15843,N_15851);
or U16180 (N_16180,N_15880,N_15990);
nor U16181 (N_16181,N_15783,N_15767);
nor U16182 (N_16182,N_15898,N_15823);
nor U16183 (N_16183,N_15911,N_15963);
and U16184 (N_16184,N_15754,N_15872);
or U16185 (N_16185,N_15751,N_15982);
and U16186 (N_16186,N_15991,N_15851);
xnor U16187 (N_16187,N_15826,N_15938);
or U16188 (N_16188,N_15817,N_15795);
xor U16189 (N_16189,N_15917,N_15936);
and U16190 (N_16190,N_15994,N_15807);
nor U16191 (N_16191,N_15903,N_15877);
xnor U16192 (N_16192,N_15813,N_15777);
nor U16193 (N_16193,N_15820,N_15963);
or U16194 (N_16194,N_15760,N_15786);
xnor U16195 (N_16195,N_15984,N_15835);
nor U16196 (N_16196,N_15975,N_15811);
nor U16197 (N_16197,N_15806,N_15950);
nor U16198 (N_16198,N_15920,N_15761);
nand U16199 (N_16199,N_15975,N_15935);
or U16200 (N_16200,N_15777,N_15821);
nor U16201 (N_16201,N_15801,N_15859);
nor U16202 (N_16202,N_15992,N_15801);
or U16203 (N_16203,N_15896,N_15801);
nor U16204 (N_16204,N_15867,N_15869);
nand U16205 (N_16205,N_15818,N_15871);
nor U16206 (N_16206,N_15770,N_15760);
xnor U16207 (N_16207,N_15862,N_15969);
xor U16208 (N_16208,N_15826,N_15783);
and U16209 (N_16209,N_15931,N_15777);
or U16210 (N_16210,N_15753,N_15841);
or U16211 (N_16211,N_15825,N_15882);
nor U16212 (N_16212,N_15779,N_15990);
nor U16213 (N_16213,N_15948,N_15863);
or U16214 (N_16214,N_15983,N_15777);
and U16215 (N_16215,N_15985,N_15922);
xnor U16216 (N_16216,N_15950,N_15910);
xnor U16217 (N_16217,N_15909,N_15820);
xnor U16218 (N_16218,N_15903,N_15801);
xor U16219 (N_16219,N_15790,N_15999);
xor U16220 (N_16220,N_15795,N_15874);
nand U16221 (N_16221,N_15820,N_15797);
or U16222 (N_16222,N_15887,N_15925);
nand U16223 (N_16223,N_15873,N_15806);
or U16224 (N_16224,N_15859,N_15950);
xnor U16225 (N_16225,N_15762,N_15949);
xor U16226 (N_16226,N_15827,N_15811);
and U16227 (N_16227,N_15881,N_15811);
nand U16228 (N_16228,N_15832,N_15836);
xnor U16229 (N_16229,N_15755,N_15832);
nor U16230 (N_16230,N_15998,N_15868);
nor U16231 (N_16231,N_15781,N_15770);
xnor U16232 (N_16232,N_15965,N_15885);
nand U16233 (N_16233,N_15910,N_15906);
nand U16234 (N_16234,N_15927,N_15839);
xor U16235 (N_16235,N_15974,N_15988);
and U16236 (N_16236,N_15908,N_15857);
nand U16237 (N_16237,N_15977,N_15787);
or U16238 (N_16238,N_15770,N_15946);
nand U16239 (N_16239,N_15978,N_15876);
or U16240 (N_16240,N_15938,N_15815);
xor U16241 (N_16241,N_15980,N_15983);
nor U16242 (N_16242,N_15939,N_15785);
nand U16243 (N_16243,N_15890,N_15948);
and U16244 (N_16244,N_15822,N_15816);
or U16245 (N_16245,N_15971,N_15808);
nor U16246 (N_16246,N_15774,N_15902);
and U16247 (N_16247,N_15851,N_15990);
nor U16248 (N_16248,N_15989,N_15961);
nor U16249 (N_16249,N_15857,N_15919);
and U16250 (N_16250,N_16027,N_16029);
nor U16251 (N_16251,N_16100,N_16043);
and U16252 (N_16252,N_16007,N_16168);
nand U16253 (N_16253,N_16159,N_16119);
nor U16254 (N_16254,N_16115,N_16012);
and U16255 (N_16255,N_16000,N_16062);
and U16256 (N_16256,N_16203,N_16073);
nor U16257 (N_16257,N_16191,N_16136);
and U16258 (N_16258,N_16145,N_16020);
nand U16259 (N_16259,N_16064,N_16197);
or U16260 (N_16260,N_16188,N_16044);
or U16261 (N_16261,N_16167,N_16211);
or U16262 (N_16262,N_16098,N_16139);
or U16263 (N_16263,N_16005,N_16118);
nor U16264 (N_16264,N_16134,N_16083);
or U16265 (N_16265,N_16017,N_16034);
or U16266 (N_16266,N_16143,N_16013);
nor U16267 (N_16267,N_16156,N_16111);
nor U16268 (N_16268,N_16063,N_16080);
nor U16269 (N_16269,N_16117,N_16028);
nor U16270 (N_16270,N_16233,N_16165);
nand U16271 (N_16271,N_16045,N_16190);
or U16272 (N_16272,N_16201,N_16177);
xnor U16273 (N_16273,N_16133,N_16169);
xor U16274 (N_16274,N_16171,N_16040);
xor U16275 (N_16275,N_16014,N_16228);
or U16276 (N_16276,N_16230,N_16052);
nand U16277 (N_16277,N_16222,N_16079);
or U16278 (N_16278,N_16137,N_16086);
or U16279 (N_16279,N_16219,N_16008);
or U16280 (N_16280,N_16113,N_16204);
or U16281 (N_16281,N_16002,N_16241);
nor U16282 (N_16282,N_16174,N_16009);
xnor U16283 (N_16283,N_16180,N_16221);
xor U16284 (N_16284,N_16006,N_16061);
nor U16285 (N_16285,N_16185,N_16108);
xor U16286 (N_16286,N_16172,N_16106);
and U16287 (N_16287,N_16128,N_16198);
and U16288 (N_16288,N_16181,N_16056);
and U16289 (N_16289,N_16032,N_16011);
nor U16290 (N_16290,N_16127,N_16076);
nor U16291 (N_16291,N_16199,N_16232);
and U16292 (N_16292,N_16166,N_16178);
xnor U16293 (N_16293,N_16231,N_16109);
nor U16294 (N_16294,N_16060,N_16225);
nand U16295 (N_16295,N_16025,N_16140);
nand U16296 (N_16296,N_16175,N_16132);
nand U16297 (N_16297,N_16154,N_16249);
and U16298 (N_16298,N_16068,N_16024);
or U16299 (N_16299,N_16092,N_16051);
xor U16300 (N_16300,N_16224,N_16066);
and U16301 (N_16301,N_16164,N_16196);
and U16302 (N_16302,N_16081,N_16200);
or U16303 (N_16303,N_16184,N_16220);
or U16304 (N_16304,N_16194,N_16049);
nand U16305 (N_16305,N_16215,N_16202);
nand U16306 (N_16306,N_16142,N_16094);
nand U16307 (N_16307,N_16039,N_16138);
nor U16308 (N_16308,N_16170,N_16097);
xnor U16309 (N_16309,N_16212,N_16223);
and U16310 (N_16310,N_16041,N_16089);
and U16311 (N_16311,N_16072,N_16207);
or U16312 (N_16312,N_16157,N_16120);
or U16313 (N_16313,N_16019,N_16144);
nand U16314 (N_16314,N_16016,N_16148);
nor U16315 (N_16315,N_16248,N_16004);
xor U16316 (N_16316,N_16218,N_16090);
xor U16317 (N_16317,N_16071,N_16242);
xnor U16318 (N_16318,N_16240,N_16229);
nand U16319 (N_16319,N_16161,N_16130);
nor U16320 (N_16320,N_16046,N_16114);
or U16321 (N_16321,N_16216,N_16077);
nand U16322 (N_16322,N_16050,N_16176);
xor U16323 (N_16323,N_16226,N_16037);
nor U16324 (N_16324,N_16234,N_16010);
nor U16325 (N_16325,N_16205,N_16055);
nand U16326 (N_16326,N_16206,N_16182);
nor U16327 (N_16327,N_16179,N_16239);
xor U16328 (N_16328,N_16173,N_16151);
xnor U16329 (N_16329,N_16087,N_16163);
nor U16330 (N_16330,N_16131,N_16158);
nand U16331 (N_16331,N_16030,N_16186);
xor U16332 (N_16332,N_16074,N_16059);
nand U16333 (N_16333,N_16075,N_16147);
or U16334 (N_16334,N_16247,N_16053);
or U16335 (N_16335,N_16146,N_16112);
nor U16336 (N_16336,N_16069,N_16105);
xnor U16337 (N_16337,N_16036,N_16085);
or U16338 (N_16338,N_16195,N_16054);
nor U16339 (N_16339,N_16244,N_16135);
nor U16340 (N_16340,N_16217,N_16023);
or U16341 (N_16341,N_16235,N_16123);
nor U16342 (N_16342,N_16096,N_16018);
xnor U16343 (N_16343,N_16084,N_16057);
xor U16344 (N_16344,N_16088,N_16033);
nand U16345 (N_16345,N_16125,N_16035);
nor U16346 (N_16346,N_16124,N_16214);
or U16347 (N_16347,N_16107,N_16078);
nor U16348 (N_16348,N_16001,N_16091);
nand U16349 (N_16349,N_16149,N_16187);
and U16350 (N_16350,N_16038,N_16189);
or U16351 (N_16351,N_16110,N_16208);
and U16352 (N_16352,N_16237,N_16104);
nand U16353 (N_16353,N_16093,N_16129);
and U16354 (N_16354,N_16193,N_16238);
nor U16355 (N_16355,N_16015,N_16192);
nand U16356 (N_16356,N_16070,N_16003);
nor U16357 (N_16357,N_16152,N_16102);
nor U16358 (N_16358,N_16126,N_16243);
xor U16359 (N_16359,N_16183,N_16162);
or U16360 (N_16360,N_16141,N_16095);
or U16361 (N_16361,N_16021,N_16031);
nor U16362 (N_16362,N_16082,N_16103);
and U16363 (N_16363,N_16099,N_16042);
and U16364 (N_16364,N_16246,N_16121);
and U16365 (N_16365,N_16022,N_16160);
nand U16366 (N_16366,N_16210,N_16048);
xor U16367 (N_16367,N_16122,N_16101);
or U16368 (N_16368,N_16047,N_16209);
xnor U16369 (N_16369,N_16153,N_16067);
nand U16370 (N_16370,N_16065,N_16236);
or U16371 (N_16371,N_16213,N_16245);
and U16372 (N_16372,N_16150,N_16058);
and U16373 (N_16373,N_16227,N_16026);
nor U16374 (N_16374,N_16155,N_16116);
nand U16375 (N_16375,N_16234,N_16081);
or U16376 (N_16376,N_16142,N_16038);
nor U16377 (N_16377,N_16206,N_16219);
and U16378 (N_16378,N_16008,N_16073);
and U16379 (N_16379,N_16007,N_16031);
xnor U16380 (N_16380,N_16231,N_16178);
or U16381 (N_16381,N_16142,N_16015);
nand U16382 (N_16382,N_16002,N_16161);
or U16383 (N_16383,N_16227,N_16203);
and U16384 (N_16384,N_16249,N_16239);
and U16385 (N_16385,N_16094,N_16131);
nor U16386 (N_16386,N_16058,N_16181);
or U16387 (N_16387,N_16216,N_16132);
and U16388 (N_16388,N_16160,N_16115);
nor U16389 (N_16389,N_16120,N_16153);
nor U16390 (N_16390,N_16134,N_16241);
xnor U16391 (N_16391,N_16034,N_16163);
nor U16392 (N_16392,N_16102,N_16002);
xor U16393 (N_16393,N_16207,N_16003);
nor U16394 (N_16394,N_16148,N_16172);
xor U16395 (N_16395,N_16118,N_16094);
nor U16396 (N_16396,N_16220,N_16173);
xnor U16397 (N_16397,N_16032,N_16133);
nand U16398 (N_16398,N_16201,N_16073);
nor U16399 (N_16399,N_16210,N_16177);
xnor U16400 (N_16400,N_16072,N_16115);
xnor U16401 (N_16401,N_16127,N_16047);
nor U16402 (N_16402,N_16050,N_16056);
or U16403 (N_16403,N_16101,N_16008);
xor U16404 (N_16404,N_16029,N_16066);
nand U16405 (N_16405,N_16238,N_16127);
nand U16406 (N_16406,N_16120,N_16194);
nand U16407 (N_16407,N_16005,N_16223);
nand U16408 (N_16408,N_16234,N_16121);
nor U16409 (N_16409,N_16138,N_16185);
nand U16410 (N_16410,N_16061,N_16077);
and U16411 (N_16411,N_16211,N_16124);
xnor U16412 (N_16412,N_16177,N_16187);
xnor U16413 (N_16413,N_16031,N_16134);
or U16414 (N_16414,N_16036,N_16091);
nor U16415 (N_16415,N_16202,N_16001);
and U16416 (N_16416,N_16034,N_16190);
or U16417 (N_16417,N_16076,N_16072);
nor U16418 (N_16418,N_16114,N_16031);
or U16419 (N_16419,N_16248,N_16169);
and U16420 (N_16420,N_16143,N_16133);
or U16421 (N_16421,N_16019,N_16054);
and U16422 (N_16422,N_16037,N_16026);
nand U16423 (N_16423,N_16016,N_16178);
nor U16424 (N_16424,N_16238,N_16175);
and U16425 (N_16425,N_16154,N_16230);
or U16426 (N_16426,N_16162,N_16091);
and U16427 (N_16427,N_16179,N_16082);
and U16428 (N_16428,N_16013,N_16082);
nor U16429 (N_16429,N_16152,N_16132);
or U16430 (N_16430,N_16215,N_16142);
or U16431 (N_16431,N_16151,N_16138);
and U16432 (N_16432,N_16131,N_16223);
or U16433 (N_16433,N_16244,N_16205);
xor U16434 (N_16434,N_16199,N_16225);
and U16435 (N_16435,N_16196,N_16074);
or U16436 (N_16436,N_16058,N_16013);
or U16437 (N_16437,N_16011,N_16180);
and U16438 (N_16438,N_16224,N_16020);
nor U16439 (N_16439,N_16079,N_16009);
or U16440 (N_16440,N_16241,N_16223);
nand U16441 (N_16441,N_16183,N_16052);
xnor U16442 (N_16442,N_16036,N_16142);
and U16443 (N_16443,N_16109,N_16206);
and U16444 (N_16444,N_16068,N_16150);
and U16445 (N_16445,N_16144,N_16139);
xor U16446 (N_16446,N_16187,N_16091);
nand U16447 (N_16447,N_16201,N_16021);
nand U16448 (N_16448,N_16219,N_16180);
xor U16449 (N_16449,N_16053,N_16070);
nor U16450 (N_16450,N_16088,N_16144);
xor U16451 (N_16451,N_16228,N_16157);
and U16452 (N_16452,N_16209,N_16031);
xor U16453 (N_16453,N_16175,N_16037);
xnor U16454 (N_16454,N_16043,N_16151);
nand U16455 (N_16455,N_16220,N_16131);
and U16456 (N_16456,N_16218,N_16204);
nand U16457 (N_16457,N_16021,N_16192);
nand U16458 (N_16458,N_16133,N_16175);
nand U16459 (N_16459,N_16074,N_16199);
or U16460 (N_16460,N_16238,N_16182);
or U16461 (N_16461,N_16048,N_16092);
and U16462 (N_16462,N_16114,N_16166);
nand U16463 (N_16463,N_16031,N_16177);
nand U16464 (N_16464,N_16099,N_16034);
and U16465 (N_16465,N_16067,N_16229);
nor U16466 (N_16466,N_16051,N_16203);
nor U16467 (N_16467,N_16013,N_16050);
nor U16468 (N_16468,N_16165,N_16220);
xor U16469 (N_16469,N_16179,N_16222);
nand U16470 (N_16470,N_16008,N_16051);
xnor U16471 (N_16471,N_16178,N_16149);
and U16472 (N_16472,N_16117,N_16096);
and U16473 (N_16473,N_16179,N_16107);
nor U16474 (N_16474,N_16204,N_16239);
nand U16475 (N_16475,N_16158,N_16128);
or U16476 (N_16476,N_16237,N_16149);
nand U16477 (N_16477,N_16211,N_16084);
and U16478 (N_16478,N_16221,N_16121);
nand U16479 (N_16479,N_16136,N_16078);
or U16480 (N_16480,N_16071,N_16062);
and U16481 (N_16481,N_16245,N_16218);
nor U16482 (N_16482,N_16236,N_16020);
and U16483 (N_16483,N_16189,N_16222);
nand U16484 (N_16484,N_16100,N_16150);
nand U16485 (N_16485,N_16053,N_16003);
nand U16486 (N_16486,N_16076,N_16175);
or U16487 (N_16487,N_16189,N_16076);
nand U16488 (N_16488,N_16044,N_16164);
nand U16489 (N_16489,N_16084,N_16065);
nor U16490 (N_16490,N_16212,N_16203);
nor U16491 (N_16491,N_16160,N_16065);
nand U16492 (N_16492,N_16132,N_16191);
xnor U16493 (N_16493,N_16195,N_16190);
or U16494 (N_16494,N_16136,N_16086);
xnor U16495 (N_16495,N_16187,N_16136);
or U16496 (N_16496,N_16011,N_16064);
xor U16497 (N_16497,N_16200,N_16176);
xor U16498 (N_16498,N_16247,N_16120);
xor U16499 (N_16499,N_16167,N_16053);
and U16500 (N_16500,N_16421,N_16436);
xor U16501 (N_16501,N_16452,N_16416);
nor U16502 (N_16502,N_16438,N_16498);
xor U16503 (N_16503,N_16310,N_16256);
or U16504 (N_16504,N_16384,N_16311);
xnor U16505 (N_16505,N_16455,N_16497);
and U16506 (N_16506,N_16378,N_16426);
or U16507 (N_16507,N_16399,N_16465);
xnor U16508 (N_16508,N_16411,N_16295);
and U16509 (N_16509,N_16484,N_16440);
nand U16510 (N_16510,N_16451,N_16418);
or U16511 (N_16511,N_16284,N_16280);
and U16512 (N_16512,N_16406,N_16366);
nor U16513 (N_16513,N_16373,N_16352);
nor U16514 (N_16514,N_16315,N_16439);
and U16515 (N_16515,N_16359,N_16414);
nor U16516 (N_16516,N_16413,N_16273);
nand U16517 (N_16517,N_16463,N_16345);
nand U16518 (N_16518,N_16294,N_16492);
nand U16519 (N_16519,N_16347,N_16391);
xnor U16520 (N_16520,N_16475,N_16265);
nor U16521 (N_16521,N_16319,N_16410);
xnor U16522 (N_16522,N_16253,N_16389);
nor U16523 (N_16523,N_16376,N_16289);
and U16524 (N_16524,N_16478,N_16431);
and U16525 (N_16525,N_16393,N_16292);
nand U16526 (N_16526,N_16458,N_16488);
nor U16527 (N_16527,N_16453,N_16272);
xor U16528 (N_16528,N_16277,N_16403);
nor U16529 (N_16529,N_16472,N_16367);
xor U16530 (N_16530,N_16355,N_16344);
nor U16531 (N_16531,N_16369,N_16486);
nand U16532 (N_16532,N_16285,N_16258);
nand U16533 (N_16533,N_16398,N_16381);
nor U16534 (N_16534,N_16377,N_16473);
or U16535 (N_16535,N_16270,N_16288);
nand U16536 (N_16536,N_16457,N_16481);
and U16537 (N_16537,N_16379,N_16456);
xor U16538 (N_16538,N_16309,N_16263);
and U16539 (N_16539,N_16477,N_16420);
nand U16540 (N_16540,N_16482,N_16314);
nor U16541 (N_16541,N_16450,N_16323);
or U16542 (N_16542,N_16428,N_16474);
and U16543 (N_16543,N_16363,N_16286);
nand U16544 (N_16544,N_16464,N_16491);
xor U16545 (N_16545,N_16275,N_16358);
nand U16546 (N_16546,N_16490,N_16330);
nor U16547 (N_16547,N_16297,N_16301);
xnor U16548 (N_16548,N_16415,N_16307);
xor U16549 (N_16549,N_16287,N_16268);
or U16550 (N_16550,N_16448,N_16365);
nand U16551 (N_16551,N_16326,N_16437);
nor U16552 (N_16552,N_16255,N_16350);
or U16553 (N_16553,N_16296,N_16282);
nand U16554 (N_16554,N_16269,N_16495);
nand U16555 (N_16555,N_16308,N_16400);
or U16556 (N_16556,N_16254,N_16349);
nand U16557 (N_16557,N_16338,N_16290);
nand U16558 (N_16558,N_16383,N_16252);
xor U16559 (N_16559,N_16250,N_16298);
and U16560 (N_16560,N_16405,N_16329);
xnor U16561 (N_16561,N_16435,N_16446);
and U16562 (N_16562,N_16317,N_16407);
and U16563 (N_16563,N_16479,N_16404);
nand U16564 (N_16564,N_16336,N_16499);
nor U16565 (N_16565,N_16483,N_16466);
and U16566 (N_16566,N_16362,N_16444);
and U16567 (N_16567,N_16274,N_16493);
or U16568 (N_16568,N_16434,N_16401);
nor U16569 (N_16569,N_16364,N_16468);
and U16570 (N_16570,N_16300,N_16412);
xnor U16571 (N_16571,N_16306,N_16348);
nand U16572 (N_16572,N_16324,N_16433);
nor U16573 (N_16573,N_16283,N_16331);
or U16574 (N_16574,N_16343,N_16467);
xnor U16575 (N_16575,N_16494,N_16312);
xnor U16576 (N_16576,N_16386,N_16341);
nand U16577 (N_16577,N_16346,N_16432);
nand U16578 (N_16578,N_16469,N_16325);
nand U16579 (N_16579,N_16271,N_16470);
and U16580 (N_16580,N_16264,N_16356);
nor U16581 (N_16581,N_16302,N_16380);
nor U16582 (N_16582,N_16460,N_16441);
nand U16583 (N_16583,N_16368,N_16257);
or U16584 (N_16584,N_16396,N_16462);
nor U16585 (N_16585,N_16388,N_16417);
and U16586 (N_16586,N_16332,N_16423);
or U16587 (N_16587,N_16392,N_16461);
xor U16588 (N_16588,N_16370,N_16279);
nand U16589 (N_16589,N_16454,N_16335);
or U16590 (N_16590,N_16328,N_16259);
nor U16591 (N_16591,N_16291,N_16459);
nand U16592 (N_16592,N_16442,N_16471);
or U16593 (N_16593,N_16251,N_16327);
xnor U16594 (N_16594,N_16267,N_16293);
nor U16595 (N_16595,N_16430,N_16374);
xor U16596 (N_16596,N_16419,N_16449);
and U16597 (N_16597,N_16402,N_16382);
and U16598 (N_16598,N_16337,N_16371);
nor U16599 (N_16599,N_16443,N_16360);
nor U16600 (N_16600,N_16260,N_16489);
nor U16601 (N_16601,N_16276,N_16333);
and U16602 (N_16602,N_16390,N_16357);
nor U16603 (N_16603,N_16429,N_16305);
nor U16604 (N_16604,N_16278,N_16375);
xnor U16605 (N_16605,N_16316,N_16487);
nor U16606 (N_16606,N_16409,N_16427);
nor U16607 (N_16607,N_16320,N_16422);
and U16608 (N_16608,N_16299,N_16340);
or U16609 (N_16609,N_16361,N_16281);
nand U16610 (N_16610,N_16321,N_16339);
and U16611 (N_16611,N_16262,N_16424);
and U16612 (N_16612,N_16397,N_16322);
or U16613 (N_16613,N_16445,N_16354);
xnor U16614 (N_16614,N_16480,N_16266);
nand U16615 (N_16615,N_16318,N_16342);
or U16616 (N_16616,N_16353,N_16408);
xor U16617 (N_16617,N_16447,N_16485);
nand U16618 (N_16618,N_16387,N_16496);
or U16619 (N_16619,N_16313,N_16303);
nand U16620 (N_16620,N_16425,N_16385);
and U16621 (N_16621,N_16261,N_16351);
and U16622 (N_16622,N_16394,N_16476);
nor U16623 (N_16623,N_16304,N_16372);
nor U16624 (N_16624,N_16334,N_16395);
and U16625 (N_16625,N_16314,N_16387);
or U16626 (N_16626,N_16347,N_16421);
or U16627 (N_16627,N_16381,N_16361);
nor U16628 (N_16628,N_16260,N_16454);
or U16629 (N_16629,N_16486,N_16252);
and U16630 (N_16630,N_16292,N_16437);
nand U16631 (N_16631,N_16276,N_16363);
and U16632 (N_16632,N_16406,N_16265);
xor U16633 (N_16633,N_16470,N_16309);
nor U16634 (N_16634,N_16463,N_16276);
xor U16635 (N_16635,N_16463,N_16437);
nand U16636 (N_16636,N_16354,N_16367);
xnor U16637 (N_16637,N_16328,N_16470);
xor U16638 (N_16638,N_16490,N_16273);
and U16639 (N_16639,N_16300,N_16266);
nand U16640 (N_16640,N_16483,N_16469);
nor U16641 (N_16641,N_16392,N_16266);
and U16642 (N_16642,N_16394,N_16405);
xnor U16643 (N_16643,N_16292,N_16352);
nor U16644 (N_16644,N_16319,N_16255);
or U16645 (N_16645,N_16279,N_16254);
or U16646 (N_16646,N_16278,N_16269);
nand U16647 (N_16647,N_16362,N_16395);
or U16648 (N_16648,N_16464,N_16420);
nor U16649 (N_16649,N_16383,N_16475);
nor U16650 (N_16650,N_16464,N_16281);
nor U16651 (N_16651,N_16268,N_16475);
and U16652 (N_16652,N_16480,N_16332);
and U16653 (N_16653,N_16368,N_16376);
or U16654 (N_16654,N_16479,N_16396);
nor U16655 (N_16655,N_16489,N_16252);
and U16656 (N_16656,N_16271,N_16413);
or U16657 (N_16657,N_16355,N_16457);
or U16658 (N_16658,N_16442,N_16322);
or U16659 (N_16659,N_16323,N_16352);
and U16660 (N_16660,N_16415,N_16437);
xor U16661 (N_16661,N_16492,N_16339);
or U16662 (N_16662,N_16339,N_16310);
nand U16663 (N_16663,N_16425,N_16414);
and U16664 (N_16664,N_16411,N_16441);
nand U16665 (N_16665,N_16451,N_16496);
nand U16666 (N_16666,N_16324,N_16269);
and U16667 (N_16667,N_16253,N_16411);
xnor U16668 (N_16668,N_16304,N_16343);
nor U16669 (N_16669,N_16331,N_16318);
xor U16670 (N_16670,N_16335,N_16386);
nor U16671 (N_16671,N_16383,N_16404);
nand U16672 (N_16672,N_16313,N_16419);
nand U16673 (N_16673,N_16292,N_16439);
and U16674 (N_16674,N_16433,N_16264);
nor U16675 (N_16675,N_16374,N_16440);
xnor U16676 (N_16676,N_16393,N_16269);
and U16677 (N_16677,N_16395,N_16498);
xor U16678 (N_16678,N_16349,N_16260);
and U16679 (N_16679,N_16314,N_16363);
nand U16680 (N_16680,N_16358,N_16337);
xnor U16681 (N_16681,N_16257,N_16454);
xnor U16682 (N_16682,N_16382,N_16360);
xnor U16683 (N_16683,N_16471,N_16324);
nand U16684 (N_16684,N_16411,N_16261);
and U16685 (N_16685,N_16385,N_16376);
or U16686 (N_16686,N_16490,N_16282);
or U16687 (N_16687,N_16397,N_16254);
or U16688 (N_16688,N_16412,N_16457);
nor U16689 (N_16689,N_16272,N_16489);
nor U16690 (N_16690,N_16272,N_16348);
nand U16691 (N_16691,N_16254,N_16263);
nor U16692 (N_16692,N_16318,N_16293);
xnor U16693 (N_16693,N_16369,N_16495);
xor U16694 (N_16694,N_16284,N_16441);
xor U16695 (N_16695,N_16495,N_16318);
and U16696 (N_16696,N_16325,N_16464);
xnor U16697 (N_16697,N_16444,N_16483);
xnor U16698 (N_16698,N_16359,N_16319);
and U16699 (N_16699,N_16466,N_16343);
nor U16700 (N_16700,N_16496,N_16407);
xnor U16701 (N_16701,N_16309,N_16252);
xor U16702 (N_16702,N_16377,N_16443);
nor U16703 (N_16703,N_16392,N_16314);
and U16704 (N_16704,N_16462,N_16271);
xnor U16705 (N_16705,N_16270,N_16463);
nand U16706 (N_16706,N_16498,N_16436);
or U16707 (N_16707,N_16317,N_16303);
and U16708 (N_16708,N_16269,N_16494);
xor U16709 (N_16709,N_16493,N_16400);
and U16710 (N_16710,N_16478,N_16493);
xor U16711 (N_16711,N_16311,N_16309);
nor U16712 (N_16712,N_16332,N_16355);
or U16713 (N_16713,N_16254,N_16251);
and U16714 (N_16714,N_16389,N_16420);
and U16715 (N_16715,N_16326,N_16383);
nor U16716 (N_16716,N_16263,N_16440);
nor U16717 (N_16717,N_16413,N_16442);
nor U16718 (N_16718,N_16464,N_16374);
nand U16719 (N_16719,N_16454,N_16409);
or U16720 (N_16720,N_16491,N_16263);
nor U16721 (N_16721,N_16468,N_16286);
and U16722 (N_16722,N_16461,N_16424);
nor U16723 (N_16723,N_16292,N_16396);
xor U16724 (N_16724,N_16294,N_16297);
nor U16725 (N_16725,N_16326,N_16281);
nor U16726 (N_16726,N_16421,N_16309);
xor U16727 (N_16727,N_16446,N_16402);
nor U16728 (N_16728,N_16437,N_16390);
or U16729 (N_16729,N_16366,N_16487);
nand U16730 (N_16730,N_16437,N_16479);
nor U16731 (N_16731,N_16447,N_16365);
and U16732 (N_16732,N_16450,N_16476);
xnor U16733 (N_16733,N_16400,N_16371);
or U16734 (N_16734,N_16407,N_16321);
and U16735 (N_16735,N_16421,N_16296);
and U16736 (N_16736,N_16452,N_16307);
nor U16737 (N_16737,N_16386,N_16374);
nor U16738 (N_16738,N_16250,N_16368);
or U16739 (N_16739,N_16456,N_16346);
nand U16740 (N_16740,N_16469,N_16390);
nor U16741 (N_16741,N_16472,N_16294);
or U16742 (N_16742,N_16358,N_16426);
or U16743 (N_16743,N_16357,N_16404);
xnor U16744 (N_16744,N_16347,N_16424);
nand U16745 (N_16745,N_16271,N_16302);
nand U16746 (N_16746,N_16449,N_16297);
nor U16747 (N_16747,N_16361,N_16252);
nand U16748 (N_16748,N_16267,N_16349);
or U16749 (N_16749,N_16413,N_16408);
nor U16750 (N_16750,N_16507,N_16682);
nand U16751 (N_16751,N_16544,N_16749);
and U16752 (N_16752,N_16596,N_16742);
nor U16753 (N_16753,N_16524,N_16611);
nor U16754 (N_16754,N_16741,N_16689);
or U16755 (N_16755,N_16565,N_16679);
xnor U16756 (N_16756,N_16558,N_16718);
nand U16757 (N_16757,N_16716,N_16663);
and U16758 (N_16758,N_16639,N_16502);
nor U16759 (N_16759,N_16549,N_16748);
and U16760 (N_16760,N_16560,N_16568);
nand U16761 (N_16761,N_16669,N_16736);
nand U16762 (N_16762,N_16548,N_16569);
nor U16763 (N_16763,N_16539,N_16523);
xor U16764 (N_16764,N_16729,N_16527);
or U16765 (N_16765,N_16661,N_16651);
nand U16766 (N_16766,N_16590,N_16747);
or U16767 (N_16767,N_16552,N_16723);
nand U16768 (N_16768,N_16583,N_16664);
or U16769 (N_16769,N_16694,N_16585);
and U16770 (N_16770,N_16619,N_16654);
or U16771 (N_16771,N_16739,N_16638);
and U16772 (N_16772,N_16719,N_16541);
xnor U16773 (N_16773,N_16600,N_16695);
xor U16774 (N_16774,N_16522,N_16599);
xor U16775 (N_16775,N_16563,N_16645);
xor U16776 (N_16776,N_16746,N_16530);
xor U16777 (N_16777,N_16637,N_16588);
or U16778 (N_16778,N_16531,N_16674);
nor U16779 (N_16779,N_16553,N_16697);
and U16780 (N_16780,N_16728,N_16510);
nand U16781 (N_16781,N_16618,N_16547);
nand U16782 (N_16782,N_16644,N_16567);
nand U16783 (N_16783,N_16575,N_16594);
nor U16784 (N_16784,N_16744,N_16589);
xnor U16785 (N_16785,N_16666,N_16528);
nand U16786 (N_16786,N_16630,N_16631);
nor U16787 (N_16787,N_16622,N_16655);
and U16788 (N_16788,N_16628,N_16701);
and U16789 (N_16789,N_16702,N_16572);
nand U16790 (N_16790,N_16658,N_16513);
and U16791 (N_16791,N_16705,N_16571);
nor U16792 (N_16792,N_16505,N_16721);
or U16793 (N_16793,N_16678,N_16598);
xor U16794 (N_16794,N_16681,N_16613);
nor U16795 (N_16795,N_16557,N_16667);
and U16796 (N_16796,N_16595,N_16508);
nor U16797 (N_16797,N_16672,N_16730);
xnor U16798 (N_16798,N_16545,N_16546);
or U16799 (N_16799,N_16511,N_16738);
nor U16800 (N_16800,N_16532,N_16727);
and U16801 (N_16801,N_16710,N_16625);
nand U16802 (N_16802,N_16709,N_16680);
and U16803 (N_16803,N_16616,N_16743);
nor U16804 (N_16804,N_16609,N_16538);
or U16805 (N_16805,N_16632,N_16602);
nor U16806 (N_16806,N_16706,N_16635);
or U16807 (N_16807,N_16647,N_16636);
xor U16808 (N_16808,N_16670,N_16501);
nand U16809 (N_16809,N_16684,N_16659);
and U16810 (N_16810,N_16521,N_16581);
and U16811 (N_16811,N_16686,N_16733);
and U16812 (N_16812,N_16580,N_16601);
and U16813 (N_16813,N_16506,N_16612);
nor U16814 (N_16814,N_16559,N_16693);
and U16815 (N_16815,N_16649,N_16641);
nand U16816 (N_16816,N_16561,N_16656);
nor U16817 (N_16817,N_16665,N_16592);
nor U16818 (N_16818,N_16725,N_16621);
or U16819 (N_16819,N_16711,N_16677);
nor U16820 (N_16820,N_16662,N_16717);
xnor U16821 (N_16821,N_16700,N_16518);
or U16822 (N_16822,N_16550,N_16608);
nor U16823 (N_16823,N_16629,N_16529);
xor U16824 (N_16824,N_16543,N_16564);
nor U16825 (N_16825,N_16503,N_16657);
nor U16826 (N_16826,N_16692,N_16675);
xnor U16827 (N_16827,N_16646,N_16615);
nor U16828 (N_16828,N_16626,N_16707);
and U16829 (N_16829,N_16703,N_16516);
and U16830 (N_16830,N_16542,N_16556);
or U16831 (N_16831,N_16708,N_16577);
nor U16832 (N_16832,N_16554,N_16734);
nor U16833 (N_16833,N_16597,N_16668);
and U16834 (N_16834,N_16555,N_16520);
xnor U16835 (N_16835,N_16606,N_16573);
or U16836 (N_16836,N_16525,N_16652);
and U16837 (N_16837,N_16737,N_16724);
nand U16838 (N_16838,N_16683,N_16740);
and U16839 (N_16839,N_16515,N_16673);
xor U16840 (N_16840,N_16610,N_16620);
xor U16841 (N_16841,N_16614,N_16648);
nor U16842 (N_16842,N_16704,N_16714);
nand U16843 (N_16843,N_16535,N_16690);
and U16844 (N_16844,N_16720,N_16688);
and U16845 (N_16845,N_16562,N_16514);
and U16846 (N_16846,N_16582,N_16698);
nor U16847 (N_16847,N_16526,N_16536);
and U16848 (N_16848,N_16603,N_16745);
or U16849 (N_16849,N_16533,N_16712);
xor U16850 (N_16850,N_16579,N_16537);
or U16851 (N_16851,N_16500,N_16591);
or U16852 (N_16852,N_16576,N_16570);
and U16853 (N_16853,N_16715,N_16691);
and U16854 (N_16854,N_16512,N_16699);
nand U16855 (N_16855,N_16584,N_16551);
and U16856 (N_16856,N_16650,N_16634);
nand U16857 (N_16857,N_16696,N_16633);
and U16858 (N_16858,N_16587,N_16726);
and U16859 (N_16859,N_16578,N_16713);
xor U16860 (N_16860,N_16517,N_16640);
or U16861 (N_16861,N_16593,N_16732);
nand U16862 (N_16862,N_16586,N_16605);
xor U16863 (N_16863,N_16735,N_16540);
xnor U16864 (N_16864,N_16627,N_16671);
and U16865 (N_16865,N_16624,N_16534);
and U16866 (N_16866,N_16722,N_16623);
or U16867 (N_16867,N_16685,N_16676);
and U16868 (N_16868,N_16519,N_16604);
nand U16869 (N_16869,N_16574,N_16617);
or U16870 (N_16870,N_16653,N_16642);
and U16871 (N_16871,N_16643,N_16504);
nand U16872 (N_16872,N_16509,N_16607);
nand U16873 (N_16873,N_16566,N_16660);
xnor U16874 (N_16874,N_16687,N_16731);
nor U16875 (N_16875,N_16518,N_16644);
xor U16876 (N_16876,N_16727,N_16681);
and U16877 (N_16877,N_16567,N_16540);
or U16878 (N_16878,N_16735,N_16618);
xnor U16879 (N_16879,N_16706,N_16674);
nand U16880 (N_16880,N_16630,N_16554);
xnor U16881 (N_16881,N_16720,N_16669);
and U16882 (N_16882,N_16689,N_16711);
nor U16883 (N_16883,N_16643,N_16530);
or U16884 (N_16884,N_16575,N_16645);
or U16885 (N_16885,N_16509,N_16533);
and U16886 (N_16886,N_16636,N_16651);
nand U16887 (N_16887,N_16614,N_16702);
xor U16888 (N_16888,N_16565,N_16627);
xnor U16889 (N_16889,N_16620,N_16687);
nor U16890 (N_16890,N_16667,N_16610);
nand U16891 (N_16891,N_16605,N_16741);
xnor U16892 (N_16892,N_16671,N_16673);
or U16893 (N_16893,N_16690,N_16526);
nor U16894 (N_16894,N_16568,N_16526);
xor U16895 (N_16895,N_16725,N_16690);
nand U16896 (N_16896,N_16534,N_16584);
nand U16897 (N_16897,N_16613,N_16733);
xor U16898 (N_16898,N_16662,N_16515);
and U16899 (N_16899,N_16551,N_16605);
nand U16900 (N_16900,N_16637,N_16556);
xor U16901 (N_16901,N_16714,N_16567);
nand U16902 (N_16902,N_16744,N_16730);
and U16903 (N_16903,N_16646,N_16621);
nand U16904 (N_16904,N_16547,N_16606);
nor U16905 (N_16905,N_16536,N_16530);
or U16906 (N_16906,N_16740,N_16730);
nor U16907 (N_16907,N_16642,N_16630);
or U16908 (N_16908,N_16671,N_16529);
xor U16909 (N_16909,N_16728,N_16726);
or U16910 (N_16910,N_16501,N_16619);
or U16911 (N_16911,N_16515,N_16668);
nand U16912 (N_16912,N_16650,N_16681);
nand U16913 (N_16913,N_16693,N_16696);
nor U16914 (N_16914,N_16649,N_16578);
and U16915 (N_16915,N_16697,N_16548);
and U16916 (N_16916,N_16716,N_16545);
and U16917 (N_16917,N_16560,N_16588);
or U16918 (N_16918,N_16502,N_16598);
nand U16919 (N_16919,N_16527,N_16628);
or U16920 (N_16920,N_16611,N_16724);
nor U16921 (N_16921,N_16563,N_16693);
nor U16922 (N_16922,N_16620,N_16674);
or U16923 (N_16923,N_16602,N_16578);
nor U16924 (N_16924,N_16548,N_16573);
nand U16925 (N_16925,N_16587,N_16549);
nor U16926 (N_16926,N_16562,N_16689);
nor U16927 (N_16927,N_16592,N_16512);
nor U16928 (N_16928,N_16513,N_16535);
and U16929 (N_16929,N_16682,N_16616);
or U16930 (N_16930,N_16642,N_16566);
nand U16931 (N_16931,N_16709,N_16612);
or U16932 (N_16932,N_16634,N_16598);
nand U16933 (N_16933,N_16625,N_16682);
nand U16934 (N_16934,N_16513,N_16590);
nor U16935 (N_16935,N_16602,N_16633);
or U16936 (N_16936,N_16604,N_16642);
and U16937 (N_16937,N_16641,N_16684);
xnor U16938 (N_16938,N_16672,N_16596);
nand U16939 (N_16939,N_16676,N_16517);
xnor U16940 (N_16940,N_16735,N_16665);
xnor U16941 (N_16941,N_16607,N_16672);
and U16942 (N_16942,N_16558,N_16600);
nor U16943 (N_16943,N_16686,N_16645);
nand U16944 (N_16944,N_16513,N_16659);
or U16945 (N_16945,N_16539,N_16615);
and U16946 (N_16946,N_16563,N_16551);
nor U16947 (N_16947,N_16741,N_16686);
nor U16948 (N_16948,N_16593,N_16540);
nand U16949 (N_16949,N_16634,N_16737);
nor U16950 (N_16950,N_16745,N_16669);
and U16951 (N_16951,N_16551,N_16673);
xnor U16952 (N_16952,N_16513,N_16533);
nand U16953 (N_16953,N_16701,N_16566);
nor U16954 (N_16954,N_16602,N_16542);
and U16955 (N_16955,N_16661,N_16579);
xor U16956 (N_16956,N_16657,N_16541);
and U16957 (N_16957,N_16685,N_16621);
and U16958 (N_16958,N_16505,N_16588);
nor U16959 (N_16959,N_16729,N_16664);
or U16960 (N_16960,N_16659,N_16545);
nor U16961 (N_16961,N_16692,N_16589);
nand U16962 (N_16962,N_16631,N_16619);
nand U16963 (N_16963,N_16565,N_16603);
nand U16964 (N_16964,N_16626,N_16698);
nor U16965 (N_16965,N_16622,N_16513);
nor U16966 (N_16966,N_16559,N_16519);
nor U16967 (N_16967,N_16605,N_16738);
nor U16968 (N_16968,N_16626,N_16617);
and U16969 (N_16969,N_16596,N_16603);
xor U16970 (N_16970,N_16525,N_16674);
or U16971 (N_16971,N_16609,N_16655);
nor U16972 (N_16972,N_16619,N_16553);
nand U16973 (N_16973,N_16522,N_16503);
nand U16974 (N_16974,N_16679,N_16671);
or U16975 (N_16975,N_16519,N_16732);
nor U16976 (N_16976,N_16746,N_16707);
or U16977 (N_16977,N_16547,N_16623);
nand U16978 (N_16978,N_16677,N_16582);
nor U16979 (N_16979,N_16695,N_16622);
or U16980 (N_16980,N_16519,N_16628);
and U16981 (N_16981,N_16716,N_16734);
and U16982 (N_16982,N_16551,N_16568);
nor U16983 (N_16983,N_16550,N_16595);
nor U16984 (N_16984,N_16636,N_16564);
nand U16985 (N_16985,N_16507,N_16630);
and U16986 (N_16986,N_16706,N_16531);
or U16987 (N_16987,N_16534,N_16620);
and U16988 (N_16988,N_16650,N_16577);
nor U16989 (N_16989,N_16538,N_16583);
nand U16990 (N_16990,N_16519,N_16537);
nor U16991 (N_16991,N_16655,N_16581);
xnor U16992 (N_16992,N_16531,N_16539);
and U16993 (N_16993,N_16564,N_16529);
xnor U16994 (N_16994,N_16523,N_16659);
xnor U16995 (N_16995,N_16668,N_16679);
nor U16996 (N_16996,N_16680,N_16565);
nand U16997 (N_16997,N_16660,N_16721);
nor U16998 (N_16998,N_16703,N_16579);
nand U16999 (N_16999,N_16504,N_16597);
or U17000 (N_17000,N_16932,N_16902);
and U17001 (N_17001,N_16883,N_16763);
nor U17002 (N_17002,N_16781,N_16813);
xnor U17003 (N_17003,N_16957,N_16821);
nor U17004 (N_17004,N_16916,N_16770);
or U17005 (N_17005,N_16989,N_16981);
and U17006 (N_17006,N_16839,N_16840);
xor U17007 (N_17007,N_16882,N_16992);
or U17008 (N_17008,N_16941,N_16944);
and U17009 (N_17009,N_16885,N_16884);
nand U17010 (N_17010,N_16983,N_16774);
or U17011 (N_17011,N_16999,N_16857);
xor U17012 (N_17012,N_16986,N_16845);
or U17013 (N_17013,N_16935,N_16893);
xnor U17014 (N_17014,N_16961,N_16812);
nand U17015 (N_17015,N_16755,N_16985);
xor U17016 (N_17016,N_16925,N_16933);
nand U17017 (N_17017,N_16834,N_16830);
or U17018 (N_17018,N_16759,N_16750);
nor U17019 (N_17019,N_16807,N_16841);
nor U17020 (N_17020,N_16888,N_16842);
nand U17021 (N_17021,N_16877,N_16822);
xor U17022 (N_17022,N_16849,N_16868);
nand U17023 (N_17023,N_16817,N_16936);
and U17024 (N_17024,N_16769,N_16804);
xor U17025 (N_17025,N_16931,N_16897);
xnor U17026 (N_17026,N_16905,N_16785);
xor U17027 (N_17027,N_16896,N_16790);
and U17028 (N_17028,N_16930,N_16901);
and U17029 (N_17029,N_16940,N_16850);
xnor U17030 (N_17030,N_16824,N_16838);
or U17031 (N_17031,N_16767,N_16778);
xnor U17032 (N_17032,N_16818,N_16918);
or U17033 (N_17033,N_16797,N_16972);
and U17034 (N_17034,N_16776,N_16870);
xnor U17035 (N_17035,N_16964,N_16793);
or U17036 (N_17036,N_16924,N_16831);
xnor U17037 (N_17037,N_16965,N_16805);
xnor U17038 (N_17038,N_16955,N_16779);
or U17039 (N_17039,N_16846,N_16996);
nand U17040 (N_17040,N_16786,N_16806);
or U17041 (N_17041,N_16894,N_16973);
xor U17042 (N_17042,N_16809,N_16851);
and U17043 (N_17043,N_16919,N_16907);
xnor U17044 (N_17044,N_16945,N_16802);
nor U17045 (N_17045,N_16795,N_16903);
and U17046 (N_17046,N_16867,N_16782);
nand U17047 (N_17047,N_16803,N_16967);
or U17048 (N_17048,N_16844,N_16752);
nor U17049 (N_17049,N_16953,N_16939);
xnor U17050 (N_17050,N_16856,N_16980);
nand U17051 (N_17051,N_16993,N_16796);
or U17052 (N_17052,N_16764,N_16861);
nor U17053 (N_17053,N_16995,N_16835);
xnor U17054 (N_17054,N_16757,N_16971);
and U17055 (N_17055,N_16801,N_16761);
nand U17056 (N_17056,N_16946,N_16966);
nor U17057 (N_17057,N_16784,N_16880);
nor U17058 (N_17058,N_16852,N_16917);
nor U17059 (N_17059,N_16900,N_16768);
nand U17060 (N_17060,N_16810,N_16753);
nand U17061 (N_17061,N_16928,N_16780);
and U17062 (N_17062,N_16891,N_16811);
nand U17063 (N_17063,N_16873,N_16938);
nor U17064 (N_17064,N_16923,N_16827);
or U17065 (N_17065,N_16843,N_16816);
or U17066 (N_17066,N_16799,N_16862);
xnor U17067 (N_17067,N_16765,N_16832);
xor U17068 (N_17068,N_16829,N_16828);
or U17069 (N_17069,N_16998,N_16871);
nand U17070 (N_17070,N_16977,N_16798);
nor U17071 (N_17071,N_16988,N_16920);
nor U17072 (N_17072,N_16848,N_16866);
and U17073 (N_17073,N_16773,N_16886);
nor U17074 (N_17074,N_16875,N_16970);
nor U17075 (N_17075,N_16911,N_16826);
xor U17076 (N_17076,N_16899,N_16974);
nor U17077 (N_17077,N_16775,N_16820);
and U17078 (N_17078,N_16895,N_16978);
or U17079 (N_17079,N_16951,N_16959);
or U17080 (N_17080,N_16864,N_16890);
nand U17081 (N_17081,N_16836,N_16892);
nor U17082 (N_17082,N_16969,N_16760);
or U17083 (N_17083,N_16791,N_16934);
xor U17084 (N_17084,N_16863,N_16756);
xnor U17085 (N_17085,N_16976,N_16984);
nand U17086 (N_17086,N_16968,N_16777);
nor U17087 (N_17087,N_16975,N_16858);
nor U17088 (N_17088,N_16913,N_16869);
nand U17089 (N_17089,N_16954,N_16956);
nand U17090 (N_17090,N_16979,N_16906);
xnor U17091 (N_17091,N_16787,N_16952);
nor U17092 (N_17092,N_16825,N_16929);
nor U17093 (N_17093,N_16963,N_16758);
nand U17094 (N_17094,N_16889,N_16990);
nand U17095 (N_17095,N_16908,N_16909);
xnor U17096 (N_17096,N_16833,N_16879);
and U17097 (N_17097,N_16878,N_16927);
nand U17098 (N_17098,N_16942,N_16859);
nor U17099 (N_17099,N_16815,N_16860);
and U17100 (N_17100,N_16960,N_16997);
xor U17101 (N_17101,N_16887,N_16947);
or U17102 (N_17102,N_16987,N_16881);
nor U17103 (N_17103,N_16994,N_16950);
or U17104 (N_17104,N_16962,N_16921);
and U17105 (N_17105,N_16794,N_16754);
or U17106 (N_17106,N_16937,N_16783);
nor U17107 (N_17107,N_16949,N_16800);
and U17108 (N_17108,N_16865,N_16872);
nor U17109 (N_17109,N_16874,N_16847);
or U17110 (N_17110,N_16789,N_16814);
or U17111 (N_17111,N_16922,N_16958);
nor U17112 (N_17112,N_16808,N_16751);
and U17113 (N_17113,N_16912,N_16876);
nand U17114 (N_17114,N_16898,N_16792);
xnor U17115 (N_17115,N_16904,N_16982);
nand U17116 (N_17116,N_16766,N_16772);
xnor U17117 (N_17117,N_16914,N_16948);
and U17118 (N_17118,N_16910,N_16823);
nand U17119 (N_17119,N_16771,N_16762);
xnor U17120 (N_17120,N_16788,N_16991);
nor U17121 (N_17121,N_16926,N_16853);
nor U17122 (N_17122,N_16837,N_16915);
nand U17123 (N_17123,N_16854,N_16819);
or U17124 (N_17124,N_16943,N_16855);
and U17125 (N_17125,N_16833,N_16785);
and U17126 (N_17126,N_16936,N_16901);
nor U17127 (N_17127,N_16949,N_16902);
nand U17128 (N_17128,N_16842,N_16929);
nor U17129 (N_17129,N_16857,N_16775);
nor U17130 (N_17130,N_16954,N_16779);
nand U17131 (N_17131,N_16916,N_16965);
or U17132 (N_17132,N_16830,N_16881);
and U17133 (N_17133,N_16769,N_16855);
xor U17134 (N_17134,N_16937,N_16947);
nor U17135 (N_17135,N_16790,N_16918);
or U17136 (N_17136,N_16860,N_16921);
nand U17137 (N_17137,N_16762,N_16835);
and U17138 (N_17138,N_16946,N_16978);
xnor U17139 (N_17139,N_16996,N_16901);
nor U17140 (N_17140,N_16987,N_16968);
nor U17141 (N_17141,N_16792,N_16903);
xor U17142 (N_17142,N_16883,N_16798);
or U17143 (N_17143,N_16763,N_16855);
xor U17144 (N_17144,N_16850,N_16999);
xnor U17145 (N_17145,N_16879,N_16969);
or U17146 (N_17146,N_16943,N_16929);
nor U17147 (N_17147,N_16862,N_16945);
or U17148 (N_17148,N_16942,N_16804);
and U17149 (N_17149,N_16896,N_16940);
and U17150 (N_17150,N_16964,N_16832);
and U17151 (N_17151,N_16870,N_16940);
nand U17152 (N_17152,N_16755,N_16901);
and U17153 (N_17153,N_16991,N_16778);
nand U17154 (N_17154,N_16830,N_16915);
nand U17155 (N_17155,N_16896,N_16861);
xnor U17156 (N_17156,N_16825,N_16761);
nand U17157 (N_17157,N_16785,N_16998);
nor U17158 (N_17158,N_16838,N_16900);
and U17159 (N_17159,N_16848,N_16755);
and U17160 (N_17160,N_16950,N_16954);
nand U17161 (N_17161,N_16974,N_16757);
nor U17162 (N_17162,N_16857,N_16928);
xnor U17163 (N_17163,N_16805,N_16979);
and U17164 (N_17164,N_16810,N_16836);
xnor U17165 (N_17165,N_16848,N_16780);
or U17166 (N_17166,N_16973,N_16888);
or U17167 (N_17167,N_16860,N_16783);
nor U17168 (N_17168,N_16849,N_16777);
nor U17169 (N_17169,N_16940,N_16768);
or U17170 (N_17170,N_16858,N_16846);
nand U17171 (N_17171,N_16832,N_16951);
nor U17172 (N_17172,N_16942,N_16754);
nand U17173 (N_17173,N_16791,N_16984);
or U17174 (N_17174,N_16827,N_16991);
nand U17175 (N_17175,N_16755,N_16876);
xor U17176 (N_17176,N_16865,N_16763);
xor U17177 (N_17177,N_16849,N_16953);
nand U17178 (N_17178,N_16976,N_16943);
or U17179 (N_17179,N_16756,N_16891);
nand U17180 (N_17180,N_16898,N_16823);
nor U17181 (N_17181,N_16793,N_16847);
nand U17182 (N_17182,N_16831,N_16807);
and U17183 (N_17183,N_16919,N_16894);
nand U17184 (N_17184,N_16775,N_16842);
nand U17185 (N_17185,N_16967,N_16981);
nand U17186 (N_17186,N_16923,N_16943);
xnor U17187 (N_17187,N_16958,N_16918);
xor U17188 (N_17188,N_16770,N_16938);
nor U17189 (N_17189,N_16974,N_16788);
and U17190 (N_17190,N_16995,N_16894);
xor U17191 (N_17191,N_16777,N_16847);
xor U17192 (N_17192,N_16780,N_16924);
xor U17193 (N_17193,N_16913,N_16767);
nand U17194 (N_17194,N_16833,N_16761);
nor U17195 (N_17195,N_16877,N_16920);
nand U17196 (N_17196,N_16854,N_16774);
and U17197 (N_17197,N_16887,N_16980);
xor U17198 (N_17198,N_16787,N_16880);
nor U17199 (N_17199,N_16976,N_16909);
nor U17200 (N_17200,N_16900,N_16955);
and U17201 (N_17201,N_16752,N_16801);
or U17202 (N_17202,N_16986,N_16913);
nand U17203 (N_17203,N_16930,N_16840);
nand U17204 (N_17204,N_16927,N_16790);
nand U17205 (N_17205,N_16870,N_16815);
nor U17206 (N_17206,N_16873,N_16763);
nor U17207 (N_17207,N_16907,N_16786);
xnor U17208 (N_17208,N_16863,N_16753);
nand U17209 (N_17209,N_16789,N_16911);
and U17210 (N_17210,N_16903,N_16939);
and U17211 (N_17211,N_16786,N_16927);
nor U17212 (N_17212,N_16919,N_16805);
xnor U17213 (N_17213,N_16938,N_16950);
nor U17214 (N_17214,N_16774,N_16841);
or U17215 (N_17215,N_16798,N_16845);
xnor U17216 (N_17216,N_16829,N_16988);
and U17217 (N_17217,N_16762,N_16862);
and U17218 (N_17218,N_16854,N_16979);
nand U17219 (N_17219,N_16993,N_16959);
nor U17220 (N_17220,N_16764,N_16881);
xor U17221 (N_17221,N_16803,N_16951);
nand U17222 (N_17222,N_16759,N_16780);
and U17223 (N_17223,N_16978,N_16815);
and U17224 (N_17224,N_16993,N_16928);
nor U17225 (N_17225,N_16757,N_16950);
and U17226 (N_17226,N_16889,N_16786);
and U17227 (N_17227,N_16949,N_16942);
xnor U17228 (N_17228,N_16988,N_16918);
or U17229 (N_17229,N_16786,N_16928);
xnor U17230 (N_17230,N_16771,N_16892);
and U17231 (N_17231,N_16763,N_16779);
nor U17232 (N_17232,N_16966,N_16915);
nand U17233 (N_17233,N_16885,N_16994);
and U17234 (N_17234,N_16919,N_16923);
nand U17235 (N_17235,N_16795,N_16951);
xnor U17236 (N_17236,N_16875,N_16785);
xor U17237 (N_17237,N_16821,N_16989);
xor U17238 (N_17238,N_16880,N_16830);
or U17239 (N_17239,N_16863,N_16805);
and U17240 (N_17240,N_16941,N_16882);
xnor U17241 (N_17241,N_16772,N_16858);
or U17242 (N_17242,N_16836,N_16834);
xor U17243 (N_17243,N_16945,N_16803);
or U17244 (N_17244,N_16862,N_16895);
nand U17245 (N_17245,N_16958,N_16945);
xor U17246 (N_17246,N_16894,N_16786);
or U17247 (N_17247,N_16841,N_16784);
nand U17248 (N_17248,N_16941,N_16851);
and U17249 (N_17249,N_16989,N_16908);
and U17250 (N_17250,N_17075,N_17080);
nand U17251 (N_17251,N_17015,N_17153);
or U17252 (N_17252,N_17127,N_17025);
nor U17253 (N_17253,N_17161,N_17020);
nor U17254 (N_17254,N_17057,N_17234);
and U17255 (N_17255,N_17196,N_17164);
or U17256 (N_17256,N_17206,N_17100);
xor U17257 (N_17257,N_17160,N_17069);
nand U17258 (N_17258,N_17115,N_17066);
or U17259 (N_17259,N_17007,N_17105);
nor U17260 (N_17260,N_17035,N_17013);
xor U17261 (N_17261,N_17119,N_17023);
and U17262 (N_17262,N_17139,N_17144);
nand U17263 (N_17263,N_17245,N_17223);
xnor U17264 (N_17264,N_17097,N_17049);
nor U17265 (N_17265,N_17113,N_17209);
or U17266 (N_17266,N_17215,N_17064);
or U17267 (N_17267,N_17212,N_17017);
nand U17268 (N_17268,N_17034,N_17031);
or U17269 (N_17269,N_17026,N_17051);
xnor U17270 (N_17270,N_17148,N_17094);
nand U17271 (N_17271,N_17016,N_17074);
nand U17272 (N_17272,N_17237,N_17201);
xnor U17273 (N_17273,N_17226,N_17089);
nand U17274 (N_17274,N_17087,N_17041);
nand U17275 (N_17275,N_17042,N_17009);
nand U17276 (N_17276,N_17043,N_17036);
and U17277 (N_17277,N_17242,N_17134);
xor U17278 (N_17278,N_17152,N_17118);
or U17279 (N_17279,N_17176,N_17207);
nor U17280 (N_17280,N_17214,N_17005);
and U17281 (N_17281,N_17168,N_17175);
or U17282 (N_17282,N_17155,N_17181);
nand U17283 (N_17283,N_17233,N_17059);
or U17284 (N_17284,N_17142,N_17056);
nand U17285 (N_17285,N_17117,N_17194);
nand U17286 (N_17286,N_17170,N_17159);
nor U17287 (N_17287,N_17240,N_17053);
and U17288 (N_17288,N_17030,N_17129);
and U17289 (N_17289,N_17203,N_17140);
and U17290 (N_17290,N_17073,N_17241);
nor U17291 (N_17291,N_17172,N_17027);
nor U17292 (N_17292,N_17228,N_17093);
and U17293 (N_17293,N_17112,N_17072);
xnor U17294 (N_17294,N_17179,N_17230);
xnor U17295 (N_17295,N_17191,N_17090);
nor U17296 (N_17296,N_17038,N_17067);
and U17297 (N_17297,N_17183,N_17040);
and U17298 (N_17298,N_17138,N_17244);
nand U17299 (N_17299,N_17116,N_17008);
or U17300 (N_17300,N_17032,N_17149);
nand U17301 (N_17301,N_17156,N_17218);
nand U17302 (N_17302,N_17098,N_17182);
and U17303 (N_17303,N_17126,N_17227);
nand U17304 (N_17304,N_17178,N_17143);
or U17305 (N_17305,N_17239,N_17079);
xor U17306 (N_17306,N_17039,N_17063);
nand U17307 (N_17307,N_17232,N_17174);
nand U17308 (N_17308,N_17185,N_17166);
xor U17309 (N_17309,N_17150,N_17095);
xor U17310 (N_17310,N_17052,N_17222);
xnor U17311 (N_17311,N_17060,N_17199);
and U17312 (N_17312,N_17123,N_17165);
nand U17313 (N_17313,N_17044,N_17107);
xor U17314 (N_17314,N_17022,N_17157);
or U17315 (N_17315,N_17188,N_17121);
and U17316 (N_17316,N_17106,N_17248);
and U17317 (N_17317,N_17229,N_17122);
or U17318 (N_17318,N_17109,N_17128);
nand U17319 (N_17319,N_17103,N_17208);
and U17320 (N_17320,N_17077,N_17102);
and U17321 (N_17321,N_17202,N_17180);
nor U17322 (N_17322,N_17101,N_17224);
and U17323 (N_17323,N_17210,N_17083);
or U17324 (N_17324,N_17088,N_17146);
or U17325 (N_17325,N_17192,N_17243);
nor U17326 (N_17326,N_17000,N_17220);
xor U17327 (N_17327,N_17186,N_17058);
nand U17328 (N_17328,N_17213,N_17195);
xnor U17329 (N_17329,N_17033,N_17200);
nand U17330 (N_17330,N_17046,N_17193);
or U17331 (N_17331,N_17154,N_17014);
xor U17332 (N_17332,N_17091,N_17189);
nor U17333 (N_17333,N_17028,N_17238);
nor U17334 (N_17334,N_17187,N_17068);
nor U17335 (N_17335,N_17133,N_17130);
nor U17336 (N_17336,N_17198,N_17171);
or U17337 (N_17337,N_17114,N_17082);
or U17338 (N_17338,N_17120,N_17135);
nand U17339 (N_17339,N_17048,N_17003);
nand U17340 (N_17340,N_17211,N_17132);
or U17341 (N_17341,N_17084,N_17055);
xor U17342 (N_17342,N_17177,N_17184);
nor U17343 (N_17343,N_17071,N_17024);
or U17344 (N_17344,N_17006,N_17151);
or U17345 (N_17345,N_17225,N_17001);
and U17346 (N_17346,N_17221,N_17125);
xnor U17347 (N_17347,N_17141,N_17037);
xor U17348 (N_17348,N_17104,N_17145);
nor U17349 (N_17349,N_17099,N_17197);
and U17350 (N_17350,N_17205,N_17158);
and U17351 (N_17351,N_17147,N_17061);
nand U17352 (N_17352,N_17002,N_17047);
nand U17353 (N_17353,N_17219,N_17054);
or U17354 (N_17354,N_17011,N_17092);
nor U17355 (N_17355,N_17076,N_17162);
and U17356 (N_17356,N_17246,N_17167);
nor U17357 (N_17357,N_17012,N_17163);
xnor U17358 (N_17358,N_17085,N_17086);
and U17359 (N_17359,N_17029,N_17216);
xor U17360 (N_17360,N_17173,N_17070);
nand U17361 (N_17361,N_17236,N_17190);
nor U17362 (N_17362,N_17204,N_17065);
xor U17363 (N_17363,N_17169,N_17096);
and U17364 (N_17364,N_17050,N_17249);
or U17365 (N_17365,N_17110,N_17131);
nor U17366 (N_17366,N_17018,N_17247);
and U17367 (N_17367,N_17235,N_17137);
or U17368 (N_17368,N_17019,N_17124);
or U17369 (N_17369,N_17062,N_17078);
or U17370 (N_17370,N_17004,N_17108);
nand U17371 (N_17371,N_17231,N_17111);
nor U17372 (N_17372,N_17081,N_17010);
or U17373 (N_17373,N_17021,N_17217);
xnor U17374 (N_17374,N_17045,N_17136);
or U17375 (N_17375,N_17237,N_17027);
and U17376 (N_17376,N_17148,N_17136);
and U17377 (N_17377,N_17022,N_17070);
xnor U17378 (N_17378,N_17203,N_17182);
and U17379 (N_17379,N_17070,N_17075);
nand U17380 (N_17380,N_17016,N_17062);
and U17381 (N_17381,N_17038,N_17245);
or U17382 (N_17382,N_17110,N_17249);
and U17383 (N_17383,N_17095,N_17040);
xor U17384 (N_17384,N_17175,N_17030);
nand U17385 (N_17385,N_17067,N_17013);
and U17386 (N_17386,N_17187,N_17000);
xor U17387 (N_17387,N_17214,N_17130);
xor U17388 (N_17388,N_17024,N_17205);
nor U17389 (N_17389,N_17214,N_17204);
or U17390 (N_17390,N_17016,N_17050);
and U17391 (N_17391,N_17183,N_17238);
nor U17392 (N_17392,N_17099,N_17042);
nor U17393 (N_17393,N_17157,N_17126);
nor U17394 (N_17394,N_17038,N_17156);
and U17395 (N_17395,N_17248,N_17220);
nand U17396 (N_17396,N_17143,N_17021);
nor U17397 (N_17397,N_17043,N_17224);
or U17398 (N_17398,N_17234,N_17183);
and U17399 (N_17399,N_17154,N_17005);
nor U17400 (N_17400,N_17095,N_17240);
nand U17401 (N_17401,N_17081,N_17204);
or U17402 (N_17402,N_17175,N_17210);
xnor U17403 (N_17403,N_17022,N_17076);
or U17404 (N_17404,N_17184,N_17168);
nor U17405 (N_17405,N_17220,N_17067);
and U17406 (N_17406,N_17234,N_17189);
nor U17407 (N_17407,N_17061,N_17219);
nor U17408 (N_17408,N_17155,N_17005);
or U17409 (N_17409,N_17185,N_17129);
nor U17410 (N_17410,N_17084,N_17043);
nand U17411 (N_17411,N_17096,N_17227);
xnor U17412 (N_17412,N_17093,N_17217);
and U17413 (N_17413,N_17249,N_17106);
nor U17414 (N_17414,N_17014,N_17107);
nand U17415 (N_17415,N_17234,N_17204);
nor U17416 (N_17416,N_17024,N_17236);
and U17417 (N_17417,N_17035,N_17221);
xnor U17418 (N_17418,N_17204,N_17121);
nand U17419 (N_17419,N_17132,N_17040);
or U17420 (N_17420,N_17041,N_17049);
xor U17421 (N_17421,N_17048,N_17204);
xor U17422 (N_17422,N_17104,N_17128);
and U17423 (N_17423,N_17055,N_17156);
and U17424 (N_17424,N_17061,N_17064);
nand U17425 (N_17425,N_17174,N_17113);
nand U17426 (N_17426,N_17171,N_17024);
xnor U17427 (N_17427,N_17102,N_17020);
or U17428 (N_17428,N_17070,N_17155);
nand U17429 (N_17429,N_17111,N_17055);
nand U17430 (N_17430,N_17147,N_17047);
nor U17431 (N_17431,N_17246,N_17020);
nand U17432 (N_17432,N_17234,N_17198);
or U17433 (N_17433,N_17117,N_17000);
xor U17434 (N_17434,N_17198,N_17001);
nand U17435 (N_17435,N_17101,N_17045);
or U17436 (N_17436,N_17246,N_17226);
and U17437 (N_17437,N_17141,N_17140);
and U17438 (N_17438,N_17132,N_17152);
or U17439 (N_17439,N_17051,N_17182);
xor U17440 (N_17440,N_17150,N_17233);
xnor U17441 (N_17441,N_17121,N_17089);
nor U17442 (N_17442,N_17073,N_17219);
nand U17443 (N_17443,N_17038,N_17124);
nand U17444 (N_17444,N_17028,N_17184);
nand U17445 (N_17445,N_17223,N_17004);
nor U17446 (N_17446,N_17175,N_17156);
nor U17447 (N_17447,N_17138,N_17032);
and U17448 (N_17448,N_17225,N_17093);
and U17449 (N_17449,N_17043,N_17183);
or U17450 (N_17450,N_17212,N_17098);
and U17451 (N_17451,N_17202,N_17212);
and U17452 (N_17452,N_17059,N_17084);
xnor U17453 (N_17453,N_17188,N_17216);
and U17454 (N_17454,N_17095,N_17201);
and U17455 (N_17455,N_17225,N_17199);
xnor U17456 (N_17456,N_17000,N_17166);
and U17457 (N_17457,N_17219,N_17195);
nand U17458 (N_17458,N_17059,N_17220);
nor U17459 (N_17459,N_17066,N_17112);
xor U17460 (N_17460,N_17187,N_17069);
and U17461 (N_17461,N_17107,N_17178);
nand U17462 (N_17462,N_17002,N_17229);
and U17463 (N_17463,N_17112,N_17058);
xor U17464 (N_17464,N_17118,N_17073);
and U17465 (N_17465,N_17193,N_17013);
xor U17466 (N_17466,N_17044,N_17235);
and U17467 (N_17467,N_17152,N_17106);
nor U17468 (N_17468,N_17129,N_17167);
or U17469 (N_17469,N_17233,N_17082);
xor U17470 (N_17470,N_17231,N_17246);
nor U17471 (N_17471,N_17148,N_17242);
xnor U17472 (N_17472,N_17064,N_17216);
or U17473 (N_17473,N_17095,N_17167);
nor U17474 (N_17474,N_17039,N_17064);
and U17475 (N_17475,N_17054,N_17233);
and U17476 (N_17476,N_17109,N_17102);
nor U17477 (N_17477,N_17075,N_17015);
and U17478 (N_17478,N_17179,N_17129);
nand U17479 (N_17479,N_17089,N_17244);
or U17480 (N_17480,N_17064,N_17102);
nand U17481 (N_17481,N_17113,N_17155);
and U17482 (N_17482,N_17240,N_17126);
nand U17483 (N_17483,N_17061,N_17014);
nand U17484 (N_17484,N_17147,N_17149);
nor U17485 (N_17485,N_17014,N_17184);
or U17486 (N_17486,N_17155,N_17078);
or U17487 (N_17487,N_17037,N_17130);
nor U17488 (N_17488,N_17104,N_17163);
nand U17489 (N_17489,N_17073,N_17084);
or U17490 (N_17490,N_17030,N_17001);
nor U17491 (N_17491,N_17174,N_17154);
nand U17492 (N_17492,N_17058,N_17075);
or U17493 (N_17493,N_17134,N_17110);
and U17494 (N_17494,N_17066,N_17155);
nor U17495 (N_17495,N_17187,N_17116);
nor U17496 (N_17496,N_17240,N_17161);
nor U17497 (N_17497,N_17013,N_17014);
nand U17498 (N_17498,N_17166,N_17120);
xor U17499 (N_17499,N_17028,N_17207);
xnor U17500 (N_17500,N_17455,N_17406);
nor U17501 (N_17501,N_17302,N_17373);
or U17502 (N_17502,N_17471,N_17399);
and U17503 (N_17503,N_17462,N_17267);
or U17504 (N_17504,N_17374,N_17338);
or U17505 (N_17505,N_17423,N_17270);
or U17506 (N_17506,N_17320,N_17494);
nand U17507 (N_17507,N_17253,N_17358);
or U17508 (N_17508,N_17314,N_17475);
nand U17509 (N_17509,N_17484,N_17491);
nand U17510 (N_17510,N_17478,N_17271);
xnor U17511 (N_17511,N_17480,N_17301);
nand U17512 (N_17512,N_17367,N_17312);
and U17513 (N_17513,N_17427,N_17284);
nand U17514 (N_17514,N_17305,N_17357);
xnor U17515 (N_17515,N_17313,N_17274);
nor U17516 (N_17516,N_17332,N_17479);
or U17517 (N_17517,N_17420,N_17465);
nor U17518 (N_17518,N_17261,N_17459);
nand U17519 (N_17519,N_17397,N_17372);
nand U17520 (N_17520,N_17456,N_17496);
xnor U17521 (N_17521,N_17366,N_17251);
or U17522 (N_17522,N_17381,N_17498);
nor U17523 (N_17523,N_17371,N_17341);
nor U17524 (N_17524,N_17388,N_17375);
xnor U17525 (N_17525,N_17452,N_17428);
and U17526 (N_17526,N_17453,N_17395);
xnor U17527 (N_17527,N_17266,N_17383);
or U17528 (N_17528,N_17382,N_17443);
xnor U17529 (N_17529,N_17264,N_17359);
and U17530 (N_17530,N_17461,N_17269);
nand U17531 (N_17531,N_17447,N_17281);
and U17532 (N_17532,N_17396,N_17370);
or U17533 (N_17533,N_17265,N_17310);
or U17534 (N_17534,N_17450,N_17356);
nand U17535 (N_17535,N_17262,N_17430);
nand U17536 (N_17536,N_17368,N_17328);
and U17537 (N_17537,N_17365,N_17460);
nand U17538 (N_17538,N_17432,N_17492);
xnor U17539 (N_17539,N_17387,N_17353);
nor U17540 (N_17540,N_17355,N_17385);
and U17541 (N_17541,N_17250,N_17445);
nor U17542 (N_17542,N_17437,N_17409);
and U17543 (N_17543,N_17340,N_17325);
nor U17544 (N_17544,N_17438,N_17369);
nand U17545 (N_17545,N_17477,N_17327);
nand U17546 (N_17546,N_17280,N_17490);
nor U17547 (N_17547,N_17434,N_17431);
nand U17548 (N_17548,N_17362,N_17417);
xor U17549 (N_17549,N_17364,N_17348);
xnor U17550 (N_17550,N_17335,N_17411);
nand U17551 (N_17551,N_17260,N_17408);
nand U17552 (N_17552,N_17293,N_17457);
xnor U17553 (N_17553,N_17287,N_17345);
nor U17554 (N_17554,N_17289,N_17354);
nor U17555 (N_17555,N_17435,N_17404);
nor U17556 (N_17556,N_17499,N_17346);
nand U17557 (N_17557,N_17441,N_17489);
nor U17558 (N_17558,N_17292,N_17323);
nor U17559 (N_17559,N_17485,N_17268);
and U17560 (N_17560,N_17278,N_17318);
or U17561 (N_17561,N_17403,N_17418);
and U17562 (N_17562,N_17259,N_17321);
nand U17563 (N_17563,N_17306,N_17497);
xor U17564 (N_17564,N_17415,N_17483);
or U17565 (N_17565,N_17444,N_17472);
nand U17566 (N_17566,N_17424,N_17466);
nor U17567 (N_17567,N_17446,N_17386);
nand U17568 (N_17568,N_17339,N_17413);
nor U17569 (N_17569,N_17300,N_17482);
and U17570 (N_17570,N_17330,N_17277);
xnor U17571 (N_17571,N_17326,N_17350);
and U17572 (N_17572,N_17273,N_17394);
xnor U17573 (N_17573,N_17487,N_17285);
and U17574 (N_17574,N_17425,N_17351);
nor U17575 (N_17575,N_17481,N_17263);
nor U17576 (N_17576,N_17298,N_17393);
and U17577 (N_17577,N_17282,N_17333);
xor U17578 (N_17578,N_17276,N_17454);
or U17579 (N_17579,N_17275,N_17296);
and U17580 (N_17580,N_17493,N_17464);
or U17581 (N_17581,N_17402,N_17334);
and U17582 (N_17582,N_17421,N_17324);
or U17583 (N_17583,N_17342,N_17468);
xor U17584 (N_17584,N_17319,N_17436);
nand U17585 (N_17585,N_17288,N_17467);
nor U17586 (N_17586,N_17476,N_17449);
xnor U17587 (N_17587,N_17458,N_17309);
nand U17588 (N_17588,N_17389,N_17422);
or U17589 (N_17589,N_17448,N_17294);
nor U17590 (N_17590,N_17295,N_17390);
nand U17591 (N_17591,N_17255,N_17398);
nand U17592 (N_17592,N_17470,N_17401);
and U17593 (N_17593,N_17469,N_17360);
nor U17594 (N_17594,N_17376,N_17400);
nand U17595 (N_17595,N_17344,N_17258);
or U17596 (N_17596,N_17315,N_17405);
xor U17597 (N_17597,N_17363,N_17286);
nor U17598 (N_17598,N_17426,N_17451);
or U17599 (N_17599,N_17317,N_17307);
nor U17600 (N_17600,N_17429,N_17407);
xnor U17601 (N_17601,N_17392,N_17349);
and U17602 (N_17602,N_17463,N_17290);
nand U17603 (N_17603,N_17257,N_17486);
xor U17604 (N_17604,N_17256,N_17322);
nand U17605 (N_17605,N_17303,N_17384);
xor U17606 (N_17606,N_17433,N_17361);
xor U17607 (N_17607,N_17329,N_17316);
and U17608 (N_17608,N_17252,N_17419);
nor U17609 (N_17609,N_17304,N_17380);
and U17610 (N_17610,N_17412,N_17308);
nor U17611 (N_17611,N_17378,N_17347);
or U17612 (N_17612,N_17299,N_17336);
nand U17613 (N_17613,N_17331,N_17495);
and U17614 (N_17614,N_17410,N_17379);
nand U17615 (N_17615,N_17473,N_17474);
xnor U17616 (N_17616,N_17291,N_17297);
or U17617 (N_17617,N_17416,N_17377);
or U17618 (N_17618,N_17442,N_17311);
nor U17619 (N_17619,N_17440,N_17279);
or U17620 (N_17620,N_17272,N_17337);
xnor U17621 (N_17621,N_17283,N_17488);
and U17622 (N_17622,N_17352,N_17391);
xnor U17623 (N_17623,N_17254,N_17414);
xor U17624 (N_17624,N_17439,N_17343);
or U17625 (N_17625,N_17346,N_17311);
nand U17626 (N_17626,N_17364,N_17282);
and U17627 (N_17627,N_17371,N_17461);
xor U17628 (N_17628,N_17425,N_17329);
and U17629 (N_17629,N_17410,N_17312);
or U17630 (N_17630,N_17426,N_17286);
nand U17631 (N_17631,N_17350,N_17475);
nand U17632 (N_17632,N_17267,N_17456);
or U17633 (N_17633,N_17354,N_17368);
nand U17634 (N_17634,N_17313,N_17256);
nand U17635 (N_17635,N_17330,N_17427);
nor U17636 (N_17636,N_17337,N_17483);
and U17637 (N_17637,N_17274,N_17403);
xor U17638 (N_17638,N_17382,N_17426);
and U17639 (N_17639,N_17468,N_17414);
and U17640 (N_17640,N_17420,N_17447);
xor U17641 (N_17641,N_17258,N_17480);
nand U17642 (N_17642,N_17394,N_17415);
xnor U17643 (N_17643,N_17405,N_17391);
nor U17644 (N_17644,N_17449,N_17388);
and U17645 (N_17645,N_17344,N_17283);
or U17646 (N_17646,N_17383,N_17324);
xor U17647 (N_17647,N_17324,N_17297);
nand U17648 (N_17648,N_17405,N_17488);
and U17649 (N_17649,N_17462,N_17402);
nand U17650 (N_17650,N_17307,N_17457);
nor U17651 (N_17651,N_17495,N_17499);
nand U17652 (N_17652,N_17298,N_17357);
or U17653 (N_17653,N_17380,N_17267);
nand U17654 (N_17654,N_17469,N_17476);
and U17655 (N_17655,N_17377,N_17381);
nand U17656 (N_17656,N_17464,N_17323);
and U17657 (N_17657,N_17373,N_17325);
xor U17658 (N_17658,N_17354,N_17351);
nand U17659 (N_17659,N_17332,N_17366);
and U17660 (N_17660,N_17343,N_17456);
xor U17661 (N_17661,N_17259,N_17387);
and U17662 (N_17662,N_17316,N_17299);
nor U17663 (N_17663,N_17463,N_17404);
or U17664 (N_17664,N_17289,N_17271);
xor U17665 (N_17665,N_17440,N_17314);
and U17666 (N_17666,N_17364,N_17492);
xor U17667 (N_17667,N_17255,N_17292);
nand U17668 (N_17668,N_17281,N_17368);
nor U17669 (N_17669,N_17280,N_17353);
xor U17670 (N_17670,N_17328,N_17258);
nor U17671 (N_17671,N_17293,N_17436);
or U17672 (N_17672,N_17435,N_17340);
xnor U17673 (N_17673,N_17264,N_17374);
or U17674 (N_17674,N_17418,N_17267);
and U17675 (N_17675,N_17475,N_17455);
and U17676 (N_17676,N_17254,N_17463);
xor U17677 (N_17677,N_17338,N_17404);
or U17678 (N_17678,N_17369,N_17424);
nand U17679 (N_17679,N_17361,N_17322);
xnor U17680 (N_17680,N_17467,N_17327);
nand U17681 (N_17681,N_17285,N_17431);
and U17682 (N_17682,N_17419,N_17260);
nand U17683 (N_17683,N_17263,N_17477);
nor U17684 (N_17684,N_17424,N_17426);
nand U17685 (N_17685,N_17387,N_17497);
xnor U17686 (N_17686,N_17316,N_17382);
or U17687 (N_17687,N_17410,N_17298);
xor U17688 (N_17688,N_17328,N_17276);
nand U17689 (N_17689,N_17445,N_17464);
or U17690 (N_17690,N_17323,N_17302);
nor U17691 (N_17691,N_17279,N_17469);
nand U17692 (N_17692,N_17317,N_17332);
xnor U17693 (N_17693,N_17418,N_17408);
and U17694 (N_17694,N_17401,N_17286);
xnor U17695 (N_17695,N_17311,N_17350);
and U17696 (N_17696,N_17384,N_17334);
and U17697 (N_17697,N_17348,N_17375);
nand U17698 (N_17698,N_17367,N_17297);
or U17699 (N_17699,N_17365,N_17407);
and U17700 (N_17700,N_17308,N_17421);
xor U17701 (N_17701,N_17463,N_17294);
xnor U17702 (N_17702,N_17388,N_17269);
xor U17703 (N_17703,N_17360,N_17364);
nor U17704 (N_17704,N_17426,N_17258);
xor U17705 (N_17705,N_17434,N_17488);
nand U17706 (N_17706,N_17340,N_17351);
and U17707 (N_17707,N_17264,N_17369);
nand U17708 (N_17708,N_17296,N_17425);
xnor U17709 (N_17709,N_17461,N_17494);
nor U17710 (N_17710,N_17418,N_17485);
nand U17711 (N_17711,N_17358,N_17433);
nand U17712 (N_17712,N_17321,N_17472);
or U17713 (N_17713,N_17342,N_17261);
nor U17714 (N_17714,N_17307,N_17424);
or U17715 (N_17715,N_17360,N_17351);
nor U17716 (N_17716,N_17264,N_17436);
nor U17717 (N_17717,N_17304,N_17251);
or U17718 (N_17718,N_17487,N_17253);
nor U17719 (N_17719,N_17353,N_17342);
or U17720 (N_17720,N_17407,N_17462);
and U17721 (N_17721,N_17261,N_17322);
or U17722 (N_17722,N_17363,N_17406);
xnor U17723 (N_17723,N_17470,N_17372);
xor U17724 (N_17724,N_17266,N_17260);
xnor U17725 (N_17725,N_17268,N_17330);
and U17726 (N_17726,N_17486,N_17373);
xor U17727 (N_17727,N_17357,N_17352);
and U17728 (N_17728,N_17469,N_17274);
or U17729 (N_17729,N_17316,N_17373);
nor U17730 (N_17730,N_17475,N_17433);
nand U17731 (N_17731,N_17422,N_17342);
and U17732 (N_17732,N_17462,N_17448);
and U17733 (N_17733,N_17402,N_17322);
and U17734 (N_17734,N_17297,N_17276);
nor U17735 (N_17735,N_17358,N_17396);
nand U17736 (N_17736,N_17272,N_17265);
nand U17737 (N_17737,N_17276,N_17420);
and U17738 (N_17738,N_17348,N_17448);
or U17739 (N_17739,N_17439,N_17374);
or U17740 (N_17740,N_17313,N_17360);
nor U17741 (N_17741,N_17290,N_17265);
or U17742 (N_17742,N_17477,N_17373);
and U17743 (N_17743,N_17351,N_17412);
xor U17744 (N_17744,N_17330,N_17401);
and U17745 (N_17745,N_17380,N_17340);
nor U17746 (N_17746,N_17406,N_17387);
xnor U17747 (N_17747,N_17350,N_17309);
nand U17748 (N_17748,N_17456,N_17412);
nor U17749 (N_17749,N_17339,N_17369);
xor U17750 (N_17750,N_17727,N_17564);
and U17751 (N_17751,N_17618,N_17623);
and U17752 (N_17752,N_17560,N_17744);
nor U17753 (N_17753,N_17590,N_17638);
and U17754 (N_17754,N_17717,N_17655);
nand U17755 (N_17755,N_17624,N_17559);
and U17756 (N_17756,N_17606,N_17679);
and U17757 (N_17757,N_17563,N_17531);
nor U17758 (N_17758,N_17574,N_17724);
and U17759 (N_17759,N_17696,N_17729);
and U17760 (N_17760,N_17736,N_17709);
nand U17761 (N_17761,N_17621,N_17682);
nand U17762 (N_17762,N_17680,N_17613);
and U17763 (N_17763,N_17636,N_17523);
xor U17764 (N_17764,N_17708,N_17582);
and U17765 (N_17765,N_17675,N_17627);
nand U17766 (N_17766,N_17516,N_17702);
xor U17767 (N_17767,N_17601,N_17630);
or U17768 (N_17768,N_17572,N_17551);
or U17769 (N_17769,N_17690,N_17747);
or U17770 (N_17770,N_17643,N_17584);
nor U17771 (N_17771,N_17605,N_17598);
and U17772 (N_17772,N_17625,N_17700);
nor U17773 (N_17773,N_17664,N_17652);
or U17774 (N_17774,N_17528,N_17715);
nand U17775 (N_17775,N_17555,N_17656);
nand U17776 (N_17776,N_17588,N_17710);
xor U17777 (N_17777,N_17683,N_17549);
nor U17778 (N_17778,N_17622,N_17739);
or U17779 (N_17779,N_17703,N_17616);
and U17780 (N_17780,N_17681,N_17641);
nand U17781 (N_17781,N_17697,N_17562);
and U17782 (N_17782,N_17721,N_17501);
xnor U17783 (N_17783,N_17527,N_17662);
nor U17784 (N_17784,N_17650,N_17629);
and U17785 (N_17785,N_17500,N_17665);
xnor U17786 (N_17786,N_17547,N_17670);
nand U17787 (N_17787,N_17597,N_17612);
xnor U17788 (N_17788,N_17737,N_17692);
nand U17789 (N_17789,N_17689,N_17694);
or U17790 (N_17790,N_17723,N_17586);
or U17791 (N_17791,N_17746,N_17544);
and U17792 (N_17792,N_17719,N_17515);
and U17793 (N_17793,N_17631,N_17611);
nand U17794 (N_17794,N_17735,N_17732);
or U17795 (N_17795,N_17568,N_17554);
nor U17796 (N_17796,N_17647,N_17540);
nand U17797 (N_17797,N_17740,N_17570);
nor U17798 (N_17798,N_17529,N_17640);
nor U17799 (N_17799,N_17706,N_17573);
xnor U17800 (N_17800,N_17645,N_17599);
and U17801 (N_17801,N_17649,N_17698);
nand U17802 (N_17802,N_17669,N_17566);
or U17803 (N_17803,N_17507,N_17628);
xnor U17804 (N_17804,N_17594,N_17632);
nor U17805 (N_17805,N_17660,N_17579);
or U17806 (N_17806,N_17575,N_17561);
or U17807 (N_17807,N_17541,N_17672);
nor U17808 (N_17808,N_17593,N_17514);
or U17809 (N_17809,N_17667,N_17596);
or U17810 (N_17810,N_17704,N_17522);
nand U17811 (N_17811,N_17651,N_17684);
or U17812 (N_17812,N_17589,N_17535);
or U17813 (N_17813,N_17580,N_17609);
nand U17814 (N_17814,N_17626,N_17550);
or U17815 (N_17815,N_17646,N_17674);
xnor U17816 (N_17816,N_17745,N_17686);
or U17817 (N_17817,N_17707,N_17539);
or U17818 (N_17818,N_17663,N_17509);
nand U17819 (N_17819,N_17637,N_17654);
or U17820 (N_17820,N_17533,N_17603);
and U17821 (N_17821,N_17571,N_17639);
or U17822 (N_17822,N_17595,N_17602);
and U17823 (N_17823,N_17688,N_17720);
or U17824 (N_17824,N_17748,N_17693);
nor U17825 (N_17825,N_17600,N_17502);
and U17826 (N_17826,N_17699,N_17587);
or U17827 (N_17827,N_17543,N_17614);
nand U17828 (N_17828,N_17733,N_17526);
nand U17829 (N_17829,N_17743,N_17685);
xor U17830 (N_17830,N_17749,N_17545);
nor U17831 (N_17831,N_17635,N_17725);
or U17832 (N_17832,N_17673,N_17519);
nor U17833 (N_17833,N_17512,N_17565);
or U17834 (N_17834,N_17716,N_17648);
xnor U17835 (N_17835,N_17532,N_17581);
nand U17836 (N_17836,N_17546,N_17726);
xor U17837 (N_17837,N_17558,N_17511);
and U17838 (N_17838,N_17569,N_17661);
xnor U17839 (N_17839,N_17666,N_17542);
or U17840 (N_17840,N_17712,N_17634);
nand U17841 (N_17841,N_17508,N_17518);
and U17842 (N_17842,N_17521,N_17695);
xnor U17843 (N_17843,N_17676,N_17678);
or U17844 (N_17844,N_17520,N_17615);
or U17845 (N_17845,N_17538,N_17738);
nand U17846 (N_17846,N_17671,N_17705);
and U17847 (N_17847,N_17687,N_17557);
nand U17848 (N_17848,N_17536,N_17503);
nand U17849 (N_17849,N_17517,N_17510);
nand U17850 (N_17850,N_17734,N_17701);
xor U17851 (N_17851,N_17718,N_17607);
and U17852 (N_17852,N_17653,N_17513);
xor U17853 (N_17853,N_17530,N_17644);
or U17854 (N_17854,N_17576,N_17730);
nor U17855 (N_17855,N_17567,N_17577);
and U17856 (N_17856,N_17619,N_17583);
nand U17857 (N_17857,N_17556,N_17659);
nand U17858 (N_17858,N_17534,N_17608);
nor U17859 (N_17859,N_17691,N_17525);
or U17860 (N_17860,N_17592,N_17610);
or U17861 (N_17861,N_17617,N_17677);
nor U17862 (N_17862,N_17591,N_17578);
nor U17863 (N_17863,N_17506,N_17657);
or U17864 (N_17864,N_17668,N_17553);
or U17865 (N_17865,N_17731,N_17620);
or U17866 (N_17866,N_17742,N_17504);
and U17867 (N_17867,N_17524,N_17552);
nand U17868 (N_17868,N_17633,N_17714);
xor U17869 (N_17869,N_17741,N_17658);
nand U17870 (N_17870,N_17548,N_17604);
or U17871 (N_17871,N_17505,N_17642);
xor U17872 (N_17872,N_17585,N_17722);
or U17873 (N_17873,N_17728,N_17713);
or U17874 (N_17874,N_17537,N_17711);
nand U17875 (N_17875,N_17691,N_17601);
nand U17876 (N_17876,N_17731,N_17625);
xor U17877 (N_17877,N_17536,N_17742);
nand U17878 (N_17878,N_17606,N_17534);
nor U17879 (N_17879,N_17710,N_17528);
and U17880 (N_17880,N_17601,N_17509);
and U17881 (N_17881,N_17558,N_17614);
xor U17882 (N_17882,N_17579,N_17552);
nor U17883 (N_17883,N_17663,N_17592);
nor U17884 (N_17884,N_17557,N_17583);
nand U17885 (N_17885,N_17549,N_17681);
nand U17886 (N_17886,N_17566,N_17560);
or U17887 (N_17887,N_17628,N_17634);
nor U17888 (N_17888,N_17548,N_17653);
xnor U17889 (N_17889,N_17749,N_17672);
and U17890 (N_17890,N_17502,N_17561);
xnor U17891 (N_17891,N_17500,N_17727);
xnor U17892 (N_17892,N_17609,N_17579);
nand U17893 (N_17893,N_17732,N_17710);
and U17894 (N_17894,N_17705,N_17593);
xnor U17895 (N_17895,N_17646,N_17699);
nor U17896 (N_17896,N_17705,N_17636);
nand U17897 (N_17897,N_17584,N_17676);
and U17898 (N_17898,N_17530,N_17712);
nand U17899 (N_17899,N_17701,N_17539);
nor U17900 (N_17900,N_17550,N_17523);
and U17901 (N_17901,N_17631,N_17682);
or U17902 (N_17902,N_17519,N_17602);
nor U17903 (N_17903,N_17622,N_17533);
nor U17904 (N_17904,N_17742,N_17552);
nand U17905 (N_17905,N_17594,N_17719);
and U17906 (N_17906,N_17534,N_17516);
or U17907 (N_17907,N_17567,N_17500);
nand U17908 (N_17908,N_17722,N_17685);
or U17909 (N_17909,N_17672,N_17732);
nand U17910 (N_17910,N_17552,N_17572);
or U17911 (N_17911,N_17670,N_17659);
xor U17912 (N_17912,N_17646,N_17581);
nor U17913 (N_17913,N_17727,N_17621);
and U17914 (N_17914,N_17550,N_17503);
or U17915 (N_17915,N_17715,N_17716);
or U17916 (N_17916,N_17563,N_17637);
nand U17917 (N_17917,N_17733,N_17628);
nor U17918 (N_17918,N_17734,N_17700);
nor U17919 (N_17919,N_17627,N_17597);
xnor U17920 (N_17920,N_17741,N_17732);
or U17921 (N_17921,N_17563,N_17522);
or U17922 (N_17922,N_17500,N_17611);
nand U17923 (N_17923,N_17673,N_17562);
nand U17924 (N_17924,N_17533,N_17566);
or U17925 (N_17925,N_17621,N_17570);
and U17926 (N_17926,N_17721,N_17599);
nor U17927 (N_17927,N_17623,N_17720);
xnor U17928 (N_17928,N_17714,N_17645);
nand U17929 (N_17929,N_17623,N_17583);
nand U17930 (N_17930,N_17614,N_17738);
nand U17931 (N_17931,N_17584,N_17695);
xnor U17932 (N_17932,N_17741,N_17647);
xnor U17933 (N_17933,N_17537,N_17651);
nor U17934 (N_17934,N_17596,N_17692);
or U17935 (N_17935,N_17614,N_17668);
xnor U17936 (N_17936,N_17703,N_17550);
nand U17937 (N_17937,N_17713,N_17595);
xor U17938 (N_17938,N_17747,N_17556);
xor U17939 (N_17939,N_17501,N_17609);
nand U17940 (N_17940,N_17725,N_17675);
xnor U17941 (N_17941,N_17544,N_17668);
nand U17942 (N_17942,N_17682,N_17737);
or U17943 (N_17943,N_17744,N_17555);
xor U17944 (N_17944,N_17620,N_17598);
nor U17945 (N_17945,N_17519,N_17718);
and U17946 (N_17946,N_17658,N_17570);
nand U17947 (N_17947,N_17660,N_17639);
or U17948 (N_17948,N_17577,N_17723);
nor U17949 (N_17949,N_17626,N_17596);
nand U17950 (N_17950,N_17578,N_17631);
nor U17951 (N_17951,N_17675,N_17748);
and U17952 (N_17952,N_17706,N_17687);
or U17953 (N_17953,N_17501,N_17743);
or U17954 (N_17954,N_17676,N_17695);
xnor U17955 (N_17955,N_17675,N_17710);
nor U17956 (N_17956,N_17613,N_17596);
xor U17957 (N_17957,N_17726,N_17725);
and U17958 (N_17958,N_17589,N_17727);
or U17959 (N_17959,N_17524,N_17706);
and U17960 (N_17960,N_17551,N_17544);
nor U17961 (N_17961,N_17505,N_17541);
or U17962 (N_17962,N_17510,N_17568);
or U17963 (N_17963,N_17554,N_17677);
or U17964 (N_17964,N_17677,N_17540);
or U17965 (N_17965,N_17541,N_17684);
and U17966 (N_17966,N_17650,N_17579);
nor U17967 (N_17967,N_17691,N_17573);
nor U17968 (N_17968,N_17732,N_17516);
nor U17969 (N_17969,N_17723,N_17564);
and U17970 (N_17970,N_17624,N_17693);
nand U17971 (N_17971,N_17598,N_17580);
nand U17972 (N_17972,N_17660,N_17572);
nor U17973 (N_17973,N_17594,N_17713);
or U17974 (N_17974,N_17681,N_17735);
or U17975 (N_17975,N_17689,N_17624);
or U17976 (N_17976,N_17639,N_17691);
and U17977 (N_17977,N_17546,N_17695);
and U17978 (N_17978,N_17619,N_17553);
xor U17979 (N_17979,N_17546,N_17542);
or U17980 (N_17980,N_17574,N_17737);
or U17981 (N_17981,N_17509,N_17673);
and U17982 (N_17982,N_17596,N_17606);
nand U17983 (N_17983,N_17729,N_17523);
nor U17984 (N_17984,N_17711,N_17635);
xor U17985 (N_17985,N_17541,N_17655);
xor U17986 (N_17986,N_17729,N_17594);
or U17987 (N_17987,N_17672,N_17711);
or U17988 (N_17988,N_17577,N_17728);
nor U17989 (N_17989,N_17592,N_17702);
xor U17990 (N_17990,N_17513,N_17710);
or U17991 (N_17991,N_17652,N_17656);
xor U17992 (N_17992,N_17542,N_17527);
nor U17993 (N_17993,N_17581,N_17514);
and U17994 (N_17994,N_17596,N_17674);
or U17995 (N_17995,N_17697,N_17522);
nor U17996 (N_17996,N_17700,N_17580);
xor U17997 (N_17997,N_17725,N_17590);
nor U17998 (N_17998,N_17536,N_17502);
xnor U17999 (N_17999,N_17689,N_17501);
and U18000 (N_18000,N_17982,N_17828);
and U18001 (N_18001,N_17841,N_17784);
xor U18002 (N_18002,N_17955,N_17879);
or U18003 (N_18003,N_17781,N_17911);
nand U18004 (N_18004,N_17752,N_17948);
xor U18005 (N_18005,N_17882,N_17874);
and U18006 (N_18006,N_17860,N_17919);
and U18007 (N_18007,N_17968,N_17931);
and U18008 (N_18008,N_17960,N_17765);
xnor U18009 (N_18009,N_17913,N_17839);
or U18010 (N_18010,N_17909,N_17923);
and U18011 (N_18011,N_17887,N_17917);
xor U18012 (N_18012,N_17946,N_17949);
and U18013 (N_18013,N_17844,N_17893);
and U18014 (N_18014,N_17975,N_17997);
and U18015 (N_18015,N_17869,N_17876);
and U18016 (N_18016,N_17832,N_17936);
xnor U18017 (N_18017,N_17950,N_17932);
or U18018 (N_18018,N_17782,N_17957);
and U18019 (N_18019,N_17827,N_17958);
xnor U18020 (N_18020,N_17941,N_17978);
xor U18021 (N_18021,N_17868,N_17811);
or U18022 (N_18022,N_17859,N_17863);
xor U18023 (N_18023,N_17956,N_17902);
and U18024 (N_18024,N_17779,N_17865);
or U18025 (N_18025,N_17812,N_17980);
xor U18026 (N_18026,N_17750,N_17773);
nor U18027 (N_18027,N_17878,N_17954);
and U18028 (N_18028,N_17891,N_17915);
nor U18029 (N_18029,N_17979,N_17873);
or U18030 (N_18030,N_17764,N_17988);
nand U18031 (N_18031,N_17774,N_17961);
xnor U18032 (N_18032,N_17989,N_17758);
nor U18033 (N_18033,N_17904,N_17757);
and U18034 (N_18034,N_17830,N_17974);
or U18035 (N_18035,N_17787,N_17751);
or U18036 (N_18036,N_17938,N_17759);
and U18037 (N_18037,N_17761,N_17835);
xnor U18038 (N_18038,N_17867,N_17994);
nor U18039 (N_18039,N_17918,N_17846);
and U18040 (N_18040,N_17984,N_17944);
xnor U18041 (N_18041,N_17840,N_17864);
nand U18042 (N_18042,N_17836,N_17753);
nor U18043 (N_18043,N_17940,N_17854);
xnor U18044 (N_18044,N_17888,N_17924);
nand U18045 (N_18045,N_17807,N_17837);
and U18046 (N_18046,N_17772,N_17763);
xnor U18047 (N_18047,N_17780,N_17770);
and U18048 (N_18048,N_17826,N_17922);
nand U18049 (N_18049,N_17755,N_17767);
nor U18050 (N_18050,N_17991,N_17792);
xnor U18051 (N_18051,N_17806,N_17999);
and U18052 (N_18052,N_17793,N_17816);
nor U18053 (N_18053,N_17791,N_17762);
or U18054 (N_18054,N_17908,N_17995);
nor U18055 (N_18055,N_17848,N_17894);
and U18056 (N_18056,N_17800,N_17905);
xor U18057 (N_18057,N_17834,N_17886);
and U18058 (N_18058,N_17880,N_17829);
or U18059 (N_18059,N_17756,N_17766);
nor U18060 (N_18060,N_17921,N_17771);
nand U18061 (N_18061,N_17953,N_17866);
or U18062 (N_18062,N_17945,N_17900);
xor U18063 (N_18063,N_17783,N_17809);
nand U18064 (N_18064,N_17799,N_17796);
nand U18065 (N_18065,N_17855,N_17943);
or U18066 (N_18066,N_17778,N_17817);
or U18067 (N_18067,N_17754,N_17852);
nand U18068 (N_18068,N_17805,N_17804);
xor U18069 (N_18069,N_17933,N_17898);
and U18070 (N_18070,N_17910,N_17903);
or U18071 (N_18071,N_17897,N_17843);
or U18072 (N_18072,N_17976,N_17973);
nor U18073 (N_18073,N_17883,N_17824);
or U18074 (N_18074,N_17896,N_17937);
nor U18075 (N_18075,N_17930,N_17785);
nand U18076 (N_18076,N_17769,N_17890);
nand U18077 (N_18077,N_17987,N_17986);
or U18078 (N_18078,N_17998,N_17907);
or U18079 (N_18079,N_17990,N_17971);
or U18080 (N_18080,N_17858,N_17789);
or U18081 (N_18081,N_17916,N_17985);
xor U18082 (N_18082,N_17795,N_17966);
and U18083 (N_18083,N_17821,N_17925);
nor U18084 (N_18084,N_17962,N_17967);
xnor U18085 (N_18085,N_17776,N_17853);
nor U18086 (N_18086,N_17920,N_17798);
or U18087 (N_18087,N_17808,N_17881);
or U18088 (N_18088,N_17872,N_17803);
xor U18089 (N_18089,N_17768,N_17815);
nor U18090 (N_18090,N_17951,N_17856);
xnor U18091 (N_18091,N_17845,N_17877);
xor U18092 (N_18092,N_17777,N_17810);
and U18093 (N_18093,N_17790,N_17901);
xor U18094 (N_18094,N_17788,N_17794);
and U18095 (N_18095,N_17814,N_17942);
xor U18096 (N_18096,N_17786,N_17849);
and U18097 (N_18097,N_17927,N_17851);
or U18098 (N_18098,N_17965,N_17947);
nand U18099 (N_18099,N_17939,N_17802);
or U18100 (N_18100,N_17914,N_17822);
and U18101 (N_18101,N_17972,N_17838);
nand U18102 (N_18102,N_17963,N_17825);
and U18103 (N_18103,N_17833,N_17797);
xnor U18104 (N_18104,N_17875,N_17906);
or U18105 (N_18105,N_17823,N_17934);
or U18106 (N_18106,N_17885,N_17964);
xnor U18107 (N_18107,N_17760,N_17977);
or U18108 (N_18108,N_17935,N_17818);
and U18109 (N_18109,N_17969,N_17970);
nor U18110 (N_18110,N_17959,N_17847);
nand U18111 (N_18111,N_17993,N_17899);
nand U18112 (N_18112,N_17850,N_17861);
nand U18113 (N_18113,N_17912,N_17820);
and U18114 (N_18114,N_17813,N_17996);
nor U18115 (N_18115,N_17871,N_17926);
nand U18116 (N_18116,N_17895,N_17801);
or U18117 (N_18117,N_17870,N_17819);
and U18118 (N_18118,N_17884,N_17983);
xnor U18119 (N_18119,N_17929,N_17775);
and U18120 (N_18120,N_17889,N_17892);
nor U18121 (N_18121,N_17842,N_17981);
xnor U18122 (N_18122,N_17952,N_17857);
and U18123 (N_18123,N_17928,N_17862);
or U18124 (N_18124,N_17831,N_17992);
and U18125 (N_18125,N_17774,N_17770);
and U18126 (N_18126,N_17843,N_17982);
or U18127 (N_18127,N_17860,N_17902);
and U18128 (N_18128,N_17973,N_17850);
and U18129 (N_18129,N_17771,N_17867);
or U18130 (N_18130,N_17964,N_17781);
and U18131 (N_18131,N_17774,N_17798);
xor U18132 (N_18132,N_17813,N_17868);
or U18133 (N_18133,N_17916,N_17978);
nand U18134 (N_18134,N_17847,N_17895);
xor U18135 (N_18135,N_17949,N_17929);
or U18136 (N_18136,N_17787,N_17851);
nor U18137 (N_18137,N_17856,N_17919);
xnor U18138 (N_18138,N_17768,N_17854);
or U18139 (N_18139,N_17760,N_17879);
xnor U18140 (N_18140,N_17929,N_17861);
or U18141 (N_18141,N_17828,N_17974);
nor U18142 (N_18142,N_17937,N_17947);
or U18143 (N_18143,N_17988,N_17908);
or U18144 (N_18144,N_17802,N_17908);
and U18145 (N_18145,N_17781,N_17917);
or U18146 (N_18146,N_17981,N_17755);
nand U18147 (N_18147,N_17824,N_17948);
or U18148 (N_18148,N_17799,N_17900);
xnor U18149 (N_18149,N_17943,N_17763);
nand U18150 (N_18150,N_17908,N_17965);
nand U18151 (N_18151,N_17982,N_17767);
and U18152 (N_18152,N_17830,N_17807);
and U18153 (N_18153,N_17917,N_17857);
and U18154 (N_18154,N_17926,N_17994);
nor U18155 (N_18155,N_17996,N_17778);
or U18156 (N_18156,N_17827,N_17954);
and U18157 (N_18157,N_17974,N_17924);
nor U18158 (N_18158,N_17788,N_17853);
nor U18159 (N_18159,N_17938,N_17843);
and U18160 (N_18160,N_17869,N_17858);
or U18161 (N_18161,N_17783,N_17768);
nor U18162 (N_18162,N_17754,N_17793);
nor U18163 (N_18163,N_17955,N_17999);
or U18164 (N_18164,N_17813,N_17956);
xor U18165 (N_18165,N_17958,N_17876);
xnor U18166 (N_18166,N_17810,N_17982);
or U18167 (N_18167,N_17929,N_17767);
xor U18168 (N_18168,N_17805,N_17838);
xor U18169 (N_18169,N_17994,N_17938);
xor U18170 (N_18170,N_17935,N_17971);
nor U18171 (N_18171,N_17883,N_17793);
nor U18172 (N_18172,N_17807,N_17760);
xnor U18173 (N_18173,N_17841,N_17821);
or U18174 (N_18174,N_17965,N_17857);
or U18175 (N_18175,N_17877,N_17944);
xor U18176 (N_18176,N_17982,N_17951);
xor U18177 (N_18177,N_17788,N_17984);
or U18178 (N_18178,N_17989,N_17926);
or U18179 (N_18179,N_17976,N_17846);
nor U18180 (N_18180,N_17824,N_17892);
nor U18181 (N_18181,N_17777,N_17949);
nor U18182 (N_18182,N_17903,N_17943);
or U18183 (N_18183,N_17851,N_17823);
and U18184 (N_18184,N_17803,N_17952);
xnor U18185 (N_18185,N_17837,N_17846);
nor U18186 (N_18186,N_17811,N_17875);
and U18187 (N_18187,N_17879,N_17916);
xnor U18188 (N_18188,N_17800,N_17972);
nand U18189 (N_18189,N_17969,N_17856);
nand U18190 (N_18190,N_17956,N_17900);
and U18191 (N_18191,N_17825,N_17805);
nor U18192 (N_18192,N_17870,N_17791);
or U18193 (N_18193,N_17982,N_17942);
or U18194 (N_18194,N_17946,N_17977);
nor U18195 (N_18195,N_17768,N_17931);
and U18196 (N_18196,N_17751,N_17884);
or U18197 (N_18197,N_17775,N_17908);
xor U18198 (N_18198,N_17798,N_17966);
and U18199 (N_18199,N_17906,N_17762);
nor U18200 (N_18200,N_17934,N_17870);
nand U18201 (N_18201,N_17920,N_17938);
xor U18202 (N_18202,N_17943,N_17929);
nor U18203 (N_18203,N_17950,N_17963);
and U18204 (N_18204,N_17868,N_17898);
nand U18205 (N_18205,N_17797,N_17994);
or U18206 (N_18206,N_17768,N_17801);
nor U18207 (N_18207,N_17819,N_17825);
or U18208 (N_18208,N_17906,N_17944);
or U18209 (N_18209,N_17915,N_17841);
xnor U18210 (N_18210,N_17831,N_17937);
or U18211 (N_18211,N_17786,N_17870);
nor U18212 (N_18212,N_17888,N_17842);
and U18213 (N_18213,N_17921,N_17855);
nand U18214 (N_18214,N_17776,N_17765);
nand U18215 (N_18215,N_17903,N_17803);
nand U18216 (N_18216,N_17894,N_17878);
xnor U18217 (N_18217,N_17904,N_17791);
or U18218 (N_18218,N_17753,N_17966);
xnor U18219 (N_18219,N_17870,N_17811);
or U18220 (N_18220,N_17943,N_17761);
and U18221 (N_18221,N_17895,N_17850);
nand U18222 (N_18222,N_17934,N_17905);
or U18223 (N_18223,N_17766,N_17842);
or U18224 (N_18224,N_17837,N_17804);
and U18225 (N_18225,N_17868,N_17788);
nand U18226 (N_18226,N_17821,N_17853);
nor U18227 (N_18227,N_17880,N_17877);
and U18228 (N_18228,N_17800,N_17962);
xor U18229 (N_18229,N_17841,N_17953);
nand U18230 (N_18230,N_17877,N_17810);
nor U18231 (N_18231,N_17994,N_17838);
and U18232 (N_18232,N_17869,N_17804);
nand U18233 (N_18233,N_17782,N_17830);
xnor U18234 (N_18234,N_17764,N_17858);
or U18235 (N_18235,N_17985,N_17952);
nand U18236 (N_18236,N_17822,N_17793);
xor U18237 (N_18237,N_17848,N_17892);
nor U18238 (N_18238,N_17896,N_17959);
nor U18239 (N_18239,N_17878,N_17801);
nor U18240 (N_18240,N_17872,N_17787);
and U18241 (N_18241,N_17956,N_17927);
nand U18242 (N_18242,N_17929,N_17757);
xnor U18243 (N_18243,N_17836,N_17799);
xor U18244 (N_18244,N_17812,N_17770);
xor U18245 (N_18245,N_17894,N_17896);
nor U18246 (N_18246,N_17799,N_17944);
or U18247 (N_18247,N_17979,N_17913);
and U18248 (N_18248,N_17846,N_17869);
and U18249 (N_18249,N_17791,N_17786);
nor U18250 (N_18250,N_18168,N_18007);
and U18251 (N_18251,N_18009,N_18178);
or U18252 (N_18252,N_18030,N_18187);
xor U18253 (N_18253,N_18025,N_18125);
and U18254 (N_18254,N_18219,N_18065);
nand U18255 (N_18255,N_18183,N_18026);
nor U18256 (N_18256,N_18239,N_18121);
and U18257 (N_18257,N_18217,N_18015);
xnor U18258 (N_18258,N_18222,N_18218);
nand U18259 (N_18259,N_18014,N_18016);
and U18260 (N_18260,N_18197,N_18024);
nor U18261 (N_18261,N_18001,N_18203);
nor U18262 (N_18262,N_18116,N_18227);
xnor U18263 (N_18263,N_18027,N_18127);
xnor U18264 (N_18264,N_18237,N_18072);
nor U18265 (N_18265,N_18152,N_18108);
xnor U18266 (N_18266,N_18191,N_18079);
nor U18267 (N_18267,N_18155,N_18151);
or U18268 (N_18268,N_18171,N_18149);
nor U18269 (N_18269,N_18081,N_18164);
nand U18270 (N_18270,N_18226,N_18051);
or U18271 (N_18271,N_18002,N_18068);
xor U18272 (N_18272,N_18229,N_18181);
or U18273 (N_18273,N_18193,N_18052);
or U18274 (N_18274,N_18141,N_18192);
nor U18275 (N_18275,N_18048,N_18156);
nor U18276 (N_18276,N_18120,N_18209);
nand U18277 (N_18277,N_18163,N_18180);
nor U18278 (N_18278,N_18160,N_18131);
or U18279 (N_18279,N_18088,N_18043);
and U18280 (N_18280,N_18240,N_18049);
xnor U18281 (N_18281,N_18169,N_18008);
nor U18282 (N_18282,N_18038,N_18235);
and U18283 (N_18283,N_18135,N_18147);
or U18284 (N_18284,N_18221,N_18159);
nand U18285 (N_18285,N_18101,N_18073);
xnor U18286 (N_18286,N_18000,N_18039);
nand U18287 (N_18287,N_18084,N_18078);
nor U18288 (N_18288,N_18115,N_18211);
xnor U18289 (N_18289,N_18182,N_18041);
or U18290 (N_18290,N_18003,N_18213);
nor U18291 (N_18291,N_18104,N_18242);
nor U18292 (N_18292,N_18053,N_18050);
xor U18293 (N_18293,N_18139,N_18200);
nor U18294 (N_18294,N_18035,N_18148);
nand U18295 (N_18295,N_18154,N_18106);
nand U18296 (N_18296,N_18208,N_18214);
xor U18297 (N_18297,N_18201,N_18165);
or U18298 (N_18298,N_18249,N_18013);
or U18299 (N_18299,N_18138,N_18080);
nor U18300 (N_18300,N_18145,N_18146);
and U18301 (N_18301,N_18188,N_18062);
and U18302 (N_18302,N_18074,N_18196);
or U18303 (N_18303,N_18109,N_18118);
and U18304 (N_18304,N_18224,N_18021);
xnor U18305 (N_18305,N_18114,N_18132);
nor U18306 (N_18306,N_18045,N_18179);
or U18307 (N_18307,N_18018,N_18100);
nor U18308 (N_18308,N_18142,N_18020);
xor U18309 (N_18309,N_18089,N_18085);
nand U18310 (N_18310,N_18158,N_18011);
nand U18311 (N_18311,N_18238,N_18096);
and U18312 (N_18312,N_18059,N_18103);
nand U18313 (N_18313,N_18199,N_18105);
nand U18314 (N_18314,N_18090,N_18093);
and U18315 (N_18315,N_18150,N_18184);
nand U18316 (N_18316,N_18231,N_18205);
nor U18317 (N_18317,N_18243,N_18069);
and U18318 (N_18318,N_18206,N_18056);
nor U18319 (N_18319,N_18212,N_18128);
nand U18320 (N_18320,N_18225,N_18006);
nand U18321 (N_18321,N_18143,N_18233);
xor U18322 (N_18322,N_18004,N_18244);
and U18323 (N_18323,N_18210,N_18070);
or U18324 (N_18324,N_18023,N_18173);
xor U18325 (N_18325,N_18012,N_18195);
nand U18326 (N_18326,N_18130,N_18055);
and U18327 (N_18327,N_18044,N_18019);
and U18328 (N_18328,N_18058,N_18134);
nor U18329 (N_18329,N_18246,N_18063);
or U18330 (N_18330,N_18133,N_18034);
or U18331 (N_18331,N_18102,N_18232);
nor U18332 (N_18332,N_18247,N_18112);
xnor U18333 (N_18333,N_18060,N_18144);
xor U18334 (N_18334,N_18075,N_18234);
or U18335 (N_18335,N_18174,N_18033);
and U18336 (N_18336,N_18046,N_18129);
or U18337 (N_18337,N_18136,N_18198);
nand U18338 (N_18338,N_18066,N_18057);
nor U18339 (N_18339,N_18153,N_18177);
nor U18340 (N_18340,N_18175,N_18029);
nand U18341 (N_18341,N_18017,N_18220);
xnor U18342 (N_18342,N_18124,N_18086);
xor U18343 (N_18343,N_18216,N_18094);
nand U18344 (N_18344,N_18037,N_18157);
nor U18345 (N_18345,N_18137,N_18228);
nand U18346 (N_18346,N_18236,N_18167);
or U18347 (N_18347,N_18166,N_18241);
nor U18348 (N_18348,N_18185,N_18083);
and U18349 (N_18349,N_18189,N_18176);
xor U18350 (N_18350,N_18061,N_18202);
and U18351 (N_18351,N_18162,N_18194);
nor U18352 (N_18352,N_18190,N_18036);
nor U18353 (N_18353,N_18032,N_18067);
nor U18354 (N_18354,N_18170,N_18126);
or U18355 (N_18355,N_18064,N_18161);
and U18356 (N_18356,N_18119,N_18113);
or U18357 (N_18357,N_18215,N_18054);
and U18358 (N_18358,N_18140,N_18117);
and U18359 (N_18359,N_18022,N_18091);
nor U18360 (N_18360,N_18095,N_18087);
nand U18361 (N_18361,N_18110,N_18097);
xnor U18362 (N_18362,N_18040,N_18107);
nor U18363 (N_18363,N_18071,N_18099);
xor U18364 (N_18364,N_18076,N_18082);
xor U18365 (N_18365,N_18092,N_18123);
nor U18366 (N_18366,N_18248,N_18031);
nand U18367 (N_18367,N_18077,N_18122);
nand U18368 (N_18368,N_18207,N_18028);
nand U18369 (N_18369,N_18186,N_18230);
xnor U18370 (N_18370,N_18245,N_18223);
nor U18371 (N_18371,N_18098,N_18010);
or U18372 (N_18372,N_18047,N_18042);
xor U18373 (N_18373,N_18204,N_18172);
and U18374 (N_18374,N_18005,N_18111);
nand U18375 (N_18375,N_18123,N_18215);
nor U18376 (N_18376,N_18162,N_18189);
nor U18377 (N_18377,N_18235,N_18042);
and U18378 (N_18378,N_18035,N_18009);
nand U18379 (N_18379,N_18220,N_18074);
or U18380 (N_18380,N_18225,N_18240);
xor U18381 (N_18381,N_18132,N_18074);
nand U18382 (N_18382,N_18065,N_18224);
xnor U18383 (N_18383,N_18210,N_18224);
nor U18384 (N_18384,N_18121,N_18114);
or U18385 (N_18385,N_18121,N_18089);
and U18386 (N_18386,N_18237,N_18109);
and U18387 (N_18387,N_18186,N_18031);
or U18388 (N_18388,N_18205,N_18218);
nand U18389 (N_18389,N_18090,N_18139);
xnor U18390 (N_18390,N_18147,N_18059);
nor U18391 (N_18391,N_18075,N_18138);
xor U18392 (N_18392,N_18128,N_18247);
and U18393 (N_18393,N_18123,N_18046);
nor U18394 (N_18394,N_18050,N_18175);
nor U18395 (N_18395,N_18192,N_18105);
nor U18396 (N_18396,N_18110,N_18131);
xor U18397 (N_18397,N_18057,N_18038);
or U18398 (N_18398,N_18080,N_18021);
nand U18399 (N_18399,N_18206,N_18021);
or U18400 (N_18400,N_18041,N_18130);
xor U18401 (N_18401,N_18015,N_18095);
nor U18402 (N_18402,N_18123,N_18249);
xor U18403 (N_18403,N_18193,N_18077);
nor U18404 (N_18404,N_18106,N_18192);
nand U18405 (N_18405,N_18033,N_18081);
and U18406 (N_18406,N_18170,N_18006);
and U18407 (N_18407,N_18099,N_18083);
nand U18408 (N_18408,N_18185,N_18169);
xor U18409 (N_18409,N_18070,N_18139);
and U18410 (N_18410,N_18024,N_18016);
nand U18411 (N_18411,N_18225,N_18000);
xor U18412 (N_18412,N_18091,N_18196);
and U18413 (N_18413,N_18243,N_18162);
and U18414 (N_18414,N_18150,N_18045);
nor U18415 (N_18415,N_18128,N_18036);
or U18416 (N_18416,N_18058,N_18127);
or U18417 (N_18417,N_18195,N_18037);
xor U18418 (N_18418,N_18156,N_18227);
or U18419 (N_18419,N_18053,N_18230);
xor U18420 (N_18420,N_18218,N_18234);
or U18421 (N_18421,N_18032,N_18234);
xnor U18422 (N_18422,N_18224,N_18032);
and U18423 (N_18423,N_18226,N_18080);
or U18424 (N_18424,N_18027,N_18234);
or U18425 (N_18425,N_18066,N_18085);
nor U18426 (N_18426,N_18233,N_18176);
or U18427 (N_18427,N_18126,N_18033);
nor U18428 (N_18428,N_18026,N_18087);
or U18429 (N_18429,N_18247,N_18217);
or U18430 (N_18430,N_18228,N_18033);
xnor U18431 (N_18431,N_18156,N_18193);
xor U18432 (N_18432,N_18113,N_18225);
or U18433 (N_18433,N_18230,N_18201);
xor U18434 (N_18434,N_18119,N_18024);
nand U18435 (N_18435,N_18216,N_18111);
and U18436 (N_18436,N_18146,N_18022);
or U18437 (N_18437,N_18030,N_18233);
nand U18438 (N_18438,N_18148,N_18074);
or U18439 (N_18439,N_18091,N_18239);
nor U18440 (N_18440,N_18132,N_18077);
xor U18441 (N_18441,N_18050,N_18038);
nand U18442 (N_18442,N_18104,N_18065);
xnor U18443 (N_18443,N_18144,N_18110);
nor U18444 (N_18444,N_18028,N_18023);
or U18445 (N_18445,N_18092,N_18229);
nand U18446 (N_18446,N_18092,N_18100);
nor U18447 (N_18447,N_18044,N_18159);
nor U18448 (N_18448,N_18031,N_18222);
or U18449 (N_18449,N_18068,N_18217);
or U18450 (N_18450,N_18049,N_18206);
nand U18451 (N_18451,N_18156,N_18057);
nor U18452 (N_18452,N_18142,N_18217);
or U18453 (N_18453,N_18182,N_18109);
nor U18454 (N_18454,N_18068,N_18219);
and U18455 (N_18455,N_18202,N_18002);
nand U18456 (N_18456,N_18000,N_18010);
xor U18457 (N_18457,N_18233,N_18183);
xnor U18458 (N_18458,N_18126,N_18128);
nor U18459 (N_18459,N_18237,N_18171);
nand U18460 (N_18460,N_18196,N_18044);
nand U18461 (N_18461,N_18174,N_18085);
or U18462 (N_18462,N_18210,N_18241);
nor U18463 (N_18463,N_18024,N_18187);
or U18464 (N_18464,N_18069,N_18150);
xor U18465 (N_18465,N_18225,N_18101);
nor U18466 (N_18466,N_18134,N_18021);
xnor U18467 (N_18467,N_18098,N_18093);
and U18468 (N_18468,N_18109,N_18078);
nand U18469 (N_18469,N_18192,N_18013);
and U18470 (N_18470,N_18183,N_18100);
xnor U18471 (N_18471,N_18177,N_18235);
nor U18472 (N_18472,N_18176,N_18135);
nand U18473 (N_18473,N_18210,N_18163);
or U18474 (N_18474,N_18130,N_18176);
nor U18475 (N_18475,N_18129,N_18127);
or U18476 (N_18476,N_18196,N_18097);
nor U18477 (N_18477,N_18071,N_18123);
xnor U18478 (N_18478,N_18175,N_18128);
nand U18479 (N_18479,N_18075,N_18091);
or U18480 (N_18480,N_18073,N_18017);
xor U18481 (N_18481,N_18054,N_18185);
nand U18482 (N_18482,N_18092,N_18213);
or U18483 (N_18483,N_18049,N_18210);
or U18484 (N_18484,N_18091,N_18113);
nor U18485 (N_18485,N_18240,N_18231);
nor U18486 (N_18486,N_18010,N_18051);
nor U18487 (N_18487,N_18223,N_18139);
or U18488 (N_18488,N_18004,N_18053);
or U18489 (N_18489,N_18081,N_18020);
or U18490 (N_18490,N_18122,N_18181);
nor U18491 (N_18491,N_18160,N_18031);
nor U18492 (N_18492,N_18123,N_18081);
and U18493 (N_18493,N_18176,N_18181);
nand U18494 (N_18494,N_18147,N_18177);
and U18495 (N_18495,N_18003,N_18091);
and U18496 (N_18496,N_18239,N_18146);
xor U18497 (N_18497,N_18193,N_18013);
and U18498 (N_18498,N_18211,N_18163);
xor U18499 (N_18499,N_18200,N_18030);
nor U18500 (N_18500,N_18413,N_18475);
or U18501 (N_18501,N_18493,N_18452);
nand U18502 (N_18502,N_18395,N_18321);
nand U18503 (N_18503,N_18444,N_18343);
or U18504 (N_18504,N_18341,N_18455);
or U18505 (N_18505,N_18316,N_18358);
or U18506 (N_18506,N_18253,N_18370);
xor U18507 (N_18507,N_18438,N_18274);
nor U18508 (N_18508,N_18404,N_18350);
or U18509 (N_18509,N_18342,N_18313);
or U18510 (N_18510,N_18406,N_18305);
and U18511 (N_18511,N_18340,N_18448);
xnor U18512 (N_18512,N_18257,N_18458);
or U18513 (N_18513,N_18272,N_18380);
or U18514 (N_18514,N_18471,N_18351);
or U18515 (N_18515,N_18287,N_18259);
and U18516 (N_18516,N_18388,N_18472);
or U18517 (N_18517,N_18385,N_18330);
and U18518 (N_18518,N_18394,N_18386);
nor U18519 (N_18519,N_18379,N_18424);
and U18520 (N_18520,N_18466,N_18401);
nand U18521 (N_18521,N_18271,N_18353);
or U18522 (N_18522,N_18348,N_18312);
nor U18523 (N_18523,N_18415,N_18267);
and U18524 (N_18524,N_18450,N_18322);
xnor U18525 (N_18525,N_18431,N_18467);
xor U18526 (N_18526,N_18295,N_18464);
nor U18527 (N_18527,N_18275,N_18279);
xor U18528 (N_18528,N_18364,N_18479);
nor U18529 (N_18529,N_18308,N_18282);
and U18530 (N_18530,N_18426,N_18349);
or U18531 (N_18531,N_18473,N_18463);
or U18532 (N_18532,N_18266,N_18314);
or U18533 (N_18533,N_18390,N_18293);
and U18534 (N_18534,N_18446,N_18262);
or U18535 (N_18535,N_18260,N_18344);
xnor U18536 (N_18536,N_18252,N_18309);
nand U18537 (N_18537,N_18373,N_18442);
xnor U18538 (N_18538,N_18420,N_18317);
xor U18539 (N_18539,N_18368,N_18276);
or U18540 (N_18540,N_18382,N_18427);
xor U18541 (N_18541,N_18434,N_18294);
nand U18542 (N_18542,N_18410,N_18497);
or U18543 (N_18543,N_18453,N_18425);
xnor U18544 (N_18544,N_18255,N_18430);
or U18545 (N_18545,N_18359,N_18355);
xor U18546 (N_18546,N_18481,N_18469);
xnor U18547 (N_18547,N_18254,N_18303);
nand U18548 (N_18548,N_18311,N_18422);
and U18549 (N_18549,N_18407,N_18457);
xor U18550 (N_18550,N_18449,N_18398);
nand U18551 (N_18551,N_18286,N_18374);
xnor U18552 (N_18552,N_18357,N_18432);
and U18553 (N_18553,N_18423,N_18402);
and U18554 (N_18554,N_18494,N_18456);
nand U18555 (N_18555,N_18334,N_18400);
nor U18556 (N_18556,N_18387,N_18347);
xnor U18557 (N_18557,N_18338,N_18483);
nor U18558 (N_18558,N_18482,N_18278);
xnor U18559 (N_18559,N_18478,N_18315);
nand U18560 (N_18560,N_18320,N_18288);
nor U18561 (N_18561,N_18470,N_18412);
or U18562 (N_18562,N_18496,N_18462);
xnor U18563 (N_18563,N_18263,N_18346);
nor U18564 (N_18564,N_18325,N_18437);
or U18565 (N_18565,N_18391,N_18264);
nor U18566 (N_18566,N_18433,N_18290);
xnor U18567 (N_18567,N_18332,N_18445);
and U18568 (N_18568,N_18440,N_18337);
xor U18569 (N_18569,N_18280,N_18299);
xnor U18570 (N_18570,N_18258,N_18488);
nor U18571 (N_18571,N_18414,N_18285);
xor U18572 (N_18572,N_18283,N_18459);
nand U18573 (N_18573,N_18384,N_18339);
nor U18574 (N_18574,N_18490,N_18408);
nor U18575 (N_18575,N_18250,N_18298);
or U18576 (N_18576,N_18327,N_18381);
xnor U18577 (N_18577,N_18273,N_18292);
or U18578 (N_18578,N_18416,N_18336);
nor U18579 (N_18579,N_18492,N_18329);
and U18580 (N_18580,N_18435,N_18465);
xnor U18581 (N_18581,N_18460,N_18461);
and U18582 (N_18582,N_18405,N_18306);
nor U18583 (N_18583,N_18474,N_18477);
or U18584 (N_18584,N_18403,N_18360);
or U18585 (N_18585,N_18451,N_18326);
xor U18586 (N_18586,N_18447,N_18269);
nand U18587 (N_18587,N_18439,N_18376);
or U18588 (N_18588,N_18399,N_18251);
nand U18589 (N_18589,N_18480,N_18454);
and U18590 (N_18590,N_18369,N_18281);
and U18591 (N_18591,N_18307,N_18345);
nor U18592 (N_18592,N_18277,N_18378);
nand U18593 (N_18593,N_18371,N_18396);
nand U18594 (N_18594,N_18495,N_18383);
xor U18595 (N_18595,N_18367,N_18261);
or U18596 (N_18596,N_18323,N_18485);
and U18597 (N_18597,N_18491,N_18476);
and U18598 (N_18598,N_18468,N_18256);
nor U18599 (N_18599,N_18304,N_18409);
nand U18600 (N_18600,N_18310,N_18328);
nor U18601 (N_18601,N_18361,N_18429);
or U18602 (N_18602,N_18421,N_18411);
or U18603 (N_18603,N_18289,N_18441);
nand U18604 (N_18604,N_18375,N_18397);
and U18605 (N_18605,N_18291,N_18319);
nor U18606 (N_18606,N_18302,N_18365);
and U18607 (N_18607,N_18333,N_18352);
and U18608 (N_18608,N_18268,N_18265);
nor U18609 (N_18609,N_18366,N_18284);
and U18610 (N_18610,N_18362,N_18331);
nand U18611 (N_18611,N_18428,N_18363);
and U18612 (N_18612,N_18498,N_18300);
nand U18613 (N_18613,N_18487,N_18489);
and U18614 (N_18614,N_18324,N_18389);
or U18615 (N_18615,N_18301,N_18377);
nand U18616 (N_18616,N_18499,N_18484);
and U18617 (N_18617,N_18356,N_18335);
xor U18618 (N_18618,N_18296,N_18372);
and U18619 (N_18619,N_18392,N_18436);
and U18620 (N_18620,N_18270,N_18297);
xnor U18621 (N_18621,N_18418,N_18443);
xnor U18622 (N_18622,N_18417,N_18393);
and U18623 (N_18623,N_18419,N_18318);
and U18624 (N_18624,N_18354,N_18486);
xor U18625 (N_18625,N_18495,N_18443);
nand U18626 (N_18626,N_18419,N_18399);
or U18627 (N_18627,N_18464,N_18259);
nor U18628 (N_18628,N_18469,N_18486);
xnor U18629 (N_18629,N_18350,N_18483);
and U18630 (N_18630,N_18479,N_18455);
or U18631 (N_18631,N_18424,N_18481);
or U18632 (N_18632,N_18408,N_18365);
and U18633 (N_18633,N_18332,N_18404);
nand U18634 (N_18634,N_18366,N_18378);
nor U18635 (N_18635,N_18442,N_18297);
and U18636 (N_18636,N_18491,N_18271);
or U18637 (N_18637,N_18308,N_18318);
nand U18638 (N_18638,N_18368,N_18337);
nor U18639 (N_18639,N_18389,N_18483);
nand U18640 (N_18640,N_18257,N_18379);
xor U18641 (N_18641,N_18342,N_18392);
nor U18642 (N_18642,N_18357,N_18271);
and U18643 (N_18643,N_18273,N_18436);
xnor U18644 (N_18644,N_18414,N_18429);
and U18645 (N_18645,N_18425,N_18395);
xnor U18646 (N_18646,N_18423,N_18427);
or U18647 (N_18647,N_18488,N_18423);
nand U18648 (N_18648,N_18399,N_18458);
nand U18649 (N_18649,N_18452,N_18387);
nand U18650 (N_18650,N_18372,N_18252);
xnor U18651 (N_18651,N_18276,N_18436);
and U18652 (N_18652,N_18394,N_18339);
nand U18653 (N_18653,N_18372,N_18277);
xnor U18654 (N_18654,N_18383,N_18268);
nor U18655 (N_18655,N_18277,N_18345);
nand U18656 (N_18656,N_18463,N_18295);
nor U18657 (N_18657,N_18362,N_18269);
and U18658 (N_18658,N_18310,N_18251);
and U18659 (N_18659,N_18485,N_18378);
nand U18660 (N_18660,N_18353,N_18435);
nand U18661 (N_18661,N_18449,N_18458);
nor U18662 (N_18662,N_18424,N_18301);
nand U18663 (N_18663,N_18338,N_18422);
and U18664 (N_18664,N_18440,N_18476);
xor U18665 (N_18665,N_18452,N_18295);
xnor U18666 (N_18666,N_18337,N_18283);
or U18667 (N_18667,N_18301,N_18479);
nand U18668 (N_18668,N_18260,N_18490);
and U18669 (N_18669,N_18436,N_18261);
nand U18670 (N_18670,N_18470,N_18424);
and U18671 (N_18671,N_18407,N_18448);
nand U18672 (N_18672,N_18422,N_18465);
xor U18673 (N_18673,N_18324,N_18390);
and U18674 (N_18674,N_18440,N_18444);
and U18675 (N_18675,N_18279,N_18284);
xor U18676 (N_18676,N_18306,N_18453);
or U18677 (N_18677,N_18440,N_18335);
nand U18678 (N_18678,N_18275,N_18314);
nand U18679 (N_18679,N_18494,N_18477);
and U18680 (N_18680,N_18409,N_18382);
xor U18681 (N_18681,N_18341,N_18362);
and U18682 (N_18682,N_18379,N_18444);
and U18683 (N_18683,N_18352,N_18353);
and U18684 (N_18684,N_18487,N_18403);
and U18685 (N_18685,N_18499,N_18401);
xor U18686 (N_18686,N_18456,N_18466);
nor U18687 (N_18687,N_18468,N_18447);
nand U18688 (N_18688,N_18461,N_18392);
and U18689 (N_18689,N_18380,N_18339);
nand U18690 (N_18690,N_18252,N_18351);
nand U18691 (N_18691,N_18385,N_18435);
and U18692 (N_18692,N_18467,N_18475);
or U18693 (N_18693,N_18334,N_18316);
or U18694 (N_18694,N_18300,N_18427);
nor U18695 (N_18695,N_18382,N_18476);
and U18696 (N_18696,N_18379,N_18463);
nand U18697 (N_18697,N_18411,N_18392);
and U18698 (N_18698,N_18260,N_18434);
nand U18699 (N_18699,N_18395,N_18485);
xnor U18700 (N_18700,N_18359,N_18282);
and U18701 (N_18701,N_18339,N_18391);
or U18702 (N_18702,N_18272,N_18414);
xor U18703 (N_18703,N_18384,N_18471);
and U18704 (N_18704,N_18277,N_18267);
or U18705 (N_18705,N_18301,N_18481);
xor U18706 (N_18706,N_18285,N_18299);
and U18707 (N_18707,N_18485,N_18272);
and U18708 (N_18708,N_18279,N_18363);
nor U18709 (N_18709,N_18330,N_18476);
and U18710 (N_18710,N_18498,N_18428);
or U18711 (N_18711,N_18460,N_18298);
xor U18712 (N_18712,N_18409,N_18481);
and U18713 (N_18713,N_18476,N_18297);
or U18714 (N_18714,N_18495,N_18483);
and U18715 (N_18715,N_18330,N_18279);
nand U18716 (N_18716,N_18397,N_18448);
nor U18717 (N_18717,N_18345,N_18406);
and U18718 (N_18718,N_18382,N_18332);
nand U18719 (N_18719,N_18483,N_18308);
xor U18720 (N_18720,N_18356,N_18386);
or U18721 (N_18721,N_18320,N_18392);
and U18722 (N_18722,N_18474,N_18432);
or U18723 (N_18723,N_18472,N_18469);
xnor U18724 (N_18724,N_18467,N_18412);
xor U18725 (N_18725,N_18352,N_18260);
nor U18726 (N_18726,N_18311,N_18361);
nor U18727 (N_18727,N_18473,N_18355);
nor U18728 (N_18728,N_18252,N_18350);
xor U18729 (N_18729,N_18316,N_18466);
nand U18730 (N_18730,N_18299,N_18411);
nand U18731 (N_18731,N_18383,N_18422);
xor U18732 (N_18732,N_18278,N_18384);
or U18733 (N_18733,N_18463,N_18402);
and U18734 (N_18734,N_18329,N_18459);
xnor U18735 (N_18735,N_18400,N_18345);
or U18736 (N_18736,N_18457,N_18354);
and U18737 (N_18737,N_18274,N_18253);
and U18738 (N_18738,N_18405,N_18253);
or U18739 (N_18739,N_18327,N_18429);
nand U18740 (N_18740,N_18384,N_18416);
xor U18741 (N_18741,N_18357,N_18369);
xor U18742 (N_18742,N_18423,N_18496);
or U18743 (N_18743,N_18294,N_18383);
nor U18744 (N_18744,N_18490,N_18323);
nor U18745 (N_18745,N_18323,N_18318);
xor U18746 (N_18746,N_18459,N_18267);
and U18747 (N_18747,N_18251,N_18360);
or U18748 (N_18748,N_18459,N_18284);
and U18749 (N_18749,N_18292,N_18442);
nand U18750 (N_18750,N_18661,N_18679);
nand U18751 (N_18751,N_18580,N_18716);
nand U18752 (N_18752,N_18549,N_18595);
or U18753 (N_18753,N_18564,N_18546);
or U18754 (N_18754,N_18592,N_18677);
xnor U18755 (N_18755,N_18641,N_18730);
nor U18756 (N_18756,N_18618,N_18525);
nand U18757 (N_18757,N_18587,N_18512);
nand U18758 (N_18758,N_18509,N_18579);
nor U18759 (N_18759,N_18640,N_18605);
xnor U18760 (N_18760,N_18566,N_18573);
nand U18761 (N_18761,N_18675,N_18617);
or U18762 (N_18762,N_18547,N_18646);
or U18763 (N_18763,N_18740,N_18598);
nand U18764 (N_18764,N_18621,N_18583);
xnor U18765 (N_18765,N_18505,N_18542);
or U18766 (N_18766,N_18556,N_18541);
nor U18767 (N_18767,N_18515,N_18520);
nor U18768 (N_18768,N_18739,N_18528);
or U18769 (N_18769,N_18523,N_18500);
or U18770 (N_18770,N_18553,N_18636);
xor U18771 (N_18771,N_18666,N_18539);
nor U18772 (N_18772,N_18672,N_18674);
nand U18773 (N_18773,N_18722,N_18550);
nand U18774 (N_18774,N_18729,N_18518);
nor U18775 (N_18775,N_18662,N_18634);
or U18776 (N_18776,N_18604,N_18723);
xnor U18777 (N_18777,N_18514,N_18551);
xor U18778 (N_18778,N_18517,N_18684);
nand U18779 (N_18779,N_18545,N_18726);
xor U18780 (N_18780,N_18559,N_18657);
xnor U18781 (N_18781,N_18511,N_18608);
nand U18782 (N_18782,N_18561,N_18733);
xnor U18783 (N_18783,N_18645,N_18651);
nor U18784 (N_18784,N_18575,N_18609);
and U18785 (N_18785,N_18629,N_18676);
and U18786 (N_18786,N_18698,N_18708);
nor U18787 (N_18787,N_18715,N_18630);
xor U18788 (N_18788,N_18707,N_18597);
xor U18789 (N_18789,N_18537,N_18526);
nor U18790 (N_18790,N_18601,N_18536);
nand U18791 (N_18791,N_18508,N_18714);
or U18792 (N_18792,N_18710,N_18721);
xnor U18793 (N_18793,N_18567,N_18521);
or U18794 (N_18794,N_18560,N_18504);
xnor U18795 (N_18795,N_18577,N_18652);
nand U18796 (N_18796,N_18650,N_18535);
or U18797 (N_18797,N_18642,N_18664);
and U18798 (N_18798,N_18683,N_18571);
nor U18799 (N_18799,N_18728,N_18513);
and U18800 (N_18800,N_18585,N_18736);
and U18801 (N_18801,N_18614,N_18705);
xnor U18802 (N_18802,N_18665,N_18709);
and U18803 (N_18803,N_18582,N_18531);
and U18804 (N_18804,N_18746,N_18519);
nand U18805 (N_18805,N_18685,N_18590);
nor U18806 (N_18806,N_18578,N_18678);
nand U18807 (N_18807,N_18735,N_18704);
and U18808 (N_18808,N_18693,N_18731);
nand U18809 (N_18809,N_18743,N_18501);
nand U18810 (N_18810,N_18615,N_18668);
or U18811 (N_18811,N_18638,N_18687);
and U18812 (N_18812,N_18622,N_18619);
or U18813 (N_18813,N_18529,N_18607);
or U18814 (N_18814,N_18570,N_18748);
nand U18815 (N_18815,N_18524,N_18647);
and U18816 (N_18816,N_18682,N_18548);
xnor U18817 (N_18817,N_18565,N_18725);
xor U18818 (N_18818,N_18691,N_18702);
xnor U18819 (N_18819,N_18612,N_18544);
nor U18820 (N_18820,N_18727,N_18599);
or U18821 (N_18821,N_18703,N_18562);
or U18822 (N_18822,N_18658,N_18533);
nand U18823 (N_18823,N_18749,N_18538);
nand U18824 (N_18824,N_18649,N_18572);
nor U18825 (N_18825,N_18686,N_18510);
nor U18826 (N_18826,N_18569,N_18620);
and U18827 (N_18827,N_18534,N_18695);
or U18828 (N_18828,N_18680,N_18611);
and U18829 (N_18829,N_18563,N_18540);
nand U18830 (N_18830,N_18610,N_18643);
nand U18831 (N_18831,N_18530,N_18644);
xor U18832 (N_18832,N_18655,N_18712);
nor U18833 (N_18833,N_18744,N_18692);
nor U18834 (N_18834,N_18626,N_18606);
xnor U18835 (N_18835,N_18660,N_18696);
xor U18836 (N_18836,N_18631,N_18713);
nand U18837 (N_18837,N_18557,N_18616);
or U18838 (N_18838,N_18737,N_18742);
or U18839 (N_18839,N_18625,N_18745);
or U18840 (N_18840,N_18593,N_18613);
nand U18841 (N_18841,N_18635,N_18669);
nor U18842 (N_18842,N_18552,N_18656);
xnor U18843 (N_18843,N_18706,N_18673);
nor U18844 (N_18844,N_18558,N_18663);
or U18845 (N_18845,N_18738,N_18516);
or U18846 (N_18846,N_18697,N_18532);
nor U18847 (N_18847,N_18554,N_18522);
and U18848 (N_18848,N_18591,N_18589);
nor U18849 (N_18849,N_18568,N_18717);
or U18850 (N_18850,N_18711,N_18628);
or U18851 (N_18851,N_18602,N_18701);
or U18852 (N_18852,N_18603,N_18724);
and U18853 (N_18853,N_18718,N_18690);
nand U18854 (N_18854,N_18581,N_18596);
xor U18855 (N_18855,N_18624,N_18633);
nand U18856 (N_18856,N_18506,N_18623);
xor U18857 (N_18857,N_18659,N_18637);
xor U18858 (N_18858,N_18586,N_18600);
and U18859 (N_18859,N_18502,N_18555);
nand U18860 (N_18860,N_18574,N_18694);
and U18861 (N_18861,N_18588,N_18747);
nor U18862 (N_18862,N_18507,N_18667);
or U18863 (N_18863,N_18741,N_18699);
xnor U18864 (N_18864,N_18653,N_18732);
nor U18865 (N_18865,N_18639,N_18627);
xor U18866 (N_18866,N_18543,N_18594);
xnor U18867 (N_18867,N_18670,N_18503);
nor U18868 (N_18868,N_18734,N_18648);
and U18869 (N_18869,N_18671,N_18654);
or U18870 (N_18870,N_18689,N_18720);
nand U18871 (N_18871,N_18576,N_18700);
xor U18872 (N_18872,N_18584,N_18719);
and U18873 (N_18873,N_18527,N_18632);
and U18874 (N_18874,N_18688,N_18681);
nor U18875 (N_18875,N_18550,N_18538);
nor U18876 (N_18876,N_18667,N_18585);
nand U18877 (N_18877,N_18649,N_18599);
nand U18878 (N_18878,N_18697,N_18549);
nand U18879 (N_18879,N_18509,N_18703);
xor U18880 (N_18880,N_18552,N_18551);
and U18881 (N_18881,N_18713,N_18524);
nor U18882 (N_18882,N_18698,N_18563);
nand U18883 (N_18883,N_18628,N_18575);
and U18884 (N_18884,N_18708,N_18648);
and U18885 (N_18885,N_18510,N_18511);
xor U18886 (N_18886,N_18595,N_18618);
nor U18887 (N_18887,N_18527,N_18618);
nand U18888 (N_18888,N_18572,N_18577);
and U18889 (N_18889,N_18690,N_18655);
nor U18890 (N_18890,N_18595,N_18667);
xor U18891 (N_18891,N_18718,N_18632);
and U18892 (N_18892,N_18629,N_18677);
nor U18893 (N_18893,N_18519,N_18706);
and U18894 (N_18894,N_18554,N_18671);
or U18895 (N_18895,N_18626,N_18635);
and U18896 (N_18896,N_18501,N_18716);
xnor U18897 (N_18897,N_18545,N_18530);
and U18898 (N_18898,N_18741,N_18603);
nor U18899 (N_18899,N_18630,N_18644);
xor U18900 (N_18900,N_18533,N_18709);
and U18901 (N_18901,N_18698,N_18540);
xnor U18902 (N_18902,N_18501,N_18580);
xnor U18903 (N_18903,N_18709,N_18720);
and U18904 (N_18904,N_18536,N_18613);
xnor U18905 (N_18905,N_18563,N_18659);
xnor U18906 (N_18906,N_18578,N_18533);
nand U18907 (N_18907,N_18705,N_18748);
and U18908 (N_18908,N_18635,N_18506);
and U18909 (N_18909,N_18507,N_18746);
nor U18910 (N_18910,N_18716,N_18630);
xnor U18911 (N_18911,N_18535,N_18646);
and U18912 (N_18912,N_18565,N_18687);
xnor U18913 (N_18913,N_18722,N_18515);
xnor U18914 (N_18914,N_18623,N_18576);
xnor U18915 (N_18915,N_18717,N_18519);
and U18916 (N_18916,N_18505,N_18678);
nor U18917 (N_18917,N_18512,N_18710);
and U18918 (N_18918,N_18674,N_18738);
or U18919 (N_18919,N_18727,N_18724);
and U18920 (N_18920,N_18585,N_18524);
or U18921 (N_18921,N_18541,N_18610);
or U18922 (N_18922,N_18504,N_18615);
xor U18923 (N_18923,N_18714,N_18717);
xor U18924 (N_18924,N_18643,N_18535);
xnor U18925 (N_18925,N_18667,N_18695);
and U18926 (N_18926,N_18637,N_18624);
or U18927 (N_18927,N_18502,N_18661);
nand U18928 (N_18928,N_18508,N_18516);
and U18929 (N_18929,N_18544,N_18632);
and U18930 (N_18930,N_18728,N_18555);
xor U18931 (N_18931,N_18564,N_18643);
nor U18932 (N_18932,N_18607,N_18634);
and U18933 (N_18933,N_18728,N_18528);
nor U18934 (N_18934,N_18505,N_18720);
xnor U18935 (N_18935,N_18530,N_18677);
xor U18936 (N_18936,N_18507,N_18655);
or U18937 (N_18937,N_18554,N_18706);
nor U18938 (N_18938,N_18580,N_18509);
nand U18939 (N_18939,N_18501,N_18569);
nor U18940 (N_18940,N_18537,N_18635);
nand U18941 (N_18941,N_18724,N_18646);
nor U18942 (N_18942,N_18650,N_18633);
and U18943 (N_18943,N_18687,N_18528);
and U18944 (N_18944,N_18581,N_18510);
or U18945 (N_18945,N_18520,N_18634);
or U18946 (N_18946,N_18599,N_18657);
and U18947 (N_18947,N_18526,N_18574);
and U18948 (N_18948,N_18663,N_18680);
nand U18949 (N_18949,N_18537,N_18553);
and U18950 (N_18950,N_18531,N_18646);
and U18951 (N_18951,N_18718,N_18680);
and U18952 (N_18952,N_18582,N_18645);
xnor U18953 (N_18953,N_18732,N_18627);
nor U18954 (N_18954,N_18737,N_18646);
or U18955 (N_18955,N_18717,N_18575);
nor U18956 (N_18956,N_18635,N_18620);
nand U18957 (N_18957,N_18575,N_18714);
xnor U18958 (N_18958,N_18578,N_18623);
nand U18959 (N_18959,N_18679,N_18516);
and U18960 (N_18960,N_18627,N_18551);
and U18961 (N_18961,N_18577,N_18704);
nor U18962 (N_18962,N_18630,N_18597);
xnor U18963 (N_18963,N_18609,N_18516);
nor U18964 (N_18964,N_18574,N_18663);
nand U18965 (N_18965,N_18629,N_18527);
and U18966 (N_18966,N_18703,N_18664);
xor U18967 (N_18967,N_18697,N_18641);
nand U18968 (N_18968,N_18613,N_18620);
nand U18969 (N_18969,N_18583,N_18572);
and U18970 (N_18970,N_18688,N_18526);
or U18971 (N_18971,N_18566,N_18636);
or U18972 (N_18972,N_18586,N_18547);
nor U18973 (N_18973,N_18533,N_18745);
nand U18974 (N_18974,N_18587,N_18634);
or U18975 (N_18975,N_18696,N_18680);
xor U18976 (N_18976,N_18749,N_18713);
or U18977 (N_18977,N_18501,N_18572);
and U18978 (N_18978,N_18523,N_18537);
nor U18979 (N_18979,N_18628,N_18629);
or U18980 (N_18980,N_18598,N_18550);
nor U18981 (N_18981,N_18748,N_18512);
or U18982 (N_18982,N_18749,N_18524);
xor U18983 (N_18983,N_18608,N_18741);
and U18984 (N_18984,N_18604,N_18521);
nand U18985 (N_18985,N_18749,N_18614);
or U18986 (N_18986,N_18596,N_18572);
xor U18987 (N_18987,N_18647,N_18729);
or U18988 (N_18988,N_18552,N_18542);
xor U18989 (N_18989,N_18634,N_18597);
nand U18990 (N_18990,N_18536,N_18608);
nor U18991 (N_18991,N_18545,N_18632);
or U18992 (N_18992,N_18745,N_18627);
and U18993 (N_18993,N_18559,N_18683);
nor U18994 (N_18994,N_18550,N_18583);
nand U18995 (N_18995,N_18618,N_18647);
or U18996 (N_18996,N_18660,N_18723);
nand U18997 (N_18997,N_18528,N_18529);
nor U18998 (N_18998,N_18526,N_18681);
nand U18999 (N_18999,N_18631,N_18607);
nor U19000 (N_19000,N_18774,N_18750);
nor U19001 (N_19001,N_18822,N_18961);
xor U19002 (N_19002,N_18809,N_18925);
or U19003 (N_19003,N_18869,N_18895);
xnor U19004 (N_19004,N_18969,N_18871);
nand U19005 (N_19005,N_18883,N_18981);
nand U19006 (N_19006,N_18975,N_18841);
nand U19007 (N_19007,N_18863,N_18986);
nand U19008 (N_19008,N_18773,N_18897);
nand U19009 (N_19009,N_18766,N_18872);
xor U19010 (N_19010,N_18876,N_18970);
and U19011 (N_19011,N_18962,N_18782);
and U19012 (N_19012,N_18932,N_18966);
and U19013 (N_19013,N_18976,N_18920);
or U19014 (N_19014,N_18789,N_18830);
or U19015 (N_19015,N_18855,N_18794);
or U19016 (N_19016,N_18887,N_18952);
xor U19017 (N_19017,N_18921,N_18938);
and U19018 (N_19018,N_18817,N_18781);
and U19019 (N_19019,N_18989,N_18980);
xnor U19020 (N_19020,N_18946,N_18849);
and U19021 (N_19021,N_18873,N_18957);
or U19022 (N_19022,N_18967,N_18999);
xor U19023 (N_19023,N_18800,N_18803);
xnor U19024 (N_19024,N_18922,N_18909);
and U19025 (N_19025,N_18763,N_18901);
or U19026 (N_19026,N_18868,N_18959);
nand U19027 (N_19027,N_18972,N_18791);
nand U19028 (N_19028,N_18918,N_18813);
nor U19029 (N_19029,N_18812,N_18941);
nor U19030 (N_19030,N_18998,N_18971);
nor U19031 (N_19031,N_18963,N_18808);
xnor U19032 (N_19032,N_18974,N_18891);
or U19033 (N_19033,N_18879,N_18842);
xor U19034 (N_19034,N_18765,N_18839);
nor U19035 (N_19035,N_18751,N_18825);
and U19036 (N_19036,N_18914,N_18984);
or U19037 (N_19037,N_18934,N_18771);
nand U19038 (N_19038,N_18913,N_18881);
nand U19039 (N_19039,N_18835,N_18964);
and U19040 (N_19040,N_18831,N_18995);
nand U19041 (N_19041,N_18997,N_18906);
or U19042 (N_19042,N_18933,N_18875);
and U19043 (N_19043,N_18755,N_18858);
and U19044 (N_19044,N_18878,N_18910);
xor U19045 (N_19045,N_18810,N_18856);
xnor U19046 (N_19046,N_18805,N_18983);
or U19047 (N_19047,N_18760,N_18821);
nor U19048 (N_19048,N_18786,N_18958);
nor U19049 (N_19049,N_18754,N_18767);
xor U19050 (N_19050,N_18993,N_18844);
or U19051 (N_19051,N_18948,N_18768);
nor U19052 (N_19052,N_18899,N_18757);
and U19053 (N_19053,N_18907,N_18874);
and U19054 (N_19054,N_18864,N_18775);
nor U19055 (N_19055,N_18834,N_18988);
nand U19056 (N_19056,N_18956,N_18778);
nor U19057 (N_19057,N_18930,N_18860);
xor U19058 (N_19058,N_18912,N_18811);
nor U19059 (N_19059,N_18911,N_18951);
nor U19060 (N_19060,N_18954,N_18823);
xnor U19061 (N_19061,N_18886,N_18840);
xor U19062 (N_19062,N_18788,N_18937);
or U19063 (N_19063,N_18836,N_18824);
nor U19064 (N_19064,N_18926,N_18904);
nor U19065 (N_19065,N_18792,N_18795);
nor U19066 (N_19066,N_18882,N_18939);
xnor U19067 (N_19067,N_18853,N_18862);
nand U19068 (N_19068,N_18947,N_18870);
or U19069 (N_19069,N_18780,N_18827);
or U19070 (N_19070,N_18770,N_18761);
nor U19071 (N_19071,N_18776,N_18806);
and U19072 (N_19072,N_18854,N_18960);
nor U19073 (N_19073,N_18815,N_18769);
nand U19074 (N_19074,N_18866,N_18777);
xnor U19075 (N_19075,N_18919,N_18950);
or U19076 (N_19076,N_18838,N_18846);
or U19077 (N_19077,N_18987,N_18793);
nor U19078 (N_19078,N_18851,N_18804);
nand U19079 (N_19079,N_18807,N_18826);
and U19080 (N_19080,N_18785,N_18845);
and U19081 (N_19081,N_18936,N_18790);
and U19082 (N_19082,N_18880,N_18942);
xnor U19083 (N_19083,N_18990,N_18928);
nand U19084 (N_19084,N_18814,N_18867);
or U19085 (N_19085,N_18977,N_18759);
xnor U19086 (N_19086,N_18892,N_18985);
or U19087 (N_19087,N_18762,N_18848);
and U19088 (N_19088,N_18923,N_18888);
and U19089 (N_19089,N_18833,N_18752);
nand U19090 (N_19090,N_18852,N_18784);
nand U19091 (N_19091,N_18978,N_18973);
nand U19092 (N_19092,N_18829,N_18968);
nor U19093 (N_19093,N_18865,N_18756);
and U19094 (N_19094,N_18787,N_18982);
and U19095 (N_19095,N_18884,N_18955);
nor U19096 (N_19096,N_18949,N_18935);
and U19097 (N_19097,N_18931,N_18905);
nor U19098 (N_19098,N_18953,N_18944);
or U19099 (N_19099,N_18850,N_18991);
xnor U19100 (N_19100,N_18828,N_18843);
nand U19101 (N_19101,N_18772,N_18885);
nor U19102 (N_19102,N_18796,N_18861);
nor U19103 (N_19103,N_18898,N_18797);
nand U19104 (N_19104,N_18832,N_18816);
xnor U19105 (N_19105,N_18819,N_18798);
nor U19106 (N_19106,N_18753,N_18758);
xor U19107 (N_19107,N_18908,N_18992);
xor U19108 (N_19108,N_18818,N_18799);
nand U19109 (N_19109,N_18802,N_18857);
nor U19110 (N_19110,N_18943,N_18820);
xnor U19111 (N_19111,N_18924,N_18917);
xor U19112 (N_19112,N_18801,N_18915);
nand U19113 (N_19113,N_18894,N_18877);
or U19114 (N_19114,N_18893,N_18900);
and U19115 (N_19115,N_18890,N_18979);
nor U19116 (N_19116,N_18847,N_18945);
nor U19117 (N_19117,N_18837,N_18764);
xor U19118 (N_19118,N_18927,N_18994);
nand U19119 (N_19119,N_18779,N_18896);
or U19120 (N_19120,N_18916,N_18783);
nand U19121 (N_19121,N_18940,N_18965);
xnor U19122 (N_19122,N_18996,N_18903);
nand U19123 (N_19123,N_18902,N_18889);
nor U19124 (N_19124,N_18929,N_18859);
and U19125 (N_19125,N_18978,N_18824);
and U19126 (N_19126,N_18836,N_18855);
nand U19127 (N_19127,N_18952,N_18784);
xnor U19128 (N_19128,N_18963,N_18801);
and U19129 (N_19129,N_18939,N_18854);
or U19130 (N_19130,N_18755,N_18799);
and U19131 (N_19131,N_18882,N_18960);
nor U19132 (N_19132,N_18788,N_18948);
xnor U19133 (N_19133,N_18767,N_18912);
or U19134 (N_19134,N_18915,N_18864);
nand U19135 (N_19135,N_18775,N_18964);
xnor U19136 (N_19136,N_18755,N_18786);
or U19137 (N_19137,N_18818,N_18951);
and U19138 (N_19138,N_18948,N_18781);
nand U19139 (N_19139,N_18891,N_18874);
xor U19140 (N_19140,N_18892,N_18880);
xor U19141 (N_19141,N_18838,N_18911);
xnor U19142 (N_19142,N_18782,N_18929);
xor U19143 (N_19143,N_18802,N_18772);
and U19144 (N_19144,N_18937,N_18793);
nor U19145 (N_19145,N_18793,N_18870);
nor U19146 (N_19146,N_18771,N_18864);
or U19147 (N_19147,N_18854,N_18890);
or U19148 (N_19148,N_18844,N_18829);
nand U19149 (N_19149,N_18888,N_18993);
xor U19150 (N_19150,N_18981,N_18755);
and U19151 (N_19151,N_18772,N_18969);
xor U19152 (N_19152,N_18759,N_18831);
or U19153 (N_19153,N_18858,N_18846);
nor U19154 (N_19154,N_18786,N_18990);
nand U19155 (N_19155,N_18825,N_18959);
xor U19156 (N_19156,N_18869,N_18941);
and U19157 (N_19157,N_18927,N_18792);
xor U19158 (N_19158,N_18850,N_18796);
nand U19159 (N_19159,N_18965,N_18795);
and U19160 (N_19160,N_18860,N_18813);
or U19161 (N_19161,N_18825,N_18755);
xor U19162 (N_19162,N_18850,N_18762);
nand U19163 (N_19163,N_18916,N_18763);
or U19164 (N_19164,N_18865,N_18956);
nor U19165 (N_19165,N_18981,N_18816);
xnor U19166 (N_19166,N_18941,N_18825);
nor U19167 (N_19167,N_18849,N_18877);
nand U19168 (N_19168,N_18898,N_18752);
or U19169 (N_19169,N_18782,N_18914);
or U19170 (N_19170,N_18770,N_18880);
or U19171 (N_19171,N_18760,N_18878);
nor U19172 (N_19172,N_18896,N_18832);
nand U19173 (N_19173,N_18774,N_18807);
nor U19174 (N_19174,N_18962,N_18750);
xor U19175 (N_19175,N_18862,N_18936);
nand U19176 (N_19176,N_18831,N_18753);
nor U19177 (N_19177,N_18837,N_18873);
nand U19178 (N_19178,N_18997,N_18911);
nand U19179 (N_19179,N_18857,N_18908);
and U19180 (N_19180,N_18958,N_18904);
nor U19181 (N_19181,N_18789,N_18997);
and U19182 (N_19182,N_18966,N_18823);
xnor U19183 (N_19183,N_18771,N_18779);
and U19184 (N_19184,N_18988,N_18795);
or U19185 (N_19185,N_18878,N_18772);
nand U19186 (N_19186,N_18961,N_18995);
xor U19187 (N_19187,N_18993,N_18848);
xnor U19188 (N_19188,N_18819,N_18801);
or U19189 (N_19189,N_18983,N_18899);
and U19190 (N_19190,N_18870,N_18756);
nand U19191 (N_19191,N_18906,N_18975);
xor U19192 (N_19192,N_18799,N_18801);
nand U19193 (N_19193,N_18885,N_18862);
xnor U19194 (N_19194,N_18927,N_18915);
nor U19195 (N_19195,N_18898,N_18853);
and U19196 (N_19196,N_18971,N_18815);
nand U19197 (N_19197,N_18787,N_18863);
nor U19198 (N_19198,N_18918,N_18815);
nor U19199 (N_19199,N_18772,N_18862);
and U19200 (N_19200,N_18787,N_18881);
or U19201 (N_19201,N_18793,N_18984);
xnor U19202 (N_19202,N_18840,N_18821);
nor U19203 (N_19203,N_18776,N_18853);
nor U19204 (N_19204,N_18943,N_18897);
or U19205 (N_19205,N_18778,N_18948);
nor U19206 (N_19206,N_18874,N_18796);
nor U19207 (N_19207,N_18882,N_18772);
nor U19208 (N_19208,N_18966,N_18775);
or U19209 (N_19209,N_18777,N_18842);
and U19210 (N_19210,N_18904,N_18848);
nor U19211 (N_19211,N_18899,N_18827);
or U19212 (N_19212,N_18758,N_18901);
nand U19213 (N_19213,N_18954,N_18826);
nand U19214 (N_19214,N_18994,N_18969);
or U19215 (N_19215,N_18757,N_18978);
nand U19216 (N_19216,N_18830,N_18952);
nor U19217 (N_19217,N_18981,N_18884);
xnor U19218 (N_19218,N_18960,N_18959);
xnor U19219 (N_19219,N_18841,N_18810);
nand U19220 (N_19220,N_18999,N_18830);
or U19221 (N_19221,N_18794,N_18758);
nand U19222 (N_19222,N_18920,N_18786);
nor U19223 (N_19223,N_18859,N_18898);
nand U19224 (N_19224,N_18939,N_18873);
nor U19225 (N_19225,N_18762,N_18993);
and U19226 (N_19226,N_18990,N_18805);
and U19227 (N_19227,N_18853,N_18871);
nand U19228 (N_19228,N_18822,N_18894);
nor U19229 (N_19229,N_18752,N_18901);
or U19230 (N_19230,N_18870,N_18882);
nand U19231 (N_19231,N_18954,N_18808);
xor U19232 (N_19232,N_18868,N_18753);
nor U19233 (N_19233,N_18909,N_18794);
nand U19234 (N_19234,N_18794,N_18757);
and U19235 (N_19235,N_18834,N_18995);
nor U19236 (N_19236,N_18882,N_18861);
nand U19237 (N_19237,N_18811,N_18857);
nor U19238 (N_19238,N_18813,N_18931);
nand U19239 (N_19239,N_18964,N_18761);
and U19240 (N_19240,N_18988,N_18936);
xor U19241 (N_19241,N_18886,N_18899);
nor U19242 (N_19242,N_18933,N_18848);
or U19243 (N_19243,N_18849,N_18785);
and U19244 (N_19244,N_18822,N_18885);
nand U19245 (N_19245,N_18792,N_18999);
and U19246 (N_19246,N_18823,N_18833);
xor U19247 (N_19247,N_18846,N_18954);
nand U19248 (N_19248,N_18969,N_18902);
nor U19249 (N_19249,N_18929,N_18767);
xor U19250 (N_19250,N_19090,N_19074);
xor U19251 (N_19251,N_19193,N_19106);
xor U19252 (N_19252,N_19033,N_19232);
or U19253 (N_19253,N_19249,N_19105);
or U19254 (N_19254,N_19145,N_19054);
or U19255 (N_19255,N_19121,N_19247);
or U19256 (N_19256,N_19198,N_19234);
nand U19257 (N_19257,N_19125,N_19191);
nand U19258 (N_19258,N_19036,N_19155);
and U19259 (N_19259,N_19181,N_19117);
or U19260 (N_19260,N_19133,N_19050);
nor U19261 (N_19261,N_19079,N_19116);
or U19262 (N_19262,N_19171,N_19114);
or U19263 (N_19263,N_19215,N_19008);
nor U19264 (N_19264,N_19246,N_19183);
xor U19265 (N_19265,N_19158,N_19217);
or U19266 (N_19266,N_19150,N_19059);
nand U19267 (N_19267,N_19203,N_19209);
and U19268 (N_19268,N_19082,N_19045);
or U19269 (N_19269,N_19066,N_19061);
xor U19270 (N_19270,N_19113,N_19207);
xor U19271 (N_19271,N_19248,N_19179);
and U19272 (N_19272,N_19161,N_19039);
or U19273 (N_19273,N_19123,N_19241);
and U19274 (N_19274,N_19076,N_19119);
or U19275 (N_19275,N_19086,N_19068);
nand U19276 (N_19276,N_19128,N_19065);
nor U19277 (N_19277,N_19185,N_19176);
and U19278 (N_19278,N_19233,N_19013);
xnor U19279 (N_19279,N_19174,N_19043);
nand U19280 (N_19280,N_19235,N_19137);
xor U19281 (N_19281,N_19002,N_19195);
and U19282 (N_19282,N_19188,N_19189);
or U19283 (N_19283,N_19136,N_19101);
xnor U19284 (N_19284,N_19146,N_19243);
or U19285 (N_19285,N_19078,N_19032);
nor U19286 (N_19286,N_19242,N_19108);
xnor U19287 (N_19287,N_19055,N_19093);
xnor U19288 (N_19288,N_19028,N_19058);
nand U19289 (N_19289,N_19091,N_19115);
nand U19290 (N_19290,N_19141,N_19223);
and U19291 (N_19291,N_19163,N_19003);
or U19292 (N_19292,N_19026,N_19044);
nand U19293 (N_19293,N_19199,N_19154);
or U19294 (N_19294,N_19147,N_19164);
and U19295 (N_19295,N_19231,N_19130);
nor U19296 (N_19296,N_19047,N_19238);
or U19297 (N_19297,N_19149,N_19087);
and U19298 (N_19298,N_19111,N_19110);
nor U19299 (N_19299,N_19206,N_19042);
or U19300 (N_19300,N_19201,N_19120);
nand U19301 (N_19301,N_19020,N_19099);
and U19302 (N_19302,N_19041,N_19196);
nand U19303 (N_19303,N_19228,N_19175);
or U19304 (N_19304,N_19227,N_19162);
nand U19305 (N_19305,N_19152,N_19027);
nand U19306 (N_19306,N_19070,N_19073);
and U19307 (N_19307,N_19011,N_19103);
nand U19308 (N_19308,N_19034,N_19208);
nand U19309 (N_19309,N_19052,N_19134);
and U19310 (N_19310,N_19048,N_19069);
xnor U19311 (N_19311,N_19014,N_19166);
or U19312 (N_19312,N_19138,N_19022);
nand U19313 (N_19313,N_19132,N_19104);
nand U19314 (N_19314,N_19029,N_19053);
or U19315 (N_19315,N_19040,N_19015);
or U19316 (N_19316,N_19085,N_19124);
or U19317 (N_19317,N_19063,N_19010);
nand U19318 (N_19318,N_19165,N_19127);
and U19319 (N_19319,N_19216,N_19172);
or U19320 (N_19320,N_19060,N_19211);
nand U19321 (N_19321,N_19094,N_19005);
xnor U19322 (N_19322,N_19214,N_19126);
nor U19323 (N_19323,N_19023,N_19038);
xnor U19324 (N_19324,N_19031,N_19072);
or U19325 (N_19325,N_19156,N_19169);
or U19326 (N_19326,N_19064,N_19177);
and U19327 (N_19327,N_19129,N_19239);
xor U19328 (N_19328,N_19122,N_19009);
nand U19329 (N_19329,N_19098,N_19212);
or U19330 (N_19330,N_19092,N_19109);
nand U19331 (N_19331,N_19144,N_19037);
or U19332 (N_19332,N_19197,N_19017);
and U19333 (N_19333,N_19019,N_19240);
and U19334 (N_19334,N_19100,N_19056);
nand U19335 (N_19335,N_19244,N_19218);
nand U19336 (N_19336,N_19096,N_19186);
nand U19337 (N_19337,N_19148,N_19024);
xnor U19338 (N_19338,N_19071,N_19219);
or U19339 (N_19339,N_19001,N_19077);
xor U19340 (N_19340,N_19160,N_19012);
and U19341 (N_19341,N_19205,N_19213);
or U19342 (N_19342,N_19187,N_19221);
xor U19343 (N_19343,N_19200,N_19139);
and U19344 (N_19344,N_19194,N_19245);
nand U19345 (N_19345,N_19229,N_19102);
nand U19346 (N_19346,N_19088,N_19180);
and U19347 (N_19347,N_19112,N_19151);
or U19348 (N_19348,N_19168,N_19159);
nor U19349 (N_19349,N_19049,N_19153);
xnor U19350 (N_19350,N_19220,N_19083);
nor U19351 (N_19351,N_19167,N_19226);
xnor U19352 (N_19352,N_19182,N_19084);
or U19353 (N_19353,N_19000,N_19173);
or U19354 (N_19354,N_19006,N_19192);
nand U19355 (N_19355,N_19202,N_19142);
nor U19356 (N_19356,N_19007,N_19143);
and U19357 (N_19357,N_19157,N_19131);
nand U19358 (N_19358,N_19080,N_19075);
nor U19359 (N_19359,N_19204,N_19097);
and U19360 (N_19360,N_19081,N_19135);
nand U19361 (N_19361,N_19178,N_19046);
nor U19362 (N_19362,N_19237,N_19107);
nand U19363 (N_19363,N_19230,N_19051);
nand U19364 (N_19364,N_19089,N_19140);
nand U19365 (N_19365,N_19225,N_19118);
and U19366 (N_19366,N_19030,N_19224);
nor U19367 (N_19367,N_19016,N_19170);
or U19368 (N_19368,N_19095,N_19236);
xnor U19369 (N_19369,N_19018,N_19057);
nor U19370 (N_19370,N_19210,N_19021);
or U19371 (N_19371,N_19004,N_19035);
xor U19372 (N_19372,N_19067,N_19062);
xor U19373 (N_19373,N_19222,N_19190);
nor U19374 (N_19374,N_19184,N_19025);
nand U19375 (N_19375,N_19210,N_19145);
and U19376 (N_19376,N_19144,N_19151);
or U19377 (N_19377,N_19193,N_19003);
and U19378 (N_19378,N_19036,N_19201);
nand U19379 (N_19379,N_19031,N_19035);
nand U19380 (N_19380,N_19173,N_19091);
or U19381 (N_19381,N_19030,N_19199);
and U19382 (N_19382,N_19011,N_19022);
nor U19383 (N_19383,N_19068,N_19231);
and U19384 (N_19384,N_19081,N_19071);
nor U19385 (N_19385,N_19219,N_19191);
xor U19386 (N_19386,N_19204,N_19223);
xnor U19387 (N_19387,N_19062,N_19154);
or U19388 (N_19388,N_19125,N_19169);
xnor U19389 (N_19389,N_19123,N_19215);
or U19390 (N_19390,N_19225,N_19039);
xnor U19391 (N_19391,N_19109,N_19189);
nor U19392 (N_19392,N_19016,N_19022);
xor U19393 (N_19393,N_19217,N_19007);
xor U19394 (N_19394,N_19162,N_19107);
nand U19395 (N_19395,N_19135,N_19097);
nor U19396 (N_19396,N_19126,N_19248);
or U19397 (N_19397,N_19006,N_19208);
or U19398 (N_19398,N_19072,N_19146);
nand U19399 (N_19399,N_19153,N_19126);
nand U19400 (N_19400,N_19119,N_19148);
nor U19401 (N_19401,N_19088,N_19053);
nand U19402 (N_19402,N_19117,N_19068);
xor U19403 (N_19403,N_19015,N_19091);
nand U19404 (N_19404,N_19084,N_19059);
xor U19405 (N_19405,N_19049,N_19174);
nand U19406 (N_19406,N_19141,N_19025);
and U19407 (N_19407,N_19050,N_19078);
or U19408 (N_19408,N_19052,N_19179);
xnor U19409 (N_19409,N_19083,N_19014);
xnor U19410 (N_19410,N_19165,N_19086);
xor U19411 (N_19411,N_19075,N_19238);
or U19412 (N_19412,N_19146,N_19054);
and U19413 (N_19413,N_19225,N_19156);
and U19414 (N_19414,N_19068,N_19131);
nand U19415 (N_19415,N_19238,N_19017);
nand U19416 (N_19416,N_19199,N_19206);
and U19417 (N_19417,N_19092,N_19058);
or U19418 (N_19418,N_19018,N_19021);
nor U19419 (N_19419,N_19147,N_19052);
or U19420 (N_19420,N_19184,N_19162);
nor U19421 (N_19421,N_19040,N_19240);
or U19422 (N_19422,N_19222,N_19129);
xor U19423 (N_19423,N_19212,N_19234);
or U19424 (N_19424,N_19212,N_19123);
and U19425 (N_19425,N_19067,N_19071);
nor U19426 (N_19426,N_19095,N_19115);
or U19427 (N_19427,N_19190,N_19012);
or U19428 (N_19428,N_19196,N_19017);
xor U19429 (N_19429,N_19228,N_19111);
and U19430 (N_19430,N_19130,N_19079);
nand U19431 (N_19431,N_19123,N_19196);
or U19432 (N_19432,N_19035,N_19050);
xnor U19433 (N_19433,N_19199,N_19161);
xor U19434 (N_19434,N_19057,N_19100);
and U19435 (N_19435,N_19187,N_19084);
nor U19436 (N_19436,N_19107,N_19016);
nand U19437 (N_19437,N_19021,N_19013);
nand U19438 (N_19438,N_19019,N_19053);
xor U19439 (N_19439,N_19173,N_19085);
xnor U19440 (N_19440,N_19077,N_19045);
and U19441 (N_19441,N_19095,N_19019);
and U19442 (N_19442,N_19069,N_19170);
or U19443 (N_19443,N_19011,N_19241);
nor U19444 (N_19444,N_19037,N_19005);
xor U19445 (N_19445,N_19209,N_19213);
nor U19446 (N_19446,N_19033,N_19202);
nand U19447 (N_19447,N_19135,N_19032);
nor U19448 (N_19448,N_19080,N_19129);
nor U19449 (N_19449,N_19085,N_19060);
and U19450 (N_19450,N_19217,N_19238);
or U19451 (N_19451,N_19007,N_19083);
or U19452 (N_19452,N_19113,N_19158);
nor U19453 (N_19453,N_19061,N_19015);
and U19454 (N_19454,N_19107,N_19189);
and U19455 (N_19455,N_19203,N_19161);
or U19456 (N_19456,N_19144,N_19028);
and U19457 (N_19457,N_19065,N_19070);
xor U19458 (N_19458,N_19085,N_19237);
and U19459 (N_19459,N_19143,N_19081);
or U19460 (N_19460,N_19054,N_19044);
or U19461 (N_19461,N_19018,N_19161);
or U19462 (N_19462,N_19139,N_19009);
or U19463 (N_19463,N_19223,N_19187);
nand U19464 (N_19464,N_19054,N_19224);
xor U19465 (N_19465,N_19081,N_19039);
and U19466 (N_19466,N_19235,N_19027);
nand U19467 (N_19467,N_19070,N_19197);
nor U19468 (N_19468,N_19213,N_19187);
nor U19469 (N_19469,N_19122,N_19186);
and U19470 (N_19470,N_19017,N_19148);
xnor U19471 (N_19471,N_19132,N_19231);
xnor U19472 (N_19472,N_19227,N_19009);
or U19473 (N_19473,N_19130,N_19135);
nand U19474 (N_19474,N_19046,N_19154);
or U19475 (N_19475,N_19096,N_19004);
nand U19476 (N_19476,N_19082,N_19124);
nand U19477 (N_19477,N_19221,N_19228);
xor U19478 (N_19478,N_19025,N_19046);
nor U19479 (N_19479,N_19176,N_19137);
nand U19480 (N_19480,N_19141,N_19117);
xor U19481 (N_19481,N_19135,N_19144);
or U19482 (N_19482,N_19180,N_19085);
xor U19483 (N_19483,N_19249,N_19157);
nor U19484 (N_19484,N_19157,N_19110);
and U19485 (N_19485,N_19097,N_19110);
or U19486 (N_19486,N_19115,N_19139);
nand U19487 (N_19487,N_19045,N_19246);
xor U19488 (N_19488,N_19184,N_19047);
nand U19489 (N_19489,N_19111,N_19065);
or U19490 (N_19490,N_19090,N_19190);
or U19491 (N_19491,N_19013,N_19097);
nand U19492 (N_19492,N_19061,N_19004);
or U19493 (N_19493,N_19249,N_19190);
xor U19494 (N_19494,N_19055,N_19127);
and U19495 (N_19495,N_19246,N_19188);
xnor U19496 (N_19496,N_19218,N_19241);
or U19497 (N_19497,N_19042,N_19240);
and U19498 (N_19498,N_19060,N_19240);
or U19499 (N_19499,N_19012,N_19197);
and U19500 (N_19500,N_19308,N_19337);
nand U19501 (N_19501,N_19346,N_19285);
xnor U19502 (N_19502,N_19262,N_19446);
or U19503 (N_19503,N_19378,N_19351);
nor U19504 (N_19504,N_19282,N_19472);
xnor U19505 (N_19505,N_19408,N_19368);
or U19506 (N_19506,N_19321,N_19499);
xnor U19507 (N_19507,N_19402,N_19302);
and U19508 (N_19508,N_19300,N_19470);
and U19509 (N_19509,N_19333,N_19461);
nor U19510 (N_19510,N_19314,N_19443);
nand U19511 (N_19511,N_19498,N_19289);
or U19512 (N_19512,N_19264,N_19339);
nand U19513 (N_19513,N_19383,N_19418);
or U19514 (N_19514,N_19374,N_19288);
and U19515 (N_19515,N_19331,N_19329);
nor U19516 (N_19516,N_19370,N_19404);
or U19517 (N_19517,N_19482,N_19440);
and U19518 (N_19518,N_19409,N_19423);
or U19519 (N_19519,N_19493,N_19497);
nor U19520 (N_19520,N_19371,N_19388);
or U19521 (N_19521,N_19400,N_19324);
and U19522 (N_19522,N_19478,N_19367);
and U19523 (N_19523,N_19291,N_19407);
or U19524 (N_19524,N_19306,N_19369);
xnor U19525 (N_19525,N_19492,N_19458);
nor U19526 (N_19526,N_19355,N_19392);
nor U19527 (N_19527,N_19454,N_19428);
xor U19528 (N_19528,N_19310,N_19257);
nor U19529 (N_19529,N_19307,N_19320);
nand U19530 (N_19530,N_19496,N_19462);
nand U19531 (N_19531,N_19365,N_19403);
or U19532 (N_19532,N_19382,N_19277);
or U19533 (N_19533,N_19421,N_19338);
and U19534 (N_19534,N_19348,N_19340);
or U19535 (N_19535,N_19384,N_19305);
nor U19536 (N_19536,N_19299,N_19397);
or U19537 (N_19537,N_19444,N_19457);
nor U19538 (N_19538,N_19366,N_19459);
or U19539 (N_19539,N_19406,N_19380);
nor U19540 (N_19540,N_19350,N_19318);
or U19541 (N_19541,N_19389,N_19381);
xor U19542 (N_19542,N_19281,N_19431);
and U19543 (N_19543,N_19327,N_19263);
or U19544 (N_19544,N_19480,N_19469);
and U19545 (N_19545,N_19463,N_19445);
and U19546 (N_19546,N_19342,N_19358);
nor U19547 (N_19547,N_19332,N_19417);
nor U19548 (N_19548,N_19487,N_19419);
and U19549 (N_19549,N_19414,N_19483);
and U19550 (N_19550,N_19272,N_19271);
nor U19551 (N_19551,N_19259,N_19319);
nor U19552 (N_19552,N_19393,N_19465);
xor U19553 (N_19553,N_19375,N_19343);
nor U19554 (N_19554,N_19356,N_19481);
and U19555 (N_19555,N_19441,N_19447);
xor U19556 (N_19556,N_19387,N_19398);
or U19557 (N_19557,N_19325,N_19449);
or U19558 (N_19558,N_19364,N_19335);
and U19559 (N_19559,N_19316,N_19292);
or U19560 (N_19560,N_19296,N_19376);
nor U19561 (N_19561,N_19347,N_19456);
and U19562 (N_19562,N_19494,N_19274);
nand U19563 (N_19563,N_19294,N_19438);
nor U19564 (N_19564,N_19468,N_19424);
nor U19565 (N_19565,N_19390,N_19266);
nor U19566 (N_19566,N_19298,N_19442);
and U19567 (N_19567,N_19477,N_19427);
nand U19568 (N_19568,N_19295,N_19280);
and U19569 (N_19569,N_19261,N_19251);
and U19570 (N_19570,N_19467,N_19315);
nor U19571 (N_19571,N_19437,N_19475);
or U19572 (N_19572,N_19432,N_19373);
nand U19573 (N_19573,N_19391,N_19297);
and U19574 (N_19574,N_19253,N_19405);
or U19575 (N_19575,N_19354,N_19385);
and U19576 (N_19576,N_19476,N_19270);
nand U19577 (N_19577,N_19488,N_19490);
nand U19578 (N_19578,N_19326,N_19401);
or U19579 (N_19579,N_19450,N_19312);
nor U19580 (N_19580,N_19435,N_19386);
nor U19581 (N_19581,N_19453,N_19474);
xnor U19582 (N_19582,N_19452,N_19439);
xor U19583 (N_19583,N_19466,N_19413);
or U19584 (N_19584,N_19426,N_19267);
xor U19585 (N_19585,N_19359,N_19479);
nor U19586 (N_19586,N_19283,N_19352);
xor U19587 (N_19587,N_19471,N_19254);
and U19588 (N_19588,N_19394,N_19303);
xnor U19589 (N_19589,N_19276,N_19265);
and U19590 (N_19590,N_19293,N_19491);
or U19591 (N_19591,N_19420,N_19396);
nor U19592 (N_19592,N_19345,N_19361);
nor U19593 (N_19593,N_19379,N_19433);
nor U19594 (N_19594,N_19464,N_19323);
or U19595 (N_19595,N_19313,N_19422);
nor U19596 (N_19596,N_19485,N_19455);
xor U19597 (N_19597,N_19322,N_19328);
or U19598 (N_19598,N_19436,N_19410);
nor U19599 (N_19599,N_19416,N_19256);
nand U19600 (N_19600,N_19360,N_19304);
nor U19601 (N_19601,N_19399,N_19344);
nor U19602 (N_19602,N_19495,N_19317);
nand U19603 (N_19603,N_19448,N_19309);
or U19604 (N_19604,N_19434,N_19363);
and U19605 (N_19605,N_19279,N_19415);
xor U19606 (N_19606,N_19334,N_19460);
or U19607 (N_19607,N_19430,N_19425);
or U19608 (N_19608,N_19269,N_19412);
xor U19609 (N_19609,N_19311,N_19372);
and U19610 (N_19610,N_19290,N_19486);
or U19611 (N_19611,N_19252,N_19362);
and U19612 (N_19612,N_19273,N_19395);
or U19613 (N_19613,N_19286,N_19341);
xnor U19614 (N_19614,N_19301,N_19473);
nand U19615 (N_19615,N_19275,N_19357);
or U19616 (N_19616,N_19284,N_19268);
nand U19617 (N_19617,N_19255,N_19258);
and U19618 (N_19618,N_19353,N_19349);
and U19619 (N_19619,N_19336,N_19411);
nor U19620 (N_19620,N_19489,N_19260);
and U19621 (N_19621,N_19377,N_19287);
and U19622 (N_19622,N_19429,N_19278);
nand U19623 (N_19623,N_19250,N_19484);
xor U19624 (N_19624,N_19451,N_19330);
or U19625 (N_19625,N_19412,N_19458);
nand U19626 (N_19626,N_19421,N_19477);
xnor U19627 (N_19627,N_19474,N_19317);
xor U19628 (N_19628,N_19452,N_19311);
xor U19629 (N_19629,N_19314,N_19297);
or U19630 (N_19630,N_19366,N_19277);
xor U19631 (N_19631,N_19385,N_19445);
nand U19632 (N_19632,N_19455,N_19439);
xor U19633 (N_19633,N_19373,N_19453);
or U19634 (N_19634,N_19410,N_19385);
and U19635 (N_19635,N_19355,N_19494);
xnor U19636 (N_19636,N_19385,N_19392);
or U19637 (N_19637,N_19359,N_19470);
and U19638 (N_19638,N_19250,N_19493);
nor U19639 (N_19639,N_19391,N_19267);
and U19640 (N_19640,N_19323,N_19286);
nor U19641 (N_19641,N_19310,N_19419);
nor U19642 (N_19642,N_19499,N_19327);
or U19643 (N_19643,N_19253,N_19472);
or U19644 (N_19644,N_19343,N_19294);
xnor U19645 (N_19645,N_19378,N_19420);
or U19646 (N_19646,N_19452,N_19433);
nand U19647 (N_19647,N_19449,N_19406);
or U19648 (N_19648,N_19309,N_19487);
or U19649 (N_19649,N_19484,N_19314);
and U19650 (N_19650,N_19338,N_19344);
nand U19651 (N_19651,N_19317,N_19409);
nor U19652 (N_19652,N_19298,N_19263);
or U19653 (N_19653,N_19318,N_19259);
or U19654 (N_19654,N_19425,N_19435);
and U19655 (N_19655,N_19356,N_19478);
xnor U19656 (N_19656,N_19352,N_19270);
or U19657 (N_19657,N_19453,N_19406);
xor U19658 (N_19658,N_19497,N_19495);
or U19659 (N_19659,N_19318,N_19347);
and U19660 (N_19660,N_19472,N_19328);
or U19661 (N_19661,N_19357,N_19336);
nand U19662 (N_19662,N_19276,N_19495);
or U19663 (N_19663,N_19325,N_19495);
nand U19664 (N_19664,N_19447,N_19402);
xor U19665 (N_19665,N_19447,N_19493);
nand U19666 (N_19666,N_19317,N_19346);
and U19667 (N_19667,N_19455,N_19402);
nor U19668 (N_19668,N_19351,N_19436);
nand U19669 (N_19669,N_19476,N_19301);
or U19670 (N_19670,N_19293,N_19454);
and U19671 (N_19671,N_19276,N_19417);
nand U19672 (N_19672,N_19437,N_19446);
xnor U19673 (N_19673,N_19387,N_19370);
xnor U19674 (N_19674,N_19267,N_19335);
nor U19675 (N_19675,N_19436,N_19345);
nor U19676 (N_19676,N_19411,N_19299);
nor U19677 (N_19677,N_19311,N_19342);
nor U19678 (N_19678,N_19358,N_19491);
nand U19679 (N_19679,N_19409,N_19424);
nand U19680 (N_19680,N_19359,N_19289);
or U19681 (N_19681,N_19351,N_19289);
nand U19682 (N_19682,N_19269,N_19383);
xor U19683 (N_19683,N_19291,N_19261);
or U19684 (N_19684,N_19453,N_19401);
and U19685 (N_19685,N_19484,N_19441);
nand U19686 (N_19686,N_19405,N_19349);
and U19687 (N_19687,N_19254,N_19408);
nor U19688 (N_19688,N_19400,N_19430);
nor U19689 (N_19689,N_19366,N_19370);
nor U19690 (N_19690,N_19376,N_19320);
nor U19691 (N_19691,N_19321,N_19428);
or U19692 (N_19692,N_19387,N_19336);
nand U19693 (N_19693,N_19495,N_19395);
and U19694 (N_19694,N_19274,N_19258);
and U19695 (N_19695,N_19478,N_19291);
nand U19696 (N_19696,N_19476,N_19394);
and U19697 (N_19697,N_19403,N_19402);
and U19698 (N_19698,N_19294,N_19338);
xnor U19699 (N_19699,N_19459,N_19268);
xor U19700 (N_19700,N_19329,N_19279);
nor U19701 (N_19701,N_19472,N_19283);
and U19702 (N_19702,N_19268,N_19405);
nand U19703 (N_19703,N_19437,N_19380);
nand U19704 (N_19704,N_19446,N_19393);
nand U19705 (N_19705,N_19367,N_19433);
xor U19706 (N_19706,N_19478,N_19380);
and U19707 (N_19707,N_19459,N_19275);
nand U19708 (N_19708,N_19359,N_19324);
xor U19709 (N_19709,N_19334,N_19286);
xnor U19710 (N_19710,N_19312,N_19492);
nor U19711 (N_19711,N_19450,N_19385);
xor U19712 (N_19712,N_19409,N_19290);
nand U19713 (N_19713,N_19408,N_19309);
nand U19714 (N_19714,N_19380,N_19486);
or U19715 (N_19715,N_19498,N_19367);
or U19716 (N_19716,N_19377,N_19499);
or U19717 (N_19717,N_19408,N_19318);
and U19718 (N_19718,N_19411,N_19322);
nor U19719 (N_19719,N_19427,N_19491);
and U19720 (N_19720,N_19437,N_19324);
xor U19721 (N_19721,N_19440,N_19344);
nor U19722 (N_19722,N_19322,N_19356);
and U19723 (N_19723,N_19455,N_19445);
xnor U19724 (N_19724,N_19368,N_19485);
nand U19725 (N_19725,N_19279,N_19367);
or U19726 (N_19726,N_19338,N_19477);
nand U19727 (N_19727,N_19263,N_19470);
or U19728 (N_19728,N_19366,N_19349);
nor U19729 (N_19729,N_19458,N_19434);
xor U19730 (N_19730,N_19483,N_19339);
nand U19731 (N_19731,N_19264,N_19458);
nand U19732 (N_19732,N_19255,N_19342);
nand U19733 (N_19733,N_19370,N_19292);
xor U19734 (N_19734,N_19498,N_19376);
nand U19735 (N_19735,N_19327,N_19257);
nor U19736 (N_19736,N_19257,N_19320);
nand U19737 (N_19737,N_19444,N_19330);
nand U19738 (N_19738,N_19332,N_19264);
xnor U19739 (N_19739,N_19280,N_19272);
and U19740 (N_19740,N_19331,N_19320);
xor U19741 (N_19741,N_19348,N_19487);
and U19742 (N_19742,N_19336,N_19363);
xnor U19743 (N_19743,N_19427,N_19256);
or U19744 (N_19744,N_19459,N_19255);
and U19745 (N_19745,N_19265,N_19476);
or U19746 (N_19746,N_19440,N_19323);
and U19747 (N_19747,N_19432,N_19262);
and U19748 (N_19748,N_19311,N_19373);
xor U19749 (N_19749,N_19292,N_19415);
nor U19750 (N_19750,N_19656,N_19644);
nor U19751 (N_19751,N_19734,N_19675);
nor U19752 (N_19752,N_19683,N_19715);
or U19753 (N_19753,N_19698,N_19645);
nor U19754 (N_19754,N_19539,N_19604);
and U19755 (N_19755,N_19592,N_19540);
nand U19756 (N_19756,N_19635,N_19639);
or U19757 (N_19757,N_19659,N_19705);
or U19758 (N_19758,N_19718,N_19717);
nor U19759 (N_19759,N_19682,N_19519);
or U19760 (N_19760,N_19513,N_19660);
and U19761 (N_19761,N_19522,N_19702);
and U19762 (N_19762,N_19652,N_19509);
and U19763 (N_19763,N_19706,N_19551);
and U19764 (N_19764,N_19614,N_19613);
or U19765 (N_19765,N_19628,N_19575);
and U19766 (N_19766,N_19684,N_19500);
xor U19767 (N_19767,N_19603,N_19646);
nor U19768 (N_19768,N_19507,N_19609);
nor U19769 (N_19769,N_19531,N_19523);
or U19770 (N_19770,N_19633,N_19739);
xor U19771 (N_19771,N_19640,N_19524);
nor U19772 (N_19772,N_19710,N_19593);
nand U19773 (N_19773,N_19689,N_19668);
nand U19774 (N_19774,N_19571,N_19587);
xor U19775 (N_19775,N_19733,N_19663);
nor U19776 (N_19776,N_19653,N_19737);
nand U19777 (N_19777,N_19590,N_19637);
and U19778 (N_19778,N_19745,N_19561);
nand U19779 (N_19779,N_19729,N_19529);
xnor U19780 (N_19780,N_19517,N_19709);
nand U19781 (N_19781,N_19670,N_19708);
nand U19782 (N_19782,N_19548,N_19699);
nand U19783 (N_19783,N_19649,N_19555);
and U19784 (N_19784,N_19501,N_19605);
or U19785 (N_19785,N_19667,N_19748);
and U19786 (N_19786,N_19558,N_19695);
and U19787 (N_19787,N_19552,N_19615);
and U19788 (N_19788,N_19678,N_19679);
or U19789 (N_19789,N_19620,N_19665);
nor U19790 (N_19790,N_19688,N_19725);
or U19791 (N_19791,N_19606,N_19572);
nor U19792 (N_19792,N_19677,N_19621);
and U19793 (N_19793,N_19731,N_19631);
nand U19794 (N_19794,N_19619,N_19657);
nand U19795 (N_19795,N_19690,N_19582);
nand U19796 (N_19796,N_19610,N_19693);
and U19797 (N_19797,N_19505,N_19636);
or U19798 (N_19798,N_19586,N_19749);
nor U19799 (N_19799,N_19630,N_19553);
and U19800 (N_19800,N_19602,N_19594);
and U19801 (N_19801,N_19579,N_19691);
nand U19802 (N_19802,N_19697,N_19658);
nand U19803 (N_19803,N_19574,N_19588);
xnor U19804 (N_19804,N_19578,N_19632);
nor U19805 (N_19805,N_19744,N_19550);
xnor U19806 (N_19806,N_19671,N_19617);
nand U19807 (N_19807,N_19542,N_19591);
nand U19808 (N_19808,N_19589,N_19694);
and U19809 (N_19809,N_19511,N_19712);
nand U19810 (N_19810,N_19692,N_19597);
xnor U19811 (N_19811,N_19685,N_19662);
xnor U19812 (N_19812,N_19612,N_19726);
and U19813 (N_19813,N_19711,N_19673);
or U19814 (N_19814,N_19518,N_19506);
nand U19815 (N_19815,N_19563,N_19568);
and U19816 (N_19816,N_19720,N_19525);
nor U19817 (N_19817,N_19598,N_19569);
nor U19818 (N_19818,N_19573,N_19638);
or U19819 (N_19819,N_19520,N_19567);
xnor U19820 (N_19820,N_19623,N_19565);
nand U19821 (N_19821,N_19504,N_19716);
nor U19822 (N_19822,N_19560,N_19508);
and U19823 (N_19823,N_19747,N_19728);
xnor U19824 (N_19824,N_19641,N_19719);
nor U19825 (N_19825,N_19510,N_19562);
xnor U19826 (N_19826,N_19544,N_19611);
nor U19827 (N_19827,N_19743,N_19625);
or U19828 (N_19828,N_19554,N_19580);
and U19829 (N_19829,N_19650,N_19576);
and U19830 (N_19830,N_19532,N_19541);
and U19831 (N_19831,N_19585,N_19686);
nor U19832 (N_19832,N_19647,N_19700);
nor U19833 (N_19833,N_19570,N_19627);
xor U19834 (N_19834,N_19543,N_19687);
xor U19835 (N_19835,N_19556,N_19669);
xnor U19836 (N_19836,N_19723,N_19629);
nand U19837 (N_19837,N_19584,N_19526);
or U19838 (N_19838,N_19701,N_19714);
nand U19839 (N_19839,N_19537,N_19600);
and U19840 (N_19840,N_19740,N_19549);
xnor U19841 (N_19841,N_19648,N_19727);
nand U19842 (N_19842,N_19742,N_19672);
and U19843 (N_19843,N_19557,N_19704);
nand U19844 (N_19844,N_19547,N_19713);
or U19845 (N_19845,N_19502,N_19696);
xor U19846 (N_19846,N_19622,N_19595);
or U19847 (N_19847,N_19528,N_19746);
nor U19848 (N_19848,N_19536,N_19661);
xor U19849 (N_19849,N_19626,N_19516);
nand U19850 (N_19850,N_19616,N_19607);
xor U19851 (N_19851,N_19608,N_19642);
nand U19852 (N_19852,N_19559,N_19732);
nor U19853 (N_19853,N_19530,N_19533);
nor U19854 (N_19854,N_19666,N_19722);
xor U19855 (N_19855,N_19703,N_19564);
xor U19856 (N_19856,N_19724,N_19545);
or U19857 (N_19857,N_19674,N_19681);
xnor U19858 (N_19858,N_19735,N_19654);
nand U19859 (N_19859,N_19546,N_19521);
nand U19860 (N_19860,N_19515,N_19664);
nor U19861 (N_19861,N_19514,N_19721);
or U19862 (N_19862,N_19577,N_19651);
nor U19863 (N_19863,N_19643,N_19618);
nor U19864 (N_19864,N_19601,N_19707);
or U19865 (N_19865,N_19538,N_19634);
nand U19866 (N_19866,N_19527,N_19736);
nor U19867 (N_19867,N_19624,N_19655);
or U19868 (N_19868,N_19581,N_19680);
or U19869 (N_19869,N_19596,N_19741);
nand U19870 (N_19870,N_19738,N_19503);
nor U19871 (N_19871,N_19534,N_19566);
xor U19872 (N_19872,N_19730,N_19599);
or U19873 (N_19873,N_19535,N_19676);
nor U19874 (N_19874,N_19583,N_19512);
or U19875 (N_19875,N_19606,N_19643);
nand U19876 (N_19876,N_19573,N_19616);
or U19877 (N_19877,N_19592,N_19706);
nor U19878 (N_19878,N_19513,N_19723);
xnor U19879 (N_19879,N_19691,N_19660);
xnor U19880 (N_19880,N_19537,N_19555);
nor U19881 (N_19881,N_19510,N_19633);
or U19882 (N_19882,N_19728,N_19735);
or U19883 (N_19883,N_19560,N_19537);
nor U19884 (N_19884,N_19577,N_19540);
and U19885 (N_19885,N_19525,N_19746);
or U19886 (N_19886,N_19558,N_19619);
nor U19887 (N_19887,N_19552,N_19504);
or U19888 (N_19888,N_19715,N_19529);
nor U19889 (N_19889,N_19544,N_19527);
or U19890 (N_19890,N_19598,N_19641);
or U19891 (N_19891,N_19507,N_19640);
xor U19892 (N_19892,N_19545,N_19687);
or U19893 (N_19893,N_19693,N_19631);
or U19894 (N_19894,N_19670,N_19719);
and U19895 (N_19895,N_19613,N_19715);
nor U19896 (N_19896,N_19561,N_19570);
and U19897 (N_19897,N_19641,N_19748);
nand U19898 (N_19898,N_19725,N_19689);
xnor U19899 (N_19899,N_19746,N_19567);
nor U19900 (N_19900,N_19609,N_19672);
nand U19901 (N_19901,N_19625,N_19581);
and U19902 (N_19902,N_19739,N_19622);
nor U19903 (N_19903,N_19727,N_19693);
or U19904 (N_19904,N_19707,N_19548);
nand U19905 (N_19905,N_19582,N_19566);
xor U19906 (N_19906,N_19500,N_19566);
nand U19907 (N_19907,N_19749,N_19591);
or U19908 (N_19908,N_19660,N_19740);
xor U19909 (N_19909,N_19690,N_19505);
xor U19910 (N_19910,N_19587,N_19509);
and U19911 (N_19911,N_19703,N_19505);
nor U19912 (N_19912,N_19724,N_19697);
nor U19913 (N_19913,N_19745,N_19524);
nand U19914 (N_19914,N_19566,N_19570);
and U19915 (N_19915,N_19744,N_19535);
and U19916 (N_19916,N_19718,N_19510);
and U19917 (N_19917,N_19538,N_19650);
nand U19918 (N_19918,N_19607,N_19579);
xor U19919 (N_19919,N_19655,N_19746);
or U19920 (N_19920,N_19663,N_19633);
nand U19921 (N_19921,N_19510,N_19594);
and U19922 (N_19922,N_19595,N_19592);
nor U19923 (N_19923,N_19534,N_19621);
and U19924 (N_19924,N_19699,N_19547);
xor U19925 (N_19925,N_19517,N_19669);
nor U19926 (N_19926,N_19735,N_19571);
and U19927 (N_19927,N_19504,N_19625);
or U19928 (N_19928,N_19589,N_19656);
nor U19929 (N_19929,N_19662,N_19545);
or U19930 (N_19930,N_19576,N_19622);
and U19931 (N_19931,N_19640,N_19628);
or U19932 (N_19932,N_19586,N_19631);
nand U19933 (N_19933,N_19522,N_19505);
nor U19934 (N_19934,N_19661,N_19658);
nand U19935 (N_19935,N_19646,N_19668);
nor U19936 (N_19936,N_19562,N_19736);
or U19937 (N_19937,N_19657,N_19505);
nor U19938 (N_19938,N_19508,N_19641);
nand U19939 (N_19939,N_19739,N_19512);
nand U19940 (N_19940,N_19548,N_19581);
xnor U19941 (N_19941,N_19569,N_19501);
nor U19942 (N_19942,N_19726,N_19569);
nand U19943 (N_19943,N_19746,N_19540);
xor U19944 (N_19944,N_19582,N_19613);
nand U19945 (N_19945,N_19601,N_19635);
xor U19946 (N_19946,N_19574,N_19709);
and U19947 (N_19947,N_19603,N_19608);
nand U19948 (N_19948,N_19518,N_19566);
nand U19949 (N_19949,N_19626,N_19655);
and U19950 (N_19950,N_19616,N_19644);
nor U19951 (N_19951,N_19644,N_19518);
or U19952 (N_19952,N_19591,N_19510);
nor U19953 (N_19953,N_19508,N_19696);
nor U19954 (N_19954,N_19713,N_19647);
nor U19955 (N_19955,N_19718,N_19689);
xor U19956 (N_19956,N_19561,N_19579);
nand U19957 (N_19957,N_19714,N_19681);
xor U19958 (N_19958,N_19515,N_19698);
nand U19959 (N_19959,N_19670,N_19573);
xnor U19960 (N_19960,N_19523,N_19598);
or U19961 (N_19961,N_19510,N_19507);
nand U19962 (N_19962,N_19659,N_19687);
or U19963 (N_19963,N_19578,N_19618);
or U19964 (N_19964,N_19660,N_19546);
nor U19965 (N_19965,N_19612,N_19696);
xnor U19966 (N_19966,N_19633,N_19677);
xnor U19967 (N_19967,N_19537,N_19616);
nand U19968 (N_19968,N_19651,N_19555);
nor U19969 (N_19969,N_19631,N_19746);
xor U19970 (N_19970,N_19554,N_19725);
xnor U19971 (N_19971,N_19727,N_19657);
and U19972 (N_19972,N_19653,N_19700);
nand U19973 (N_19973,N_19704,N_19625);
nor U19974 (N_19974,N_19566,N_19748);
or U19975 (N_19975,N_19722,N_19713);
and U19976 (N_19976,N_19714,N_19610);
nor U19977 (N_19977,N_19538,N_19607);
nor U19978 (N_19978,N_19741,N_19735);
xor U19979 (N_19979,N_19603,N_19588);
nor U19980 (N_19980,N_19686,N_19625);
or U19981 (N_19981,N_19742,N_19587);
and U19982 (N_19982,N_19718,N_19745);
and U19983 (N_19983,N_19606,N_19503);
or U19984 (N_19984,N_19732,N_19529);
xnor U19985 (N_19985,N_19676,N_19529);
nand U19986 (N_19986,N_19675,N_19709);
nor U19987 (N_19987,N_19530,N_19547);
xor U19988 (N_19988,N_19573,N_19675);
xnor U19989 (N_19989,N_19749,N_19744);
nor U19990 (N_19990,N_19612,N_19741);
and U19991 (N_19991,N_19564,N_19540);
nor U19992 (N_19992,N_19704,N_19577);
nand U19993 (N_19993,N_19501,N_19683);
or U19994 (N_19994,N_19515,N_19704);
nor U19995 (N_19995,N_19544,N_19605);
or U19996 (N_19996,N_19637,N_19585);
xor U19997 (N_19997,N_19622,N_19675);
xnor U19998 (N_19998,N_19675,N_19641);
or U19999 (N_19999,N_19509,N_19718);
and U20000 (N_20000,N_19792,N_19787);
nand U20001 (N_20001,N_19901,N_19931);
xor U20002 (N_20002,N_19948,N_19842);
or U20003 (N_20003,N_19875,N_19885);
or U20004 (N_20004,N_19850,N_19848);
nor U20005 (N_20005,N_19811,N_19785);
nand U20006 (N_20006,N_19945,N_19813);
and U20007 (N_20007,N_19908,N_19896);
nor U20008 (N_20008,N_19804,N_19976);
nand U20009 (N_20009,N_19796,N_19956);
and U20010 (N_20010,N_19946,N_19910);
or U20011 (N_20011,N_19849,N_19751);
and U20012 (N_20012,N_19835,N_19970);
and U20013 (N_20013,N_19791,N_19822);
or U20014 (N_20014,N_19797,N_19987);
nand U20015 (N_20015,N_19868,N_19851);
or U20016 (N_20016,N_19788,N_19997);
xor U20017 (N_20017,N_19925,N_19818);
xor U20018 (N_20018,N_19795,N_19876);
nand U20019 (N_20019,N_19895,N_19936);
or U20020 (N_20020,N_19864,N_19886);
nand U20021 (N_20021,N_19857,N_19771);
or U20022 (N_20022,N_19928,N_19847);
nor U20023 (N_20023,N_19985,N_19753);
or U20024 (N_20024,N_19855,N_19974);
nor U20025 (N_20025,N_19762,N_19951);
and U20026 (N_20026,N_19932,N_19924);
nor U20027 (N_20027,N_19937,N_19756);
or U20028 (N_20028,N_19870,N_19975);
and U20029 (N_20029,N_19860,N_19774);
or U20030 (N_20030,N_19831,N_19898);
xnor U20031 (N_20031,N_19942,N_19890);
and U20032 (N_20032,N_19790,N_19866);
xnor U20033 (N_20033,N_19917,N_19869);
xnor U20034 (N_20034,N_19837,N_19763);
nand U20035 (N_20035,N_19834,N_19793);
nor U20036 (N_20036,N_19957,N_19999);
or U20037 (N_20037,N_19798,N_19877);
nand U20038 (N_20038,N_19752,N_19784);
xor U20039 (N_20039,N_19960,N_19879);
nor U20040 (N_20040,N_19930,N_19803);
xnor U20041 (N_20041,N_19812,N_19907);
or U20042 (N_20042,N_19846,N_19884);
nor U20043 (N_20043,N_19983,N_19794);
or U20044 (N_20044,N_19909,N_19825);
and U20045 (N_20045,N_19950,N_19780);
and U20046 (N_20046,N_19827,N_19750);
xnor U20047 (N_20047,N_19783,N_19772);
nand U20048 (N_20048,N_19961,N_19761);
nor U20049 (N_20049,N_19754,N_19921);
and U20050 (N_20050,N_19773,N_19897);
nand U20051 (N_20051,N_19964,N_19820);
or U20052 (N_20052,N_19807,N_19990);
xor U20053 (N_20053,N_19767,N_19802);
nor U20054 (N_20054,N_19839,N_19986);
nand U20055 (N_20055,N_19843,N_19815);
or U20056 (N_20056,N_19996,N_19968);
nor U20057 (N_20057,N_19880,N_19903);
and U20058 (N_20058,N_19938,N_19963);
nand U20059 (N_20059,N_19862,N_19891);
nor U20060 (N_20060,N_19958,N_19845);
nand U20061 (N_20061,N_19899,N_19915);
or U20062 (N_20062,N_19760,N_19840);
and U20063 (N_20063,N_19881,N_19995);
nor U20064 (N_20064,N_19782,N_19806);
xor U20065 (N_20065,N_19977,N_19918);
or U20066 (N_20066,N_19856,N_19994);
nor U20067 (N_20067,N_19894,N_19878);
or U20068 (N_20068,N_19913,N_19757);
xnor U20069 (N_20069,N_19872,N_19863);
or U20070 (N_20070,N_19959,N_19759);
nand U20071 (N_20071,N_19765,N_19858);
or U20072 (N_20072,N_19984,N_19871);
nand U20073 (N_20073,N_19799,N_19832);
or U20074 (N_20074,N_19883,N_19982);
or U20075 (N_20075,N_19989,N_19919);
and U20076 (N_20076,N_19852,N_19992);
and U20077 (N_20077,N_19888,N_19904);
nand U20078 (N_20078,N_19927,N_19844);
xnor U20079 (N_20079,N_19865,N_19978);
and U20080 (N_20080,N_19819,N_19912);
nand U20081 (N_20081,N_19941,N_19949);
nand U20082 (N_20082,N_19926,N_19777);
nor U20083 (N_20083,N_19944,N_19882);
and U20084 (N_20084,N_19867,N_19892);
nor U20085 (N_20085,N_19824,N_19965);
nor U20086 (N_20086,N_19947,N_19768);
nand U20087 (N_20087,N_19991,N_19922);
or U20088 (N_20088,N_19955,N_19972);
nand U20089 (N_20089,N_19810,N_19821);
xor U20090 (N_20090,N_19755,N_19778);
or U20091 (N_20091,N_19828,N_19800);
nor U20092 (N_20092,N_19873,N_19902);
or U20093 (N_20093,N_19830,N_19966);
nor U20094 (N_20094,N_19770,N_19816);
and U20095 (N_20095,N_19900,N_19838);
or U20096 (N_20096,N_19859,N_19853);
and U20097 (N_20097,N_19833,N_19998);
and U20098 (N_20098,N_19943,N_19789);
or U20099 (N_20099,N_19980,N_19779);
xor U20100 (N_20100,N_19934,N_19893);
nand U20101 (N_20101,N_19973,N_19988);
nor U20102 (N_20102,N_19939,N_19935);
nand U20103 (N_20103,N_19823,N_19962);
or U20104 (N_20104,N_19874,N_19916);
nor U20105 (N_20105,N_19764,N_19775);
xor U20106 (N_20106,N_19836,N_19952);
nand U20107 (N_20107,N_19905,N_19841);
xor U20108 (N_20108,N_19817,N_19954);
or U20109 (N_20109,N_19906,N_19933);
or U20110 (N_20110,N_19786,N_19776);
or U20111 (N_20111,N_19887,N_19809);
xor U20112 (N_20112,N_19758,N_19923);
xor U20113 (N_20113,N_19993,N_19889);
nand U20114 (N_20114,N_19861,N_19981);
nor U20115 (N_20115,N_19808,N_19805);
nor U20116 (N_20116,N_19914,N_19929);
xnor U20117 (N_20117,N_19829,N_19826);
or U20118 (N_20118,N_19769,N_19979);
xor U20119 (N_20119,N_19971,N_19814);
and U20120 (N_20120,N_19801,N_19940);
nor U20121 (N_20121,N_19854,N_19911);
and U20122 (N_20122,N_19969,N_19967);
nor U20123 (N_20123,N_19781,N_19766);
and U20124 (N_20124,N_19920,N_19953);
xor U20125 (N_20125,N_19892,N_19775);
xor U20126 (N_20126,N_19885,N_19825);
xor U20127 (N_20127,N_19921,N_19750);
or U20128 (N_20128,N_19835,N_19780);
or U20129 (N_20129,N_19896,N_19857);
and U20130 (N_20130,N_19920,N_19935);
or U20131 (N_20131,N_19889,N_19833);
nand U20132 (N_20132,N_19971,N_19829);
xnor U20133 (N_20133,N_19952,N_19809);
xor U20134 (N_20134,N_19928,N_19837);
or U20135 (N_20135,N_19884,N_19906);
or U20136 (N_20136,N_19866,N_19887);
and U20137 (N_20137,N_19883,N_19968);
or U20138 (N_20138,N_19787,N_19898);
nor U20139 (N_20139,N_19787,N_19800);
or U20140 (N_20140,N_19778,N_19829);
and U20141 (N_20141,N_19822,N_19783);
nand U20142 (N_20142,N_19771,N_19777);
nand U20143 (N_20143,N_19856,N_19963);
xnor U20144 (N_20144,N_19995,N_19992);
nand U20145 (N_20145,N_19970,N_19799);
nor U20146 (N_20146,N_19756,N_19989);
xnor U20147 (N_20147,N_19808,N_19991);
xor U20148 (N_20148,N_19869,N_19776);
or U20149 (N_20149,N_19904,N_19968);
nor U20150 (N_20150,N_19963,N_19936);
and U20151 (N_20151,N_19848,N_19948);
nand U20152 (N_20152,N_19956,N_19968);
or U20153 (N_20153,N_19969,N_19784);
and U20154 (N_20154,N_19840,N_19845);
nor U20155 (N_20155,N_19841,N_19984);
nor U20156 (N_20156,N_19940,N_19912);
or U20157 (N_20157,N_19832,N_19892);
xnor U20158 (N_20158,N_19920,N_19799);
nand U20159 (N_20159,N_19810,N_19932);
xnor U20160 (N_20160,N_19771,N_19823);
nor U20161 (N_20161,N_19916,N_19786);
nand U20162 (N_20162,N_19863,N_19769);
nor U20163 (N_20163,N_19851,N_19847);
nand U20164 (N_20164,N_19821,N_19976);
or U20165 (N_20165,N_19876,N_19866);
nand U20166 (N_20166,N_19881,N_19920);
nor U20167 (N_20167,N_19895,N_19969);
xor U20168 (N_20168,N_19981,N_19904);
nor U20169 (N_20169,N_19973,N_19941);
nor U20170 (N_20170,N_19891,N_19974);
nor U20171 (N_20171,N_19822,N_19762);
xor U20172 (N_20172,N_19789,N_19900);
nand U20173 (N_20173,N_19783,N_19777);
nor U20174 (N_20174,N_19894,N_19781);
xor U20175 (N_20175,N_19841,N_19947);
or U20176 (N_20176,N_19788,N_19799);
nor U20177 (N_20177,N_19954,N_19983);
and U20178 (N_20178,N_19990,N_19858);
nand U20179 (N_20179,N_19858,N_19931);
or U20180 (N_20180,N_19912,N_19799);
nor U20181 (N_20181,N_19918,N_19947);
nor U20182 (N_20182,N_19955,N_19855);
nor U20183 (N_20183,N_19886,N_19881);
nor U20184 (N_20184,N_19991,N_19894);
nand U20185 (N_20185,N_19990,N_19973);
nor U20186 (N_20186,N_19881,N_19955);
xnor U20187 (N_20187,N_19761,N_19809);
or U20188 (N_20188,N_19871,N_19847);
nor U20189 (N_20189,N_19784,N_19904);
nor U20190 (N_20190,N_19875,N_19933);
nand U20191 (N_20191,N_19939,N_19781);
xor U20192 (N_20192,N_19872,N_19993);
nand U20193 (N_20193,N_19768,N_19853);
nand U20194 (N_20194,N_19805,N_19765);
or U20195 (N_20195,N_19948,N_19928);
or U20196 (N_20196,N_19801,N_19927);
and U20197 (N_20197,N_19799,N_19935);
or U20198 (N_20198,N_19974,N_19842);
xor U20199 (N_20199,N_19984,N_19773);
xnor U20200 (N_20200,N_19760,N_19868);
xnor U20201 (N_20201,N_19891,N_19819);
and U20202 (N_20202,N_19910,N_19985);
nor U20203 (N_20203,N_19786,N_19891);
nor U20204 (N_20204,N_19869,N_19928);
nand U20205 (N_20205,N_19957,N_19914);
and U20206 (N_20206,N_19776,N_19986);
nor U20207 (N_20207,N_19777,N_19912);
nand U20208 (N_20208,N_19944,N_19821);
nand U20209 (N_20209,N_19865,N_19982);
nor U20210 (N_20210,N_19777,N_19969);
and U20211 (N_20211,N_19823,N_19929);
xnor U20212 (N_20212,N_19976,N_19965);
nor U20213 (N_20213,N_19957,N_19855);
nor U20214 (N_20214,N_19788,N_19970);
or U20215 (N_20215,N_19818,N_19857);
xor U20216 (N_20216,N_19868,N_19958);
or U20217 (N_20217,N_19912,N_19836);
nor U20218 (N_20218,N_19775,N_19861);
or U20219 (N_20219,N_19982,N_19769);
nor U20220 (N_20220,N_19846,N_19800);
nor U20221 (N_20221,N_19857,N_19850);
and U20222 (N_20222,N_19931,N_19750);
nor U20223 (N_20223,N_19908,N_19846);
or U20224 (N_20224,N_19970,N_19965);
nor U20225 (N_20225,N_19982,N_19770);
nand U20226 (N_20226,N_19820,N_19802);
or U20227 (N_20227,N_19922,N_19917);
or U20228 (N_20228,N_19861,N_19907);
xnor U20229 (N_20229,N_19945,N_19958);
or U20230 (N_20230,N_19758,N_19958);
or U20231 (N_20231,N_19942,N_19850);
nand U20232 (N_20232,N_19765,N_19875);
nor U20233 (N_20233,N_19874,N_19987);
nor U20234 (N_20234,N_19847,N_19804);
or U20235 (N_20235,N_19882,N_19943);
nand U20236 (N_20236,N_19947,N_19920);
nand U20237 (N_20237,N_19968,N_19795);
or U20238 (N_20238,N_19943,N_19942);
xnor U20239 (N_20239,N_19933,N_19947);
nor U20240 (N_20240,N_19959,N_19801);
xnor U20241 (N_20241,N_19993,N_19999);
nor U20242 (N_20242,N_19895,N_19784);
nor U20243 (N_20243,N_19818,N_19826);
xnor U20244 (N_20244,N_19798,N_19767);
nand U20245 (N_20245,N_19781,N_19848);
or U20246 (N_20246,N_19968,N_19891);
nand U20247 (N_20247,N_19788,N_19789);
or U20248 (N_20248,N_19799,N_19960);
xnor U20249 (N_20249,N_19791,N_19878);
or U20250 (N_20250,N_20124,N_20051);
nand U20251 (N_20251,N_20138,N_20232);
and U20252 (N_20252,N_20147,N_20167);
or U20253 (N_20253,N_20210,N_20021);
and U20254 (N_20254,N_20187,N_20110);
and U20255 (N_20255,N_20205,N_20047);
or U20256 (N_20256,N_20086,N_20134);
xor U20257 (N_20257,N_20125,N_20236);
nor U20258 (N_20258,N_20239,N_20193);
or U20259 (N_20259,N_20074,N_20178);
and U20260 (N_20260,N_20230,N_20028);
xor U20261 (N_20261,N_20226,N_20234);
nand U20262 (N_20262,N_20188,N_20161);
or U20263 (N_20263,N_20235,N_20029);
nand U20264 (N_20264,N_20071,N_20034);
or U20265 (N_20265,N_20065,N_20093);
xor U20266 (N_20266,N_20160,N_20139);
nand U20267 (N_20267,N_20246,N_20092);
and U20268 (N_20268,N_20038,N_20245);
or U20269 (N_20269,N_20105,N_20208);
nand U20270 (N_20270,N_20025,N_20127);
and U20271 (N_20271,N_20128,N_20222);
nand U20272 (N_20272,N_20227,N_20219);
nor U20273 (N_20273,N_20087,N_20101);
nor U20274 (N_20274,N_20249,N_20141);
or U20275 (N_20275,N_20043,N_20217);
or U20276 (N_20276,N_20094,N_20243);
or U20277 (N_20277,N_20162,N_20069);
nand U20278 (N_20278,N_20186,N_20073);
nand U20279 (N_20279,N_20011,N_20149);
or U20280 (N_20280,N_20185,N_20015);
nand U20281 (N_20281,N_20221,N_20129);
xor U20282 (N_20282,N_20152,N_20049);
and U20283 (N_20283,N_20153,N_20126);
or U20284 (N_20284,N_20039,N_20197);
nand U20285 (N_20285,N_20096,N_20137);
nor U20286 (N_20286,N_20248,N_20118);
and U20287 (N_20287,N_20023,N_20064);
nor U20288 (N_20288,N_20136,N_20080);
xnor U20289 (N_20289,N_20056,N_20014);
or U20290 (N_20290,N_20077,N_20201);
xnor U20291 (N_20291,N_20184,N_20117);
nor U20292 (N_20292,N_20055,N_20169);
and U20293 (N_20293,N_20111,N_20133);
and U20294 (N_20294,N_20224,N_20240);
xor U20295 (N_20295,N_20022,N_20102);
xor U20296 (N_20296,N_20106,N_20066);
nor U20297 (N_20297,N_20070,N_20183);
or U20298 (N_20298,N_20109,N_20067);
nor U20299 (N_20299,N_20114,N_20050);
xor U20300 (N_20300,N_20084,N_20179);
and U20301 (N_20301,N_20012,N_20171);
and U20302 (N_20302,N_20196,N_20181);
xor U20303 (N_20303,N_20182,N_20061);
nand U20304 (N_20304,N_20079,N_20059);
xnor U20305 (N_20305,N_20044,N_20082);
and U20306 (N_20306,N_20237,N_20078);
nand U20307 (N_20307,N_20207,N_20215);
nand U20308 (N_20308,N_20058,N_20233);
and U20309 (N_20309,N_20003,N_20089);
nand U20310 (N_20310,N_20004,N_20030);
xor U20311 (N_20311,N_20140,N_20241);
nand U20312 (N_20312,N_20036,N_20040);
nor U20313 (N_20313,N_20116,N_20091);
nand U20314 (N_20314,N_20006,N_20026);
xnor U20315 (N_20315,N_20228,N_20143);
nand U20316 (N_20316,N_20142,N_20033);
and U20317 (N_20317,N_20103,N_20214);
nor U20318 (N_20318,N_20148,N_20062);
and U20319 (N_20319,N_20122,N_20045);
or U20320 (N_20320,N_20017,N_20155);
and U20321 (N_20321,N_20032,N_20075);
nand U20322 (N_20322,N_20198,N_20041);
xor U20323 (N_20323,N_20027,N_20001);
xor U20324 (N_20324,N_20060,N_20154);
xnor U20325 (N_20325,N_20192,N_20002);
or U20326 (N_20326,N_20159,N_20115);
nand U20327 (N_20327,N_20173,N_20156);
xnor U20328 (N_20328,N_20081,N_20174);
or U20329 (N_20329,N_20010,N_20048);
or U20330 (N_20330,N_20054,N_20016);
nand U20331 (N_20331,N_20019,N_20037);
and U20332 (N_20332,N_20212,N_20083);
nor U20333 (N_20333,N_20009,N_20053);
xnor U20334 (N_20334,N_20052,N_20238);
and U20335 (N_20335,N_20031,N_20170);
or U20336 (N_20336,N_20172,N_20144);
nor U20337 (N_20337,N_20220,N_20225);
and U20338 (N_20338,N_20199,N_20042);
nand U20339 (N_20339,N_20200,N_20145);
xor U20340 (N_20340,N_20191,N_20131);
nor U20341 (N_20341,N_20113,N_20218);
nand U20342 (N_20342,N_20008,N_20132);
and U20343 (N_20343,N_20164,N_20104);
xor U20344 (N_20344,N_20206,N_20046);
nand U20345 (N_20345,N_20189,N_20216);
nand U20346 (N_20346,N_20203,N_20085);
or U20347 (N_20347,N_20165,N_20146);
or U20348 (N_20348,N_20135,N_20112);
xor U20349 (N_20349,N_20000,N_20202);
xor U20350 (N_20350,N_20098,N_20204);
xnor U20351 (N_20351,N_20119,N_20211);
nor U20352 (N_20352,N_20005,N_20057);
or U20353 (N_20353,N_20013,N_20018);
nor U20354 (N_20354,N_20175,N_20108);
nand U20355 (N_20355,N_20024,N_20123);
and U20356 (N_20356,N_20097,N_20242);
and U20357 (N_20357,N_20020,N_20072);
or U20358 (N_20358,N_20076,N_20090);
or U20359 (N_20359,N_20068,N_20130);
nor U20360 (N_20360,N_20120,N_20035);
nand U20361 (N_20361,N_20176,N_20223);
or U20362 (N_20362,N_20194,N_20121);
or U20363 (N_20363,N_20177,N_20095);
xnor U20364 (N_20364,N_20168,N_20209);
xnor U20365 (N_20365,N_20151,N_20244);
or U20366 (N_20366,N_20163,N_20063);
xor U20367 (N_20367,N_20158,N_20213);
or U20368 (N_20368,N_20180,N_20157);
xnor U20369 (N_20369,N_20229,N_20150);
and U20370 (N_20370,N_20099,N_20190);
nor U20371 (N_20371,N_20100,N_20088);
and U20372 (N_20372,N_20247,N_20107);
nor U20373 (N_20373,N_20195,N_20231);
nand U20374 (N_20374,N_20166,N_20007);
nor U20375 (N_20375,N_20065,N_20183);
nor U20376 (N_20376,N_20065,N_20227);
xnor U20377 (N_20377,N_20203,N_20158);
and U20378 (N_20378,N_20153,N_20183);
nor U20379 (N_20379,N_20219,N_20243);
xnor U20380 (N_20380,N_20039,N_20145);
nand U20381 (N_20381,N_20003,N_20056);
nand U20382 (N_20382,N_20014,N_20145);
nor U20383 (N_20383,N_20115,N_20126);
and U20384 (N_20384,N_20178,N_20004);
xor U20385 (N_20385,N_20062,N_20189);
or U20386 (N_20386,N_20000,N_20078);
or U20387 (N_20387,N_20082,N_20161);
and U20388 (N_20388,N_20113,N_20093);
nor U20389 (N_20389,N_20079,N_20167);
and U20390 (N_20390,N_20118,N_20066);
and U20391 (N_20391,N_20194,N_20028);
xnor U20392 (N_20392,N_20074,N_20038);
nor U20393 (N_20393,N_20024,N_20040);
or U20394 (N_20394,N_20146,N_20163);
and U20395 (N_20395,N_20006,N_20222);
xor U20396 (N_20396,N_20058,N_20147);
nand U20397 (N_20397,N_20106,N_20190);
or U20398 (N_20398,N_20141,N_20248);
or U20399 (N_20399,N_20164,N_20090);
or U20400 (N_20400,N_20075,N_20027);
nand U20401 (N_20401,N_20114,N_20236);
xnor U20402 (N_20402,N_20055,N_20217);
xor U20403 (N_20403,N_20061,N_20185);
nand U20404 (N_20404,N_20156,N_20088);
xor U20405 (N_20405,N_20153,N_20135);
nand U20406 (N_20406,N_20070,N_20062);
nand U20407 (N_20407,N_20088,N_20233);
nor U20408 (N_20408,N_20229,N_20178);
nor U20409 (N_20409,N_20200,N_20134);
and U20410 (N_20410,N_20151,N_20018);
or U20411 (N_20411,N_20219,N_20052);
or U20412 (N_20412,N_20130,N_20073);
xnor U20413 (N_20413,N_20021,N_20058);
xor U20414 (N_20414,N_20103,N_20038);
or U20415 (N_20415,N_20066,N_20183);
nor U20416 (N_20416,N_20053,N_20200);
nand U20417 (N_20417,N_20216,N_20248);
nor U20418 (N_20418,N_20178,N_20144);
nand U20419 (N_20419,N_20021,N_20104);
nor U20420 (N_20420,N_20110,N_20214);
or U20421 (N_20421,N_20045,N_20001);
or U20422 (N_20422,N_20000,N_20043);
nand U20423 (N_20423,N_20238,N_20094);
nand U20424 (N_20424,N_20108,N_20232);
or U20425 (N_20425,N_20111,N_20024);
nand U20426 (N_20426,N_20184,N_20066);
nand U20427 (N_20427,N_20011,N_20178);
xnor U20428 (N_20428,N_20075,N_20109);
and U20429 (N_20429,N_20122,N_20249);
nand U20430 (N_20430,N_20042,N_20097);
nor U20431 (N_20431,N_20226,N_20034);
and U20432 (N_20432,N_20226,N_20003);
xor U20433 (N_20433,N_20011,N_20029);
or U20434 (N_20434,N_20023,N_20052);
and U20435 (N_20435,N_20244,N_20236);
and U20436 (N_20436,N_20146,N_20034);
or U20437 (N_20437,N_20145,N_20079);
xor U20438 (N_20438,N_20072,N_20144);
or U20439 (N_20439,N_20195,N_20058);
nand U20440 (N_20440,N_20037,N_20084);
and U20441 (N_20441,N_20133,N_20094);
nand U20442 (N_20442,N_20201,N_20065);
nor U20443 (N_20443,N_20099,N_20103);
nor U20444 (N_20444,N_20087,N_20030);
or U20445 (N_20445,N_20188,N_20137);
nor U20446 (N_20446,N_20021,N_20125);
or U20447 (N_20447,N_20001,N_20185);
or U20448 (N_20448,N_20062,N_20077);
xor U20449 (N_20449,N_20168,N_20221);
nor U20450 (N_20450,N_20011,N_20021);
or U20451 (N_20451,N_20200,N_20197);
nand U20452 (N_20452,N_20187,N_20073);
xor U20453 (N_20453,N_20021,N_20176);
nand U20454 (N_20454,N_20217,N_20181);
and U20455 (N_20455,N_20125,N_20121);
and U20456 (N_20456,N_20169,N_20030);
nand U20457 (N_20457,N_20132,N_20131);
nand U20458 (N_20458,N_20223,N_20148);
nand U20459 (N_20459,N_20038,N_20169);
xnor U20460 (N_20460,N_20159,N_20201);
nand U20461 (N_20461,N_20111,N_20229);
and U20462 (N_20462,N_20115,N_20048);
or U20463 (N_20463,N_20068,N_20139);
xor U20464 (N_20464,N_20133,N_20134);
nor U20465 (N_20465,N_20237,N_20248);
xnor U20466 (N_20466,N_20089,N_20188);
xor U20467 (N_20467,N_20070,N_20052);
and U20468 (N_20468,N_20177,N_20049);
or U20469 (N_20469,N_20061,N_20035);
or U20470 (N_20470,N_20235,N_20159);
and U20471 (N_20471,N_20110,N_20234);
nor U20472 (N_20472,N_20154,N_20004);
nor U20473 (N_20473,N_20143,N_20200);
nand U20474 (N_20474,N_20134,N_20071);
or U20475 (N_20475,N_20141,N_20191);
xor U20476 (N_20476,N_20069,N_20225);
or U20477 (N_20477,N_20077,N_20204);
and U20478 (N_20478,N_20063,N_20157);
nand U20479 (N_20479,N_20125,N_20135);
nor U20480 (N_20480,N_20122,N_20141);
nand U20481 (N_20481,N_20118,N_20111);
nand U20482 (N_20482,N_20193,N_20014);
nor U20483 (N_20483,N_20009,N_20035);
xor U20484 (N_20484,N_20215,N_20001);
and U20485 (N_20485,N_20014,N_20016);
nor U20486 (N_20486,N_20153,N_20019);
nor U20487 (N_20487,N_20186,N_20195);
xnor U20488 (N_20488,N_20090,N_20136);
and U20489 (N_20489,N_20159,N_20049);
nor U20490 (N_20490,N_20070,N_20248);
nand U20491 (N_20491,N_20076,N_20026);
and U20492 (N_20492,N_20244,N_20072);
nor U20493 (N_20493,N_20217,N_20170);
nand U20494 (N_20494,N_20158,N_20081);
xor U20495 (N_20495,N_20131,N_20009);
nor U20496 (N_20496,N_20118,N_20017);
nor U20497 (N_20497,N_20239,N_20147);
xor U20498 (N_20498,N_20112,N_20199);
and U20499 (N_20499,N_20087,N_20163);
and U20500 (N_20500,N_20416,N_20377);
nand U20501 (N_20501,N_20456,N_20452);
or U20502 (N_20502,N_20408,N_20251);
nor U20503 (N_20503,N_20401,N_20438);
nor U20504 (N_20504,N_20369,N_20422);
nor U20505 (N_20505,N_20261,N_20449);
or U20506 (N_20506,N_20287,N_20361);
nand U20507 (N_20507,N_20352,N_20492);
or U20508 (N_20508,N_20347,N_20292);
nand U20509 (N_20509,N_20488,N_20411);
nand U20510 (N_20510,N_20354,N_20450);
and U20511 (N_20511,N_20472,N_20406);
and U20512 (N_20512,N_20447,N_20436);
and U20513 (N_20513,N_20274,N_20433);
nor U20514 (N_20514,N_20388,N_20439);
and U20515 (N_20515,N_20442,N_20282);
nor U20516 (N_20516,N_20493,N_20262);
nor U20517 (N_20517,N_20276,N_20333);
nor U20518 (N_20518,N_20288,N_20353);
nand U20519 (N_20519,N_20463,N_20397);
nor U20520 (N_20520,N_20336,N_20345);
or U20521 (N_20521,N_20289,N_20253);
and U20522 (N_20522,N_20327,N_20317);
nor U20523 (N_20523,N_20443,N_20350);
xor U20524 (N_20524,N_20476,N_20432);
nor U20525 (N_20525,N_20268,N_20480);
or U20526 (N_20526,N_20426,N_20373);
and U20527 (N_20527,N_20475,N_20425);
nand U20528 (N_20528,N_20257,N_20330);
nand U20529 (N_20529,N_20474,N_20338);
and U20530 (N_20530,N_20356,N_20269);
nand U20531 (N_20531,N_20371,N_20351);
nand U20532 (N_20532,N_20305,N_20363);
and U20533 (N_20533,N_20477,N_20465);
nand U20534 (N_20534,N_20483,N_20491);
nand U20535 (N_20535,N_20484,N_20300);
and U20536 (N_20536,N_20283,N_20277);
or U20537 (N_20537,N_20427,N_20271);
and U20538 (N_20538,N_20420,N_20295);
nor U20539 (N_20539,N_20360,N_20340);
and U20540 (N_20540,N_20368,N_20323);
nand U20541 (N_20541,N_20322,N_20272);
xnor U20542 (N_20542,N_20342,N_20429);
xor U20543 (N_20543,N_20349,N_20306);
xor U20544 (N_20544,N_20309,N_20403);
or U20545 (N_20545,N_20421,N_20281);
xor U20546 (N_20546,N_20417,N_20307);
xor U20547 (N_20547,N_20355,N_20337);
and U20548 (N_20548,N_20339,N_20486);
nand U20549 (N_20549,N_20409,N_20490);
nand U20550 (N_20550,N_20376,N_20335);
xnor U20551 (N_20551,N_20441,N_20326);
xor U20552 (N_20552,N_20428,N_20348);
xnor U20553 (N_20553,N_20263,N_20407);
nand U20554 (N_20554,N_20270,N_20334);
or U20555 (N_20555,N_20259,N_20479);
nor U20556 (N_20556,N_20423,N_20460);
or U20557 (N_20557,N_20255,N_20386);
xnor U20558 (N_20558,N_20390,N_20294);
and U20559 (N_20559,N_20412,N_20383);
xnor U20560 (N_20560,N_20310,N_20487);
xnor U20561 (N_20561,N_20466,N_20458);
or U20562 (N_20562,N_20256,N_20446);
nand U20563 (N_20563,N_20316,N_20258);
nand U20564 (N_20564,N_20343,N_20324);
and U20565 (N_20565,N_20481,N_20329);
nor U20566 (N_20566,N_20328,N_20318);
nor U20567 (N_20567,N_20413,N_20320);
nand U20568 (N_20568,N_20430,N_20284);
nor U20569 (N_20569,N_20489,N_20457);
nor U20570 (N_20570,N_20266,N_20332);
xor U20571 (N_20571,N_20496,N_20357);
and U20572 (N_20572,N_20293,N_20385);
or U20573 (N_20573,N_20391,N_20437);
nand U20574 (N_20574,N_20264,N_20308);
and U20575 (N_20575,N_20344,N_20455);
and U20576 (N_20576,N_20359,N_20459);
nand U20577 (N_20577,N_20393,N_20431);
or U20578 (N_20578,N_20331,N_20302);
or U20579 (N_20579,N_20448,N_20499);
nor U20580 (N_20580,N_20372,N_20346);
xor U20581 (N_20581,N_20498,N_20473);
xnor U20582 (N_20582,N_20313,N_20399);
xor U20583 (N_20583,N_20415,N_20396);
or U20584 (N_20584,N_20392,N_20410);
and U20585 (N_20585,N_20404,N_20445);
or U20586 (N_20586,N_20303,N_20440);
nor U20587 (N_20587,N_20285,N_20453);
xnor U20588 (N_20588,N_20312,N_20485);
xnor U20589 (N_20589,N_20379,N_20497);
and U20590 (N_20590,N_20341,N_20434);
xnor U20591 (N_20591,N_20250,N_20389);
or U20592 (N_20592,N_20435,N_20362);
xor U20593 (N_20593,N_20400,N_20319);
or U20594 (N_20594,N_20315,N_20286);
and U20595 (N_20595,N_20384,N_20298);
nand U20596 (N_20596,N_20367,N_20311);
nand U20597 (N_20597,N_20380,N_20358);
or U20598 (N_20598,N_20444,N_20402);
and U20599 (N_20599,N_20419,N_20414);
or U20600 (N_20600,N_20275,N_20494);
nor U20601 (N_20601,N_20304,N_20290);
nor U20602 (N_20602,N_20321,N_20365);
or U20603 (N_20603,N_20297,N_20387);
xor U20604 (N_20604,N_20394,N_20418);
or U20605 (N_20605,N_20299,N_20462);
nor U20606 (N_20606,N_20469,N_20482);
nand U20607 (N_20607,N_20382,N_20364);
and U20608 (N_20608,N_20375,N_20314);
or U20609 (N_20609,N_20467,N_20398);
xor U20610 (N_20610,N_20252,N_20291);
and U20611 (N_20611,N_20495,N_20374);
and U20612 (N_20612,N_20325,N_20454);
nand U20613 (N_20613,N_20267,N_20461);
or U20614 (N_20614,N_20405,N_20468);
and U20615 (N_20615,N_20279,N_20265);
and U20616 (N_20616,N_20378,N_20278);
or U20617 (N_20617,N_20451,N_20370);
nor U20618 (N_20618,N_20470,N_20273);
nor U20619 (N_20619,N_20296,N_20254);
nand U20620 (N_20620,N_20280,N_20424);
nor U20621 (N_20621,N_20366,N_20395);
or U20622 (N_20622,N_20301,N_20478);
and U20623 (N_20623,N_20260,N_20464);
xor U20624 (N_20624,N_20471,N_20381);
or U20625 (N_20625,N_20344,N_20373);
nand U20626 (N_20626,N_20261,N_20291);
nor U20627 (N_20627,N_20416,N_20351);
nand U20628 (N_20628,N_20458,N_20477);
nand U20629 (N_20629,N_20296,N_20353);
nand U20630 (N_20630,N_20351,N_20347);
xnor U20631 (N_20631,N_20397,N_20400);
or U20632 (N_20632,N_20366,N_20290);
nand U20633 (N_20633,N_20338,N_20376);
nand U20634 (N_20634,N_20348,N_20400);
and U20635 (N_20635,N_20376,N_20331);
nor U20636 (N_20636,N_20416,N_20331);
xor U20637 (N_20637,N_20337,N_20491);
and U20638 (N_20638,N_20408,N_20489);
and U20639 (N_20639,N_20320,N_20338);
nand U20640 (N_20640,N_20440,N_20412);
nor U20641 (N_20641,N_20414,N_20467);
or U20642 (N_20642,N_20467,N_20444);
and U20643 (N_20643,N_20456,N_20422);
and U20644 (N_20644,N_20346,N_20420);
xor U20645 (N_20645,N_20403,N_20414);
or U20646 (N_20646,N_20317,N_20499);
xnor U20647 (N_20647,N_20307,N_20251);
nor U20648 (N_20648,N_20275,N_20364);
or U20649 (N_20649,N_20336,N_20296);
nor U20650 (N_20650,N_20350,N_20476);
nor U20651 (N_20651,N_20282,N_20265);
nand U20652 (N_20652,N_20299,N_20327);
and U20653 (N_20653,N_20276,N_20265);
or U20654 (N_20654,N_20417,N_20467);
or U20655 (N_20655,N_20315,N_20294);
or U20656 (N_20656,N_20341,N_20274);
xnor U20657 (N_20657,N_20306,N_20297);
and U20658 (N_20658,N_20427,N_20328);
nor U20659 (N_20659,N_20316,N_20434);
or U20660 (N_20660,N_20273,N_20307);
xor U20661 (N_20661,N_20494,N_20479);
nand U20662 (N_20662,N_20310,N_20425);
and U20663 (N_20663,N_20446,N_20362);
or U20664 (N_20664,N_20485,N_20349);
nor U20665 (N_20665,N_20442,N_20406);
xnor U20666 (N_20666,N_20300,N_20383);
xor U20667 (N_20667,N_20314,N_20350);
or U20668 (N_20668,N_20324,N_20264);
or U20669 (N_20669,N_20447,N_20370);
or U20670 (N_20670,N_20379,N_20385);
and U20671 (N_20671,N_20379,N_20271);
nand U20672 (N_20672,N_20381,N_20286);
and U20673 (N_20673,N_20274,N_20335);
and U20674 (N_20674,N_20344,N_20264);
nand U20675 (N_20675,N_20460,N_20287);
nor U20676 (N_20676,N_20444,N_20316);
and U20677 (N_20677,N_20481,N_20402);
nand U20678 (N_20678,N_20388,N_20293);
nor U20679 (N_20679,N_20279,N_20311);
nand U20680 (N_20680,N_20436,N_20431);
nor U20681 (N_20681,N_20480,N_20256);
xnor U20682 (N_20682,N_20352,N_20462);
and U20683 (N_20683,N_20394,N_20355);
or U20684 (N_20684,N_20459,N_20273);
nor U20685 (N_20685,N_20269,N_20256);
nand U20686 (N_20686,N_20408,N_20422);
or U20687 (N_20687,N_20454,N_20498);
and U20688 (N_20688,N_20299,N_20350);
nor U20689 (N_20689,N_20408,N_20477);
and U20690 (N_20690,N_20292,N_20492);
nand U20691 (N_20691,N_20438,N_20336);
xor U20692 (N_20692,N_20373,N_20465);
nor U20693 (N_20693,N_20499,N_20406);
nor U20694 (N_20694,N_20392,N_20378);
or U20695 (N_20695,N_20379,N_20254);
xor U20696 (N_20696,N_20410,N_20447);
xnor U20697 (N_20697,N_20483,N_20438);
or U20698 (N_20698,N_20276,N_20301);
and U20699 (N_20699,N_20370,N_20422);
and U20700 (N_20700,N_20416,N_20463);
nand U20701 (N_20701,N_20436,N_20394);
xnor U20702 (N_20702,N_20465,N_20353);
and U20703 (N_20703,N_20285,N_20303);
or U20704 (N_20704,N_20492,N_20466);
nor U20705 (N_20705,N_20262,N_20304);
xor U20706 (N_20706,N_20410,N_20340);
or U20707 (N_20707,N_20285,N_20487);
nand U20708 (N_20708,N_20444,N_20491);
and U20709 (N_20709,N_20273,N_20435);
or U20710 (N_20710,N_20260,N_20342);
xor U20711 (N_20711,N_20341,N_20400);
and U20712 (N_20712,N_20420,N_20318);
xor U20713 (N_20713,N_20445,N_20328);
or U20714 (N_20714,N_20346,N_20337);
xor U20715 (N_20715,N_20302,N_20467);
xor U20716 (N_20716,N_20450,N_20499);
or U20717 (N_20717,N_20269,N_20413);
nand U20718 (N_20718,N_20417,N_20486);
and U20719 (N_20719,N_20357,N_20278);
xnor U20720 (N_20720,N_20318,N_20376);
nor U20721 (N_20721,N_20293,N_20396);
and U20722 (N_20722,N_20498,N_20415);
nor U20723 (N_20723,N_20464,N_20305);
nor U20724 (N_20724,N_20452,N_20326);
and U20725 (N_20725,N_20462,N_20458);
nor U20726 (N_20726,N_20267,N_20329);
xnor U20727 (N_20727,N_20252,N_20381);
xor U20728 (N_20728,N_20387,N_20363);
nand U20729 (N_20729,N_20374,N_20296);
xor U20730 (N_20730,N_20321,N_20385);
and U20731 (N_20731,N_20499,N_20307);
and U20732 (N_20732,N_20319,N_20266);
or U20733 (N_20733,N_20260,N_20453);
and U20734 (N_20734,N_20476,N_20404);
and U20735 (N_20735,N_20422,N_20381);
nand U20736 (N_20736,N_20325,N_20311);
nor U20737 (N_20737,N_20314,N_20281);
nand U20738 (N_20738,N_20313,N_20366);
and U20739 (N_20739,N_20295,N_20492);
xnor U20740 (N_20740,N_20460,N_20305);
nor U20741 (N_20741,N_20461,N_20334);
nand U20742 (N_20742,N_20295,N_20441);
or U20743 (N_20743,N_20331,N_20289);
xor U20744 (N_20744,N_20304,N_20347);
nor U20745 (N_20745,N_20289,N_20290);
or U20746 (N_20746,N_20263,N_20449);
nor U20747 (N_20747,N_20465,N_20253);
or U20748 (N_20748,N_20407,N_20351);
or U20749 (N_20749,N_20344,N_20391);
or U20750 (N_20750,N_20652,N_20578);
or U20751 (N_20751,N_20564,N_20732);
nor U20752 (N_20752,N_20500,N_20534);
or U20753 (N_20753,N_20747,N_20645);
nand U20754 (N_20754,N_20643,N_20686);
or U20755 (N_20755,N_20667,N_20581);
or U20756 (N_20756,N_20600,N_20687);
xor U20757 (N_20757,N_20634,N_20622);
nor U20758 (N_20758,N_20748,N_20642);
or U20759 (N_20759,N_20736,N_20721);
and U20760 (N_20760,N_20665,N_20654);
nor U20761 (N_20761,N_20726,N_20513);
nor U20762 (N_20762,N_20720,N_20633);
and U20763 (N_20763,N_20698,N_20606);
nand U20764 (N_20764,N_20683,N_20524);
and U20765 (N_20765,N_20708,N_20531);
xor U20766 (N_20766,N_20532,N_20505);
xnor U20767 (N_20767,N_20678,N_20657);
and U20768 (N_20768,N_20680,N_20696);
and U20769 (N_20769,N_20653,N_20663);
nor U20770 (N_20770,N_20681,N_20662);
nor U20771 (N_20771,N_20685,N_20629);
and U20772 (N_20772,N_20504,N_20515);
xor U20773 (N_20773,N_20547,N_20517);
and U20774 (N_20774,N_20546,N_20553);
or U20775 (N_20775,N_20670,N_20635);
nand U20776 (N_20776,N_20571,N_20527);
nand U20777 (N_20777,N_20522,N_20697);
xor U20778 (N_20778,N_20742,N_20668);
nor U20779 (N_20779,N_20567,N_20511);
xnor U20780 (N_20780,N_20743,N_20577);
and U20781 (N_20781,N_20509,N_20576);
nor U20782 (N_20782,N_20684,N_20514);
or U20783 (N_20783,N_20714,N_20636);
or U20784 (N_20784,N_20519,N_20614);
and U20785 (N_20785,N_20554,N_20594);
or U20786 (N_20786,N_20692,N_20619);
xor U20787 (N_20787,N_20722,N_20529);
nand U20788 (N_20788,N_20583,N_20612);
nor U20789 (N_20789,N_20566,N_20701);
xnor U20790 (N_20790,N_20510,N_20664);
xor U20791 (N_20791,N_20521,N_20580);
or U20792 (N_20792,N_20723,N_20711);
or U20793 (N_20793,N_20725,N_20617);
xor U20794 (N_20794,N_20674,N_20604);
xnor U20795 (N_20795,N_20618,N_20733);
nor U20796 (N_20796,N_20632,N_20609);
nor U20797 (N_20797,N_20535,N_20691);
nor U20798 (N_20798,N_20630,N_20512);
and U20799 (N_20799,N_20506,N_20565);
nor U20800 (N_20800,N_20658,N_20563);
and U20801 (N_20801,N_20693,N_20501);
nand U20802 (N_20802,N_20699,N_20575);
and U20803 (N_20803,N_20560,N_20637);
and U20804 (N_20804,N_20682,N_20608);
xnor U20805 (N_20805,N_20562,N_20555);
nand U20806 (N_20806,N_20556,N_20741);
or U20807 (N_20807,N_20628,N_20574);
nand U20808 (N_20808,N_20552,N_20688);
and U20809 (N_20809,N_20666,N_20738);
and U20810 (N_20810,N_20620,N_20702);
and U20811 (N_20811,N_20719,N_20689);
and U20812 (N_20812,N_20536,N_20705);
xnor U20813 (N_20813,N_20558,N_20650);
xor U20814 (N_20814,N_20731,N_20585);
and U20815 (N_20815,N_20729,N_20543);
xor U20816 (N_20816,N_20605,N_20598);
xor U20817 (N_20817,N_20737,N_20727);
and U20818 (N_20818,N_20623,N_20542);
nor U20819 (N_20819,N_20710,N_20525);
nand U20820 (N_20820,N_20610,N_20584);
xor U20821 (N_20821,N_20621,N_20545);
and U20822 (N_20822,N_20707,N_20713);
or U20823 (N_20823,N_20591,N_20669);
nand U20824 (N_20824,N_20728,N_20588);
or U20825 (N_20825,N_20596,N_20656);
nor U20826 (N_20826,N_20589,N_20603);
xor U20827 (N_20827,N_20661,N_20508);
or U20828 (N_20828,N_20744,N_20539);
xnor U20829 (N_20829,N_20557,N_20526);
or U20830 (N_20830,N_20549,N_20695);
or U20831 (N_20831,N_20587,N_20651);
and U20832 (N_20832,N_20572,N_20616);
nand U20833 (N_20833,N_20538,N_20700);
nor U20834 (N_20834,N_20615,N_20551);
nor U20835 (N_20835,N_20735,N_20715);
nand U20836 (N_20836,N_20592,N_20520);
nor U20837 (N_20837,N_20749,N_20746);
and U20838 (N_20838,N_20679,N_20640);
xor U20839 (N_20839,N_20627,N_20646);
or U20840 (N_20840,N_20694,N_20582);
nor U20841 (N_20841,N_20676,N_20595);
nor U20842 (N_20842,N_20639,N_20641);
and U20843 (N_20843,N_20659,N_20590);
or U20844 (N_20844,N_20660,N_20631);
nand U20845 (N_20845,N_20671,N_20550);
nor U20846 (N_20846,N_20673,N_20611);
xor U20847 (N_20847,N_20706,N_20734);
nand U20848 (N_20848,N_20613,N_20644);
and U20849 (N_20849,N_20625,N_20607);
nand U20850 (N_20850,N_20724,N_20675);
or U20851 (N_20851,N_20507,N_20739);
nor U20852 (N_20852,N_20709,N_20648);
and U20853 (N_20853,N_20533,N_20569);
xnor U20854 (N_20854,N_20599,N_20677);
or U20855 (N_20855,N_20544,N_20561);
or U20856 (N_20856,N_20540,N_20537);
xnor U20857 (N_20857,N_20638,N_20672);
nor U20858 (N_20858,N_20649,N_20716);
or U20859 (N_20859,N_20559,N_20745);
and U20860 (N_20860,N_20528,N_20573);
and U20861 (N_20861,N_20690,N_20597);
xnor U20862 (N_20862,N_20602,N_20518);
xnor U20863 (N_20863,N_20655,N_20718);
or U20864 (N_20864,N_20704,N_20717);
and U20865 (N_20865,N_20624,N_20548);
nor U20866 (N_20866,N_20647,N_20579);
xor U20867 (N_20867,N_20530,N_20730);
and U20868 (N_20868,N_20516,N_20503);
nor U20869 (N_20869,N_20568,N_20626);
or U20870 (N_20870,N_20601,N_20703);
nand U20871 (N_20871,N_20502,N_20570);
xnor U20872 (N_20872,N_20593,N_20523);
and U20873 (N_20873,N_20712,N_20586);
nand U20874 (N_20874,N_20740,N_20541);
nor U20875 (N_20875,N_20732,N_20696);
or U20876 (N_20876,N_20541,N_20542);
nor U20877 (N_20877,N_20560,N_20734);
nand U20878 (N_20878,N_20545,N_20524);
and U20879 (N_20879,N_20652,N_20503);
nor U20880 (N_20880,N_20659,N_20600);
nor U20881 (N_20881,N_20739,N_20535);
or U20882 (N_20882,N_20682,N_20610);
or U20883 (N_20883,N_20737,N_20649);
or U20884 (N_20884,N_20737,N_20606);
nor U20885 (N_20885,N_20685,N_20655);
or U20886 (N_20886,N_20696,N_20500);
nor U20887 (N_20887,N_20511,N_20689);
xor U20888 (N_20888,N_20700,N_20549);
or U20889 (N_20889,N_20521,N_20732);
nor U20890 (N_20890,N_20583,N_20642);
or U20891 (N_20891,N_20736,N_20595);
and U20892 (N_20892,N_20610,N_20748);
and U20893 (N_20893,N_20603,N_20654);
or U20894 (N_20894,N_20703,N_20535);
xor U20895 (N_20895,N_20692,N_20570);
nand U20896 (N_20896,N_20513,N_20501);
or U20897 (N_20897,N_20591,N_20630);
or U20898 (N_20898,N_20609,N_20582);
nor U20899 (N_20899,N_20693,N_20650);
nor U20900 (N_20900,N_20555,N_20665);
nor U20901 (N_20901,N_20633,N_20606);
nand U20902 (N_20902,N_20599,N_20719);
and U20903 (N_20903,N_20735,N_20617);
xor U20904 (N_20904,N_20575,N_20656);
and U20905 (N_20905,N_20674,N_20598);
nand U20906 (N_20906,N_20650,N_20697);
nand U20907 (N_20907,N_20608,N_20526);
nor U20908 (N_20908,N_20638,N_20701);
or U20909 (N_20909,N_20561,N_20610);
xnor U20910 (N_20910,N_20735,N_20508);
nand U20911 (N_20911,N_20652,N_20687);
nand U20912 (N_20912,N_20741,N_20553);
nand U20913 (N_20913,N_20504,N_20744);
or U20914 (N_20914,N_20583,N_20689);
nor U20915 (N_20915,N_20539,N_20581);
nand U20916 (N_20916,N_20701,N_20677);
nor U20917 (N_20917,N_20718,N_20653);
nor U20918 (N_20918,N_20560,N_20639);
nand U20919 (N_20919,N_20690,N_20666);
nor U20920 (N_20920,N_20653,N_20511);
or U20921 (N_20921,N_20602,N_20749);
nor U20922 (N_20922,N_20546,N_20550);
or U20923 (N_20923,N_20526,N_20685);
nor U20924 (N_20924,N_20669,N_20705);
or U20925 (N_20925,N_20504,N_20613);
or U20926 (N_20926,N_20638,N_20719);
or U20927 (N_20927,N_20589,N_20601);
xor U20928 (N_20928,N_20594,N_20625);
and U20929 (N_20929,N_20585,N_20653);
or U20930 (N_20930,N_20648,N_20723);
nand U20931 (N_20931,N_20645,N_20526);
nand U20932 (N_20932,N_20598,N_20626);
nor U20933 (N_20933,N_20512,N_20744);
xor U20934 (N_20934,N_20608,N_20618);
or U20935 (N_20935,N_20734,N_20710);
nand U20936 (N_20936,N_20585,N_20713);
nand U20937 (N_20937,N_20679,N_20601);
nand U20938 (N_20938,N_20591,N_20713);
and U20939 (N_20939,N_20593,N_20598);
and U20940 (N_20940,N_20651,N_20517);
nor U20941 (N_20941,N_20717,N_20581);
and U20942 (N_20942,N_20742,N_20589);
and U20943 (N_20943,N_20683,N_20657);
and U20944 (N_20944,N_20633,N_20569);
and U20945 (N_20945,N_20530,N_20604);
and U20946 (N_20946,N_20615,N_20670);
and U20947 (N_20947,N_20557,N_20611);
and U20948 (N_20948,N_20702,N_20743);
and U20949 (N_20949,N_20504,N_20592);
nor U20950 (N_20950,N_20562,N_20729);
nand U20951 (N_20951,N_20671,N_20661);
nor U20952 (N_20952,N_20542,N_20528);
or U20953 (N_20953,N_20612,N_20728);
and U20954 (N_20954,N_20561,N_20719);
and U20955 (N_20955,N_20615,N_20586);
nand U20956 (N_20956,N_20710,N_20721);
nand U20957 (N_20957,N_20685,N_20502);
and U20958 (N_20958,N_20704,N_20658);
or U20959 (N_20959,N_20728,N_20724);
or U20960 (N_20960,N_20566,N_20606);
and U20961 (N_20961,N_20744,N_20704);
nor U20962 (N_20962,N_20684,N_20660);
xnor U20963 (N_20963,N_20547,N_20578);
nand U20964 (N_20964,N_20542,N_20693);
xnor U20965 (N_20965,N_20626,N_20733);
and U20966 (N_20966,N_20573,N_20589);
nor U20967 (N_20967,N_20705,N_20730);
or U20968 (N_20968,N_20507,N_20509);
or U20969 (N_20969,N_20576,N_20739);
nor U20970 (N_20970,N_20659,N_20680);
nor U20971 (N_20971,N_20504,N_20517);
or U20972 (N_20972,N_20651,N_20518);
nor U20973 (N_20973,N_20522,N_20581);
and U20974 (N_20974,N_20532,N_20673);
or U20975 (N_20975,N_20597,N_20604);
and U20976 (N_20976,N_20598,N_20689);
nor U20977 (N_20977,N_20600,N_20648);
and U20978 (N_20978,N_20583,N_20688);
nor U20979 (N_20979,N_20502,N_20503);
and U20980 (N_20980,N_20699,N_20565);
and U20981 (N_20981,N_20662,N_20658);
nor U20982 (N_20982,N_20585,N_20598);
xnor U20983 (N_20983,N_20712,N_20620);
or U20984 (N_20984,N_20728,N_20654);
xor U20985 (N_20985,N_20706,N_20595);
or U20986 (N_20986,N_20541,N_20620);
and U20987 (N_20987,N_20645,N_20517);
and U20988 (N_20988,N_20559,N_20670);
xnor U20989 (N_20989,N_20574,N_20712);
nor U20990 (N_20990,N_20717,N_20742);
and U20991 (N_20991,N_20665,N_20684);
and U20992 (N_20992,N_20669,N_20728);
or U20993 (N_20993,N_20543,N_20706);
xnor U20994 (N_20994,N_20663,N_20519);
xor U20995 (N_20995,N_20569,N_20541);
nor U20996 (N_20996,N_20577,N_20575);
and U20997 (N_20997,N_20616,N_20542);
nand U20998 (N_20998,N_20613,N_20505);
nand U20999 (N_20999,N_20618,N_20547);
nand U21000 (N_21000,N_20932,N_20915);
nor U21001 (N_21001,N_20966,N_20789);
and U21002 (N_21002,N_20767,N_20862);
nand U21003 (N_21003,N_20810,N_20913);
xnor U21004 (N_21004,N_20931,N_20845);
or U21005 (N_21005,N_20909,N_20800);
nor U21006 (N_21006,N_20930,N_20993);
or U21007 (N_21007,N_20837,N_20847);
nand U21008 (N_21008,N_20998,N_20826);
nor U21009 (N_21009,N_20790,N_20763);
and U21010 (N_21010,N_20924,N_20971);
xor U21011 (N_21011,N_20900,N_20921);
xnor U21012 (N_21012,N_20944,N_20755);
or U21013 (N_21013,N_20779,N_20990);
nand U21014 (N_21014,N_20877,N_20896);
and U21015 (N_21015,N_20916,N_20815);
nor U21016 (N_21016,N_20906,N_20936);
nor U21017 (N_21017,N_20866,N_20824);
nor U21018 (N_21018,N_20798,N_20761);
or U21019 (N_21019,N_20939,N_20899);
nor U21020 (N_21020,N_20927,N_20849);
and U21021 (N_21021,N_20951,N_20961);
nand U21022 (N_21022,N_20994,N_20992);
xor U21023 (N_21023,N_20928,N_20867);
or U21024 (N_21024,N_20969,N_20783);
and U21025 (N_21025,N_20912,N_20801);
xnor U21026 (N_21026,N_20859,N_20978);
nor U21027 (N_21027,N_20943,N_20781);
xor U21028 (N_21028,N_20777,N_20856);
nand U21029 (N_21029,N_20977,N_20982);
nand U21030 (N_21030,N_20773,N_20965);
and U21031 (N_21031,N_20942,N_20959);
nand U21032 (N_21032,N_20843,N_20883);
and U21033 (N_21033,N_20973,N_20769);
or U21034 (N_21034,N_20934,N_20811);
nand U21035 (N_21035,N_20898,N_20803);
nor U21036 (N_21036,N_20879,N_20980);
nand U21037 (N_21037,N_20793,N_20886);
or U21038 (N_21038,N_20870,N_20764);
nand U21039 (N_21039,N_20771,N_20937);
and U21040 (N_21040,N_20786,N_20788);
or U21041 (N_21041,N_20822,N_20825);
and U21042 (N_21042,N_20947,N_20989);
or U21043 (N_21043,N_20981,N_20950);
and U21044 (N_21044,N_20860,N_20817);
nand U21045 (N_21045,N_20920,N_20890);
nand U21046 (N_21046,N_20888,N_20938);
nand U21047 (N_21047,N_20832,N_20850);
nor U21048 (N_21048,N_20751,N_20882);
or U21049 (N_21049,N_20858,N_20857);
or U21050 (N_21050,N_20772,N_20967);
xor U21051 (N_21051,N_20794,N_20956);
or U21052 (N_21052,N_20997,N_20820);
and U21053 (N_21053,N_20902,N_20756);
nand U21054 (N_21054,N_20952,N_20754);
nand U21055 (N_21055,N_20897,N_20910);
xor U21056 (N_21056,N_20799,N_20917);
and U21057 (N_21057,N_20878,N_20809);
and U21058 (N_21058,N_20874,N_20988);
and U21059 (N_21059,N_20983,N_20962);
xnor U21060 (N_21060,N_20975,N_20923);
xor U21061 (N_21061,N_20808,N_20797);
nand U21062 (N_21062,N_20835,N_20868);
and U21063 (N_21063,N_20829,N_20972);
and U21064 (N_21064,N_20758,N_20796);
xnor U21065 (N_21065,N_20831,N_20821);
nand U21066 (N_21066,N_20833,N_20984);
nand U21067 (N_21067,N_20986,N_20871);
or U21068 (N_21068,N_20848,N_20907);
or U21069 (N_21069,N_20827,N_20949);
and U21070 (N_21070,N_20863,N_20816);
nand U21071 (N_21071,N_20855,N_20887);
nand U21072 (N_21072,N_20861,N_20834);
nor U21073 (N_21073,N_20974,N_20918);
nor U21074 (N_21074,N_20880,N_20753);
or U21075 (N_21075,N_20804,N_20881);
and U21076 (N_21076,N_20819,N_20846);
nor U21077 (N_21077,N_20894,N_20784);
or U21078 (N_21078,N_20780,N_20873);
nor U21079 (N_21079,N_20941,N_20979);
and U21080 (N_21080,N_20933,N_20991);
xor U21081 (N_21081,N_20987,N_20935);
nand U21082 (N_21082,N_20812,N_20760);
and U21083 (N_21083,N_20778,N_20964);
xnor U21084 (N_21084,N_20785,N_20791);
and U21085 (N_21085,N_20852,N_20940);
and U21086 (N_21086,N_20953,N_20818);
or U21087 (N_21087,N_20922,N_20995);
nor U21088 (N_21088,N_20851,N_20813);
nor U21089 (N_21089,N_20946,N_20814);
xor U21090 (N_21090,N_20854,N_20948);
or U21091 (N_21091,N_20872,N_20976);
nor U21092 (N_21092,N_20774,N_20752);
or U21093 (N_21093,N_20792,N_20842);
nand U21094 (N_21094,N_20963,N_20839);
xnor U21095 (N_21095,N_20806,N_20807);
nor U21096 (N_21096,N_20911,N_20840);
nand U21097 (N_21097,N_20958,N_20765);
and U21098 (N_21098,N_20823,N_20954);
nor U21099 (N_21099,N_20838,N_20955);
or U21100 (N_21100,N_20885,N_20929);
nor U21101 (N_21101,N_20768,N_20762);
nor U21102 (N_21102,N_20853,N_20892);
and U21103 (N_21103,N_20828,N_20795);
nor U21104 (N_21104,N_20901,N_20905);
nand U21105 (N_21105,N_20893,N_20970);
xor U21106 (N_21106,N_20841,N_20919);
nand U21107 (N_21107,N_20957,N_20782);
nor U21108 (N_21108,N_20914,N_20757);
nand U21109 (N_21109,N_20999,N_20750);
nor U21110 (N_21110,N_20869,N_20770);
nand U21111 (N_21111,N_20985,N_20875);
xnor U21112 (N_21112,N_20830,N_20925);
or U21113 (N_21113,N_20775,N_20996);
and U21114 (N_21114,N_20864,N_20805);
or U21115 (N_21115,N_20891,N_20759);
xor U21116 (N_21116,N_20960,N_20908);
and U21117 (N_21117,N_20904,N_20903);
xnor U21118 (N_21118,N_20884,N_20968);
and U21119 (N_21119,N_20776,N_20895);
or U21120 (N_21120,N_20876,N_20802);
xnor U21121 (N_21121,N_20865,N_20926);
or U21122 (N_21122,N_20889,N_20836);
nor U21123 (N_21123,N_20787,N_20945);
and U21124 (N_21124,N_20766,N_20844);
xor U21125 (N_21125,N_20900,N_20805);
or U21126 (N_21126,N_20954,N_20846);
and U21127 (N_21127,N_20897,N_20911);
and U21128 (N_21128,N_20903,N_20892);
or U21129 (N_21129,N_20787,N_20907);
or U21130 (N_21130,N_20991,N_20951);
and U21131 (N_21131,N_20965,N_20904);
nand U21132 (N_21132,N_20914,N_20791);
or U21133 (N_21133,N_20751,N_20986);
nand U21134 (N_21134,N_20867,N_20972);
nand U21135 (N_21135,N_20804,N_20820);
or U21136 (N_21136,N_20960,N_20804);
or U21137 (N_21137,N_20983,N_20996);
and U21138 (N_21138,N_20843,N_20812);
nor U21139 (N_21139,N_20911,N_20877);
nor U21140 (N_21140,N_20974,N_20840);
xor U21141 (N_21141,N_20850,N_20785);
nor U21142 (N_21142,N_20829,N_20954);
and U21143 (N_21143,N_20933,N_20918);
or U21144 (N_21144,N_20899,N_20945);
or U21145 (N_21145,N_20798,N_20889);
nand U21146 (N_21146,N_20921,N_20877);
xnor U21147 (N_21147,N_20764,N_20889);
nor U21148 (N_21148,N_20827,N_20931);
nand U21149 (N_21149,N_20881,N_20811);
or U21150 (N_21150,N_20863,N_20971);
or U21151 (N_21151,N_20882,N_20851);
or U21152 (N_21152,N_20750,N_20751);
nand U21153 (N_21153,N_20973,N_20980);
nor U21154 (N_21154,N_20894,N_20760);
xor U21155 (N_21155,N_20955,N_20816);
nor U21156 (N_21156,N_20797,N_20853);
or U21157 (N_21157,N_20871,N_20884);
or U21158 (N_21158,N_20800,N_20880);
nand U21159 (N_21159,N_20770,N_20976);
nor U21160 (N_21160,N_20855,N_20956);
and U21161 (N_21161,N_20789,N_20860);
nor U21162 (N_21162,N_20953,N_20857);
nand U21163 (N_21163,N_20830,N_20946);
xor U21164 (N_21164,N_20899,N_20970);
xor U21165 (N_21165,N_20938,N_20777);
xor U21166 (N_21166,N_20897,N_20905);
and U21167 (N_21167,N_20964,N_20800);
and U21168 (N_21168,N_20954,N_20953);
nand U21169 (N_21169,N_20985,N_20944);
and U21170 (N_21170,N_20956,N_20972);
or U21171 (N_21171,N_20754,N_20893);
or U21172 (N_21172,N_20916,N_20996);
nand U21173 (N_21173,N_20792,N_20953);
and U21174 (N_21174,N_20959,N_20999);
or U21175 (N_21175,N_20815,N_20819);
xor U21176 (N_21176,N_20855,N_20928);
nand U21177 (N_21177,N_20781,N_20995);
xnor U21178 (N_21178,N_20852,N_20842);
or U21179 (N_21179,N_20869,N_20764);
and U21180 (N_21180,N_20996,N_20795);
nand U21181 (N_21181,N_20757,N_20860);
or U21182 (N_21182,N_20894,N_20809);
or U21183 (N_21183,N_20821,N_20847);
or U21184 (N_21184,N_20798,N_20947);
nand U21185 (N_21185,N_20891,N_20826);
nand U21186 (N_21186,N_20760,N_20978);
nor U21187 (N_21187,N_20989,N_20939);
or U21188 (N_21188,N_20899,N_20940);
xnor U21189 (N_21189,N_20943,N_20835);
nor U21190 (N_21190,N_20778,N_20791);
nand U21191 (N_21191,N_20776,N_20919);
xnor U21192 (N_21192,N_20944,N_20878);
and U21193 (N_21193,N_20924,N_20819);
nor U21194 (N_21194,N_20976,N_20821);
nor U21195 (N_21195,N_20752,N_20951);
nand U21196 (N_21196,N_20811,N_20929);
nor U21197 (N_21197,N_20927,N_20909);
and U21198 (N_21198,N_20755,N_20965);
xnor U21199 (N_21199,N_20775,N_20816);
nand U21200 (N_21200,N_20953,N_20805);
or U21201 (N_21201,N_20792,N_20873);
or U21202 (N_21202,N_20964,N_20919);
and U21203 (N_21203,N_20859,N_20840);
and U21204 (N_21204,N_20780,N_20803);
nor U21205 (N_21205,N_20795,N_20802);
xor U21206 (N_21206,N_20833,N_20856);
xnor U21207 (N_21207,N_20848,N_20949);
or U21208 (N_21208,N_20786,N_20967);
xor U21209 (N_21209,N_20844,N_20795);
xor U21210 (N_21210,N_20995,N_20816);
or U21211 (N_21211,N_20948,N_20999);
or U21212 (N_21212,N_20804,N_20798);
nor U21213 (N_21213,N_20977,N_20909);
nor U21214 (N_21214,N_20908,N_20824);
or U21215 (N_21215,N_20759,N_20868);
xor U21216 (N_21216,N_20809,N_20976);
nor U21217 (N_21217,N_20937,N_20932);
and U21218 (N_21218,N_20850,N_20806);
nor U21219 (N_21219,N_20937,N_20848);
and U21220 (N_21220,N_20918,N_20785);
xor U21221 (N_21221,N_20775,N_20865);
xor U21222 (N_21222,N_20993,N_20863);
nor U21223 (N_21223,N_20878,N_20852);
xor U21224 (N_21224,N_20825,N_20987);
nor U21225 (N_21225,N_20987,N_20764);
xor U21226 (N_21226,N_20792,N_20991);
nand U21227 (N_21227,N_20796,N_20764);
or U21228 (N_21228,N_20991,N_20940);
xor U21229 (N_21229,N_20889,N_20920);
or U21230 (N_21230,N_20829,N_20955);
xnor U21231 (N_21231,N_20812,N_20984);
nor U21232 (N_21232,N_20755,N_20806);
nand U21233 (N_21233,N_20831,N_20942);
xor U21234 (N_21234,N_20948,N_20786);
nor U21235 (N_21235,N_20979,N_20935);
nand U21236 (N_21236,N_20856,N_20837);
or U21237 (N_21237,N_20937,N_20874);
or U21238 (N_21238,N_20866,N_20909);
nand U21239 (N_21239,N_20907,N_20949);
nand U21240 (N_21240,N_20931,N_20844);
nand U21241 (N_21241,N_20801,N_20910);
and U21242 (N_21242,N_20877,N_20958);
xnor U21243 (N_21243,N_20822,N_20864);
nor U21244 (N_21244,N_20851,N_20878);
or U21245 (N_21245,N_20981,N_20969);
and U21246 (N_21246,N_20889,N_20835);
xor U21247 (N_21247,N_20887,N_20975);
xor U21248 (N_21248,N_20881,N_20985);
xor U21249 (N_21249,N_20767,N_20991);
nand U21250 (N_21250,N_21032,N_21225);
nand U21251 (N_21251,N_21203,N_21097);
nand U21252 (N_21252,N_21040,N_21174);
and U21253 (N_21253,N_21004,N_21237);
and U21254 (N_21254,N_21012,N_21227);
xnor U21255 (N_21255,N_21199,N_21109);
xor U21256 (N_21256,N_21100,N_21164);
xor U21257 (N_21257,N_21131,N_21211);
xor U21258 (N_21258,N_21246,N_21188);
and U21259 (N_21259,N_21242,N_21221);
and U21260 (N_21260,N_21185,N_21000);
nor U21261 (N_21261,N_21103,N_21244);
xor U21262 (N_21262,N_21011,N_21057);
nand U21263 (N_21263,N_21022,N_21158);
and U21264 (N_21264,N_21133,N_21072);
nor U21265 (N_21265,N_21029,N_21023);
or U21266 (N_21266,N_21106,N_21087);
nor U21267 (N_21267,N_21105,N_21045);
nand U21268 (N_21268,N_21066,N_21206);
nand U21269 (N_21269,N_21202,N_21092);
xnor U21270 (N_21270,N_21141,N_21075);
xor U21271 (N_21271,N_21041,N_21183);
nand U21272 (N_21272,N_21049,N_21006);
nor U21273 (N_21273,N_21030,N_21217);
and U21274 (N_21274,N_21198,N_21150);
and U21275 (N_21275,N_21193,N_21140);
xnor U21276 (N_21276,N_21060,N_21191);
nor U21277 (N_21277,N_21025,N_21216);
and U21278 (N_21278,N_21107,N_21014);
nand U21279 (N_21279,N_21001,N_21058);
and U21280 (N_21280,N_21116,N_21208);
nand U21281 (N_21281,N_21228,N_21080);
xor U21282 (N_21282,N_21205,N_21148);
and U21283 (N_21283,N_21130,N_21160);
or U21284 (N_21284,N_21162,N_21010);
and U21285 (N_21285,N_21156,N_21241);
or U21286 (N_21286,N_21082,N_21240);
nor U21287 (N_21287,N_21120,N_21063);
or U21288 (N_21288,N_21077,N_21181);
xor U21289 (N_21289,N_21102,N_21219);
or U21290 (N_21290,N_21003,N_21115);
xor U21291 (N_21291,N_21220,N_21054);
and U21292 (N_21292,N_21009,N_21074);
and U21293 (N_21293,N_21236,N_21079);
and U21294 (N_21294,N_21214,N_21136);
nor U21295 (N_21295,N_21125,N_21039);
and U21296 (N_21296,N_21096,N_21065);
and U21297 (N_21297,N_21145,N_21171);
or U21298 (N_21298,N_21226,N_21161);
or U21299 (N_21299,N_21071,N_21051);
nand U21300 (N_21300,N_21117,N_21044);
nand U21301 (N_21301,N_21104,N_21248);
xor U21302 (N_21302,N_21197,N_21149);
nor U21303 (N_21303,N_21035,N_21114);
xnor U21304 (N_21304,N_21186,N_21016);
and U21305 (N_21305,N_21033,N_21031);
nor U21306 (N_21306,N_21056,N_21143);
xnor U21307 (N_21307,N_21182,N_21207);
or U21308 (N_21308,N_21084,N_21194);
xnor U21309 (N_21309,N_21245,N_21215);
and U21310 (N_21310,N_21247,N_21201);
or U21311 (N_21311,N_21052,N_21089);
and U21312 (N_21312,N_21135,N_21078);
and U21313 (N_21313,N_21166,N_21076);
and U21314 (N_21314,N_21128,N_21243);
and U21315 (N_21315,N_21083,N_21026);
xnor U21316 (N_21316,N_21134,N_21068);
xnor U21317 (N_21317,N_21213,N_21177);
and U21318 (N_21318,N_21222,N_21024);
xor U21319 (N_21319,N_21176,N_21231);
xnor U21320 (N_21320,N_21098,N_21218);
or U21321 (N_21321,N_21047,N_21094);
nor U21322 (N_21322,N_21192,N_21055);
and U21323 (N_21323,N_21053,N_21196);
nor U21324 (N_21324,N_21173,N_21007);
xnor U21325 (N_21325,N_21034,N_21157);
nor U21326 (N_21326,N_21099,N_21138);
and U21327 (N_21327,N_21209,N_21050);
xnor U21328 (N_21328,N_21005,N_21043);
xor U21329 (N_21329,N_21189,N_21200);
or U21330 (N_21330,N_21224,N_21059);
and U21331 (N_21331,N_21070,N_21190);
nor U21332 (N_21332,N_21064,N_21061);
and U21333 (N_21333,N_21165,N_21144);
and U21334 (N_21334,N_21085,N_21154);
nand U21335 (N_21335,N_21204,N_21038);
nor U21336 (N_21336,N_21081,N_21095);
nand U21337 (N_21337,N_21233,N_21238);
and U21338 (N_21338,N_21111,N_21123);
nor U21339 (N_21339,N_21110,N_21239);
nand U21340 (N_21340,N_21112,N_21013);
nand U21341 (N_21341,N_21008,N_21147);
nor U21342 (N_21342,N_21015,N_21142);
and U21343 (N_21343,N_21180,N_21178);
nand U21344 (N_21344,N_21137,N_21127);
and U21345 (N_21345,N_21170,N_21223);
nor U21346 (N_21346,N_21086,N_21113);
and U21347 (N_21347,N_21101,N_21046);
nand U21348 (N_21348,N_21187,N_21129);
or U21349 (N_21349,N_21119,N_21018);
nand U21350 (N_21350,N_21155,N_21124);
or U21351 (N_21351,N_21017,N_21027);
nand U21352 (N_21352,N_21163,N_21020);
and U21353 (N_21353,N_21172,N_21122);
nand U21354 (N_21354,N_21168,N_21184);
nor U21355 (N_21355,N_21159,N_21108);
xor U21356 (N_21356,N_21019,N_21229);
or U21357 (N_21357,N_21153,N_21152);
xor U21358 (N_21358,N_21179,N_21132);
xor U21359 (N_21359,N_21230,N_21036);
nand U21360 (N_21360,N_21037,N_21069);
nor U21361 (N_21361,N_21195,N_21169);
xnor U21362 (N_21362,N_21048,N_21028);
and U21363 (N_21363,N_21151,N_21210);
and U21364 (N_21364,N_21002,N_21088);
nand U21365 (N_21365,N_21118,N_21139);
xnor U21366 (N_21366,N_21232,N_21062);
xor U21367 (N_21367,N_21073,N_21167);
nand U21368 (N_21368,N_21021,N_21067);
xnor U21369 (N_21369,N_21146,N_21090);
xnor U21370 (N_21370,N_21212,N_21234);
or U21371 (N_21371,N_21126,N_21235);
nor U21372 (N_21372,N_21249,N_21091);
xnor U21373 (N_21373,N_21121,N_21093);
nor U21374 (N_21374,N_21042,N_21175);
or U21375 (N_21375,N_21149,N_21056);
xnor U21376 (N_21376,N_21152,N_21081);
xnor U21377 (N_21377,N_21085,N_21097);
xor U21378 (N_21378,N_21044,N_21229);
xnor U21379 (N_21379,N_21151,N_21120);
or U21380 (N_21380,N_21232,N_21149);
nor U21381 (N_21381,N_21121,N_21166);
xnor U21382 (N_21382,N_21143,N_21196);
and U21383 (N_21383,N_21172,N_21184);
and U21384 (N_21384,N_21206,N_21212);
nor U21385 (N_21385,N_21143,N_21194);
nor U21386 (N_21386,N_21120,N_21075);
xnor U21387 (N_21387,N_21061,N_21162);
xnor U21388 (N_21388,N_21056,N_21088);
nand U21389 (N_21389,N_21067,N_21000);
and U21390 (N_21390,N_21064,N_21164);
nor U21391 (N_21391,N_21038,N_21011);
and U21392 (N_21392,N_21231,N_21203);
nand U21393 (N_21393,N_21158,N_21208);
xor U21394 (N_21394,N_21003,N_21006);
and U21395 (N_21395,N_21132,N_21022);
xnor U21396 (N_21396,N_21222,N_21207);
or U21397 (N_21397,N_21140,N_21191);
and U21398 (N_21398,N_21104,N_21174);
xor U21399 (N_21399,N_21147,N_21213);
nor U21400 (N_21400,N_21222,N_21076);
and U21401 (N_21401,N_21117,N_21036);
and U21402 (N_21402,N_21037,N_21017);
and U21403 (N_21403,N_21198,N_21111);
xnor U21404 (N_21404,N_21041,N_21199);
and U21405 (N_21405,N_21057,N_21082);
nand U21406 (N_21406,N_21127,N_21085);
or U21407 (N_21407,N_21016,N_21226);
and U21408 (N_21408,N_21007,N_21120);
and U21409 (N_21409,N_21030,N_21087);
xor U21410 (N_21410,N_21113,N_21114);
nand U21411 (N_21411,N_21133,N_21040);
or U21412 (N_21412,N_21226,N_21192);
nor U21413 (N_21413,N_21203,N_21099);
and U21414 (N_21414,N_21247,N_21101);
and U21415 (N_21415,N_21041,N_21109);
or U21416 (N_21416,N_21174,N_21006);
and U21417 (N_21417,N_21010,N_21101);
or U21418 (N_21418,N_21238,N_21188);
nand U21419 (N_21419,N_21217,N_21129);
and U21420 (N_21420,N_21039,N_21206);
xor U21421 (N_21421,N_21243,N_21006);
nor U21422 (N_21422,N_21231,N_21156);
nor U21423 (N_21423,N_21157,N_21057);
xor U21424 (N_21424,N_21227,N_21078);
and U21425 (N_21425,N_21065,N_21237);
xor U21426 (N_21426,N_21052,N_21116);
nor U21427 (N_21427,N_21063,N_21065);
nand U21428 (N_21428,N_21021,N_21242);
nor U21429 (N_21429,N_21210,N_21176);
nand U21430 (N_21430,N_21233,N_21099);
or U21431 (N_21431,N_21203,N_21201);
or U21432 (N_21432,N_21246,N_21202);
xor U21433 (N_21433,N_21048,N_21235);
and U21434 (N_21434,N_21201,N_21177);
and U21435 (N_21435,N_21070,N_21165);
or U21436 (N_21436,N_21073,N_21225);
xnor U21437 (N_21437,N_21088,N_21068);
and U21438 (N_21438,N_21112,N_21179);
or U21439 (N_21439,N_21117,N_21094);
nor U21440 (N_21440,N_21200,N_21079);
nand U21441 (N_21441,N_21246,N_21128);
and U21442 (N_21442,N_21129,N_21182);
and U21443 (N_21443,N_21188,N_21070);
xor U21444 (N_21444,N_21134,N_21032);
and U21445 (N_21445,N_21028,N_21099);
nand U21446 (N_21446,N_21132,N_21016);
nand U21447 (N_21447,N_21051,N_21085);
nand U21448 (N_21448,N_21090,N_21029);
and U21449 (N_21449,N_21058,N_21200);
and U21450 (N_21450,N_21014,N_21030);
and U21451 (N_21451,N_21158,N_21143);
xor U21452 (N_21452,N_21061,N_21200);
and U21453 (N_21453,N_21021,N_21243);
or U21454 (N_21454,N_21188,N_21057);
and U21455 (N_21455,N_21239,N_21218);
or U21456 (N_21456,N_21198,N_21137);
or U21457 (N_21457,N_21241,N_21122);
xnor U21458 (N_21458,N_21141,N_21047);
nand U21459 (N_21459,N_21245,N_21230);
xnor U21460 (N_21460,N_21080,N_21179);
nand U21461 (N_21461,N_21244,N_21025);
nand U21462 (N_21462,N_21202,N_21125);
nand U21463 (N_21463,N_21051,N_21084);
nor U21464 (N_21464,N_21099,N_21022);
nand U21465 (N_21465,N_21064,N_21034);
and U21466 (N_21466,N_21072,N_21216);
xor U21467 (N_21467,N_21230,N_21097);
nor U21468 (N_21468,N_21239,N_21174);
xor U21469 (N_21469,N_21017,N_21009);
nand U21470 (N_21470,N_21172,N_21075);
and U21471 (N_21471,N_21017,N_21070);
xnor U21472 (N_21472,N_21125,N_21083);
xnor U21473 (N_21473,N_21121,N_21125);
or U21474 (N_21474,N_21099,N_21091);
xor U21475 (N_21475,N_21029,N_21219);
nand U21476 (N_21476,N_21072,N_21179);
or U21477 (N_21477,N_21046,N_21208);
nand U21478 (N_21478,N_21170,N_21221);
or U21479 (N_21479,N_21193,N_21002);
nand U21480 (N_21480,N_21161,N_21142);
and U21481 (N_21481,N_21209,N_21196);
or U21482 (N_21482,N_21214,N_21149);
and U21483 (N_21483,N_21219,N_21160);
nor U21484 (N_21484,N_21088,N_21006);
nand U21485 (N_21485,N_21041,N_21127);
nor U21486 (N_21486,N_21078,N_21048);
or U21487 (N_21487,N_21027,N_21014);
xnor U21488 (N_21488,N_21230,N_21118);
nor U21489 (N_21489,N_21089,N_21124);
and U21490 (N_21490,N_21119,N_21044);
nand U21491 (N_21491,N_21187,N_21095);
xor U21492 (N_21492,N_21121,N_21081);
xor U21493 (N_21493,N_21063,N_21035);
or U21494 (N_21494,N_21127,N_21007);
or U21495 (N_21495,N_21185,N_21240);
xor U21496 (N_21496,N_21230,N_21238);
xor U21497 (N_21497,N_21010,N_21065);
xor U21498 (N_21498,N_21202,N_21240);
nor U21499 (N_21499,N_21167,N_21081);
or U21500 (N_21500,N_21303,N_21471);
or U21501 (N_21501,N_21262,N_21289);
or U21502 (N_21502,N_21392,N_21481);
nor U21503 (N_21503,N_21445,N_21497);
xor U21504 (N_21504,N_21261,N_21333);
nand U21505 (N_21505,N_21381,N_21374);
nand U21506 (N_21506,N_21311,N_21326);
and U21507 (N_21507,N_21436,N_21335);
nand U21508 (N_21508,N_21274,N_21364);
nor U21509 (N_21509,N_21295,N_21258);
nor U21510 (N_21510,N_21293,N_21328);
nor U21511 (N_21511,N_21473,N_21412);
nor U21512 (N_21512,N_21345,N_21332);
xor U21513 (N_21513,N_21380,N_21477);
xnor U21514 (N_21514,N_21443,N_21496);
nand U21515 (N_21515,N_21306,N_21438);
nand U21516 (N_21516,N_21250,N_21309);
nor U21517 (N_21517,N_21448,N_21498);
and U21518 (N_21518,N_21367,N_21395);
or U21519 (N_21519,N_21350,N_21384);
and U21520 (N_21520,N_21279,N_21465);
nor U21521 (N_21521,N_21493,N_21483);
nand U21522 (N_21522,N_21322,N_21355);
xnor U21523 (N_21523,N_21442,N_21468);
or U21524 (N_21524,N_21296,N_21317);
xor U21525 (N_21525,N_21269,N_21329);
nor U21526 (N_21526,N_21416,N_21290);
xnor U21527 (N_21527,N_21349,N_21461);
xnor U21528 (N_21528,N_21342,N_21464);
nor U21529 (N_21529,N_21255,N_21385);
nor U21530 (N_21530,N_21469,N_21361);
nor U21531 (N_21531,N_21387,N_21418);
nand U21532 (N_21532,N_21432,N_21359);
xor U21533 (N_21533,N_21302,N_21479);
nor U21534 (N_21534,N_21456,N_21450);
or U21535 (N_21535,N_21383,N_21273);
xor U21536 (N_21536,N_21382,N_21478);
or U21537 (N_21537,N_21489,N_21260);
xnor U21538 (N_21538,N_21439,N_21449);
and U21539 (N_21539,N_21453,N_21298);
xor U21540 (N_21540,N_21429,N_21467);
xor U21541 (N_21541,N_21372,N_21271);
xor U21542 (N_21542,N_21344,N_21406);
xor U21543 (N_21543,N_21491,N_21299);
nor U21544 (N_21544,N_21370,N_21324);
nor U21545 (N_21545,N_21424,N_21422);
or U21546 (N_21546,N_21320,N_21462);
and U21547 (N_21547,N_21256,N_21259);
nor U21548 (N_21548,N_21430,N_21437);
and U21549 (N_21549,N_21401,N_21282);
xnor U21550 (N_21550,N_21321,N_21356);
nor U21551 (N_21551,N_21458,N_21411);
nand U21552 (N_21552,N_21375,N_21341);
or U21553 (N_21553,N_21492,N_21390);
nor U21554 (N_21554,N_21495,N_21407);
nand U21555 (N_21555,N_21315,N_21447);
and U21556 (N_21556,N_21423,N_21485);
or U21557 (N_21557,N_21339,N_21494);
nand U21558 (N_21558,N_21425,N_21360);
xor U21559 (N_21559,N_21454,N_21313);
nor U21560 (N_21560,N_21441,N_21314);
xnor U21561 (N_21561,N_21253,N_21263);
and U21562 (N_21562,N_21421,N_21368);
nor U21563 (N_21563,N_21354,N_21325);
nand U21564 (N_21564,N_21294,N_21460);
and U21565 (N_21565,N_21484,N_21331);
and U21566 (N_21566,N_21480,N_21376);
nor U21567 (N_21567,N_21337,N_21466);
xor U21568 (N_21568,N_21257,N_21431);
or U21569 (N_21569,N_21283,N_21347);
nor U21570 (N_21570,N_21276,N_21488);
and U21571 (N_21571,N_21292,N_21459);
nor U21572 (N_21572,N_21297,N_21300);
and U21573 (N_21573,N_21472,N_21265);
nor U21574 (N_21574,N_21386,N_21451);
nand U21575 (N_21575,N_21365,N_21266);
nor U21576 (N_21576,N_21379,N_21373);
nand U21577 (N_21577,N_21318,N_21394);
xnor U21578 (N_21578,N_21270,N_21340);
nor U21579 (N_21579,N_21363,N_21252);
and U21580 (N_21580,N_21362,N_21420);
xor U21581 (N_21581,N_21413,N_21316);
nor U21582 (N_21582,N_21474,N_21277);
or U21583 (N_21583,N_21452,N_21404);
nand U21584 (N_21584,N_21482,N_21334);
and U21585 (N_21585,N_21251,N_21399);
or U21586 (N_21586,N_21264,N_21357);
and U21587 (N_21587,N_21323,N_21396);
or U21588 (N_21588,N_21267,N_21440);
and U21589 (N_21589,N_21393,N_21338);
nor U21590 (N_21590,N_21304,N_21278);
or U21591 (N_21591,N_21410,N_21470);
and U21592 (N_21592,N_21408,N_21398);
nand U21593 (N_21593,N_21308,N_21402);
nand U21594 (N_21594,N_21352,N_21377);
xnor U21595 (N_21595,N_21280,N_21463);
xor U21596 (N_21596,N_21371,N_21284);
xor U21597 (N_21597,N_21388,N_21476);
nand U21598 (N_21598,N_21435,N_21327);
nor U21599 (N_21599,N_21285,N_21417);
nor U21600 (N_21600,N_21490,N_21455);
nand U21601 (N_21601,N_21336,N_21409);
nand U21602 (N_21602,N_21369,N_21389);
xor U21603 (N_21603,N_21428,N_21330);
xor U21604 (N_21604,N_21291,N_21310);
or U21605 (N_21605,N_21486,N_21288);
or U21606 (N_21606,N_21301,N_21378);
nor U21607 (N_21607,N_21281,N_21287);
or U21608 (N_21608,N_21254,N_21348);
nand U21609 (N_21609,N_21346,N_21343);
nand U21610 (N_21610,N_21434,N_21415);
nor U21611 (N_21611,N_21307,N_21444);
and U21612 (N_21612,N_21405,N_21457);
or U21613 (N_21613,N_21286,N_21433);
and U21614 (N_21614,N_21475,N_21426);
and U21615 (N_21615,N_21305,N_21268);
xnor U21616 (N_21616,N_21351,N_21275);
nor U21617 (N_21617,N_21353,N_21319);
nor U21618 (N_21618,N_21414,N_21487);
nor U21619 (N_21619,N_21400,N_21366);
nor U21620 (N_21620,N_21272,N_21427);
nand U21621 (N_21621,N_21419,N_21397);
or U21622 (N_21622,N_21358,N_21312);
and U21623 (N_21623,N_21446,N_21391);
nand U21624 (N_21624,N_21499,N_21403);
and U21625 (N_21625,N_21377,N_21486);
nor U21626 (N_21626,N_21269,N_21283);
or U21627 (N_21627,N_21268,N_21267);
xnor U21628 (N_21628,N_21353,N_21376);
and U21629 (N_21629,N_21340,N_21342);
or U21630 (N_21630,N_21327,N_21324);
or U21631 (N_21631,N_21295,N_21344);
nor U21632 (N_21632,N_21375,N_21371);
nand U21633 (N_21633,N_21269,N_21395);
or U21634 (N_21634,N_21402,N_21386);
nor U21635 (N_21635,N_21306,N_21358);
nor U21636 (N_21636,N_21353,N_21324);
nor U21637 (N_21637,N_21452,N_21264);
nor U21638 (N_21638,N_21472,N_21383);
and U21639 (N_21639,N_21270,N_21496);
and U21640 (N_21640,N_21411,N_21253);
nor U21641 (N_21641,N_21430,N_21369);
xnor U21642 (N_21642,N_21265,N_21359);
nand U21643 (N_21643,N_21310,N_21394);
nor U21644 (N_21644,N_21332,N_21447);
or U21645 (N_21645,N_21412,N_21324);
nor U21646 (N_21646,N_21372,N_21401);
xnor U21647 (N_21647,N_21328,N_21416);
nand U21648 (N_21648,N_21278,N_21317);
or U21649 (N_21649,N_21373,N_21492);
and U21650 (N_21650,N_21274,N_21333);
xor U21651 (N_21651,N_21416,N_21364);
nor U21652 (N_21652,N_21360,N_21391);
and U21653 (N_21653,N_21250,N_21359);
nand U21654 (N_21654,N_21316,N_21469);
nand U21655 (N_21655,N_21294,N_21281);
nor U21656 (N_21656,N_21311,N_21300);
and U21657 (N_21657,N_21386,N_21313);
or U21658 (N_21658,N_21395,N_21279);
or U21659 (N_21659,N_21312,N_21320);
or U21660 (N_21660,N_21434,N_21289);
or U21661 (N_21661,N_21333,N_21285);
nor U21662 (N_21662,N_21478,N_21450);
xnor U21663 (N_21663,N_21317,N_21497);
xor U21664 (N_21664,N_21404,N_21330);
nor U21665 (N_21665,N_21315,N_21294);
nor U21666 (N_21666,N_21317,N_21287);
nand U21667 (N_21667,N_21270,N_21398);
xnor U21668 (N_21668,N_21465,N_21475);
nand U21669 (N_21669,N_21391,N_21366);
nand U21670 (N_21670,N_21343,N_21424);
xnor U21671 (N_21671,N_21336,N_21291);
nor U21672 (N_21672,N_21333,N_21489);
xor U21673 (N_21673,N_21398,N_21314);
nor U21674 (N_21674,N_21325,N_21478);
and U21675 (N_21675,N_21281,N_21338);
nand U21676 (N_21676,N_21291,N_21366);
nand U21677 (N_21677,N_21437,N_21326);
nor U21678 (N_21678,N_21437,N_21440);
nand U21679 (N_21679,N_21483,N_21371);
nand U21680 (N_21680,N_21467,N_21299);
nor U21681 (N_21681,N_21335,N_21298);
nor U21682 (N_21682,N_21254,N_21363);
xor U21683 (N_21683,N_21324,N_21278);
nand U21684 (N_21684,N_21332,N_21251);
nand U21685 (N_21685,N_21326,N_21338);
nand U21686 (N_21686,N_21422,N_21347);
and U21687 (N_21687,N_21346,N_21292);
xnor U21688 (N_21688,N_21303,N_21475);
xnor U21689 (N_21689,N_21414,N_21323);
or U21690 (N_21690,N_21404,N_21433);
xor U21691 (N_21691,N_21316,N_21337);
and U21692 (N_21692,N_21309,N_21395);
and U21693 (N_21693,N_21495,N_21422);
nor U21694 (N_21694,N_21388,N_21316);
nor U21695 (N_21695,N_21341,N_21458);
xor U21696 (N_21696,N_21478,N_21280);
xnor U21697 (N_21697,N_21454,N_21445);
xor U21698 (N_21698,N_21467,N_21325);
and U21699 (N_21699,N_21366,N_21345);
xor U21700 (N_21700,N_21273,N_21412);
nand U21701 (N_21701,N_21480,N_21423);
or U21702 (N_21702,N_21373,N_21282);
nand U21703 (N_21703,N_21350,N_21422);
or U21704 (N_21704,N_21309,N_21319);
nor U21705 (N_21705,N_21432,N_21467);
nand U21706 (N_21706,N_21431,N_21428);
or U21707 (N_21707,N_21451,N_21394);
or U21708 (N_21708,N_21294,N_21347);
and U21709 (N_21709,N_21357,N_21339);
and U21710 (N_21710,N_21386,N_21317);
nor U21711 (N_21711,N_21359,N_21264);
nand U21712 (N_21712,N_21256,N_21369);
nand U21713 (N_21713,N_21377,N_21299);
nor U21714 (N_21714,N_21363,N_21373);
nor U21715 (N_21715,N_21308,N_21345);
nand U21716 (N_21716,N_21337,N_21291);
or U21717 (N_21717,N_21339,N_21311);
or U21718 (N_21718,N_21400,N_21488);
xor U21719 (N_21719,N_21339,N_21393);
and U21720 (N_21720,N_21487,N_21451);
nor U21721 (N_21721,N_21263,N_21467);
nand U21722 (N_21722,N_21258,N_21497);
or U21723 (N_21723,N_21287,N_21344);
and U21724 (N_21724,N_21268,N_21320);
xnor U21725 (N_21725,N_21424,N_21383);
and U21726 (N_21726,N_21254,N_21428);
nand U21727 (N_21727,N_21318,N_21303);
nand U21728 (N_21728,N_21305,N_21457);
or U21729 (N_21729,N_21419,N_21291);
and U21730 (N_21730,N_21285,N_21343);
xnor U21731 (N_21731,N_21429,N_21408);
nand U21732 (N_21732,N_21418,N_21465);
nand U21733 (N_21733,N_21462,N_21346);
xor U21734 (N_21734,N_21496,N_21456);
nor U21735 (N_21735,N_21403,N_21420);
or U21736 (N_21736,N_21331,N_21278);
or U21737 (N_21737,N_21285,N_21300);
or U21738 (N_21738,N_21368,N_21467);
or U21739 (N_21739,N_21342,N_21286);
and U21740 (N_21740,N_21365,N_21420);
nand U21741 (N_21741,N_21480,N_21476);
or U21742 (N_21742,N_21302,N_21350);
or U21743 (N_21743,N_21497,N_21254);
nand U21744 (N_21744,N_21462,N_21423);
or U21745 (N_21745,N_21291,N_21472);
nor U21746 (N_21746,N_21420,N_21458);
xor U21747 (N_21747,N_21442,N_21466);
or U21748 (N_21748,N_21306,N_21434);
and U21749 (N_21749,N_21256,N_21453);
nor U21750 (N_21750,N_21535,N_21509);
or U21751 (N_21751,N_21665,N_21693);
xor U21752 (N_21752,N_21689,N_21570);
xor U21753 (N_21753,N_21623,N_21530);
xor U21754 (N_21754,N_21562,N_21555);
and U21755 (N_21755,N_21549,N_21632);
or U21756 (N_21756,N_21634,N_21548);
nor U21757 (N_21757,N_21646,N_21576);
or U21758 (N_21758,N_21597,N_21720);
nand U21759 (N_21759,N_21622,N_21726);
nor U21760 (N_21760,N_21502,N_21711);
nand U21761 (N_21761,N_21559,N_21742);
xnor U21762 (N_21762,N_21567,N_21675);
xnor U21763 (N_21763,N_21514,N_21749);
nand U21764 (N_21764,N_21560,N_21589);
and U21765 (N_21765,N_21704,N_21640);
nand U21766 (N_21766,N_21543,N_21635);
nor U21767 (N_21767,N_21531,N_21702);
xnor U21768 (N_21768,N_21506,N_21546);
and U21769 (N_21769,N_21608,N_21563);
nor U21770 (N_21770,N_21600,N_21568);
or U21771 (N_21771,N_21554,N_21593);
nor U21772 (N_21772,N_21669,N_21721);
nand U21773 (N_21773,N_21737,N_21673);
nor U21774 (N_21774,N_21627,N_21719);
nor U21775 (N_21775,N_21588,N_21525);
nand U21776 (N_21776,N_21660,N_21591);
nor U21777 (N_21777,N_21683,N_21537);
nand U21778 (N_21778,N_21633,N_21670);
nand U21779 (N_21779,N_21504,N_21672);
nor U21780 (N_21780,N_21644,N_21636);
nand U21781 (N_21781,N_21577,N_21609);
nand U21782 (N_21782,N_21618,N_21688);
or U21783 (N_21783,N_21662,N_21557);
and U21784 (N_21784,N_21735,N_21575);
and U21785 (N_21785,N_21641,N_21579);
nor U21786 (N_21786,N_21652,N_21615);
or U21787 (N_21787,N_21629,N_21612);
and U21788 (N_21788,N_21518,N_21658);
and U21789 (N_21789,N_21678,N_21611);
nand U21790 (N_21790,N_21607,N_21651);
and U21791 (N_21791,N_21654,N_21653);
nand U21792 (N_21792,N_21690,N_21534);
and U21793 (N_21793,N_21691,N_21699);
nor U21794 (N_21794,N_21601,N_21727);
or U21795 (N_21795,N_21558,N_21692);
nor U21796 (N_21796,N_21639,N_21728);
and U21797 (N_21797,N_21657,N_21697);
nand U21798 (N_21798,N_21604,N_21648);
nor U21799 (N_21799,N_21547,N_21508);
or U21800 (N_21800,N_21666,N_21712);
and U21801 (N_21801,N_21717,N_21606);
xor U21802 (N_21802,N_21694,N_21521);
nand U21803 (N_21803,N_21541,N_21626);
xnor U21804 (N_21804,N_21650,N_21741);
nor U21805 (N_21805,N_21630,N_21723);
and U21806 (N_21806,N_21590,N_21663);
nor U21807 (N_21807,N_21625,N_21680);
xnor U21808 (N_21808,N_21709,N_21732);
nor U21809 (N_21809,N_21659,N_21681);
and U21810 (N_21810,N_21520,N_21532);
and U21811 (N_21811,N_21746,N_21605);
or U21812 (N_21812,N_21628,N_21552);
xor U21813 (N_21813,N_21507,N_21545);
or U21814 (N_21814,N_21512,N_21573);
or U21815 (N_21815,N_21667,N_21501);
nor U21816 (N_21816,N_21528,N_21592);
and U21817 (N_21817,N_21561,N_21649);
and U21818 (N_21818,N_21716,N_21700);
or U21819 (N_21819,N_21613,N_21715);
xor U21820 (N_21820,N_21682,N_21685);
nand U21821 (N_21821,N_21510,N_21610);
nand U21822 (N_21822,N_21731,N_21655);
nor U21823 (N_21823,N_21513,N_21707);
nor U21824 (N_21824,N_21744,N_21643);
and U21825 (N_21825,N_21676,N_21586);
and U21826 (N_21826,N_21522,N_21603);
and U21827 (N_21827,N_21718,N_21587);
nand U21828 (N_21828,N_21527,N_21544);
xor U21829 (N_21829,N_21743,N_21684);
nor U21830 (N_21830,N_21511,N_21701);
nand U21831 (N_21831,N_21747,N_21677);
nand U21832 (N_21832,N_21631,N_21536);
and U21833 (N_21833,N_21595,N_21569);
and U21834 (N_21834,N_21505,N_21526);
nor U21835 (N_21835,N_21637,N_21578);
or U21836 (N_21836,N_21714,N_21582);
and U21837 (N_21837,N_21733,N_21722);
or U21838 (N_21838,N_21687,N_21551);
nand U21839 (N_21839,N_21594,N_21713);
and U21840 (N_21840,N_21674,N_21724);
nand U21841 (N_21841,N_21736,N_21671);
nor U21842 (N_21842,N_21710,N_21542);
nand U21843 (N_21843,N_21642,N_21571);
nand U21844 (N_21844,N_21556,N_21647);
nand U21845 (N_21845,N_21624,N_21538);
nand U21846 (N_21846,N_21523,N_21583);
nand U21847 (N_21847,N_21550,N_21698);
xnor U21848 (N_21848,N_21503,N_21638);
nand U21849 (N_21849,N_21706,N_21739);
nand U21850 (N_21850,N_21529,N_21730);
or U21851 (N_21851,N_21585,N_21517);
nor U21852 (N_21852,N_21679,N_21664);
and U21853 (N_21853,N_21616,N_21598);
nor U21854 (N_21854,N_21519,N_21614);
nand U21855 (N_21855,N_21729,N_21533);
or U21856 (N_21856,N_21708,N_21740);
nand U21857 (N_21857,N_21553,N_21617);
or U21858 (N_21858,N_21734,N_21572);
nor U21859 (N_21859,N_21621,N_21599);
xor U21860 (N_21860,N_21738,N_21580);
and U21861 (N_21861,N_21745,N_21748);
or U21862 (N_21862,N_21565,N_21620);
nor U21863 (N_21863,N_21500,N_21703);
xor U21864 (N_21864,N_21661,N_21540);
nand U21865 (N_21865,N_21515,N_21695);
or U21866 (N_21866,N_21596,N_21539);
nand U21867 (N_21867,N_21584,N_21564);
xnor U21868 (N_21868,N_21705,N_21602);
xor U21869 (N_21869,N_21516,N_21725);
nand U21870 (N_21870,N_21645,N_21696);
or U21871 (N_21871,N_21686,N_21581);
xnor U21872 (N_21872,N_21619,N_21524);
xor U21873 (N_21873,N_21566,N_21668);
and U21874 (N_21874,N_21656,N_21574);
nand U21875 (N_21875,N_21615,N_21694);
nand U21876 (N_21876,N_21568,N_21618);
nand U21877 (N_21877,N_21658,N_21641);
nor U21878 (N_21878,N_21552,N_21692);
xor U21879 (N_21879,N_21727,N_21587);
and U21880 (N_21880,N_21546,N_21662);
or U21881 (N_21881,N_21686,N_21625);
or U21882 (N_21882,N_21550,N_21521);
nand U21883 (N_21883,N_21659,N_21620);
or U21884 (N_21884,N_21685,N_21734);
nand U21885 (N_21885,N_21522,N_21661);
xnor U21886 (N_21886,N_21662,N_21623);
or U21887 (N_21887,N_21511,N_21525);
and U21888 (N_21888,N_21703,N_21737);
or U21889 (N_21889,N_21530,N_21691);
nand U21890 (N_21890,N_21588,N_21643);
or U21891 (N_21891,N_21518,N_21707);
and U21892 (N_21892,N_21699,N_21666);
or U21893 (N_21893,N_21690,N_21500);
or U21894 (N_21894,N_21736,N_21705);
and U21895 (N_21895,N_21506,N_21735);
or U21896 (N_21896,N_21684,N_21731);
or U21897 (N_21897,N_21537,N_21568);
nand U21898 (N_21898,N_21741,N_21700);
nand U21899 (N_21899,N_21612,N_21573);
nand U21900 (N_21900,N_21627,N_21717);
or U21901 (N_21901,N_21632,N_21708);
nand U21902 (N_21902,N_21561,N_21513);
xnor U21903 (N_21903,N_21556,N_21740);
nand U21904 (N_21904,N_21642,N_21545);
or U21905 (N_21905,N_21591,N_21622);
xor U21906 (N_21906,N_21503,N_21689);
nand U21907 (N_21907,N_21674,N_21663);
nor U21908 (N_21908,N_21536,N_21514);
nand U21909 (N_21909,N_21560,N_21627);
or U21910 (N_21910,N_21579,N_21723);
or U21911 (N_21911,N_21541,N_21603);
nand U21912 (N_21912,N_21684,N_21575);
nor U21913 (N_21913,N_21522,N_21672);
nor U21914 (N_21914,N_21535,N_21572);
or U21915 (N_21915,N_21549,N_21614);
nor U21916 (N_21916,N_21528,N_21654);
nand U21917 (N_21917,N_21707,N_21722);
or U21918 (N_21918,N_21643,N_21682);
and U21919 (N_21919,N_21695,N_21619);
nand U21920 (N_21920,N_21577,N_21675);
nand U21921 (N_21921,N_21632,N_21525);
and U21922 (N_21922,N_21501,N_21563);
nor U21923 (N_21923,N_21633,N_21641);
or U21924 (N_21924,N_21666,N_21648);
or U21925 (N_21925,N_21726,N_21586);
xnor U21926 (N_21926,N_21618,N_21500);
xnor U21927 (N_21927,N_21678,N_21543);
xnor U21928 (N_21928,N_21732,N_21509);
or U21929 (N_21929,N_21519,N_21661);
nand U21930 (N_21930,N_21578,N_21727);
nor U21931 (N_21931,N_21570,N_21652);
xnor U21932 (N_21932,N_21546,N_21639);
and U21933 (N_21933,N_21673,N_21616);
nor U21934 (N_21934,N_21704,N_21631);
or U21935 (N_21935,N_21531,N_21654);
nor U21936 (N_21936,N_21574,N_21515);
or U21937 (N_21937,N_21500,N_21506);
and U21938 (N_21938,N_21545,N_21724);
nand U21939 (N_21939,N_21630,N_21523);
and U21940 (N_21940,N_21660,N_21676);
nand U21941 (N_21941,N_21556,N_21503);
and U21942 (N_21942,N_21644,N_21564);
and U21943 (N_21943,N_21505,N_21660);
nand U21944 (N_21944,N_21746,N_21594);
or U21945 (N_21945,N_21627,N_21528);
xnor U21946 (N_21946,N_21582,N_21710);
xnor U21947 (N_21947,N_21509,N_21615);
xnor U21948 (N_21948,N_21552,N_21599);
nand U21949 (N_21949,N_21500,N_21567);
xnor U21950 (N_21950,N_21509,N_21687);
nor U21951 (N_21951,N_21700,N_21633);
and U21952 (N_21952,N_21712,N_21693);
or U21953 (N_21953,N_21591,N_21736);
xor U21954 (N_21954,N_21539,N_21621);
nand U21955 (N_21955,N_21625,N_21746);
nand U21956 (N_21956,N_21669,N_21506);
and U21957 (N_21957,N_21515,N_21617);
nor U21958 (N_21958,N_21543,N_21552);
or U21959 (N_21959,N_21617,N_21696);
xnor U21960 (N_21960,N_21594,N_21738);
xor U21961 (N_21961,N_21665,N_21530);
and U21962 (N_21962,N_21675,N_21625);
nor U21963 (N_21963,N_21665,N_21514);
nor U21964 (N_21964,N_21682,N_21621);
xnor U21965 (N_21965,N_21667,N_21635);
or U21966 (N_21966,N_21745,N_21701);
nor U21967 (N_21967,N_21742,N_21706);
nor U21968 (N_21968,N_21626,N_21651);
and U21969 (N_21969,N_21631,N_21706);
and U21970 (N_21970,N_21627,N_21584);
xor U21971 (N_21971,N_21653,N_21717);
nand U21972 (N_21972,N_21556,N_21730);
xor U21973 (N_21973,N_21735,N_21607);
or U21974 (N_21974,N_21534,N_21591);
or U21975 (N_21975,N_21624,N_21738);
nand U21976 (N_21976,N_21712,N_21740);
nor U21977 (N_21977,N_21717,N_21664);
or U21978 (N_21978,N_21673,N_21747);
xor U21979 (N_21979,N_21733,N_21647);
xor U21980 (N_21980,N_21702,N_21593);
or U21981 (N_21981,N_21696,N_21618);
or U21982 (N_21982,N_21593,N_21635);
nand U21983 (N_21983,N_21624,N_21563);
and U21984 (N_21984,N_21704,N_21727);
xnor U21985 (N_21985,N_21567,N_21516);
nor U21986 (N_21986,N_21716,N_21550);
or U21987 (N_21987,N_21744,N_21677);
xor U21988 (N_21988,N_21717,N_21736);
nor U21989 (N_21989,N_21673,N_21505);
nand U21990 (N_21990,N_21660,N_21553);
nand U21991 (N_21991,N_21605,N_21515);
and U21992 (N_21992,N_21639,N_21726);
and U21993 (N_21993,N_21705,N_21655);
xnor U21994 (N_21994,N_21696,N_21681);
and U21995 (N_21995,N_21711,N_21521);
nand U21996 (N_21996,N_21516,N_21635);
xnor U21997 (N_21997,N_21707,N_21564);
and U21998 (N_21998,N_21536,N_21629);
xor U21999 (N_21999,N_21533,N_21579);
nor U22000 (N_22000,N_21833,N_21987);
or U22001 (N_22001,N_21885,N_21923);
nor U22002 (N_22002,N_21804,N_21819);
nand U22003 (N_22003,N_21775,N_21887);
nor U22004 (N_22004,N_21812,N_21818);
and U22005 (N_22005,N_21838,N_21984);
xnor U22006 (N_22006,N_21945,N_21920);
or U22007 (N_22007,N_21755,N_21814);
and U22008 (N_22008,N_21898,N_21900);
and U22009 (N_22009,N_21990,N_21928);
nor U22010 (N_22010,N_21808,N_21946);
or U22011 (N_22011,N_21758,N_21910);
or U22012 (N_22012,N_21968,N_21986);
nand U22013 (N_22013,N_21947,N_21779);
nor U22014 (N_22014,N_21974,N_21925);
nor U22015 (N_22015,N_21911,N_21913);
or U22016 (N_22016,N_21912,N_21922);
nand U22017 (N_22017,N_21853,N_21849);
nand U22018 (N_22018,N_21908,N_21877);
xor U22019 (N_22019,N_21992,N_21896);
or U22020 (N_22020,N_21862,N_21916);
or U22021 (N_22021,N_21964,N_21832);
nand U22022 (N_22022,N_21865,N_21997);
or U22023 (N_22023,N_21991,N_21800);
nor U22024 (N_22024,N_21905,N_21772);
and U22025 (N_22025,N_21753,N_21881);
xor U22026 (N_22026,N_21893,N_21999);
or U22027 (N_22027,N_21941,N_21882);
nand U22028 (N_22028,N_21939,N_21926);
xnor U22029 (N_22029,N_21759,N_21764);
nor U22030 (N_22030,N_21857,N_21914);
nor U22031 (N_22031,N_21846,N_21763);
nand U22032 (N_22032,N_21963,N_21785);
nor U22033 (N_22033,N_21762,N_21782);
or U22034 (N_22034,N_21820,N_21867);
xnor U22035 (N_22035,N_21957,N_21932);
and U22036 (N_22036,N_21767,N_21852);
and U22037 (N_22037,N_21891,N_21944);
nand U22038 (N_22038,N_21953,N_21972);
and U22039 (N_22039,N_21958,N_21949);
and U22040 (N_22040,N_21988,N_21828);
and U22041 (N_22041,N_21844,N_21869);
nand U22042 (N_22042,N_21786,N_21831);
xor U22043 (N_22043,N_21854,N_21791);
nor U22044 (N_22044,N_21927,N_21909);
nor U22045 (N_22045,N_21825,N_21821);
nor U22046 (N_22046,N_21871,N_21899);
nor U22047 (N_22047,N_21970,N_21805);
or U22048 (N_22048,N_21952,N_21792);
and U22049 (N_22049,N_21872,N_21813);
nand U22050 (N_22050,N_21858,N_21794);
xnor U22051 (N_22051,N_21904,N_21847);
and U22052 (N_22052,N_21883,N_21868);
xor U22053 (N_22053,N_21835,N_21980);
xor U22054 (N_22054,N_21864,N_21751);
or U22055 (N_22055,N_21940,N_21915);
and U22056 (N_22056,N_21770,N_21766);
or U22057 (N_22057,N_21873,N_21777);
nand U22058 (N_22058,N_21967,N_21981);
nand U22059 (N_22059,N_21757,N_21827);
nor U22060 (N_22060,N_21801,N_21894);
xnor U22061 (N_22061,N_21876,N_21760);
nor U22062 (N_22062,N_21906,N_21822);
nand U22063 (N_22063,N_21901,N_21938);
xnor U22064 (N_22064,N_21934,N_21975);
nor U22065 (N_22065,N_21917,N_21955);
and U22066 (N_22066,N_21769,N_21826);
nand U22067 (N_22067,N_21778,N_21860);
or U22068 (N_22068,N_21870,N_21982);
nand U22069 (N_22069,N_21977,N_21851);
and U22070 (N_22070,N_21810,N_21796);
xor U22071 (N_22071,N_21965,N_21836);
or U22072 (N_22072,N_21998,N_21880);
and U22073 (N_22073,N_21781,N_21929);
and U22074 (N_22074,N_21930,N_21839);
nand U22075 (N_22075,N_21790,N_21888);
or U22076 (N_22076,N_21787,N_21834);
or U22077 (N_22077,N_21850,N_21803);
and U22078 (N_22078,N_21830,N_21823);
xor U22079 (N_22079,N_21856,N_21879);
or U22080 (N_22080,N_21817,N_21948);
or U22081 (N_22081,N_21774,N_21961);
or U22082 (N_22082,N_21976,N_21993);
xnor U22083 (N_22083,N_21962,N_21837);
nand U22084 (N_22084,N_21979,N_21861);
xor U22085 (N_22085,N_21890,N_21848);
xnor U22086 (N_22086,N_21884,N_21843);
and U22087 (N_22087,N_21784,N_21985);
xnor U22088 (N_22088,N_21892,N_21902);
or U22089 (N_22089,N_21995,N_21788);
or U22090 (N_22090,N_21895,N_21969);
or U22091 (N_22091,N_21807,N_21809);
xor U22092 (N_22092,N_21989,N_21752);
and U22093 (N_22093,N_21761,N_21996);
or U22094 (N_22094,N_21933,N_21956);
nor U22095 (N_22095,N_21874,N_21776);
and U22096 (N_22096,N_21960,N_21983);
nand U22097 (N_22097,N_21966,N_21845);
nor U22098 (N_22098,N_21924,N_21875);
xor U22099 (N_22099,N_21943,N_21931);
and U22100 (N_22100,N_21771,N_21811);
nand U22101 (N_22101,N_21824,N_21780);
or U22102 (N_22102,N_21768,N_21799);
nor U22103 (N_22103,N_21841,N_21907);
nand U22104 (N_22104,N_21829,N_21863);
nor U22105 (N_22105,N_21971,N_21942);
xnor U22106 (N_22106,N_21756,N_21978);
xnor U22107 (N_22107,N_21754,N_21918);
xnor U22108 (N_22108,N_21951,N_21936);
nand U22109 (N_22109,N_21954,N_21889);
and U22110 (N_22110,N_21903,N_21950);
or U22111 (N_22111,N_21795,N_21855);
nor U22112 (N_22112,N_21797,N_21919);
or U22113 (N_22113,N_21866,N_21959);
and U22114 (N_22114,N_21789,N_21897);
and U22115 (N_22115,N_21773,N_21750);
or U22116 (N_22116,N_21802,N_21937);
xnor U22117 (N_22117,N_21886,N_21859);
nand U22118 (N_22118,N_21973,N_21815);
and U22119 (N_22119,N_21878,N_21840);
xnor U22120 (N_22120,N_21806,N_21921);
xnor U22121 (N_22121,N_21842,N_21793);
nor U22122 (N_22122,N_21935,N_21783);
nand U22123 (N_22123,N_21816,N_21994);
nor U22124 (N_22124,N_21798,N_21765);
or U22125 (N_22125,N_21914,N_21788);
and U22126 (N_22126,N_21839,N_21894);
and U22127 (N_22127,N_21972,N_21769);
xor U22128 (N_22128,N_21859,N_21765);
nor U22129 (N_22129,N_21964,N_21958);
xor U22130 (N_22130,N_21892,N_21835);
nor U22131 (N_22131,N_21907,N_21758);
and U22132 (N_22132,N_21853,N_21895);
or U22133 (N_22133,N_21907,N_21866);
xnor U22134 (N_22134,N_21750,N_21935);
xnor U22135 (N_22135,N_21940,N_21911);
nor U22136 (N_22136,N_21990,N_21938);
or U22137 (N_22137,N_21927,N_21915);
xnor U22138 (N_22138,N_21939,N_21889);
xor U22139 (N_22139,N_21855,N_21951);
nand U22140 (N_22140,N_21754,N_21873);
and U22141 (N_22141,N_21779,N_21812);
and U22142 (N_22142,N_21976,N_21839);
or U22143 (N_22143,N_21755,N_21999);
nand U22144 (N_22144,N_21784,N_21957);
nand U22145 (N_22145,N_21750,N_21877);
nand U22146 (N_22146,N_21922,N_21822);
or U22147 (N_22147,N_21991,N_21877);
and U22148 (N_22148,N_21852,N_21769);
and U22149 (N_22149,N_21766,N_21925);
nand U22150 (N_22150,N_21845,N_21848);
or U22151 (N_22151,N_21938,N_21752);
nand U22152 (N_22152,N_21844,N_21839);
and U22153 (N_22153,N_21911,N_21991);
or U22154 (N_22154,N_21750,N_21888);
nor U22155 (N_22155,N_21860,N_21979);
or U22156 (N_22156,N_21772,N_21896);
nor U22157 (N_22157,N_21994,N_21926);
nor U22158 (N_22158,N_21939,N_21973);
or U22159 (N_22159,N_21840,N_21909);
xnor U22160 (N_22160,N_21936,N_21873);
and U22161 (N_22161,N_21796,N_21824);
and U22162 (N_22162,N_21944,N_21867);
and U22163 (N_22163,N_21806,N_21765);
or U22164 (N_22164,N_21782,N_21781);
nand U22165 (N_22165,N_21825,N_21787);
nand U22166 (N_22166,N_21922,N_21925);
xnor U22167 (N_22167,N_21755,N_21993);
nand U22168 (N_22168,N_21910,N_21766);
nand U22169 (N_22169,N_21767,N_21909);
nor U22170 (N_22170,N_21921,N_21817);
nand U22171 (N_22171,N_21804,N_21779);
xor U22172 (N_22172,N_21778,N_21888);
xnor U22173 (N_22173,N_21932,N_21790);
and U22174 (N_22174,N_21941,N_21834);
and U22175 (N_22175,N_21927,N_21940);
or U22176 (N_22176,N_21780,N_21946);
xnor U22177 (N_22177,N_21836,N_21904);
nand U22178 (N_22178,N_21752,N_21988);
xnor U22179 (N_22179,N_21842,N_21880);
nand U22180 (N_22180,N_21892,N_21922);
xnor U22181 (N_22181,N_21960,N_21781);
nand U22182 (N_22182,N_21973,N_21846);
xor U22183 (N_22183,N_21800,N_21777);
xor U22184 (N_22184,N_21771,N_21991);
nor U22185 (N_22185,N_21780,N_21893);
and U22186 (N_22186,N_21838,N_21898);
nand U22187 (N_22187,N_21922,N_21828);
or U22188 (N_22188,N_21888,N_21915);
or U22189 (N_22189,N_21784,N_21813);
nor U22190 (N_22190,N_21872,N_21980);
or U22191 (N_22191,N_21954,N_21867);
and U22192 (N_22192,N_21830,N_21876);
nand U22193 (N_22193,N_21769,N_21864);
or U22194 (N_22194,N_21774,N_21912);
nand U22195 (N_22195,N_21997,N_21989);
xor U22196 (N_22196,N_21766,N_21822);
nor U22197 (N_22197,N_21822,N_21949);
or U22198 (N_22198,N_21912,N_21964);
and U22199 (N_22199,N_21927,N_21779);
or U22200 (N_22200,N_21975,N_21922);
nand U22201 (N_22201,N_21862,N_21844);
nor U22202 (N_22202,N_21892,N_21759);
or U22203 (N_22203,N_21865,N_21763);
nand U22204 (N_22204,N_21956,N_21940);
or U22205 (N_22205,N_21911,N_21837);
nor U22206 (N_22206,N_21969,N_21959);
and U22207 (N_22207,N_21899,N_21974);
xor U22208 (N_22208,N_21966,N_21780);
and U22209 (N_22209,N_21880,N_21996);
nor U22210 (N_22210,N_21867,N_21956);
nor U22211 (N_22211,N_21921,N_21952);
xnor U22212 (N_22212,N_21774,N_21826);
or U22213 (N_22213,N_21791,N_21820);
and U22214 (N_22214,N_21990,N_21893);
and U22215 (N_22215,N_21860,N_21810);
nor U22216 (N_22216,N_21987,N_21822);
and U22217 (N_22217,N_21832,N_21961);
xnor U22218 (N_22218,N_21897,N_21853);
xor U22219 (N_22219,N_21817,N_21978);
nand U22220 (N_22220,N_21871,N_21788);
nor U22221 (N_22221,N_21873,N_21943);
xnor U22222 (N_22222,N_21969,N_21953);
nand U22223 (N_22223,N_21780,N_21847);
or U22224 (N_22224,N_21985,N_21783);
nand U22225 (N_22225,N_21933,N_21803);
or U22226 (N_22226,N_21878,N_21821);
nand U22227 (N_22227,N_21793,N_21824);
nor U22228 (N_22228,N_21767,N_21879);
and U22229 (N_22229,N_21972,N_21959);
nand U22230 (N_22230,N_21835,N_21851);
nor U22231 (N_22231,N_21775,N_21852);
nand U22232 (N_22232,N_21903,N_21808);
nand U22233 (N_22233,N_21960,N_21910);
nor U22234 (N_22234,N_21874,N_21810);
or U22235 (N_22235,N_21878,N_21786);
nand U22236 (N_22236,N_21976,N_21887);
or U22237 (N_22237,N_21751,N_21893);
and U22238 (N_22238,N_21919,N_21962);
or U22239 (N_22239,N_21904,N_21834);
nor U22240 (N_22240,N_21887,N_21855);
nor U22241 (N_22241,N_21863,N_21945);
nand U22242 (N_22242,N_21863,N_21750);
xor U22243 (N_22243,N_21889,N_21935);
and U22244 (N_22244,N_21968,N_21795);
nor U22245 (N_22245,N_21932,N_21892);
and U22246 (N_22246,N_21956,N_21806);
xor U22247 (N_22247,N_21829,N_21872);
nand U22248 (N_22248,N_21943,N_21957);
nor U22249 (N_22249,N_21880,N_21993);
nor U22250 (N_22250,N_22033,N_22055);
and U22251 (N_22251,N_22019,N_22139);
xor U22252 (N_22252,N_22241,N_22085);
xor U22253 (N_22253,N_22129,N_22024);
nor U22254 (N_22254,N_22011,N_22195);
or U22255 (N_22255,N_22211,N_22018);
nand U22256 (N_22256,N_22166,N_22067);
nor U22257 (N_22257,N_22186,N_22236);
nor U22258 (N_22258,N_22091,N_22007);
nand U22259 (N_22259,N_22196,N_22042);
or U22260 (N_22260,N_22145,N_22143);
or U22261 (N_22261,N_22046,N_22012);
or U22262 (N_22262,N_22247,N_22208);
or U22263 (N_22263,N_22061,N_22179);
and U22264 (N_22264,N_22169,N_22246);
and U22265 (N_22265,N_22117,N_22095);
xnor U22266 (N_22266,N_22022,N_22128);
nand U22267 (N_22267,N_22213,N_22232);
nor U22268 (N_22268,N_22003,N_22058);
or U22269 (N_22269,N_22132,N_22131);
nand U22270 (N_22270,N_22069,N_22014);
nor U22271 (N_22271,N_22057,N_22173);
and U22272 (N_22272,N_22175,N_22001);
xnor U22273 (N_22273,N_22079,N_22048);
and U22274 (N_22274,N_22133,N_22162);
nor U22275 (N_22275,N_22080,N_22191);
nand U22276 (N_22276,N_22160,N_22201);
xor U22277 (N_22277,N_22050,N_22222);
xor U22278 (N_22278,N_22063,N_22200);
nor U22279 (N_22279,N_22218,N_22205);
or U22280 (N_22280,N_22230,N_22093);
nor U22281 (N_22281,N_22231,N_22161);
nor U22282 (N_22282,N_22141,N_22081);
nor U22283 (N_22283,N_22189,N_22113);
xor U22284 (N_22284,N_22020,N_22051);
xnor U22285 (N_22285,N_22233,N_22036);
xnor U22286 (N_22286,N_22060,N_22116);
xnor U22287 (N_22287,N_22077,N_22157);
nor U22288 (N_22288,N_22006,N_22040);
or U22289 (N_22289,N_22108,N_22065);
and U22290 (N_22290,N_22168,N_22184);
xnor U22291 (N_22291,N_22053,N_22100);
nor U22292 (N_22292,N_22068,N_22119);
or U22293 (N_22293,N_22188,N_22192);
nand U22294 (N_22294,N_22158,N_22146);
and U22295 (N_22295,N_22062,N_22176);
nor U22296 (N_22296,N_22082,N_22219);
or U22297 (N_22297,N_22167,N_22107);
nor U22298 (N_22298,N_22094,N_22045);
nand U22299 (N_22299,N_22105,N_22140);
and U22300 (N_22300,N_22228,N_22031);
or U22301 (N_22301,N_22041,N_22084);
nand U22302 (N_22302,N_22004,N_22089);
xnor U22303 (N_22303,N_22052,N_22056);
and U22304 (N_22304,N_22190,N_22049);
nand U22305 (N_22305,N_22059,N_22087);
or U22306 (N_22306,N_22227,N_22206);
nor U22307 (N_22307,N_22203,N_22183);
xnor U22308 (N_22308,N_22178,N_22248);
or U22309 (N_22309,N_22151,N_22096);
nand U22310 (N_22310,N_22245,N_22101);
or U22311 (N_22311,N_22066,N_22071);
xor U22312 (N_22312,N_22144,N_22038);
or U22313 (N_22313,N_22198,N_22090);
xor U22314 (N_22314,N_22153,N_22194);
xnor U22315 (N_22315,N_22074,N_22110);
or U22316 (N_22316,N_22037,N_22127);
and U22317 (N_22317,N_22148,N_22135);
or U22318 (N_22318,N_22075,N_22210);
or U22319 (N_22319,N_22070,N_22026);
xor U22320 (N_22320,N_22076,N_22008);
xnor U22321 (N_22321,N_22137,N_22182);
nand U22322 (N_22322,N_22244,N_22002);
nor U22323 (N_22323,N_22225,N_22152);
or U22324 (N_22324,N_22199,N_22023);
nor U22325 (N_22325,N_22083,N_22229);
and U22326 (N_22326,N_22207,N_22187);
xnor U22327 (N_22327,N_22156,N_22121);
xnor U22328 (N_22328,N_22030,N_22235);
xnor U22329 (N_22329,N_22109,N_22193);
and U22330 (N_22330,N_22044,N_22102);
xor U22331 (N_22331,N_22214,N_22138);
and U22332 (N_22332,N_22159,N_22025);
nor U22333 (N_22333,N_22134,N_22064);
or U22334 (N_22334,N_22220,N_22072);
or U22335 (N_22335,N_22249,N_22015);
or U22336 (N_22336,N_22098,N_22212);
xor U22337 (N_22337,N_22112,N_22154);
nor U22338 (N_22338,N_22185,N_22017);
nor U22339 (N_22339,N_22111,N_22122);
nand U22340 (N_22340,N_22088,N_22016);
or U22341 (N_22341,N_22039,N_22130);
xor U22342 (N_22342,N_22000,N_22177);
or U22343 (N_22343,N_22180,N_22150);
or U22344 (N_22344,N_22147,N_22005);
nor U22345 (N_22345,N_22243,N_22054);
and U22346 (N_22346,N_22027,N_22217);
or U22347 (N_22347,N_22171,N_22086);
nor U22348 (N_22348,N_22170,N_22123);
and U22349 (N_22349,N_22221,N_22240);
nor U22350 (N_22350,N_22149,N_22009);
nand U22351 (N_22351,N_22197,N_22237);
xor U22352 (N_22352,N_22029,N_22043);
xnor U22353 (N_22353,N_22032,N_22239);
nor U22354 (N_22354,N_22163,N_22073);
xor U22355 (N_22355,N_22224,N_22035);
or U22356 (N_22356,N_22013,N_22142);
or U22357 (N_22357,N_22164,N_22226);
nor U22358 (N_22358,N_22165,N_22215);
xnor U22359 (N_22359,N_22097,N_22120);
or U22360 (N_22360,N_22034,N_22115);
xnor U22361 (N_22361,N_22118,N_22126);
nand U22362 (N_22362,N_22021,N_22204);
and U22363 (N_22363,N_22125,N_22242);
and U22364 (N_22364,N_22104,N_22092);
xnor U22365 (N_22365,N_22216,N_22099);
nor U22366 (N_22366,N_22028,N_22047);
nand U22367 (N_22367,N_22078,N_22209);
xnor U22368 (N_22368,N_22202,N_22155);
or U22369 (N_22369,N_22106,N_22114);
nor U22370 (N_22370,N_22223,N_22124);
and U22371 (N_22371,N_22181,N_22234);
nor U22372 (N_22372,N_22172,N_22103);
nor U22373 (N_22373,N_22010,N_22174);
and U22374 (N_22374,N_22136,N_22238);
and U22375 (N_22375,N_22014,N_22163);
xor U22376 (N_22376,N_22012,N_22153);
xor U22377 (N_22377,N_22191,N_22178);
xnor U22378 (N_22378,N_22083,N_22234);
nor U22379 (N_22379,N_22097,N_22022);
or U22380 (N_22380,N_22031,N_22156);
or U22381 (N_22381,N_22139,N_22013);
xnor U22382 (N_22382,N_22034,N_22214);
and U22383 (N_22383,N_22189,N_22099);
and U22384 (N_22384,N_22231,N_22058);
or U22385 (N_22385,N_22018,N_22188);
nand U22386 (N_22386,N_22191,N_22179);
xor U22387 (N_22387,N_22161,N_22150);
and U22388 (N_22388,N_22035,N_22036);
or U22389 (N_22389,N_22195,N_22053);
xor U22390 (N_22390,N_22192,N_22052);
or U22391 (N_22391,N_22137,N_22040);
and U22392 (N_22392,N_22137,N_22057);
or U22393 (N_22393,N_22216,N_22205);
nor U22394 (N_22394,N_22029,N_22126);
and U22395 (N_22395,N_22181,N_22214);
xor U22396 (N_22396,N_22246,N_22174);
xor U22397 (N_22397,N_22144,N_22161);
or U22398 (N_22398,N_22079,N_22216);
and U22399 (N_22399,N_22076,N_22040);
nor U22400 (N_22400,N_22039,N_22102);
xnor U22401 (N_22401,N_22206,N_22219);
or U22402 (N_22402,N_22194,N_22100);
xnor U22403 (N_22403,N_22037,N_22093);
xor U22404 (N_22404,N_22086,N_22184);
or U22405 (N_22405,N_22087,N_22198);
nor U22406 (N_22406,N_22091,N_22019);
or U22407 (N_22407,N_22192,N_22205);
or U22408 (N_22408,N_22182,N_22186);
xnor U22409 (N_22409,N_22093,N_22153);
and U22410 (N_22410,N_22001,N_22104);
nand U22411 (N_22411,N_22215,N_22117);
and U22412 (N_22412,N_22094,N_22240);
xnor U22413 (N_22413,N_22075,N_22248);
or U22414 (N_22414,N_22101,N_22130);
xnor U22415 (N_22415,N_22102,N_22040);
and U22416 (N_22416,N_22219,N_22059);
and U22417 (N_22417,N_22178,N_22098);
xor U22418 (N_22418,N_22159,N_22070);
or U22419 (N_22419,N_22146,N_22077);
xnor U22420 (N_22420,N_22151,N_22123);
xor U22421 (N_22421,N_22066,N_22214);
and U22422 (N_22422,N_22243,N_22176);
and U22423 (N_22423,N_22075,N_22185);
xor U22424 (N_22424,N_22209,N_22035);
or U22425 (N_22425,N_22159,N_22072);
nand U22426 (N_22426,N_22057,N_22058);
nor U22427 (N_22427,N_22065,N_22144);
and U22428 (N_22428,N_22164,N_22184);
nand U22429 (N_22429,N_22012,N_22128);
xnor U22430 (N_22430,N_22122,N_22211);
nand U22431 (N_22431,N_22033,N_22129);
nor U22432 (N_22432,N_22132,N_22079);
nand U22433 (N_22433,N_22054,N_22017);
xor U22434 (N_22434,N_22168,N_22207);
xor U22435 (N_22435,N_22117,N_22086);
nor U22436 (N_22436,N_22136,N_22126);
xnor U22437 (N_22437,N_22160,N_22151);
or U22438 (N_22438,N_22176,N_22197);
and U22439 (N_22439,N_22152,N_22121);
or U22440 (N_22440,N_22142,N_22154);
or U22441 (N_22441,N_22083,N_22166);
xnor U22442 (N_22442,N_22138,N_22170);
and U22443 (N_22443,N_22216,N_22232);
nand U22444 (N_22444,N_22089,N_22126);
nand U22445 (N_22445,N_22105,N_22235);
xnor U22446 (N_22446,N_22152,N_22238);
and U22447 (N_22447,N_22132,N_22189);
or U22448 (N_22448,N_22175,N_22105);
nor U22449 (N_22449,N_22193,N_22066);
xor U22450 (N_22450,N_22067,N_22073);
xnor U22451 (N_22451,N_22216,N_22139);
or U22452 (N_22452,N_22009,N_22106);
or U22453 (N_22453,N_22097,N_22074);
nand U22454 (N_22454,N_22022,N_22082);
or U22455 (N_22455,N_22140,N_22146);
or U22456 (N_22456,N_22007,N_22062);
xor U22457 (N_22457,N_22208,N_22180);
xor U22458 (N_22458,N_22046,N_22142);
or U22459 (N_22459,N_22245,N_22124);
xnor U22460 (N_22460,N_22065,N_22134);
nor U22461 (N_22461,N_22013,N_22133);
and U22462 (N_22462,N_22247,N_22116);
and U22463 (N_22463,N_22103,N_22161);
or U22464 (N_22464,N_22100,N_22191);
and U22465 (N_22465,N_22247,N_22235);
xor U22466 (N_22466,N_22090,N_22100);
nor U22467 (N_22467,N_22188,N_22171);
xnor U22468 (N_22468,N_22191,N_22163);
and U22469 (N_22469,N_22029,N_22077);
or U22470 (N_22470,N_22192,N_22045);
nor U22471 (N_22471,N_22040,N_22227);
or U22472 (N_22472,N_22174,N_22170);
nor U22473 (N_22473,N_22062,N_22197);
nor U22474 (N_22474,N_22000,N_22189);
nor U22475 (N_22475,N_22021,N_22123);
xnor U22476 (N_22476,N_22148,N_22017);
and U22477 (N_22477,N_22068,N_22172);
nor U22478 (N_22478,N_22178,N_22182);
xnor U22479 (N_22479,N_22087,N_22171);
nor U22480 (N_22480,N_22196,N_22145);
nand U22481 (N_22481,N_22112,N_22222);
xor U22482 (N_22482,N_22064,N_22020);
nand U22483 (N_22483,N_22094,N_22146);
nand U22484 (N_22484,N_22229,N_22140);
and U22485 (N_22485,N_22069,N_22121);
nand U22486 (N_22486,N_22019,N_22006);
or U22487 (N_22487,N_22151,N_22012);
nor U22488 (N_22488,N_22047,N_22209);
nand U22489 (N_22489,N_22152,N_22167);
xor U22490 (N_22490,N_22199,N_22123);
xnor U22491 (N_22491,N_22071,N_22094);
nand U22492 (N_22492,N_22046,N_22102);
nor U22493 (N_22493,N_22059,N_22154);
xnor U22494 (N_22494,N_22085,N_22240);
nor U22495 (N_22495,N_22183,N_22046);
or U22496 (N_22496,N_22101,N_22015);
or U22497 (N_22497,N_22153,N_22098);
and U22498 (N_22498,N_22238,N_22168);
and U22499 (N_22499,N_22039,N_22191);
xnor U22500 (N_22500,N_22368,N_22260);
xor U22501 (N_22501,N_22251,N_22496);
or U22502 (N_22502,N_22495,N_22308);
nand U22503 (N_22503,N_22259,N_22432);
and U22504 (N_22504,N_22410,N_22424);
and U22505 (N_22505,N_22377,N_22345);
or U22506 (N_22506,N_22399,N_22333);
nor U22507 (N_22507,N_22394,N_22487);
nor U22508 (N_22508,N_22453,N_22463);
and U22509 (N_22509,N_22441,N_22371);
or U22510 (N_22510,N_22395,N_22253);
nor U22511 (N_22511,N_22374,N_22415);
nor U22512 (N_22512,N_22302,N_22334);
xnor U22513 (N_22513,N_22329,N_22279);
or U22514 (N_22514,N_22477,N_22484);
and U22515 (N_22515,N_22284,N_22444);
nand U22516 (N_22516,N_22330,N_22491);
and U22517 (N_22517,N_22443,N_22375);
or U22518 (N_22518,N_22266,N_22268);
or U22519 (N_22519,N_22317,N_22342);
nand U22520 (N_22520,N_22470,N_22328);
nor U22521 (N_22521,N_22250,N_22365);
or U22522 (N_22522,N_22391,N_22381);
or U22523 (N_22523,N_22425,N_22312);
nand U22524 (N_22524,N_22316,N_22256);
nand U22525 (N_22525,N_22489,N_22478);
nor U22526 (N_22526,N_22339,N_22389);
nand U22527 (N_22527,N_22386,N_22289);
xnor U22528 (N_22528,N_22303,N_22318);
and U22529 (N_22529,N_22350,N_22315);
xor U22530 (N_22530,N_22431,N_22422);
or U22531 (N_22531,N_22467,N_22497);
xnor U22532 (N_22532,N_22490,N_22382);
or U22533 (N_22533,N_22347,N_22298);
nand U22534 (N_22534,N_22255,N_22483);
xor U22535 (N_22535,N_22413,N_22384);
or U22536 (N_22536,N_22494,N_22357);
or U22537 (N_22537,N_22473,N_22421);
or U22538 (N_22538,N_22306,N_22273);
nor U22539 (N_22539,N_22323,N_22493);
xor U22540 (N_22540,N_22310,N_22403);
nand U22541 (N_22541,N_22468,N_22276);
xnor U22542 (N_22542,N_22498,N_22285);
or U22543 (N_22543,N_22355,N_22429);
nand U22544 (N_22544,N_22460,N_22362);
and U22545 (N_22545,N_22401,N_22353);
nand U22546 (N_22546,N_22331,N_22414);
and U22547 (N_22547,N_22313,N_22352);
xor U22548 (N_22548,N_22390,N_22445);
xnor U22549 (N_22549,N_22412,N_22370);
nand U22550 (N_22550,N_22332,N_22469);
nand U22551 (N_22551,N_22346,N_22461);
nor U22552 (N_22552,N_22387,N_22292);
nor U22553 (N_22553,N_22278,N_22283);
nor U22554 (N_22554,N_22397,N_22393);
and U22555 (N_22555,N_22442,N_22290);
nor U22556 (N_22556,N_22433,N_22416);
and U22557 (N_22557,N_22356,N_22499);
xor U22558 (N_22558,N_22455,N_22282);
and U22559 (N_22559,N_22417,N_22485);
xor U22560 (N_22560,N_22405,N_22309);
and U22561 (N_22561,N_22423,N_22367);
nand U22562 (N_22562,N_22411,N_22430);
nor U22563 (N_22563,N_22471,N_22379);
and U22564 (N_22564,N_22439,N_22291);
or U22565 (N_22565,N_22409,N_22407);
nor U22566 (N_22566,N_22349,N_22465);
and U22567 (N_22567,N_22435,N_22396);
or U22568 (N_22568,N_22482,N_22472);
and U22569 (N_22569,N_22277,N_22321);
xnor U22570 (N_22570,N_22456,N_22452);
or U22571 (N_22571,N_22336,N_22479);
xor U22572 (N_22572,N_22311,N_22319);
or U22573 (N_22573,N_22252,N_22359);
xor U22574 (N_22574,N_22488,N_22457);
and U22575 (N_22575,N_22449,N_22392);
xnor U22576 (N_22576,N_22344,N_22341);
xnor U22577 (N_22577,N_22327,N_22454);
or U22578 (N_22578,N_22480,N_22361);
or U22579 (N_22579,N_22300,N_22286);
nand U22580 (N_22580,N_22326,N_22301);
nor U22581 (N_22581,N_22270,N_22288);
xnor U22582 (N_22582,N_22380,N_22419);
and U22583 (N_22583,N_22481,N_22486);
and U22584 (N_22584,N_22378,N_22404);
nand U22585 (N_22585,N_22262,N_22272);
nor U22586 (N_22586,N_22281,N_22372);
xor U22587 (N_22587,N_22280,N_22335);
xor U22588 (N_22588,N_22307,N_22348);
xnor U22589 (N_22589,N_22466,N_22426);
and U22590 (N_22590,N_22462,N_22274);
xor U22591 (N_22591,N_22388,N_22299);
xor U22592 (N_22592,N_22324,N_22358);
or U22593 (N_22593,N_22383,N_22428);
or U22594 (N_22594,N_22325,N_22427);
nand U22595 (N_22595,N_22294,N_22492);
nor U22596 (N_22596,N_22475,N_22436);
nor U22597 (N_22597,N_22450,N_22265);
or U22598 (N_22598,N_22293,N_22271);
nand U22599 (N_22599,N_22287,N_22261);
and U22600 (N_22600,N_22366,N_22418);
nor U22601 (N_22601,N_22448,N_22476);
nor U22602 (N_22602,N_22464,N_22295);
nand U22603 (N_22603,N_22351,N_22474);
and U22604 (N_22604,N_22373,N_22343);
nand U22605 (N_22605,N_22451,N_22437);
xnor U22606 (N_22606,N_22254,N_22406);
nor U22607 (N_22607,N_22363,N_22269);
xor U22608 (N_22608,N_22267,N_22263);
xnor U22609 (N_22609,N_22420,N_22376);
nand U22610 (N_22610,N_22296,N_22258);
xnor U22611 (N_22611,N_22459,N_22434);
nand U22612 (N_22612,N_22297,N_22408);
xor U22613 (N_22613,N_22438,N_22402);
xor U22614 (N_22614,N_22264,N_22385);
nor U22615 (N_22615,N_22337,N_22446);
and U22616 (N_22616,N_22304,N_22354);
and U22617 (N_22617,N_22364,N_22320);
and U22618 (N_22618,N_22400,N_22340);
nor U22619 (N_22619,N_22398,N_22314);
and U22620 (N_22620,N_22305,N_22257);
and U22621 (N_22621,N_22447,N_22369);
and U22622 (N_22622,N_22322,N_22338);
nand U22623 (N_22623,N_22440,N_22275);
nand U22624 (N_22624,N_22360,N_22458);
or U22625 (N_22625,N_22264,N_22289);
nand U22626 (N_22626,N_22290,N_22260);
and U22627 (N_22627,N_22346,N_22268);
nand U22628 (N_22628,N_22338,N_22452);
or U22629 (N_22629,N_22446,N_22363);
or U22630 (N_22630,N_22333,N_22297);
or U22631 (N_22631,N_22375,N_22414);
nor U22632 (N_22632,N_22264,N_22485);
nor U22633 (N_22633,N_22469,N_22363);
nand U22634 (N_22634,N_22315,N_22346);
nand U22635 (N_22635,N_22337,N_22293);
nor U22636 (N_22636,N_22313,N_22336);
xnor U22637 (N_22637,N_22492,N_22416);
or U22638 (N_22638,N_22435,N_22327);
nor U22639 (N_22639,N_22434,N_22346);
and U22640 (N_22640,N_22272,N_22460);
xnor U22641 (N_22641,N_22289,N_22327);
xnor U22642 (N_22642,N_22339,N_22255);
nand U22643 (N_22643,N_22446,N_22309);
nor U22644 (N_22644,N_22250,N_22382);
nor U22645 (N_22645,N_22459,N_22395);
and U22646 (N_22646,N_22474,N_22383);
nor U22647 (N_22647,N_22303,N_22306);
and U22648 (N_22648,N_22333,N_22412);
nor U22649 (N_22649,N_22425,N_22333);
nand U22650 (N_22650,N_22473,N_22482);
nor U22651 (N_22651,N_22387,N_22403);
nand U22652 (N_22652,N_22498,N_22309);
nor U22653 (N_22653,N_22342,N_22336);
xnor U22654 (N_22654,N_22348,N_22413);
nand U22655 (N_22655,N_22377,N_22365);
and U22656 (N_22656,N_22396,N_22344);
nor U22657 (N_22657,N_22396,N_22250);
and U22658 (N_22658,N_22376,N_22288);
or U22659 (N_22659,N_22356,N_22402);
and U22660 (N_22660,N_22345,N_22253);
or U22661 (N_22661,N_22383,N_22495);
or U22662 (N_22662,N_22395,N_22408);
or U22663 (N_22663,N_22483,N_22411);
or U22664 (N_22664,N_22452,N_22393);
xor U22665 (N_22665,N_22399,N_22444);
nor U22666 (N_22666,N_22466,N_22300);
and U22667 (N_22667,N_22434,N_22347);
or U22668 (N_22668,N_22371,N_22395);
xnor U22669 (N_22669,N_22253,N_22291);
nor U22670 (N_22670,N_22295,N_22347);
nand U22671 (N_22671,N_22433,N_22447);
nand U22672 (N_22672,N_22393,N_22280);
or U22673 (N_22673,N_22315,N_22336);
nand U22674 (N_22674,N_22452,N_22382);
nand U22675 (N_22675,N_22373,N_22383);
xor U22676 (N_22676,N_22371,N_22390);
nand U22677 (N_22677,N_22292,N_22288);
nand U22678 (N_22678,N_22340,N_22416);
xnor U22679 (N_22679,N_22331,N_22332);
nand U22680 (N_22680,N_22341,N_22465);
and U22681 (N_22681,N_22481,N_22474);
xnor U22682 (N_22682,N_22453,N_22349);
and U22683 (N_22683,N_22448,N_22288);
xor U22684 (N_22684,N_22411,N_22449);
nor U22685 (N_22685,N_22440,N_22401);
or U22686 (N_22686,N_22310,N_22337);
xnor U22687 (N_22687,N_22435,N_22495);
and U22688 (N_22688,N_22276,N_22356);
nor U22689 (N_22689,N_22258,N_22466);
or U22690 (N_22690,N_22258,N_22393);
and U22691 (N_22691,N_22376,N_22327);
nand U22692 (N_22692,N_22289,N_22349);
or U22693 (N_22693,N_22289,N_22331);
nor U22694 (N_22694,N_22283,N_22310);
nand U22695 (N_22695,N_22280,N_22329);
and U22696 (N_22696,N_22437,N_22388);
xor U22697 (N_22697,N_22401,N_22311);
nor U22698 (N_22698,N_22305,N_22251);
nand U22699 (N_22699,N_22376,N_22285);
nand U22700 (N_22700,N_22492,N_22402);
or U22701 (N_22701,N_22385,N_22347);
nor U22702 (N_22702,N_22280,N_22486);
and U22703 (N_22703,N_22353,N_22258);
xor U22704 (N_22704,N_22390,N_22438);
nor U22705 (N_22705,N_22301,N_22401);
or U22706 (N_22706,N_22312,N_22396);
nand U22707 (N_22707,N_22306,N_22334);
or U22708 (N_22708,N_22291,N_22466);
and U22709 (N_22709,N_22300,N_22283);
nand U22710 (N_22710,N_22387,N_22299);
nand U22711 (N_22711,N_22483,N_22280);
and U22712 (N_22712,N_22417,N_22472);
and U22713 (N_22713,N_22388,N_22474);
or U22714 (N_22714,N_22445,N_22272);
xor U22715 (N_22715,N_22310,N_22424);
nor U22716 (N_22716,N_22477,N_22346);
nor U22717 (N_22717,N_22272,N_22319);
and U22718 (N_22718,N_22362,N_22280);
nor U22719 (N_22719,N_22347,N_22384);
and U22720 (N_22720,N_22279,N_22453);
nand U22721 (N_22721,N_22419,N_22387);
nor U22722 (N_22722,N_22432,N_22389);
xnor U22723 (N_22723,N_22318,N_22280);
and U22724 (N_22724,N_22336,N_22390);
xor U22725 (N_22725,N_22463,N_22494);
nand U22726 (N_22726,N_22464,N_22264);
and U22727 (N_22727,N_22335,N_22424);
nand U22728 (N_22728,N_22455,N_22382);
and U22729 (N_22729,N_22464,N_22302);
nand U22730 (N_22730,N_22298,N_22433);
nand U22731 (N_22731,N_22260,N_22329);
nand U22732 (N_22732,N_22331,N_22282);
or U22733 (N_22733,N_22276,N_22395);
nand U22734 (N_22734,N_22297,N_22252);
nor U22735 (N_22735,N_22365,N_22364);
nor U22736 (N_22736,N_22408,N_22392);
and U22737 (N_22737,N_22351,N_22313);
or U22738 (N_22738,N_22376,N_22283);
nand U22739 (N_22739,N_22322,N_22328);
and U22740 (N_22740,N_22485,N_22324);
and U22741 (N_22741,N_22339,N_22264);
xor U22742 (N_22742,N_22478,N_22340);
xnor U22743 (N_22743,N_22433,N_22319);
xor U22744 (N_22744,N_22287,N_22324);
nor U22745 (N_22745,N_22266,N_22379);
xnor U22746 (N_22746,N_22363,N_22437);
or U22747 (N_22747,N_22470,N_22435);
nand U22748 (N_22748,N_22468,N_22291);
nand U22749 (N_22749,N_22267,N_22277);
or U22750 (N_22750,N_22657,N_22592);
xor U22751 (N_22751,N_22685,N_22564);
and U22752 (N_22752,N_22598,N_22672);
and U22753 (N_22753,N_22610,N_22692);
nand U22754 (N_22754,N_22578,N_22633);
and U22755 (N_22755,N_22686,N_22509);
nand U22756 (N_22756,N_22715,N_22713);
nand U22757 (N_22757,N_22502,N_22553);
nand U22758 (N_22758,N_22611,N_22508);
nor U22759 (N_22759,N_22643,N_22644);
nand U22760 (N_22760,N_22503,N_22647);
and U22761 (N_22761,N_22655,N_22583);
nand U22762 (N_22762,N_22641,N_22595);
xor U22763 (N_22763,N_22697,N_22634);
nand U22764 (N_22764,N_22586,N_22512);
nor U22765 (N_22765,N_22582,N_22581);
or U22766 (N_22766,N_22520,N_22678);
or U22767 (N_22767,N_22673,N_22649);
xnor U22768 (N_22768,N_22566,N_22667);
nor U22769 (N_22769,N_22671,N_22711);
xor U22770 (N_22770,N_22574,N_22533);
and U22771 (N_22771,N_22620,N_22700);
nor U22772 (N_22772,N_22590,N_22603);
xnor U22773 (N_22773,N_22626,N_22628);
nor U22774 (N_22774,N_22614,N_22691);
or U22775 (N_22775,N_22573,N_22510);
or U22776 (N_22776,N_22518,N_22654);
or U22777 (N_22777,N_22524,N_22661);
xnor U22778 (N_22778,N_22571,N_22696);
or U22779 (N_22779,N_22651,N_22530);
nand U22780 (N_22780,N_22642,N_22619);
xnor U22781 (N_22781,N_22526,N_22523);
xor U22782 (N_22782,N_22679,N_22570);
nor U22783 (N_22783,N_22708,N_22561);
and U22784 (N_22784,N_22618,N_22545);
and U22785 (N_22785,N_22528,N_22727);
or U22786 (N_22786,N_22710,N_22698);
or U22787 (N_22787,N_22660,N_22638);
xnor U22788 (N_22788,N_22552,N_22741);
or U22789 (N_22789,N_22635,N_22677);
and U22790 (N_22790,N_22589,N_22615);
nand U22791 (N_22791,N_22535,N_22717);
nand U22792 (N_22792,N_22560,N_22722);
or U22793 (N_22793,N_22629,N_22605);
and U22794 (N_22794,N_22558,N_22707);
or U22795 (N_22795,N_22664,N_22748);
nor U22796 (N_22796,N_22522,N_22511);
xnor U22797 (N_22797,N_22580,N_22701);
and U22798 (N_22798,N_22714,N_22622);
nand U22799 (N_22799,N_22650,N_22540);
or U22800 (N_22800,N_22683,N_22745);
or U22801 (N_22801,N_22680,N_22551);
nor U22802 (N_22802,N_22728,N_22631);
nor U22803 (N_22803,N_22720,N_22624);
nand U22804 (N_22804,N_22705,N_22625);
nand U22805 (N_22805,N_22737,N_22519);
nand U22806 (N_22806,N_22684,N_22637);
nor U22807 (N_22807,N_22746,N_22585);
xor U22808 (N_22808,N_22501,N_22702);
nand U22809 (N_22809,N_22537,N_22703);
xor U22810 (N_22810,N_22607,N_22593);
nor U22811 (N_22811,N_22612,N_22709);
or U22812 (N_22812,N_22597,N_22645);
nand U22813 (N_22813,N_22588,N_22646);
nor U22814 (N_22814,N_22653,N_22500);
and U22815 (N_22815,N_22639,N_22565);
nand U22816 (N_22816,N_22681,N_22627);
nor U22817 (N_22817,N_22704,N_22594);
xnor U22818 (N_22818,N_22648,N_22738);
nor U22819 (N_22819,N_22517,N_22749);
xnor U22820 (N_22820,N_22587,N_22719);
or U22821 (N_22821,N_22604,N_22542);
and U22822 (N_22822,N_22576,N_22532);
or U22823 (N_22823,N_22726,N_22689);
nor U22824 (N_22824,N_22735,N_22543);
or U22825 (N_22825,N_22608,N_22544);
nand U22826 (N_22826,N_22743,N_22662);
and U22827 (N_22827,N_22538,N_22600);
nor U22828 (N_22828,N_22572,N_22623);
nor U22829 (N_22829,N_22652,N_22548);
xor U22830 (N_22830,N_22731,N_22729);
nor U22831 (N_22831,N_22670,N_22656);
xor U22832 (N_22832,N_22663,N_22632);
or U22833 (N_22833,N_22579,N_22531);
or U22834 (N_22834,N_22556,N_22695);
nand U22835 (N_22835,N_22527,N_22621);
xor U22836 (N_22836,N_22541,N_22547);
or U22837 (N_22837,N_22539,N_22546);
and U22838 (N_22838,N_22730,N_22555);
xor U22839 (N_22839,N_22721,N_22736);
and U22840 (N_22840,N_22740,N_22549);
nand U22841 (N_22841,N_22536,N_22602);
nor U22842 (N_22842,N_22723,N_22562);
and U22843 (N_22843,N_22613,N_22529);
nand U22844 (N_22844,N_22515,N_22616);
nor U22845 (N_22845,N_22668,N_22688);
and U22846 (N_22846,N_22514,N_22606);
nand U22847 (N_22847,N_22609,N_22665);
nand U22848 (N_22848,N_22567,N_22669);
xnor U22849 (N_22849,N_22747,N_22725);
and U22850 (N_22850,N_22596,N_22712);
and U22851 (N_22851,N_22563,N_22554);
xnor U22852 (N_22852,N_22682,N_22584);
nor U22853 (N_22853,N_22706,N_22666);
and U22854 (N_22854,N_22659,N_22744);
or U22855 (N_22855,N_22674,N_22599);
or U22856 (N_22856,N_22694,N_22690);
nand U22857 (N_22857,N_22630,N_22521);
nor U22858 (N_22858,N_22557,N_22534);
nor U22859 (N_22859,N_22507,N_22575);
nor U22860 (N_22860,N_22577,N_22504);
and U22861 (N_22861,N_22742,N_22568);
xnor U22862 (N_22862,N_22525,N_22601);
nand U22863 (N_22863,N_22716,N_22734);
and U22864 (N_22864,N_22676,N_22733);
nor U22865 (N_22865,N_22505,N_22617);
nand U22866 (N_22866,N_22506,N_22687);
or U22867 (N_22867,N_22516,N_22658);
or U22868 (N_22868,N_22550,N_22724);
nor U22869 (N_22869,N_22513,N_22640);
nand U22870 (N_22870,N_22732,N_22675);
and U22871 (N_22871,N_22699,N_22636);
and U22872 (N_22872,N_22693,N_22718);
xnor U22873 (N_22873,N_22739,N_22569);
and U22874 (N_22874,N_22591,N_22559);
or U22875 (N_22875,N_22685,N_22736);
or U22876 (N_22876,N_22526,N_22700);
and U22877 (N_22877,N_22549,N_22589);
xor U22878 (N_22878,N_22685,N_22672);
nor U22879 (N_22879,N_22711,N_22707);
and U22880 (N_22880,N_22561,N_22510);
and U22881 (N_22881,N_22593,N_22551);
xor U22882 (N_22882,N_22593,N_22556);
xor U22883 (N_22883,N_22651,N_22749);
nand U22884 (N_22884,N_22723,N_22572);
nand U22885 (N_22885,N_22558,N_22678);
nand U22886 (N_22886,N_22720,N_22568);
nand U22887 (N_22887,N_22640,N_22706);
xor U22888 (N_22888,N_22533,N_22683);
nand U22889 (N_22889,N_22599,N_22712);
nand U22890 (N_22890,N_22625,N_22651);
xnor U22891 (N_22891,N_22575,N_22526);
nor U22892 (N_22892,N_22564,N_22602);
nor U22893 (N_22893,N_22722,N_22614);
xor U22894 (N_22894,N_22665,N_22551);
and U22895 (N_22895,N_22686,N_22747);
xor U22896 (N_22896,N_22700,N_22661);
and U22897 (N_22897,N_22665,N_22524);
and U22898 (N_22898,N_22589,N_22686);
nor U22899 (N_22899,N_22508,N_22593);
and U22900 (N_22900,N_22612,N_22539);
nor U22901 (N_22901,N_22603,N_22548);
and U22902 (N_22902,N_22722,N_22597);
nand U22903 (N_22903,N_22655,N_22612);
or U22904 (N_22904,N_22694,N_22662);
and U22905 (N_22905,N_22611,N_22652);
xnor U22906 (N_22906,N_22559,N_22520);
nor U22907 (N_22907,N_22678,N_22592);
and U22908 (N_22908,N_22565,N_22635);
xor U22909 (N_22909,N_22617,N_22547);
or U22910 (N_22910,N_22597,N_22582);
nor U22911 (N_22911,N_22589,N_22578);
or U22912 (N_22912,N_22705,N_22708);
nor U22913 (N_22913,N_22598,N_22719);
or U22914 (N_22914,N_22673,N_22722);
nor U22915 (N_22915,N_22668,N_22659);
nor U22916 (N_22916,N_22617,N_22532);
or U22917 (N_22917,N_22526,N_22704);
and U22918 (N_22918,N_22717,N_22702);
nand U22919 (N_22919,N_22617,N_22645);
nand U22920 (N_22920,N_22591,N_22532);
and U22921 (N_22921,N_22654,N_22690);
or U22922 (N_22922,N_22595,N_22743);
nand U22923 (N_22923,N_22703,N_22501);
nand U22924 (N_22924,N_22562,N_22527);
nor U22925 (N_22925,N_22642,N_22640);
nand U22926 (N_22926,N_22561,N_22506);
or U22927 (N_22927,N_22733,N_22708);
and U22928 (N_22928,N_22705,N_22694);
xnor U22929 (N_22929,N_22664,N_22616);
xnor U22930 (N_22930,N_22725,N_22509);
or U22931 (N_22931,N_22520,N_22607);
or U22932 (N_22932,N_22524,N_22711);
and U22933 (N_22933,N_22524,N_22672);
xnor U22934 (N_22934,N_22593,N_22584);
nand U22935 (N_22935,N_22583,N_22620);
nand U22936 (N_22936,N_22727,N_22659);
or U22937 (N_22937,N_22637,N_22608);
or U22938 (N_22938,N_22701,N_22534);
xor U22939 (N_22939,N_22647,N_22704);
or U22940 (N_22940,N_22570,N_22661);
or U22941 (N_22941,N_22604,N_22590);
or U22942 (N_22942,N_22522,N_22723);
xor U22943 (N_22943,N_22593,N_22684);
xnor U22944 (N_22944,N_22515,N_22690);
nor U22945 (N_22945,N_22571,N_22541);
nand U22946 (N_22946,N_22538,N_22666);
or U22947 (N_22947,N_22743,N_22641);
nor U22948 (N_22948,N_22622,N_22535);
or U22949 (N_22949,N_22557,N_22645);
nor U22950 (N_22950,N_22629,N_22644);
or U22951 (N_22951,N_22530,N_22725);
nor U22952 (N_22952,N_22588,N_22725);
and U22953 (N_22953,N_22516,N_22571);
nor U22954 (N_22954,N_22633,N_22589);
nor U22955 (N_22955,N_22605,N_22654);
xnor U22956 (N_22956,N_22712,N_22567);
nand U22957 (N_22957,N_22715,N_22549);
or U22958 (N_22958,N_22581,N_22524);
nand U22959 (N_22959,N_22679,N_22726);
or U22960 (N_22960,N_22705,N_22525);
nand U22961 (N_22961,N_22653,N_22528);
xnor U22962 (N_22962,N_22688,N_22723);
and U22963 (N_22963,N_22647,N_22556);
and U22964 (N_22964,N_22524,N_22570);
nand U22965 (N_22965,N_22685,N_22621);
nand U22966 (N_22966,N_22683,N_22514);
nor U22967 (N_22967,N_22739,N_22683);
and U22968 (N_22968,N_22688,N_22664);
or U22969 (N_22969,N_22531,N_22694);
or U22970 (N_22970,N_22639,N_22649);
or U22971 (N_22971,N_22542,N_22504);
nor U22972 (N_22972,N_22672,N_22709);
xnor U22973 (N_22973,N_22749,N_22540);
or U22974 (N_22974,N_22524,N_22580);
xnor U22975 (N_22975,N_22644,N_22597);
nand U22976 (N_22976,N_22611,N_22661);
nand U22977 (N_22977,N_22543,N_22587);
and U22978 (N_22978,N_22508,N_22701);
nand U22979 (N_22979,N_22597,N_22654);
nand U22980 (N_22980,N_22669,N_22727);
nor U22981 (N_22981,N_22738,N_22551);
nor U22982 (N_22982,N_22536,N_22506);
or U22983 (N_22983,N_22685,N_22551);
xor U22984 (N_22984,N_22582,N_22640);
or U22985 (N_22985,N_22605,N_22661);
nor U22986 (N_22986,N_22527,N_22624);
or U22987 (N_22987,N_22576,N_22599);
xnor U22988 (N_22988,N_22647,N_22711);
or U22989 (N_22989,N_22634,N_22656);
or U22990 (N_22990,N_22687,N_22616);
xor U22991 (N_22991,N_22506,N_22510);
xnor U22992 (N_22992,N_22729,N_22610);
and U22993 (N_22993,N_22672,N_22658);
nor U22994 (N_22994,N_22672,N_22633);
nor U22995 (N_22995,N_22680,N_22619);
or U22996 (N_22996,N_22635,N_22650);
or U22997 (N_22997,N_22670,N_22591);
nor U22998 (N_22998,N_22712,N_22580);
nor U22999 (N_22999,N_22689,N_22612);
or U23000 (N_23000,N_22831,N_22960);
nand U23001 (N_23001,N_22777,N_22939);
xor U23002 (N_23002,N_22929,N_22914);
nor U23003 (N_23003,N_22856,N_22954);
and U23004 (N_23004,N_22806,N_22754);
nand U23005 (N_23005,N_22999,N_22778);
or U23006 (N_23006,N_22908,N_22752);
and U23007 (N_23007,N_22863,N_22839);
nor U23008 (N_23008,N_22901,N_22886);
nand U23009 (N_23009,N_22998,N_22773);
nand U23010 (N_23010,N_22808,N_22873);
and U23011 (N_23011,N_22834,N_22771);
xnor U23012 (N_23012,N_22865,N_22790);
nand U23013 (N_23013,N_22976,N_22857);
and U23014 (N_23014,N_22907,N_22770);
xnor U23015 (N_23015,N_22897,N_22801);
xor U23016 (N_23016,N_22995,N_22854);
nor U23017 (N_23017,N_22884,N_22896);
nor U23018 (N_23018,N_22885,N_22851);
nand U23019 (N_23019,N_22989,N_22875);
xnor U23020 (N_23020,N_22872,N_22883);
xor U23021 (N_23021,N_22799,N_22951);
nor U23022 (N_23022,N_22836,N_22924);
xnor U23023 (N_23023,N_22769,N_22877);
xor U23024 (N_23024,N_22855,N_22785);
nor U23025 (N_23025,N_22803,N_22984);
nor U23026 (N_23026,N_22940,N_22992);
and U23027 (N_23027,N_22776,N_22864);
and U23028 (N_23028,N_22842,N_22990);
nor U23029 (N_23029,N_22817,N_22833);
nand U23030 (N_23030,N_22858,N_22936);
nor U23031 (N_23031,N_22913,N_22971);
or U23032 (N_23032,N_22965,N_22973);
nor U23033 (N_23033,N_22988,N_22829);
or U23034 (N_23034,N_22893,N_22784);
nand U23035 (N_23035,N_22955,N_22802);
xnor U23036 (N_23036,N_22996,N_22755);
or U23037 (N_23037,N_22925,N_22902);
or U23038 (N_23038,N_22892,N_22757);
nor U23039 (N_23039,N_22917,N_22794);
xnor U23040 (N_23040,N_22845,N_22997);
xnor U23041 (N_23041,N_22979,N_22928);
nor U23042 (N_23042,N_22987,N_22859);
nor U23043 (N_23043,N_22958,N_22822);
and U23044 (N_23044,N_22904,N_22812);
and U23045 (N_23045,N_22821,N_22763);
nor U23046 (N_23046,N_22970,N_22753);
nor U23047 (N_23047,N_22980,N_22881);
and U23048 (N_23048,N_22948,N_22919);
and U23049 (N_23049,N_22975,N_22927);
nand U23050 (N_23050,N_22780,N_22935);
nor U23051 (N_23051,N_22759,N_22846);
or U23052 (N_23052,N_22869,N_22938);
nand U23053 (N_23053,N_22756,N_22894);
xor U23054 (N_23054,N_22926,N_22882);
and U23055 (N_23055,N_22800,N_22760);
nor U23056 (N_23056,N_22789,N_22788);
xnor U23057 (N_23057,N_22781,N_22750);
or U23058 (N_23058,N_22977,N_22792);
and U23059 (N_23059,N_22993,N_22967);
or U23060 (N_23060,N_22813,N_22941);
nand U23061 (N_23061,N_22837,N_22947);
xnor U23062 (N_23062,N_22793,N_22900);
nor U23063 (N_23063,N_22994,N_22797);
or U23064 (N_23064,N_22962,N_22815);
nand U23065 (N_23065,N_22860,N_22978);
nor U23066 (N_23066,N_22910,N_22964);
nor U23067 (N_23067,N_22816,N_22915);
xor U23068 (N_23068,N_22949,N_22923);
nand U23069 (N_23069,N_22942,N_22824);
xor U23070 (N_23070,N_22775,N_22765);
and U23071 (N_23071,N_22814,N_22787);
xnor U23072 (N_23072,N_22782,N_22844);
or U23073 (N_23073,N_22876,N_22847);
and U23074 (N_23074,N_22772,N_22943);
or U23075 (N_23075,N_22849,N_22966);
and U23076 (N_23076,N_22870,N_22868);
or U23077 (N_23077,N_22805,N_22871);
and U23078 (N_23078,N_22950,N_22874);
nor U23079 (N_23079,N_22841,N_22921);
nor U23080 (N_23080,N_22982,N_22843);
and U23081 (N_23081,N_22891,N_22823);
xor U23082 (N_23082,N_22861,N_22796);
or U23083 (N_23083,N_22768,N_22899);
or U23084 (N_23084,N_22783,N_22959);
nor U23085 (N_23085,N_22825,N_22922);
or U23086 (N_23086,N_22848,N_22903);
xnor U23087 (N_23087,N_22867,N_22911);
or U23088 (N_23088,N_22798,N_22764);
or U23089 (N_23089,N_22827,N_22887);
and U23090 (N_23090,N_22866,N_22807);
and U23091 (N_23091,N_22985,N_22878);
nor U23092 (N_23092,N_22898,N_22991);
nand U23093 (N_23093,N_22889,N_22828);
or U23094 (N_23094,N_22879,N_22767);
and U23095 (N_23095,N_22811,N_22930);
nand U23096 (N_23096,N_22952,N_22918);
xor U23097 (N_23097,N_22945,N_22786);
xor U23098 (N_23098,N_22880,N_22957);
nor U23099 (N_23099,N_22912,N_22774);
nor U23100 (N_23100,N_22826,N_22986);
nor U23101 (N_23101,N_22983,N_22830);
nor U23102 (N_23102,N_22888,N_22853);
and U23103 (N_23103,N_22818,N_22961);
and U23104 (N_23104,N_22890,N_22835);
nand U23105 (N_23105,N_22895,N_22956);
and U23106 (N_23106,N_22946,N_22981);
or U23107 (N_23107,N_22795,N_22909);
or U23108 (N_23108,N_22931,N_22791);
nor U23109 (N_23109,N_22761,N_22972);
nand U23110 (N_23110,N_22862,N_22953);
nand U23111 (N_23111,N_22934,N_22944);
and U23112 (N_23112,N_22905,N_22968);
and U23113 (N_23113,N_22932,N_22779);
and U23114 (N_23114,N_22920,N_22850);
nor U23115 (N_23115,N_22933,N_22916);
nand U23116 (N_23116,N_22751,N_22762);
and U23117 (N_23117,N_22969,N_22810);
nand U23118 (N_23118,N_22840,N_22820);
and U23119 (N_23119,N_22804,N_22832);
xnor U23120 (N_23120,N_22758,N_22838);
nand U23121 (N_23121,N_22766,N_22937);
and U23122 (N_23122,N_22906,N_22963);
and U23123 (N_23123,N_22852,N_22809);
nor U23124 (N_23124,N_22819,N_22974);
nor U23125 (N_23125,N_22863,N_22871);
nand U23126 (N_23126,N_22832,N_22880);
xor U23127 (N_23127,N_22875,N_22788);
or U23128 (N_23128,N_22769,N_22816);
nand U23129 (N_23129,N_22985,N_22996);
and U23130 (N_23130,N_22945,N_22967);
xnor U23131 (N_23131,N_22959,N_22924);
or U23132 (N_23132,N_22911,N_22779);
nor U23133 (N_23133,N_22977,N_22923);
xnor U23134 (N_23134,N_22786,N_22861);
or U23135 (N_23135,N_22937,N_22825);
nand U23136 (N_23136,N_22769,N_22899);
xor U23137 (N_23137,N_22928,N_22860);
xnor U23138 (N_23138,N_22998,N_22902);
xor U23139 (N_23139,N_22789,N_22797);
and U23140 (N_23140,N_22865,N_22829);
or U23141 (N_23141,N_22830,N_22818);
or U23142 (N_23142,N_22848,N_22931);
xor U23143 (N_23143,N_22795,N_22766);
nor U23144 (N_23144,N_22844,N_22863);
nand U23145 (N_23145,N_22887,N_22947);
and U23146 (N_23146,N_22927,N_22945);
nand U23147 (N_23147,N_22765,N_22938);
nand U23148 (N_23148,N_22928,N_22963);
nand U23149 (N_23149,N_22977,N_22814);
nand U23150 (N_23150,N_22829,N_22818);
or U23151 (N_23151,N_22811,N_22887);
nand U23152 (N_23152,N_22892,N_22941);
or U23153 (N_23153,N_22952,N_22862);
xnor U23154 (N_23154,N_22755,N_22839);
nand U23155 (N_23155,N_22844,N_22897);
nand U23156 (N_23156,N_22942,N_22940);
nand U23157 (N_23157,N_22798,N_22956);
or U23158 (N_23158,N_22766,N_22896);
and U23159 (N_23159,N_22807,N_22808);
xnor U23160 (N_23160,N_22971,N_22917);
and U23161 (N_23161,N_22809,N_22871);
nor U23162 (N_23162,N_22959,N_22871);
nand U23163 (N_23163,N_22934,N_22812);
and U23164 (N_23164,N_22771,N_22884);
and U23165 (N_23165,N_22886,N_22753);
or U23166 (N_23166,N_22775,N_22861);
or U23167 (N_23167,N_22957,N_22910);
and U23168 (N_23168,N_22763,N_22831);
and U23169 (N_23169,N_22828,N_22988);
xor U23170 (N_23170,N_22849,N_22795);
nor U23171 (N_23171,N_22772,N_22826);
nor U23172 (N_23172,N_22805,N_22869);
nand U23173 (N_23173,N_22944,N_22975);
and U23174 (N_23174,N_22926,N_22951);
nor U23175 (N_23175,N_22763,N_22958);
or U23176 (N_23176,N_22975,N_22876);
nand U23177 (N_23177,N_22972,N_22755);
and U23178 (N_23178,N_22861,N_22980);
and U23179 (N_23179,N_22840,N_22895);
or U23180 (N_23180,N_22886,N_22751);
nand U23181 (N_23181,N_22793,N_22996);
and U23182 (N_23182,N_22894,N_22865);
nor U23183 (N_23183,N_22931,N_22787);
nor U23184 (N_23184,N_22905,N_22771);
nor U23185 (N_23185,N_22902,N_22788);
xor U23186 (N_23186,N_22760,N_22825);
and U23187 (N_23187,N_22810,N_22868);
or U23188 (N_23188,N_22776,N_22848);
or U23189 (N_23189,N_22851,N_22953);
or U23190 (N_23190,N_22870,N_22954);
nor U23191 (N_23191,N_22923,N_22792);
xor U23192 (N_23192,N_22798,N_22837);
nand U23193 (N_23193,N_22857,N_22818);
nand U23194 (N_23194,N_22887,N_22837);
and U23195 (N_23195,N_22753,N_22788);
nand U23196 (N_23196,N_22891,N_22834);
or U23197 (N_23197,N_22937,N_22953);
nand U23198 (N_23198,N_22824,N_22836);
nor U23199 (N_23199,N_22780,N_22847);
or U23200 (N_23200,N_22801,N_22784);
nor U23201 (N_23201,N_22792,N_22837);
nor U23202 (N_23202,N_22804,N_22929);
nor U23203 (N_23203,N_22894,N_22810);
or U23204 (N_23204,N_22801,N_22803);
nor U23205 (N_23205,N_22912,N_22922);
or U23206 (N_23206,N_22801,N_22798);
or U23207 (N_23207,N_22912,N_22985);
nor U23208 (N_23208,N_22971,N_22864);
and U23209 (N_23209,N_22967,N_22973);
or U23210 (N_23210,N_22989,N_22903);
or U23211 (N_23211,N_22995,N_22851);
nand U23212 (N_23212,N_22822,N_22940);
or U23213 (N_23213,N_22938,N_22802);
and U23214 (N_23214,N_22846,N_22809);
xnor U23215 (N_23215,N_22846,N_22794);
xor U23216 (N_23216,N_22914,N_22942);
and U23217 (N_23217,N_22921,N_22867);
nand U23218 (N_23218,N_22921,N_22980);
or U23219 (N_23219,N_22775,N_22793);
or U23220 (N_23220,N_22980,N_22974);
nand U23221 (N_23221,N_22837,N_22803);
or U23222 (N_23222,N_22834,N_22947);
nand U23223 (N_23223,N_22993,N_22927);
nand U23224 (N_23224,N_22784,N_22816);
and U23225 (N_23225,N_22988,N_22932);
nand U23226 (N_23226,N_22840,N_22875);
nand U23227 (N_23227,N_22886,N_22772);
or U23228 (N_23228,N_22800,N_22929);
nor U23229 (N_23229,N_22864,N_22992);
xor U23230 (N_23230,N_22764,N_22827);
and U23231 (N_23231,N_22793,N_22984);
and U23232 (N_23232,N_22757,N_22891);
and U23233 (N_23233,N_22946,N_22842);
xor U23234 (N_23234,N_22828,N_22952);
xnor U23235 (N_23235,N_22940,N_22871);
xor U23236 (N_23236,N_22769,N_22814);
xor U23237 (N_23237,N_22768,N_22963);
and U23238 (N_23238,N_22812,N_22855);
and U23239 (N_23239,N_22935,N_22967);
xor U23240 (N_23240,N_22784,N_22807);
and U23241 (N_23241,N_22990,N_22794);
or U23242 (N_23242,N_22753,N_22949);
nand U23243 (N_23243,N_22770,N_22821);
xnor U23244 (N_23244,N_22928,N_22945);
xnor U23245 (N_23245,N_22865,N_22782);
xor U23246 (N_23246,N_22951,N_22804);
nand U23247 (N_23247,N_22898,N_22756);
nand U23248 (N_23248,N_22995,N_22762);
nand U23249 (N_23249,N_22862,N_22824);
and U23250 (N_23250,N_23248,N_23219);
and U23251 (N_23251,N_23040,N_23239);
or U23252 (N_23252,N_23203,N_23133);
xnor U23253 (N_23253,N_23052,N_23225);
and U23254 (N_23254,N_23087,N_23153);
or U23255 (N_23255,N_23078,N_23218);
or U23256 (N_23256,N_23084,N_23070);
nand U23257 (N_23257,N_23206,N_23011);
nand U23258 (N_23258,N_23034,N_23141);
xnor U23259 (N_23259,N_23193,N_23160);
or U23260 (N_23260,N_23191,N_23195);
nor U23261 (N_23261,N_23172,N_23100);
or U23262 (N_23262,N_23003,N_23107);
or U23263 (N_23263,N_23197,N_23104);
xnor U23264 (N_23264,N_23181,N_23146);
xnor U23265 (N_23265,N_23157,N_23132);
or U23266 (N_23266,N_23242,N_23091);
and U23267 (N_23267,N_23013,N_23051);
nor U23268 (N_23268,N_23101,N_23068);
xnor U23269 (N_23269,N_23001,N_23031);
nand U23270 (N_23270,N_23042,N_23230);
and U23271 (N_23271,N_23043,N_23095);
nor U23272 (N_23272,N_23135,N_23155);
nand U23273 (N_23273,N_23004,N_23148);
xor U23274 (N_23274,N_23074,N_23071);
xnor U23275 (N_23275,N_23030,N_23024);
or U23276 (N_23276,N_23093,N_23192);
nor U23277 (N_23277,N_23076,N_23238);
nand U23278 (N_23278,N_23039,N_23119);
nand U23279 (N_23279,N_23099,N_23180);
or U23280 (N_23280,N_23041,N_23054);
and U23281 (N_23281,N_23189,N_23023);
xnor U23282 (N_23282,N_23186,N_23077);
or U23283 (N_23283,N_23045,N_23014);
or U23284 (N_23284,N_23123,N_23231);
nand U23285 (N_23285,N_23171,N_23167);
and U23286 (N_23286,N_23179,N_23125);
xnor U23287 (N_23287,N_23130,N_23007);
or U23288 (N_23288,N_23235,N_23120);
xor U23289 (N_23289,N_23234,N_23246);
and U23290 (N_23290,N_23188,N_23217);
nor U23291 (N_23291,N_23223,N_23115);
and U23292 (N_23292,N_23144,N_23035);
or U23293 (N_23293,N_23128,N_23037);
and U23294 (N_23294,N_23194,N_23237);
xnor U23295 (N_23295,N_23117,N_23032);
xor U23296 (N_23296,N_23111,N_23010);
nor U23297 (N_23297,N_23081,N_23170);
and U23298 (N_23298,N_23088,N_23029);
nor U23299 (N_23299,N_23244,N_23102);
xnor U23300 (N_23300,N_23020,N_23106);
and U23301 (N_23301,N_23154,N_23116);
and U23302 (N_23302,N_23110,N_23137);
xnor U23303 (N_23303,N_23210,N_23075);
nor U23304 (N_23304,N_23065,N_23049);
or U23305 (N_23305,N_23131,N_23096);
or U23306 (N_23306,N_23226,N_23243);
nor U23307 (N_23307,N_23066,N_23190);
nand U23308 (N_23308,N_23050,N_23129);
and U23309 (N_23309,N_23176,N_23224);
nor U23310 (N_23310,N_23215,N_23016);
and U23311 (N_23311,N_23086,N_23134);
xor U23312 (N_23312,N_23000,N_23227);
and U23313 (N_23313,N_23199,N_23213);
nor U23314 (N_23314,N_23229,N_23178);
xnor U23315 (N_23315,N_23127,N_23205);
xnor U23316 (N_23316,N_23152,N_23187);
nand U23317 (N_23317,N_23162,N_23247);
and U23318 (N_23318,N_23151,N_23165);
nand U23319 (N_23319,N_23057,N_23241);
nand U23320 (N_23320,N_23103,N_23090);
nor U23321 (N_23321,N_23053,N_23038);
nor U23322 (N_23322,N_23113,N_23166);
or U23323 (N_23323,N_23009,N_23061);
or U23324 (N_23324,N_23184,N_23138);
nor U23325 (N_23325,N_23015,N_23198);
nor U23326 (N_23326,N_23121,N_23005);
and U23327 (N_23327,N_23240,N_23072);
or U23328 (N_23328,N_23019,N_23208);
nor U23329 (N_23329,N_23222,N_23126);
nor U23330 (N_23330,N_23025,N_23108);
xnor U23331 (N_23331,N_23082,N_23098);
or U23332 (N_23332,N_23056,N_23002);
xor U23333 (N_23333,N_23059,N_23036);
or U23334 (N_23334,N_23207,N_23033);
nand U23335 (N_23335,N_23149,N_23214);
xor U23336 (N_23336,N_23118,N_23028);
nand U23337 (N_23337,N_23147,N_23145);
nand U23338 (N_23338,N_23105,N_23047);
xnor U23339 (N_23339,N_23174,N_23067);
or U23340 (N_23340,N_23097,N_23008);
and U23341 (N_23341,N_23060,N_23046);
and U23342 (N_23342,N_23183,N_23201);
xnor U23343 (N_23343,N_23064,N_23169);
nor U23344 (N_23344,N_23143,N_23196);
xnor U23345 (N_23345,N_23221,N_23089);
or U23346 (N_23346,N_23021,N_23069);
nand U23347 (N_23347,N_23164,N_23124);
nand U23348 (N_23348,N_23185,N_23220);
xnor U23349 (N_23349,N_23112,N_23228);
nand U23350 (N_23350,N_23232,N_23158);
nand U23351 (N_23351,N_23245,N_23142);
nand U23352 (N_23352,N_23062,N_23236);
xor U23353 (N_23353,N_23017,N_23182);
xnor U23354 (N_23354,N_23048,N_23216);
nand U23355 (N_23355,N_23159,N_23055);
nand U23356 (N_23356,N_23202,N_23085);
and U23357 (N_23357,N_23211,N_23027);
nor U23358 (N_23358,N_23168,N_23079);
nor U23359 (N_23359,N_23204,N_23022);
nor U23360 (N_23360,N_23114,N_23163);
and U23361 (N_23361,N_23080,N_23139);
and U23362 (N_23362,N_23249,N_23233);
or U23363 (N_23363,N_23092,N_23200);
xnor U23364 (N_23364,N_23058,N_23150);
nor U23365 (N_23365,N_23212,N_23173);
and U23366 (N_23366,N_23161,N_23012);
nor U23367 (N_23367,N_23177,N_23006);
and U23368 (N_23368,N_23026,N_23140);
nor U23369 (N_23369,N_23044,N_23073);
and U23370 (N_23370,N_23109,N_23063);
xor U23371 (N_23371,N_23083,N_23018);
and U23372 (N_23372,N_23094,N_23209);
nor U23373 (N_23373,N_23156,N_23175);
or U23374 (N_23374,N_23122,N_23136);
nand U23375 (N_23375,N_23226,N_23233);
nand U23376 (N_23376,N_23106,N_23160);
and U23377 (N_23377,N_23080,N_23245);
or U23378 (N_23378,N_23166,N_23243);
nor U23379 (N_23379,N_23225,N_23211);
xor U23380 (N_23380,N_23119,N_23145);
xnor U23381 (N_23381,N_23087,N_23088);
nor U23382 (N_23382,N_23223,N_23140);
xor U23383 (N_23383,N_23162,N_23064);
xor U23384 (N_23384,N_23028,N_23057);
nor U23385 (N_23385,N_23208,N_23017);
nor U23386 (N_23386,N_23245,N_23163);
and U23387 (N_23387,N_23220,N_23161);
and U23388 (N_23388,N_23158,N_23034);
nand U23389 (N_23389,N_23114,N_23023);
nand U23390 (N_23390,N_23036,N_23020);
nor U23391 (N_23391,N_23241,N_23224);
or U23392 (N_23392,N_23222,N_23039);
nor U23393 (N_23393,N_23060,N_23246);
and U23394 (N_23394,N_23209,N_23247);
or U23395 (N_23395,N_23203,N_23105);
nand U23396 (N_23396,N_23068,N_23019);
nor U23397 (N_23397,N_23165,N_23157);
and U23398 (N_23398,N_23099,N_23166);
or U23399 (N_23399,N_23003,N_23246);
xnor U23400 (N_23400,N_23105,N_23197);
xor U23401 (N_23401,N_23105,N_23063);
xor U23402 (N_23402,N_23233,N_23216);
and U23403 (N_23403,N_23230,N_23185);
or U23404 (N_23404,N_23015,N_23111);
nor U23405 (N_23405,N_23130,N_23105);
xor U23406 (N_23406,N_23105,N_23091);
nor U23407 (N_23407,N_23070,N_23183);
and U23408 (N_23408,N_23224,N_23170);
xnor U23409 (N_23409,N_23105,N_23085);
and U23410 (N_23410,N_23193,N_23170);
and U23411 (N_23411,N_23049,N_23183);
or U23412 (N_23412,N_23117,N_23058);
nor U23413 (N_23413,N_23047,N_23002);
or U23414 (N_23414,N_23071,N_23042);
nand U23415 (N_23415,N_23157,N_23177);
or U23416 (N_23416,N_23103,N_23158);
and U23417 (N_23417,N_23216,N_23062);
and U23418 (N_23418,N_23090,N_23089);
nand U23419 (N_23419,N_23127,N_23230);
nor U23420 (N_23420,N_23169,N_23056);
and U23421 (N_23421,N_23207,N_23110);
xor U23422 (N_23422,N_23115,N_23090);
or U23423 (N_23423,N_23217,N_23102);
xor U23424 (N_23424,N_23165,N_23043);
or U23425 (N_23425,N_23029,N_23206);
nor U23426 (N_23426,N_23099,N_23122);
or U23427 (N_23427,N_23222,N_23228);
or U23428 (N_23428,N_23173,N_23144);
or U23429 (N_23429,N_23226,N_23140);
xor U23430 (N_23430,N_23227,N_23061);
or U23431 (N_23431,N_23185,N_23098);
nor U23432 (N_23432,N_23246,N_23215);
nand U23433 (N_23433,N_23068,N_23151);
or U23434 (N_23434,N_23105,N_23239);
and U23435 (N_23435,N_23006,N_23060);
nand U23436 (N_23436,N_23179,N_23219);
nand U23437 (N_23437,N_23033,N_23102);
or U23438 (N_23438,N_23067,N_23112);
or U23439 (N_23439,N_23109,N_23129);
xor U23440 (N_23440,N_23115,N_23067);
and U23441 (N_23441,N_23244,N_23128);
and U23442 (N_23442,N_23079,N_23107);
or U23443 (N_23443,N_23015,N_23040);
xnor U23444 (N_23444,N_23230,N_23195);
nand U23445 (N_23445,N_23006,N_23154);
nor U23446 (N_23446,N_23249,N_23172);
nor U23447 (N_23447,N_23242,N_23024);
nand U23448 (N_23448,N_23105,N_23078);
nand U23449 (N_23449,N_23118,N_23077);
or U23450 (N_23450,N_23149,N_23113);
and U23451 (N_23451,N_23202,N_23150);
nand U23452 (N_23452,N_23238,N_23103);
and U23453 (N_23453,N_23049,N_23002);
nand U23454 (N_23454,N_23000,N_23011);
and U23455 (N_23455,N_23072,N_23052);
xnor U23456 (N_23456,N_23069,N_23077);
or U23457 (N_23457,N_23239,N_23208);
nand U23458 (N_23458,N_23043,N_23020);
and U23459 (N_23459,N_23180,N_23177);
xor U23460 (N_23460,N_23064,N_23112);
nor U23461 (N_23461,N_23030,N_23035);
or U23462 (N_23462,N_23087,N_23197);
and U23463 (N_23463,N_23128,N_23044);
nand U23464 (N_23464,N_23201,N_23181);
nand U23465 (N_23465,N_23001,N_23215);
nor U23466 (N_23466,N_23109,N_23003);
xor U23467 (N_23467,N_23072,N_23234);
xnor U23468 (N_23468,N_23048,N_23113);
xor U23469 (N_23469,N_23132,N_23092);
and U23470 (N_23470,N_23153,N_23247);
and U23471 (N_23471,N_23074,N_23140);
nor U23472 (N_23472,N_23227,N_23220);
and U23473 (N_23473,N_23225,N_23040);
xor U23474 (N_23474,N_23084,N_23246);
nand U23475 (N_23475,N_23219,N_23236);
nand U23476 (N_23476,N_23225,N_23161);
nor U23477 (N_23477,N_23232,N_23206);
nand U23478 (N_23478,N_23062,N_23001);
nor U23479 (N_23479,N_23174,N_23180);
nor U23480 (N_23480,N_23091,N_23070);
xnor U23481 (N_23481,N_23154,N_23038);
and U23482 (N_23482,N_23170,N_23048);
xnor U23483 (N_23483,N_23063,N_23103);
nand U23484 (N_23484,N_23141,N_23037);
nand U23485 (N_23485,N_23044,N_23118);
and U23486 (N_23486,N_23123,N_23211);
xnor U23487 (N_23487,N_23141,N_23019);
or U23488 (N_23488,N_23058,N_23139);
nand U23489 (N_23489,N_23203,N_23233);
nand U23490 (N_23490,N_23036,N_23220);
xnor U23491 (N_23491,N_23167,N_23210);
and U23492 (N_23492,N_23175,N_23063);
and U23493 (N_23493,N_23015,N_23112);
xnor U23494 (N_23494,N_23115,N_23242);
and U23495 (N_23495,N_23008,N_23154);
nand U23496 (N_23496,N_23227,N_23036);
or U23497 (N_23497,N_23227,N_23221);
nor U23498 (N_23498,N_23189,N_23218);
xor U23499 (N_23499,N_23014,N_23077);
nand U23500 (N_23500,N_23353,N_23435);
xnor U23501 (N_23501,N_23325,N_23485);
nor U23502 (N_23502,N_23418,N_23257);
and U23503 (N_23503,N_23295,N_23357);
nand U23504 (N_23504,N_23327,N_23496);
or U23505 (N_23505,N_23271,N_23385);
xnor U23506 (N_23506,N_23263,N_23254);
and U23507 (N_23507,N_23494,N_23312);
and U23508 (N_23508,N_23472,N_23274);
nor U23509 (N_23509,N_23384,N_23448);
nand U23510 (N_23510,N_23365,N_23320);
nor U23511 (N_23511,N_23284,N_23341);
nor U23512 (N_23512,N_23497,N_23440);
xnor U23513 (N_23513,N_23446,N_23462);
and U23514 (N_23514,N_23316,N_23306);
nand U23515 (N_23515,N_23420,N_23300);
nand U23516 (N_23516,N_23350,N_23452);
xnor U23517 (N_23517,N_23348,N_23344);
and U23518 (N_23518,N_23484,N_23294);
nand U23519 (N_23519,N_23269,N_23398);
xor U23520 (N_23520,N_23467,N_23415);
or U23521 (N_23521,N_23260,N_23390);
and U23522 (N_23522,N_23423,N_23333);
or U23523 (N_23523,N_23493,N_23416);
and U23524 (N_23524,N_23377,N_23256);
and U23525 (N_23525,N_23335,N_23307);
or U23526 (N_23526,N_23308,N_23412);
xnor U23527 (N_23527,N_23417,N_23408);
and U23528 (N_23528,N_23310,N_23483);
nor U23529 (N_23529,N_23315,N_23439);
and U23530 (N_23530,N_23354,N_23381);
and U23531 (N_23531,N_23376,N_23424);
nand U23532 (N_23532,N_23375,N_23433);
and U23533 (N_23533,N_23279,N_23474);
nand U23534 (N_23534,N_23281,N_23373);
xor U23535 (N_23535,N_23414,N_23383);
xor U23536 (N_23536,N_23449,N_23473);
or U23537 (N_23537,N_23378,N_23461);
xor U23538 (N_23538,N_23498,N_23410);
and U23539 (N_23539,N_23282,N_23285);
nor U23540 (N_23540,N_23317,N_23386);
nor U23541 (N_23541,N_23491,N_23477);
nand U23542 (N_23542,N_23268,N_23459);
xor U23543 (N_23543,N_23426,N_23454);
and U23544 (N_23544,N_23468,N_23392);
nand U23545 (N_23545,N_23425,N_23442);
and U23546 (N_23546,N_23487,N_23379);
nor U23547 (N_23547,N_23321,N_23499);
or U23548 (N_23548,N_23463,N_23286);
or U23549 (N_23549,N_23305,N_23255);
nor U23550 (N_23550,N_23324,N_23358);
or U23551 (N_23551,N_23336,N_23331);
nand U23552 (N_23552,N_23409,N_23401);
and U23553 (N_23553,N_23298,N_23419);
nand U23554 (N_23554,N_23451,N_23251);
or U23555 (N_23555,N_23270,N_23480);
and U23556 (N_23556,N_23476,N_23301);
xor U23557 (N_23557,N_23492,N_23343);
nand U23558 (N_23558,N_23369,N_23431);
and U23559 (N_23559,N_23275,N_23465);
and U23560 (N_23560,N_23464,N_23391);
or U23561 (N_23561,N_23311,N_23290);
and U23562 (N_23562,N_23466,N_23323);
nor U23563 (N_23563,N_23266,N_23347);
or U23564 (N_23564,N_23460,N_23434);
nand U23565 (N_23565,N_23342,N_23261);
xor U23566 (N_23566,N_23368,N_23436);
xnor U23567 (N_23567,N_23297,N_23259);
nand U23568 (N_23568,N_23430,N_23389);
nand U23569 (N_23569,N_23490,N_23405);
nand U23570 (N_23570,N_23432,N_23455);
nor U23571 (N_23571,N_23394,N_23337);
nand U23572 (N_23572,N_23441,N_23252);
and U23573 (N_23573,N_23360,N_23338);
or U23574 (N_23574,N_23397,N_23296);
nand U23575 (N_23575,N_23422,N_23262);
or U23576 (N_23576,N_23356,N_23339);
and U23577 (N_23577,N_23469,N_23421);
or U23578 (N_23578,N_23402,N_23352);
or U23579 (N_23579,N_23444,N_23319);
nand U23580 (N_23580,N_23280,N_23453);
xnor U23581 (N_23581,N_23288,N_23488);
xnor U23582 (N_23582,N_23364,N_23314);
and U23583 (N_23583,N_23292,N_23359);
and U23584 (N_23584,N_23413,N_23481);
and U23585 (N_23585,N_23406,N_23486);
nand U23586 (N_23586,N_23318,N_23291);
xnor U23587 (N_23587,N_23407,N_23330);
or U23588 (N_23588,N_23471,N_23299);
and U23589 (N_23589,N_23277,N_23253);
or U23590 (N_23590,N_23276,N_23303);
or U23591 (N_23591,N_23404,N_23400);
nor U23592 (N_23592,N_23326,N_23478);
nor U23593 (N_23593,N_23267,N_23489);
nand U23594 (N_23594,N_23361,N_23445);
nand U23595 (N_23595,N_23427,N_23428);
or U23596 (N_23596,N_23447,N_23395);
and U23597 (N_23597,N_23374,N_23272);
and U23598 (N_23598,N_23495,N_23293);
xnor U23599 (N_23599,N_23362,N_23382);
xnor U23600 (N_23600,N_23351,N_23370);
xnor U23601 (N_23601,N_23429,N_23443);
nor U23602 (N_23602,N_23399,N_23329);
and U23603 (N_23603,N_23363,N_23265);
and U23604 (N_23604,N_23393,N_23264);
nor U23605 (N_23605,N_23283,N_23278);
and U23606 (N_23606,N_23345,N_23340);
or U23607 (N_23607,N_23387,N_23457);
or U23608 (N_23608,N_23437,N_23302);
xnor U23609 (N_23609,N_23289,N_23380);
or U23610 (N_23610,N_23479,N_23328);
nor U23611 (N_23611,N_23388,N_23438);
nand U23612 (N_23612,N_23456,N_23372);
nor U23613 (N_23613,N_23304,N_23313);
and U23614 (N_23614,N_23273,N_23458);
xnor U23615 (N_23615,N_23366,N_23475);
xnor U23616 (N_23616,N_23309,N_23470);
nand U23617 (N_23617,N_23411,N_23396);
xnor U23618 (N_23618,N_23367,N_23450);
nand U23619 (N_23619,N_23258,N_23287);
nor U23620 (N_23620,N_23334,N_23332);
and U23621 (N_23621,N_23346,N_23349);
xnor U23622 (N_23622,N_23250,N_23403);
nor U23623 (N_23623,N_23322,N_23371);
nand U23624 (N_23624,N_23355,N_23482);
nor U23625 (N_23625,N_23434,N_23376);
and U23626 (N_23626,N_23467,N_23253);
nor U23627 (N_23627,N_23267,N_23427);
or U23628 (N_23628,N_23293,N_23364);
xor U23629 (N_23629,N_23364,N_23348);
nor U23630 (N_23630,N_23394,N_23251);
xor U23631 (N_23631,N_23395,N_23427);
nor U23632 (N_23632,N_23257,N_23298);
and U23633 (N_23633,N_23336,N_23391);
nor U23634 (N_23634,N_23373,N_23260);
or U23635 (N_23635,N_23476,N_23408);
and U23636 (N_23636,N_23390,N_23333);
xor U23637 (N_23637,N_23369,N_23335);
or U23638 (N_23638,N_23379,N_23303);
or U23639 (N_23639,N_23368,N_23461);
and U23640 (N_23640,N_23290,N_23476);
xnor U23641 (N_23641,N_23425,N_23291);
or U23642 (N_23642,N_23263,N_23431);
xor U23643 (N_23643,N_23454,N_23373);
or U23644 (N_23644,N_23313,N_23468);
nand U23645 (N_23645,N_23372,N_23254);
nor U23646 (N_23646,N_23275,N_23452);
or U23647 (N_23647,N_23251,N_23414);
and U23648 (N_23648,N_23481,N_23335);
or U23649 (N_23649,N_23417,N_23490);
xnor U23650 (N_23650,N_23357,N_23420);
and U23651 (N_23651,N_23448,N_23303);
nor U23652 (N_23652,N_23431,N_23371);
nor U23653 (N_23653,N_23253,N_23278);
and U23654 (N_23654,N_23434,N_23262);
xor U23655 (N_23655,N_23354,N_23463);
nand U23656 (N_23656,N_23305,N_23262);
and U23657 (N_23657,N_23419,N_23478);
xor U23658 (N_23658,N_23363,N_23372);
nor U23659 (N_23659,N_23483,N_23498);
or U23660 (N_23660,N_23388,N_23366);
or U23661 (N_23661,N_23329,N_23380);
nor U23662 (N_23662,N_23493,N_23490);
nand U23663 (N_23663,N_23297,N_23461);
xnor U23664 (N_23664,N_23435,N_23393);
and U23665 (N_23665,N_23378,N_23262);
or U23666 (N_23666,N_23341,N_23447);
nand U23667 (N_23667,N_23479,N_23376);
xor U23668 (N_23668,N_23345,N_23395);
nand U23669 (N_23669,N_23357,N_23392);
or U23670 (N_23670,N_23367,N_23421);
nor U23671 (N_23671,N_23449,N_23261);
nor U23672 (N_23672,N_23436,N_23435);
and U23673 (N_23673,N_23303,N_23362);
xnor U23674 (N_23674,N_23349,N_23302);
nand U23675 (N_23675,N_23340,N_23265);
or U23676 (N_23676,N_23405,N_23489);
or U23677 (N_23677,N_23400,N_23328);
xor U23678 (N_23678,N_23496,N_23301);
and U23679 (N_23679,N_23425,N_23337);
and U23680 (N_23680,N_23264,N_23453);
nand U23681 (N_23681,N_23479,N_23453);
nand U23682 (N_23682,N_23398,N_23334);
xor U23683 (N_23683,N_23339,N_23365);
xor U23684 (N_23684,N_23353,N_23442);
and U23685 (N_23685,N_23497,N_23270);
nor U23686 (N_23686,N_23383,N_23432);
nand U23687 (N_23687,N_23346,N_23375);
xnor U23688 (N_23688,N_23445,N_23264);
or U23689 (N_23689,N_23473,N_23391);
and U23690 (N_23690,N_23472,N_23466);
or U23691 (N_23691,N_23308,N_23465);
and U23692 (N_23692,N_23304,N_23328);
nor U23693 (N_23693,N_23315,N_23370);
or U23694 (N_23694,N_23471,N_23286);
xor U23695 (N_23695,N_23319,N_23258);
nand U23696 (N_23696,N_23467,N_23449);
nor U23697 (N_23697,N_23493,N_23290);
nand U23698 (N_23698,N_23296,N_23408);
xnor U23699 (N_23699,N_23299,N_23369);
xnor U23700 (N_23700,N_23281,N_23447);
nand U23701 (N_23701,N_23385,N_23261);
nand U23702 (N_23702,N_23286,N_23343);
and U23703 (N_23703,N_23300,N_23392);
nor U23704 (N_23704,N_23302,N_23370);
or U23705 (N_23705,N_23377,N_23476);
nor U23706 (N_23706,N_23338,N_23306);
nor U23707 (N_23707,N_23377,N_23463);
or U23708 (N_23708,N_23300,N_23277);
and U23709 (N_23709,N_23328,N_23472);
and U23710 (N_23710,N_23484,N_23476);
or U23711 (N_23711,N_23468,N_23338);
nor U23712 (N_23712,N_23471,N_23291);
nand U23713 (N_23713,N_23454,N_23462);
nor U23714 (N_23714,N_23487,N_23391);
xor U23715 (N_23715,N_23454,N_23482);
nor U23716 (N_23716,N_23276,N_23269);
and U23717 (N_23717,N_23285,N_23395);
or U23718 (N_23718,N_23352,N_23279);
nor U23719 (N_23719,N_23333,N_23426);
xor U23720 (N_23720,N_23394,N_23482);
xor U23721 (N_23721,N_23486,N_23443);
nand U23722 (N_23722,N_23285,N_23308);
xnor U23723 (N_23723,N_23410,N_23290);
and U23724 (N_23724,N_23259,N_23294);
nor U23725 (N_23725,N_23291,N_23458);
xor U23726 (N_23726,N_23417,N_23445);
nand U23727 (N_23727,N_23495,N_23454);
xnor U23728 (N_23728,N_23446,N_23368);
nand U23729 (N_23729,N_23469,N_23442);
nor U23730 (N_23730,N_23379,N_23389);
or U23731 (N_23731,N_23271,N_23427);
or U23732 (N_23732,N_23424,N_23428);
nand U23733 (N_23733,N_23480,N_23372);
nor U23734 (N_23734,N_23299,N_23446);
nor U23735 (N_23735,N_23442,N_23373);
xor U23736 (N_23736,N_23365,N_23314);
nor U23737 (N_23737,N_23328,N_23404);
xor U23738 (N_23738,N_23379,N_23283);
xnor U23739 (N_23739,N_23386,N_23293);
or U23740 (N_23740,N_23495,N_23476);
or U23741 (N_23741,N_23313,N_23325);
or U23742 (N_23742,N_23362,N_23322);
and U23743 (N_23743,N_23325,N_23258);
nand U23744 (N_23744,N_23304,N_23262);
xnor U23745 (N_23745,N_23434,N_23302);
nand U23746 (N_23746,N_23363,N_23395);
and U23747 (N_23747,N_23418,N_23324);
nor U23748 (N_23748,N_23350,N_23274);
xor U23749 (N_23749,N_23469,N_23322);
or U23750 (N_23750,N_23542,N_23539);
xor U23751 (N_23751,N_23722,N_23674);
or U23752 (N_23752,N_23587,N_23579);
and U23753 (N_23753,N_23585,N_23618);
xnor U23754 (N_23754,N_23724,N_23550);
nor U23755 (N_23755,N_23526,N_23682);
nand U23756 (N_23756,N_23732,N_23507);
nor U23757 (N_23757,N_23731,N_23648);
xor U23758 (N_23758,N_23535,N_23555);
and U23759 (N_23759,N_23537,N_23503);
and U23760 (N_23760,N_23687,N_23529);
or U23761 (N_23761,N_23611,N_23684);
xor U23762 (N_23762,N_23737,N_23521);
and U23763 (N_23763,N_23530,N_23720);
nand U23764 (N_23764,N_23663,N_23635);
or U23765 (N_23765,N_23748,N_23514);
nand U23766 (N_23766,N_23691,N_23698);
xor U23767 (N_23767,N_23733,N_23543);
or U23768 (N_23768,N_23651,N_23710);
nor U23769 (N_23769,N_23627,N_23566);
nand U23770 (N_23770,N_23511,N_23633);
xnor U23771 (N_23771,N_23728,N_23622);
nor U23772 (N_23772,N_23640,N_23573);
and U23773 (N_23773,N_23654,N_23671);
nand U23774 (N_23774,N_23666,N_23726);
nor U23775 (N_23775,N_23609,N_23644);
xor U23776 (N_23776,N_23569,N_23749);
and U23777 (N_23777,N_23615,N_23559);
nand U23778 (N_23778,N_23567,N_23689);
nand U23779 (N_23779,N_23592,N_23641);
and U23780 (N_23780,N_23591,N_23590);
nor U23781 (N_23781,N_23582,N_23548);
xor U23782 (N_23782,N_23516,N_23744);
nor U23783 (N_23783,N_23716,N_23533);
nor U23784 (N_23784,N_23594,N_23531);
or U23785 (N_23785,N_23557,N_23700);
nand U23786 (N_23786,N_23601,N_23626);
and U23787 (N_23787,N_23576,N_23606);
nor U23788 (N_23788,N_23603,N_23657);
or U23789 (N_23789,N_23632,N_23586);
and U23790 (N_23790,N_23580,N_23670);
and U23791 (N_23791,N_23525,N_23646);
xor U23792 (N_23792,N_23575,N_23678);
and U23793 (N_23793,N_23605,N_23638);
nor U23794 (N_23794,N_23604,N_23549);
or U23795 (N_23795,N_23669,N_23699);
nor U23796 (N_23796,N_23520,N_23683);
or U23797 (N_23797,N_23564,N_23508);
xnor U23798 (N_23798,N_23563,N_23560);
nand U23799 (N_23799,N_23527,N_23505);
nand U23800 (N_23800,N_23739,N_23708);
or U23801 (N_23801,N_23634,N_23561);
and U23802 (N_23802,N_23659,N_23509);
xor U23803 (N_23803,N_23617,N_23676);
nand U23804 (N_23804,N_23723,N_23562);
or U23805 (N_23805,N_23593,N_23730);
nand U23806 (N_23806,N_23702,N_23705);
xnor U23807 (N_23807,N_23544,N_23725);
and U23808 (N_23808,N_23554,N_23685);
xnor U23809 (N_23809,N_23668,N_23565);
and U23810 (N_23810,N_23616,N_23571);
or U23811 (N_23811,N_23652,N_23597);
or U23812 (N_23812,N_23660,N_23680);
or U23813 (N_23813,N_23665,N_23653);
nand U23814 (N_23814,N_23707,N_23679);
xnor U23815 (N_23815,N_23642,N_23552);
and U23816 (N_23816,N_23528,N_23701);
or U23817 (N_23817,N_23620,N_23574);
nor U23818 (N_23818,N_23709,N_23675);
nor U23819 (N_23819,N_23547,N_23532);
or U23820 (N_23820,N_23712,N_23519);
or U23821 (N_23821,N_23694,N_23696);
nand U23822 (N_23822,N_23501,N_23738);
xor U23823 (N_23823,N_23740,N_23599);
xnor U23824 (N_23824,N_23686,N_23515);
nand U23825 (N_23825,N_23643,N_23637);
nor U23826 (N_23826,N_23598,N_23607);
and U23827 (N_23827,N_23504,N_23719);
nand U23828 (N_23828,N_23538,N_23625);
xor U23829 (N_23829,N_23619,N_23545);
nor U23830 (N_23830,N_23714,N_23517);
or U23831 (N_23831,N_23672,N_23711);
and U23832 (N_23832,N_23647,N_23715);
or U23833 (N_23833,N_23650,N_23572);
and U23834 (N_23834,N_23513,N_23727);
nor U23835 (N_23835,N_23613,N_23596);
nand U23836 (N_23836,N_23584,N_23681);
or U23837 (N_23837,N_23631,N_23536);
nor U23838 (N_23838,N_23630,N_23692);
nand U23839 (N_23839,N_23600,N_23661);
xor U23840 (N_23840,N_23610,N_23645);
nand U23841 (N_23841,N_23614,N_23734);
and U23842 (N_23842,N_23746,N_23583);
and U23843 (N_23843,N_23697,N_23664);
and U23844 (N_23844,N_23735,N_23589);
nand U23845 (N_23845,N_23729,N_23690);
nand U23846 (N_23846,N_23717,N_23523);
xor U23847 (N_23847,N_23656,N_23551);
or U23848 (N_23848,N_23741,N_23518);
and U23849 (N_23849,N_23706,N_23742);
xnor U23850 (N_23850,N_23695,N_23506);
or U23851 (N_23851,N_23568,N_23556);
or U23852 (N_23852,N_23688,N_23721);
and U23853 (N_23853,N_23588,N_23524);
and U23854 (N_23854,N_23534,N_23718);
and U23855 (N_23855,N_23655,N_23540);
or U23856 (N_23856,N_23595,N_23636);
xnor U23857 (N_23857,N_23747,N_23581);
nand U23858 (N_23858,N_23608,N_23673);
nand U23859 (N_23859,N_23745,N_23704);
or U23860 (N_23860,N_23577,N_23623);
nor U23861 (N_23861,N_23624,N_23500);
and U23862 (N_23862,N_23522,N_23649);
and U23863 (N_23863,N_23602,N_23510);
nand U23864 (N_23864,N_23621,N_23677);
nand U23865 (N_23865,N_23667,N_23553);
nor U23866 (N_23866,N_23570,N_23662);
nand U23867 (N_23867,N_23546,N_23628);
nor U23868 (N_23868,N_23736,N_23578);
nand U23869 (N_23869,N_23703,N_23612);
nand U23870 (N_23870,N_23512,N_23693);
or U23871 (N_23871,N_23541,N_23558);
and U23872 (N_23872,N_23713,N_23629);
or U23873 (N_23873,N_23658,N_23743);
xnor U23874 (N_23874,N_23639,N_23502);
nand U23875 (N_23875,N_23504,N_23741);
and U23876 (N_23876,N_23680,N_23729);
nor U23877 (N_23877,N_23698,N_23670);
and U23878 (N_23878,N_23591,N_23536);
xor U23879 (N_23879,N_23522,N_23571);
nand U23880 (N_23880,N_23603,N_23722);
or U23881 (N_23881,N_23535,N_23533);
nand U23882 (N_23882,N_23710,N_23723);
and U23883 (N_23883,N_23604,N_23670);
nand U23884 (N_23884,N_23533,N_23630);
nor U23885 (N_23885,N_23638,N_23542);
and U23886 (N_23886,N_23588,N_23591);
nand U23887 (N_23887,N_23650,N_23516);
nand U23888 (N_23888,N_23739,N_23702);
and U23889 (N_23889,N_23563,N_23564);
or U23890 (N_23890,N_23704,N_23566);
or U23891 (N_23891,N_23545,N_23596);
and U23892 (N_23892,N_23513,N_23692);
or U23893 (N_23893,N_23630,N_23535);
and U23894 (N_23894,N_23515,N_23584);
nor U23895 (N_23895,N_23569,N_23747);
or U23896 (N_23896,N_23564,N_23510);
and U23897 (N_23897,N_23551,N_23616);
nand U23898 (N_23898,N_23673,N_23719);
xnor U23899 (N_23899,N_23568,N_23704);
nand U23900 (N_23900,N_23514,N_23631);
xor U23901 (N_23901,N_23627,N_23601);
or U23902 (N_23902,N_23519,N_23534);
nor U23903 (N_23903,N_23724,N_23504);
nor U23904 (N_23904,N_23607,N_23597);
or U23905 (N_23905,N_23721,N_23572);
and U23906 (N_23906,N_23564,N_23704);
nand U23907 (N_23907,N_23514,N_23664);
or U23908 (N_23908,N_23644,N_23550);
nor U23909 (N_23909,N_23558,N_23733);
xor U23910 (N_23910,N_23691,N_23600);
and U23911 (N_23911,N_23647,N_23680);
nor U23912 (N_23912,N_23717,N_23707);
nor U23913 (N_23913,N_23507,N_23561);
and U23914 (N_23914,N_23711,N_23731);
or U23915 (N_23915,N_23664,N_23708);
or U23916 (N_23916,N_23579,N_23703);
xnor U23917 (N_23917,N_23635,N_23696);
or U23918 (N_23918,N_23611,N_23680);
nor U23919 (N_23919,N_23569,N_23718);
nor U23920 (N_23920,N_23514,N_23707);
xor U23921 (N_23921,N_23575,N_23662);
nand U23922 (N_23922,N_23741,N_23555);
xnor U23923 (N_23923,N_23617,N_23537);
and U23924 (N_23924,N_23665,N_23510);
nor U23925 (N_23925,N_23539,N_23723);
xor U23926 (N_23926,N_23695,N_23705);
nand U23927 (N_23927,N_23537,N_23507);
nand U23928 (N_23928,N_23680,N_23556);
nand U23929 (N_23929,N_23627,N_23550);
and U23930 (N_23930,N_23651,N_23655);
and U23931 (N_23931,N_23625,N_23628);
nor U23932 (N_23932,N_23625,N_23640);
and U23933 (N_23933,N_23544,N_23650);
or U23934 (N_23934,N_23725,N_23668);
nand U23935 (N_23935,N_23576,N_23588);
and U23936 (N_23936,N_23645,N_23591);
nand U23937 (N_23937,N_23731,N_23622);
xnor U23938 (N_23938,N_23651,N_23725);
and U23939 (N_23939,N_23710,N_23620);
nor U23940 (N_23940,N_23735,N_23591);
nor U23941 (N_23941,N_23530,N_23712);
xnor U23942 (N_23942,N_23508,N_23551);
or U23943 (N_23943,N_23669,N_23697);
nand U23944 (N_23944,N_23543,N_23514);
nor U23945 (N_23945,N_23676,N_23615);
nand U23946 (N_23946,N_23571,N_23647);
nand U23947 (N_23947,N_23657,N_23718);
and U23948 (N_23948,N_23544,N_23559);
xnor U23949 (N_23949,N_23560,N_23546);
and U23950 (N_23950,N_23705,N_23544);
or U23951 (N_23951,N_23674,N_23662);
and U23952 (N_23952,N_23733,N_23678);
xor U23953 (N_23953,N_23633,N_23572);
and U23954 (N_23954,N_23543,N_23745);
and U23955 (N_23955,N_23580,N_23512);
xor U23956 (N_23956,N_23735,N_23678);
nor U23957 (N_23957,N_23601,N_23693);
and U23958 (N_23958,N_23522,N_23739);
nand U23959 (N_23959,N_23632,N_23549);
nand U23960 (N_23960,N_23748,N_23659);
nand U23961 (N_23961,N_23708,N_23524);
nand U23962 (N_23962,N_23552,N_23583);
nor U23963 (N_23963,N_23556,N_23551);
xnor U23964 (N_23964,N_23707,N_23537);
xor U23965 (N_23965,N_23723,N_23606);
nand U23966 (N_23966,N_23535,N_23506);
nand U23967 (N_23967,N_23631,N_23723);
and U23968 (N_23968,N_23608,N_23612);
and U23969 (N_23969,N_23635,N_23697);
nor U23970 (N_23970,N_23597,N_23727);
nand U23971 (N_23971,N_23685,N_23578);
nor U23972 (N_23972,N_23523,N_23519);
xnor U23973 (N_23973,N_23603,N_23579);
nor U23974 (N_23974,N_23704,N_23654);
nor U23975 (N_23975,N_23559,N_23517);
nand U23976 (N_23976,N_23695,N_23710);
nor U23977 (N_23977,N_23592,N_23591);
xnor U23978 (N_23978,N_23744,N_23528);
xor U23979 (N_23979,N_23582,N_23745);
or U23980 (N_23980,N_23671,N_23658);
and U23981 (N_23981,N_23515,N_23536);
nor U23982 (N_23982,N_23611,N_23621);
and U23983 (N_23983,N_23639,N_23541);
nand U23984 (N_23984,N_23654,N_23582);
and U23985 (N_23985,N_23717,N_23654);
xor U23986 (N_23986,N_23609,N_23721);
xnor U23987 (N_23987,N_23723,N_23517);
xor U23988 (N_23988,N_23695,N_23577);
xor U23989 (N_23989,N_23588,N_23607);
or U23990 (N_23990,N_23576,N_23693);
and U23991 (N_23991,N_23675,N_23614);
nor U23992 (N_23992,N_23575,N_23723);
nand U23993 (N_23993,N_23582,N_23518);
or U23994 (N_23994,N_23591,N_23616);
nand U23995 (N_23995,N_23611,N_23528);
and U23996 (N_23996,N_23599,N_23682);
and U23997 (N_23997,N_23576,N_23522);
xnor U23998 (N_23998,N_23723,N_23648);
nor U23999 (N_23999,N_23739,N_23527);
xnor U24000 (N_24000,N_23882,N_23953);
xor U24001 (N_24001,N_23920,N_23894);
and U24002 (N_24002,N_23842,N_23936);
nor U24003 (N_24003,N_23965,N_23957);
xnor U24004 (N_24004,N_23787,N_23901);
xnor U24005 (N_24005,N_23841,N_23849);
nand U24006 (N_24006,N_23866,N_23796);
nor U24007 (N_24007,N_23880,N_23898);
xnor U24008 (N_24008,N_23973,N_23977);
and U24009 (N_24009,N_23919,N_23835);
nand U24010 (N_24010,N_23889,N_23838);
or U24011 (N_24011,N_23869,N_23964);
nand U24012 (N_24012,N_23840,N_23998);
xor U24013 (N_24013,N_23860,N_23981);
or U24014 (N_24014,N_23829,N_23974);
nand U24015 (N_24015,N_23803,N_23984);
xor U24016 (N_24016,N_23764,N_23966);
xor U24017 (N_24017,N_23995,N_23868);
and U24018 (N_24018,N_23954,N_23963);
and U24019 (N_24019,N_23767,N_23935);
nor U24020 (N_24020,N_23997,N_23991);
and U24021 (N_24021,N_23846,N_23900);
or U24022 (N_24022,N_23861,N_23929);
and U24023 (N_24023,N_23763,N_23969);
nor U24024 (N_24024,N_23923,N_23948);
xor U24025 (N_24025,N_23859,N_23983);
nor U24026 (N_24026,N_23958,N_23876);
nor U24027 (N_24027,N_23950,N_23875);
and U24028 (N_24028,N_23924,N_23938);
nor U24029 (N_24029,N_23857,N_23886);
and U24030 (N_24030,N_23858,N_23789);
nor U24031 (N_24031,N_23933,N_23776);
nor U24032 (N_24032,N_23854,N_23961);
nor U24033 (N_24033,N_23828,N_23794);
xor U24034 (N_24034,N_23836,N_23947);
nor U24035 (N_24035,N_23783,N_23941);
nor U24036 (N_24036,N_23939,N_23815);
nor U24037 (N_24037,N_23890,N_23891);
nand U24038 (N_24038,N_23855,N_23791);
nand U24039 (N_24039,N_23906,N_23999);
and U24040 (N_24040,N_23937,N_23967);
or U24041 (N_24041,N_23959,N_23793);
nand U24042 (N_24042,N_23864,N_23996);
or U24043 (N_24043,N_23975,N_23774);
nand U24044 (N_24044,N_23952,N_23820);
nor U24045 (N_24045,N_23930,N_23863);
xor U24046 (N_24046,N_23872,N_23773);
or U24047 (N_24047,N_23750,N_23944);
nand U24048 (N_24048,N_23985,N_23878);
nand U24049 (N_24049,N_23852,N_23755);
xnor U24050 (N_24050,N_23951,N_23892);
and U24051 (N_24051,N_23801,N_23753);
nor U24052 (N_24052,N_23910,N_23831);
nand U24053 (N_24053,N_23927,N_23798);
and U24054 (N_24054,N_23867,N_23821);
nand U24055 (N_24055,N_23819,N_23897);
or U24056 (N_24056,N_23822,N_23968);
or U24057 (N_24057,N_23888,N_23816);
nor U24058 (N_24058,N_23777,N_23833);
and U24059 (N_24059,N_23848,N_23903);
and U24060 (N_24060,N_23885,N_23802);
nand U24061 (N_24061,N_23871,N_23782);
and U24062 (N_24062,N_23754,N_23909);
and U24063 (N_24063,N_23980,N_23806);
and U24064 (N_24064,N_23870,N_23853);
nand U24065 (N_24065,N_23904,N_23818);
or U24066 (N_24066,N_23786,N_23770);
or U24067 (N_24067,N_23865,N_23810);
nor U24068 (N_24068,N_23784,N_23812);
nor U24069 (N_24069,N_23759,N_23987);
nand U24070 (N_24070,N_23771,N_23887);
and U24071 (N_24071,N_23814,N_23788);
nand U24072 (N_24072,N_23979,N_23781);
nor U24073 (N_24073,N_23914,N_23839);
or U24074 (N_24074,N_23921,N_23907);
or U24075 (N_24075,N_23895,N_23752);
nand U24076 (N_24076,N_23922,N_23766);
and U24077 (N_24077,N_23873,N_23915);
and U24078 (N_24078,N_23837,N_23757);
nand U24079 (N_24079,N_23808,N_23785);
or U24080 (N_24080,N_23960,N_23879);
and U24081 (N_24081,N_23918,N_23826);
nor U24082 (N_24082,N_23772,N_23899);
nand U24083 (N_24083,N_23908,N_23809);
nand U24084 (N_24084,N_23912,N_23971);
nor U24085 (N_24085,N_23905,N_23989);
or U24086 (N_24086,N_23994,N_23986);
xnor U24087 (N_24087,N_23990,N_23790);
xor U24088 (N_24088,N_23807,N_23955);
or U24089 (N_24089,N_23825,N_23800);
or U24090 (N_24090,N_23845,N_23769);
xor U24091 (N_24091,N_23843,N_23847);
or U24092 (N_24092,N_23926,N_23928);
or U24093 (N_24093,N_23834,N_23943);
xnor U24094 (N_24094,N_23942,N_23805);
xor U24095 (N_24095,N_23881,N_23976);
nand U24096 (N_24096,N_23856,N_23775);
nor U24097 (N_24097,N_23893,N_23902);
xnor U24098 (N_24098,N_23940,N_23811);
nand U24099 (N_24099,N_23911,N_23884);
nor U24100 (N_24100,N_23925,N_23945);
xnor U24101 (N_24101,N_23962,N_23896);
nor U24102 (N_24102,N_23844,N_23832);
xnor U24103 (N_24103,N_23992,N_23751);
nor U24104 (N_24104,N_23804,N_23792);
nor U24105 (N_24105,N_23913,N_23768);
nor U24106 (N_24106,N_23949,N_23779);
or U24107 (N_24107,N_23883,N_23917);
nor U24108 (N_24108,N_23824,N_23931);
and U24109 (N_24109,N_23813,N_23874);
or U24110 (N_24110,N_23982,N_23795);
nand U24111 (N_24111,N_23916,N_23850);
and U24112 (N_24112,N_23823,N_23765);
nor U24113 (N_24113,N_23956,N_23988);
xnor U24114 (N_24114,N_23827,N_23761);
nand U24115 (N_24115,N_23830,N_23934);
xor U24116 (N_24116,N_23932,N_23972);
nand U24117 (N_24117,N_23799,N_23797);
and U24118 (N_24118,N_23758,N_23817);
xnor U24119 (N_24119,N_23970,N_23862);
nor U24120 (N_24120,N_23778,N_23756);
or U24121 (N_24121,N_23993,N_23946);
and U24122 (N_24122,N_23780,N_23851);
xnor U24123 (N_24123,N_23762,N_23978);
or U24124 (N_24124,N_23877,N_23760);
nand U24125 (N_24125,N_23754,N_23971);
and U24126 (N_24126,N_23838,N_23971);
nand U24127 (N_24127,N_23918,N_23879);
nand U24128 (N_24128,N_23822,N_23764);
nand U24129 (N_24129,N_23767,N_23950);
nor U24130 (N_24130,N_23971,N_23995);
xor U24131 (N_24131,N_23973,N_23905);
nand U24132 (N_24132,N_23913,N_23952);
xor U24133 (N_24133,N_23989,N_23841);
or U24134 (N_24134,N_23908,N_23808);
nand U24135 (N_24135,N_23978,N_23754);
nor U24136 (N_24136,N_23899,N_23988);
or U24137 (N_24137,N_23853,N_23759);
xor U24138 (N_24138,N_23790,N_23785);
and U24139 (N_24139,N_23883,N_23798);
nand U24140 (N_24140,N_23911,N_23967);
nor U24141 (N_24141,N_23865,N_23760);
nand U24142 (N_24142,N_23870,N_23817);
nor U24143 (N_24143,N_23850,N_23889);
nor U24144 (N_24144,N_23917,N_23802);
and U24145 (N_24145,N_23755,N_23783);
and U24146 (N_24146,N_23758,N_23860);
nand U24147 (N_24147,N_23800,N_23762);
and U24148 (N_24148,N_23806,N_23833);
or U24149 (N_24149,N_23880,N_23995);
or U24150 (N_24150,N_23954,N_23796);
nand U24151 (N_24151,N_23819,N_23863);
nand U24152 (N_24152,N_23765,N_23857);
and U24153 (N_24153,N_23814,N_23891);
and U24154 (N_24154,N_23800,N_23873);
or U24155 (N_24155,N_23975,N_23968);
nand U24156 (N_24156,N_23942,N_23878);
nor U24157 (N_24157,N_23830,N_23832);
and U24158 (N_24158,N_23854,N_23919);
and U24159 (N_24159,N_23882,N_23836);
and U24160 (N_24160,N_23807,N_23780);
nor U24161 (N_24161,N_23862,N_23972);
xor U24162 (N_24162,N_23902,N_23775);
nand U24163 (N_24163,N_23755,N_23932);
nand U24164 (N_24164,N_23854,N_23849);
or U24165 (N_24165,N_23851,N_23836);
nor U24166 (N_24166,N_23942,N_23840);
nor U24167 (N_24167,N_23852,N_23827);
nor U24168 (N_24168,N_23752,N_23904);
xor U24169 (N_24169,N_23786,N_23798);
xnor U24170 (N_24170,N_23922,N_23760);
xnor U24171 (N_24171,N_23986,N_23764);
nor U24172 (N_24172,N_23879,N_23965);
xnor U24173 (N_24173,N_23970,N_23939);
xor U24174 (N_24174,N_23830,N_23955);
or U24175 (N_24175,N_23913,N_23757);
xnor U24176 (N_24176,N_23758,N_23857);
nand U24177 (N_24177,N_23966,N_23940);
nand U24178 (N_24178,N_23819,N_23888);
nand U24179 (N_24179,N_23938,N_23987);
and U24180 (N_24180,N_23884,N_23951);
or U24181 (N_24181,N_23899,N_23824);
nor U24182 (N_24182,N_23918,N_23843);
and U24183 (N_24183,N_23884,N_23996);
nand U24184 (N_24184,N_23900,N_23758);
or U24185 (N_24185,N_23894,N_23823);
nand U24186 (N_24186,N_23784,N_23845);
nand U24187 (N_24187,N_23786,N_23808);
xnor U24188 (N_24188,N_23884,N_23802);
nand U24189 (N_24189,N_23950,N_23858);
nand U24190 (N_24190,N_23981,N_23891);
and U24191 (N_24191,N_23803,N_23795);
xor U24192 (N_24192,N_23754,N_23774);
or U24193 (N_24193,N_23899,N_23774);
nor U24194 (N_24194,N_23904,N_23833);
and U24195 (N_24195,N_23870,N_23751);
xor U24196 (N_24196,N_23956,N_23955);
nand U24197 (N_24197,N_23986,N_23850);
xnor U24198 (N_24198,N_23908,N_23889);
nor U24199 (N_24199,N_23806,N_23908);
nand U24200 (N_24200,N_23998,N_23977);
or U24201 (N_24201,N_23912,N_23909);
or U24202 (N_24202,N_23797,N_23843);
nand U24203 (N_24203,N_23947,N_23986);
and U24204 (N_24204,N_23943,N_23798);
and U24205 (N_24205,N_23923,N_23844);
nand U24206 (N_24206,N_23988,N_23891);
xor U24207 (N_24207,N_23879,N_23771);
nor U24208 (N_24208,N_23854,N_23754);
and U24209 (N_24209,N_23823,N_23811);
nand U24210 (N_24210,N_23853,N_23920);
nand U24211 (N_24211,N_23866,N_23800);
and U24212 (N_24212,N_23776,N_23764);
nand U24213 (N_24213,N_23856,N_23822);
nand U24214 (N_24214,N_23758,N_23806);
nor U24215 (N_24215,N_23759,N_23850);
nand U24216 (N_24216,N_23998,N_23994);
xor U24217 (N_24217,N_23791,N_23777);
nand U24218 (N_24218,N_23823,N_23947);
xor U24219 (N_24219,N_23834,N_23985);
xnor U24220 (N_24220,N_23914,N_23907);
and U24221 (N_24221,N_23940,N_23991);
nor U24222 (N_24222,N_23954,N_23838);
or U24223 (N_24223,N_23790,N_23966);
and U24224 (N_24224,N_23903,N_23913);
nand U24225 (N_24225,N_23836,N_23955);
nor U24226 (N_24226,N_23803,N_23911);
or U24227 (N_24227,N_23977,N_23759);
xnor U24228 (N_24228,N_23834,N_23968);
or U24229 (N_24229,N_23921,N_23988);
nand U24230 (N_24230,N_23954,N_23829);
xor U24231 (N_24231,N_23818,N_23994);
nand U24232 (N_24232,N_23893,N_23923);
xnor U24233 (N_24233,N_23871,N_23922);
nor U24234 (N_24234,N_23940,N_23946);
nand U24235 (N_24235,N_23954,N_23952);
xor U24236 (N_24236,N_23848,N_23976);
or U24237 (N_24237,N_23775,N_23943);
and U24238 (N_24238,N_23869,N_23979);
or U24239 (N_24239,N_23998,N_23869);
or U24240 (N_24240,N_23764,N_23767);
nor U24241 (N_24241,N_23804,N_23952);
and U24242 (N_24242,N_23967,N_23898);
xnor U24243 (N_24243,N_23830,N_23839);
nor U24244 (N_24244,N_23795,N_23995);
xor U24245 (N_24245,N_23903,N_23808);
nor U24246 (N_24246,N_23826,N_23785);
nand U24247 (N_24247,N_23859,N_23799);
and U24248 (N_24248,N_23905,N_23897);
and U24249 (N_24249,N_23879,N_23804);
and U24250 (N_24250,N_24211,N_24220);
nor U24251 (N_24251,N_24031,N_24241);
or U24252 (N_24252,N_24053,N_24001);
nand U24253 (N_24253,N_24127,N_24021);
or U24254 (N_24254,N_24204,N_24023);
nor U24255 (N_24255,N_24033,N_24117);
or U24256 (N_24256,N_24179,N_24012);
nor U24257 (N_24257,N_24028,N_24199);
nor U24258 (N_24258,N_24076,N_24041);
nand U24259 (N_24259,N_24047,N_24049);
nand U24260 (N_24260,N_24232,N_24176);
xor U24261 (N_24261,N_24172,N_24135);
or U24262 (N_24262,N_24198,N_24058);
nand U24263 (N_24263,N_24158,N_24022);
or U24264 (N_24264,N_24133,N_24037);
nand U24265 (N_24265,N_24218,N_24125);
xnor U24266 (N_24266,N_24182,N_24238);
nor U24267 (N_24267,N_24234,N_24228);
nor U24268 (N_24268,N_24247,N_24036);
or U24269 (N_24269,N_24101,N_24157);
and U24270 (N_24270,N_24113,N_24161);
nor U24271 (N_24271,N_24067,N_24185);
xnor U24272 (N_24272,N_24088,N_24124);
or U24273 (N_24273,N_24075,N_24193);
and U24274 (N_24274,N_24174,N_24050);
nor U24275 (N_24275,N_24223,N_24160);
or U24276 (N_24276,N_24005,N_24108);
nor U24277 (N_24277,N_24159,N_24011);
and U24278 (N_24278,N_24120,N_24059);
nor U24279 (N_24279,N_24007,N_24191);
or U24280 (N_24280,N_24225,N_24230);
and U24281 (N_24281,N_24144,N_24136);
xor U24282 (N_24282,N_24079,N_24165);
xnor U24283 (N_24283,N_24151,N_24115);
nand U24284 (N_24284,N_24054,N_24078);
and U24285 (N_24285,N_24065,N_24095);
and U24286 (N_24286,N_24206,N_24093);
or U24287 (N_24287,N_24006,N_24083);
and U24288 (N_24288,N_24143,N_24217);
nor U24289 (N_24289,N_24129,N_24009);
nand U24290 (N_24290,N_24213,N_24014);
nor U24291 (N_24291,N_24068,N_24196);
nor U24292 (N_24292,N_24231,N_24181);
nand U24293 (N_24293,N_24072,N_24130);
xnor U24294 (N_24294,N_24192,N_24227);
and U24295 (N_24295,N_24084,N_24086);
nor U24296 (N_24296,N_24215,N_24048);
and U24297 (N_24297,N_24071,N_24186);
or U24298 (N_24298,N_24082,N_24131);
nor U24299 (N_24299,N_24178,N_24119);
nand U24300 (N_24300,N_24162,N_24187);
xnor U24301 (N_24301,N_24202,N_24121);
and U24302 (N_24302,N_24145,N_24236);
or U24303 (N_24303,N_24235,N_24122);
xor U24304 (N_24304,N_24013,N_24239);
or U24305 (N_24305,N_24141,N_24219);
xnor U24306 (N_24306,N_24132,N_24156);
nor U24307 (N_24307,N_24090,N_24189);
nor U24308 (N_24308,N_24081,N_24064);
nand U24309 (N_24309,N_24105,N_24190);
or U24310 (N_24310,N_24017,N_24044);
and U24311 (N_24311,N_24194,N_24029);
and U24312 (N_24312,N_24056,N_24224);
nor U24313 (N_24313,N_24155,N_24010);
and U24314 (N_24314,N_24094,N_24027);
and U24315 (N_24315,N_24153,N_24051);
or U24316 (N_24316,N_24074,N_24138);
xor U24317 (N_24317,N_24077,N_24098);
or U24318 (N_24318,N_24052,N_24107);
nor U24319 (N_24319,N_24140,N_24018);
nor U24320 (N_24320,N_24169,N_24139);
nand U24321 (N_24321,N_24032,N_24245);
or U24322 (N_24322,N_24055,N_24167);
xnor U24323 (N_24323,N_24016,N_24170);
xnor U24324 (N_24324,N_24175,N_24221);
nand U24325 (N_24325,N_24024,N_24216);
nor U24326 (N_24326,N_24063,N_24118);
nand U24327 (N_24327,N_24034,N_24020);
xnor U24328 (N_24328,N_24112,N_24137);
and U24329 (N_24329,N_24111,N_24104);
or U24330 (N_24330,N_24210,N_24091);
nand U24331 (N_24331,N_24146,N_24073);
or U24332 (N_24332,N_24184,N_24008);
or U24333 (N_24333,N_24102,N_24040);
nor U24334 (N_24334,N_24237,N_24026);
nor U24335 (N_24335,N_24042,N_24188);
nor U24336 (N_24336,N_24249,N_24208);
nand U24337 (N_24337,N_24103,N_24035);
nand U24338 (N_24338,N_24154,N_24000);
nor U24339 (N_24339,N_24046,N_24069);
and U24340 (N_24340,N_24123,N_24106);
xnor U24341 (N_24341,N_24148,N_24240);
or U24342 (N_24342,N_24183,N_24149);
nand U24343 (N_24343,N_24003,N_24166);
and U24344 (N_24344,N_24233,N_24180);
nor U24345 (N_24345,N_24038,N_24019);
xor U24346 (N_24346,N_24087,N_24222);
xnor U24347 (N_24347,N_24097,N_24025);
and U24348 (N_24348,N_24152,N_24168);
nor U24349 (N_24349,N_24043,N_24142);
nand U24350 (N_24350,N_24002,N_24045);
nor U24351 (N_24351,N_24116,N_24171);
nand U24352 (N_24352,N_24243,N_24147);
nor U24353 (N_24353,N_24195,N_24030);
xnor U24354 (N_24354,N_24004,N_24015);
nand U24355 (N_24355,N_24092,N_24096);
or U24356 (N_24356,N_24126,N_24246);
or U24357 (N_24357,N_24212,N_24080);
nor U24358 (N_24358,N_24200,N_24089);
or U24359 (N_24359,N_24134,N_24150);
or U24360 (N_24360,N_24163,N_24099);
xor U24361 (N_24361,N_24070,N_24066);
or U24362 (N_24362,N_24207,N_24203);
nor U24363 (N_24363,N_24057,N_24229);
nand U24364 (N_24364,N_24164,N_24205);
nor U24365 (N_24365,N_24128,N_24085);
xnor U24366 (N_24366,N_24197,N_24100);
nor U24367 (N_24367,N_24173,N_24244);
nand U24368 (N_24368,N_24248,N_24109);
xnor U24369 (N_24369,N_24242,N_24061);
nand U24370 (N_24370,N_24062,N_24209);
nand U24371 (N_24371,N_24214,N_24201);
xor U24372 (N_24372,N_24039,N_24114);
nand U24373 (N_24373,N_24060,N_24110);
or U24374 (N_24374,N_24177,N_24226);
and U24375 (N_24375,N_24111,N_24065);
nor U24376 (N_24376,N_24184,N_24079);
nor U24377 (N_24377,N_24188,N_24122);
xnor U24378 (N_24378,N_24141,N_24190);
nand U24379 (N_24379,N_24061,N_24202);
nor U24380 (N_24380,N_24081,N_24150);
or U24381 (N_24381,N_24094,N_24022);
nor U24382 (N_24382,N_24036,N_24134);
xnor U24383 (N_24383,N_24124,N_24238);
nor U24384 (N_24384,N_24208,N_24154);
and U24385 (N_24385,N_24171,N_24130);
nor U24386 (N_24386,N_24099,N_24193);
and U24387 (N_24387,N_24007,N_24117);
xnor U24388 (N_24388,N_24004,N_24168);
xor U24389 (N_24389,N_24119,N_24116);
and U24390 (N_24390,N_24037,N_24099);
and U24391 (N_24391,N_24234,N_24143);
nor U24392 (N_24392,N_24050,N_24046);
nor U24393 (N_24393,N_24113,N_24243);
and U24394 (N_24394,N_24012,N_24104);
and U24395 (N_24395,N_24036,N_24133);
nor U24396 (N_24396,N_24098,N_24112);
xnor U24397 (N_24397,N_24078,N_24200);
nand U24398 (N_24398,N_24174,N_24245);
xor U24399 (N_24399,N_24044,N_24060);
or U24400 (N_24400,N_24088,N_24153);
xor U24401 (N_24401,N_24246,N_24194);
or U24402 (N_24402,N_24049,N_24091);
or U24403 (N_24403,N_24026,N_24185);
nand U24404 (N_24404,N_24212,N_24054);
nor U24405 (N_24405,N_24210,N_24084);
xor U24406 (N_24406,N_24071,N_24249);
nor U24407 (N_24407,N_24218,N_24170);
and U24408 (N_24408,N_24111,N_24021);
nand U24409 (N_24409,N_24066,N_24166);
xor U24410 (N_24410,N_24228,N_24064);
nand U24411 (N_24411,N_24201,N_24014);
xor U24412 (N_24412,N_24050,N_24016);
or U24413 (N_24413,N_24119,N_24216);
nor U24414 (N_24414,N_24026,N_24055);
nor U24415 (N_24415,N_24126,N_24173);
xnor U24416 (N_24416,N_24170,N_24155);
nand U24417 (N_24417,N_24044,N_24019);
nand U24418 (N_24418,N_24166,N_24040);
nand U24419 (N_24419,N_24008,N_24193);
xor U24420 (N_24420,N_24148,N_24134);
and U24421 (N_24421,N_24073,N_24228);
and U24422 (N_24422,N_24133,N_24201);
or U24423 (N_24423,N_24081,N_24107);
or U24424 (N_24424,N_24018,N_24076);
xnor U24425 (N_24425,N_24146,N_24056);
or U24426 (N_24426,N_24096,N_24219);
nand U24427 (N_24427,N_24125,N_24200);
or U24428 (N_24428,N_24005,N_24152);
xnor U24429 (N_24429,N_24022,N_24183);
and U24430 (N_24430,N_24116,N_24081);
and U24431 (N_24431,N_24194,N_24137);
or U24432 (N_24432,N_24010,N_24168);
or U24433 (N_24433,N_24025,N_24086);
or U24434 (N_24434,N_24064,N_24078);
nor U24435 (N_24435,N_24242,N_24246);
nand U24436 (N_24436,N_24188,N_24125);
xnor U24437 (N_24437,N_24150,N_24042);
nor U24438 (N_24438,N_24155,N_24164);
and U24439 (N_24439,N_24145,N_24213);
xnor U24440 (N_24440,N_24214,N_24127);
xor U24441 (N_24441,N_24134,N_24246);
or U24442 (N_24442,N_24164,N_24195);
nor U24443 (N_24443,N_24190,N_24064);
xor U24444 (N_24444,N_24249,N_24205);
and U24445 (N_24445,N_24157,N_24214);
nor U24446 (N_24446,N_24101,N_24176);
and U24447 (N_24447,N_24233,N_24129);
or U24448 (N_24448,N_24034,N_24095);
nor U24449 (N_24449,N_24168,N_24073);
nand U24450 (N_24450,N_24243,N_24131);
nand U24451 (N_24451,N_24158,N_24005);
or U24452 (N_24452,N_24184,N_24009);
nor U24453 (N_24453,N_24106,N_24175);
or U24454 (N_24454,N_24174,N_24118);
or U24455 (N_24455,N_24032,N_24167);
nor U24456 (N_24456,N_24242,N_24164);
xor U24457 (N_24457,N_24153,N_24077);
nand U24458 (N_24458,N_24039,N_24056);
xor U24459 (N_24459,N_24070,N_24172);
or U24460 (N_24460,N_24069,N_24168);
nor U24461 (N_24461,N_24119,N_24031);
nor U24462 (N_24462,N_24206,N_24192);
nor U24463 (N_24463,N_24061,N_24233);
and U24464 (N_24464,N_24170,N_24046);
xor U24465 (N_24465,N_24070,N_24215);
or U24466 (N_24466,N_24128,N_24035);
nand U24467 (N_24467,N_24246,N_24162);
nand U24468 (N_24468,N_24012,N_24240);
xnor U24469 (N_24469,N_24119,N_24126);
and U24470 (N_24470,N_24212,N_24090);
or U24471 (N_24471,N_24133,N_24206);
or U24472 (N_24472,N_24221,N_24119);
nor U24473 (N_24473,N_24236,N_24021);
xnor U24474 (N_24474,N_24076,N_24164);
nor U24475 (N_24475,N_24208,N_24037);
xnor U24476 (N_24476,N_24188,N_24005);
nand U24477 (N_24477,N_24146,N_24164);
xor U24478 (N_24478,N_24189,N_24178);
and U24479 (N_24479,N_24235,N_24239);
nor U24480 (N_24480,N_24008,N_24235);
xor U24481 (N_24481,N_24210,N_24196);
or U24482 (N_24482,N_24172,N_24082);
nor U24483 (N_24483,N_24003,N_24177);
nor U24484 (N_24484,N_24006,N_24247);
xor U24485 (N_24485,N_24132,N_24034);
xnor U24486 (N_24486,N_24073,N_24244);
nand U24487 (N_24487,N_24114,N_24213);
nand U24488 (N_24488,N_24224,N_24168);
and U24489 (N_24489,N_24034,N_24051);
or U24490 (N_24490,N_24194,N_24067);
nand U24491 (N_24491,N_24163,N_24018);
xnor U24492 (N_24492,N_24088,N_24027);
xor U24493 (N_24493,N_24079,N_24022);
nand U24494 (N_24494,N_24108,N_24073);
nor U24495 (N_24495,N_24202,N_24088);
and U24496 (N_24496,N_24074,N_24087);
and U24497 (N_24497,N_24216,N_24057);
nand U24498 (N_24498,N_24160,N_24093);
nand U24499 (N_24499,N_24134,N_24183);
xnor U24500 (N_24500,N_24294,N_24489);
nand U24501 (N_24501,N_24295,N_24394);
or U24502 (N_24502,N_24466,N_24322);
and U24503 (N_24503,N_24337,N_24353);
nor U24504 (N_24504,N_24330,N_24257);
xnor U24505 (N_24505,N_24454,N_24428);
and U24506 (N_24506,N_24402,N_24306);
xor U24507 (N_24507,N_24252,N_24298);
xor U24508 (N_24508,N_24387,N_24455);
xnor U24509 (N_24509,N_24485,N_24378);
or U24510 (N_24510,N_24476,N_24366);
nor U24511 (N_24511,N_24266,N_24447);
or U24512 (N_24512,N_24432,N_24273);
and U24513 (N_24513,N_24397,N_24302);
and U24514 (N_24514,N_24376,N_24304);
xnor U24515 (N_24515,N_24349,N_24250);
nor U24516 (N_24516,N_24380,N_24461);
and U24517 (N_24517,N_24354,N_24274);
and U24518 (N_24518,N_24305,N_24281);
nand U24519 (N_24519,N_24276,N_24347);
or U24520 (N_24520,N_24443,N_24415);
and U24521 (N_24521,N_24320,N_24283);
or U24522 (N_24522,N_24311,N_24363);
or U24523 (N_24523,N_24399,N_24258);
or U24524 (N_24524,N_24297,N_24448);
xnor U24525 (N_24525,N_24496,N_24429);
and U24526 (N_24526,N_24463,N_24265);
nand U24527 (N_24527,N_24262,N_24410);
nand U24528 (N_24528,N_24420,N_24456);
or U24529 (N_24529,N_24299,N_24286);
or U24530 (N_24530,N_24260,N_24267);
nand U24531 (N_24531,N_24350,N_24417);
nand U24532 (N_24532,N_24451,N_24401);
nor U24533 (N_24533,N_24437,N_24312);
or U24534 (N_24534,N_24339,N_24405);
nand U24535 (N_24535,N_24498,N_24480);
nor U24536 (N_24536,N_24259,N_24256);
and U24537 (N_24537,N_24491,N_24255);
or U24538 (N_24538,N_24469,N_24422);
nand U24539 (N_24539,N_24470,N_24481);
xor U24540 (N_24540,N_24317,N_24418);
or U24541 (N_24541,N_24459,N_24355);
nand U24542 (N_24542,N_24453,N_24474);
nor U24543 (N_24543,N_24285,N_24413);
nand U24544 (N_24544,N_24411,N_24462);
xnor U24545 (N_24545,N_24365,N_24300);
nand U24546 (N_24546,N_24301,N_24371);
xnor U24547 (N_24547,N_24269,N_24370);
nor U24548 (N_24548,N_24490,N_24343);
nand U24549 (N_24549,N_24484,N_24479);
nor U24550 (N_24550,N_24275,N_24393);
xor U24551 (N_24551,N_24288,N_24440);
xor U24552 (N_24552,N_24319,N_24316);
xor U24553 (N_24553,N_24383,N_24385);
or U24554 (N_24554,N_24460,N_24386);
or U24555 (N_24555,N_24321,N_24403);
nand U24556 (N_24556,N_24346,N_24263);
or U24557 (N_24557,N_24293,N_24449);
or U24558 (N_24558,N_24434,N_24367);
or U24559 (N_24559,N_24360,N_24357);
and U24560 (N_24560,N_24335,N_24438);
xor U24561 (N_24561,N_24391,N_24468);
nand U24562 (N_24562,N_24442,N_24439);
nor U24563 (N_24563,N_24427,N_24436);
and U24564 (N_24564,N_24465,N_24472);
or U24565 (N_24565,N_24310,N_24356);
xor U24566 (N_24566,N_24373,N_24408);
and U24567 (N_24567,N_24426,N_24270);
nor U24568 (N_24568,N_24473,N_24328);
xnor U24569 (N_24569,N_24333,N_24336);
and U24570 (N_24570,N_24477,N_24419);
and U24571 (N_24571,N_24375,N_24493);
nand U24572 (N_24572,N_24421,N_24251);
nand U24573 (N_24573,N_24329,N_24352);
xnor U24574 (N_24574,N_24471,N_24369);
nand U24575 (N_24575,N_24326,N_24482);
and U24576 (N_24576,N_24441,N_24331);
and U24577 (N_24577,N_24342,N_24478);
and U24578 (N_24578,N_24309,N_24409);
xor U24579 (N_24579,N_24325,N_24278);
xnor U24580 (N_24580,N_24389,N_24332);
nand U24581 (N_24581,N_24396,N_24416);
and U24582 (N_24582,N_24430,N_24464);
or U24583 (N_24583,N_24398,N_24324);
and U24584 (N_24584,N_24487,N_24425);
and U24585 (N_24585,N_24338,N_24497);
or U24586 (N_24586,N_24279,N_24289);
xnor U24587 (N_24587,N_24327,N_24495);
xnor U24588 (N_24588,N_24368,N_24290);
or U24589 (N_24589,N_24435,N_24351);
nor U24590 (N_24590,N_24414,N_24431);
nand U24591 (N_24591,N_24268,N_24303);
or U24592 (N_24592,N_24340,N_24308);
and U24593 (N_24593,N_24492,N_24264);
xnor U24594 (N_24594,N_24423,N_24261);
nand U24595 (N_24595,N_24494,N_24395);
and U24596 (N_24596,N_24445,N_24483);
nor U24597 (N_24597,N_24392,N_24382);
nand U24598 (N_24598,N_24254,N_24404);
nand U24599 (N_24599,N_24424,N_24450);
xor U24600 (N_24600,N_24444,N_24284);
and U24601 (N_24601,N_24475,N_24407);
nor U24602 (N_24602,N_24307,N_24271);
xnor U24603 (N_24603,N_24318,N_24348);
xnor U24604 (N_24604,N_24334,N_24388);
or U24605 (N_24605,N_24253,N_24467);
nor U24606 (N_24606,N_24458,N_24315);
nor U24607 (N_24607,N_24296,N_24291);
and U24608 (N_24608,N_24345,N_24400);
nor U24609 (N_24609,N_24499,N_24381);
and U24610 (N_24610,N_24344,N_24282);
and U24611 (N_24611,N_24390,N_24313);
nor U24612 (N_24612,N_24374,N_24277);
and U24613 (N_24613,N_24379,N_24272);
nand U24614 (N_24614,N_24412,N_24446);
nand U24615 (N_24615,N_24323,N_24364);
and U24616 (N_24616,N_24457,N_24488);
xor U24617 (N_24617,N_24486,N_24314);
xnor U24618 (N_24618,N_24358,N_24341);
and U24619 (N_24619,N_24292,N_24280);
or U24620 (N_24620,N_24287,N_24377);
nor U24621 (N_24621,N_24406,N_24384);
nand U24622 (N_24622,N_24362,N_24372);
nor U24623 (N_24623,N_24452,N_24361);
and U24624 (N_24624,N_24433,N_24359);
nor U24625 (N_24625,N_24440,N_24339);
nand U24626 (N_24626,N_24432,N_24363);
and U24627 (N_24627,N_24322,N_24366);
or U24628 (N_24628,N_24354,N_24434);
or U24629 (N_24629,N_24384,N_24403);
xor U24630 (N_24630,N_24427,N_24455);
nor U24631 (N_24631,N_24380,N_24313);
nand U24632 (N_24632,N_24496,N_24414);
or U24633 (N_24633,N_24279,N_24364);
and U24634 (N_24634,N_24431,N_24329);
xnor U24635 (N_24635,N_24438,N_24257);
nand U24636 (N_24636,N_24488,N_24267);
and U24637 (N_24637,N_24420,N_24429);
nor U24638 (N_24638,N_24453,N_24369);
and U24639 (N_24639,N_24366,N_24317);
xnor U24640 (N_24640,N_24305,N_24251);
xor U24641 (N_24641,N_24447,N_24479);
nor U24642 (N_24642,N_24381,N_24438);
xor U24643 (N_24643,N_24370,N_24377);
nand U24644 (N_24644,N_24381,N_24437);
nand U24645 (N_24645,N_24253,N_24477);
and U24646 (N_24646,N_24433,N_24276);
nor U24647 (N_24647,N_24293,N_24416);
xor U24648 (N_24648,N_24487,N_24305);
nand U24649 (N_24649,N_24369,N_24337);
xor U24650 (N_24650,N_24402,N_24264);
xor U24651 (N_24651,N_24297,N_24368);
xnor U24652 (N_24652,N_24427,N_24274);
nand U24653 (N_24653,N_24466,N_24460);
or U24654 (N_24654,N_24333,N_24250);
nand U24655 (N_24655,N_24280,N_24494);
nor U24656 (N_24656,N_24391,N_24498);
xor U24657 (N_24657,N_24371,N_24498);
nand U24658 (N_24658,N_24364,N_24422);
nor U24659 (N_24659,N_24462,N_24268);
xnor U24660 (N_24660,N_24481,N_24291);
and U24661 (N_24661,N_24498,N_24438);
xor U24662 (N_24662,N_24400,N_24377);
xnor U24663 (N_24663,N_24454,N_24320);
and U24664 (N_24664,N_24371,N_24254);
or U24665 (N_24665,N_24459,N_24399);
nand U24666 (N_24666,N_24443,N_24493);
xor U24667 (N_24667,N_24424,N_24416);
or U24668 (N_24668,N_24335,N_24260);
and U24669 (N_24669,N_24468,N_24413);
or U24670 (N_24670,N_24405,N_24368);
nor U24671 (N_24671,N_24364,N_24298);
xor U24672 (N_24672,N_24440,N_24435);
nand U24673 (N_24673,N_24362,N_24458);
and U24674 (N_24674,N_24355,N_24280);
nand U24675 (N_24675,N_24287,N_24490);
nand U24676 (N_24676,N_24484,N_24290);
or U24677 (N_24677,N_24453,N_24307);
nand U24678 (N_24678,N_24471,N_24282);
xor U24679 (N_24679,N_24260,N_24445);
and U24680 (N_24680,N_24266,N_24340);
or U24681 (N_24681,N_24362,N_24319);
nor U24682 (N_24682,N_24467,N_24459);
nor U24683 (N_24683,N_24345,N_24418);
and U24684 (N_24684,N_24400,N_24256);
nor U24685 (N_24685,N_24368,N_24463);
or U24686 (N_24686,N_24432,N_24365);
or U24687 (N_24687,N_24369,N_24383);
or U24688 (N_24688,N_24475,N_24302);
nand U24689 (N_24689,N_24473,N_24398);
or U24690 (N_24690,N_24389,N_24453);
and U24691 (N_24691,N_24376,N_24365);
nor U24692 (N_24692,N_24400,N_24287);
xnor U24693 (N_24693,N_24450,N_24325);
or U24694 (N_24694,N_24481,N_24436);
nand U24695 (N_24695,N_24351,N_24438);
xnor U24696 (N_24696,N_24330,N_24400);
and U24697 (N_24697,N_24272,N_24277);
xor U24698 (N_24698,N_24326,N_24495);
xor U24699 (N_24699,N_24255,N_24463);
or U24700 (N_24700,N_24409,N_24450);
xnor U24701 (N_24701,N_24438,N_24312);
nor U24702 (N_24702,N_24320,N_24324);
nor U24703 (N_24703,N_24453,N_24442);
and U24704 (N_24704,N_24440,N_24266);
or U24705 (N_24705,N_24363,N_24420);
and U24706 (N_24706,N_24461,N_24267);
and U24707 (N_24707,N_24334,N_24366);
xnor U24708 (N_24708,N_24490,N_24276);
nor U24709 (N_24709,N_24335,N_24441);
nand U24710 (N_24710,N_24463,N_24402);
or U24711 (N_24711,N_24405,N_24324);
and U24712 (N_24712,N_24370,N_24335);
xnor U24713 (N_24713,N_24458,N_24489);
or U24714 (N_24714,N_24256,N_24432);
or U24715 (N_24715,N_24400,N_24475);
or U24716 (N_24716,N_24273,N_24471);
and U24717 (N_24717,N_24483,N_24407);
nor U24718 (N_24718,N_24458,N_24453);
nor U24719 (N_24719,N_24272,N_24341);
xor U24720 (N_24720,N_24384,N_24263);
and U24721 (N_24721,N_24331,N_24257);
nand U24722 (N_24722,N_24284,N_24272);
nor U24723 (N_24723,N_24442,N_24262);
or U24724 (N_24724,N_24331,N_24474);
nand U24725 (N_24725,N_24436,N_24393);
or U24726 (N_24726,N_24480,N_24304);
nand U24727 (N_24727,N_24323,N_24326);
nor U24728 (N_24728,N_24252,N_24431);
xor U24729 (N_24729,N_24288,N_24446);
xor U24730 (N_24730,N_24293,N_24418);
or U24731 (N_24731,N_24340,N_24450);
or U24732 (N_24732,N_24361,N_24436);
xor U24733 (N_24733,N_24339,N_24465);
xor U24734 (N_24734,N_24360,N_24438);
and U24735 (N_24735,N_24440,N_24282);
nor U24736 (N_24736,N_24255,N_24345);
nor U24737 (N_24737,N_24458,N_24477);
and U24738 (N_24738,N_24434,N_24427);
nor U24739 (N_24739,N_24349,N_24451);
nor U24740 (N_24740,N_24443,N_24476);
xor U24741 (N_24741,N_24375,N_24380);
xnor U24742 (N_24742,N_24266,N_24306);
xor U24743 (N_24743,N_24446,N_24470);
or U24744 (N_24744,N_24299,N_24257);
and U24745 (N_24745,N_24332,N_24376);
or U24746 (N_24746,N_24289,N_24440);
nor U24747 (N_24747,N_24322,N_24318);
nand U24748 (N_24748,N_24382,N_24412);
nor U24749 (N_24749,N_24259,N_24369);
nor U24750 (N_24750,N_24606,N_24598);
and U24751 (N_24751,N_24632,N_24633);
or U24752 (N_24752,N_24602,N_24732);
or U24753 (N_24753,N_24575,N_24704);
and U24754 (N_24754,N_24591,N_24654);
or U24755 (N_24755,N_24708,N_24748);
and U24756 (N_24756,N_24729,N_24615);
nand U24757 (N_24757,N_24600,N_24614);
or U24758 (N_24758,N_24720,N_24657);
nand U24759 (N_24759,N_24641,N_24561);
or U24760 (N_24760,N_24527,N_24722);
nand U24761 (N_24761,N_24690,N_24679);
nand U24762 (N_24762,N_24531,N_24640);
xnor U24763 (N_24763,N_24669,N_24672);
xor U24764 (N_24764,N_24659,N_24572);
nand U24765 (N_24765,N_24516,N_24656);
xnor U24766 (N_24766,N_24534,N_24581);
nor U24767 (N_24767,N_24682,N_24570);
xnor U24768 (N_24768,N_24622,N_24541);
xor U24769 (N_24769,N_24580,N_24660);
nand U24770 (N_24770,N_24565,N_24725);
xor U24771 (N_24771,N_24719,N_24674);
nor U24772 (N_24772,N_24698,N_24573);
or U24773 (N_24773,N_24515,N_24718);
nor U24774 (N_24774,N_24585,N_24529);
and U24775 (N_24775,N_24731,N_24670);
and U24776 (N_24776,N_24727,N_24624);
xor U24777 (N_24777,N_24513,N_24650);
nand U24778 (N_24778,N_24688,N_24599);
nor U24779 (N_24779,N_24611,N_24741);
nor U24780 (N_24780,N_24697,N_24685);
xor U24781 (N_24781,N_24539,N_24530);
nor U24782 (N_24782,N_24584,N_24616);
or U24783 (N_24783,N_24634,N_24740);
and U24784 (N_24784,N_24663,N_24579);
or U24785 (N_24785,N_24596,N_24746);
nand U24786 (N_24786,N_24512,N_24558);
nand U24787 (N_24787,N_24511,N_24696);
and U24788 (N_24788,N_24662,N_24522);
xor U24789 (N_24789,N_24647,N_24610);
nand U24790 (N_24790,N_24737,N_24627);
nor U24791 (N_24791,N_24566,N_24501);
xnor U24792 (N_24792,N_24604,N_24637);
and U24793 (N_24793,N_24612,N_24548);
xor U24794 (N_24794,N_24618,N_24538);
xnor U24795 (N_24795,N_24631,N_24567);
and U24796 (N_24796,N_24713,N_24597);
nor U24797 (N_24797,N_24555,N_24528);
nand U24798 (N_24798,N_24609,N_24592);
or U24799 (N_24799,N_24595,N_24687);
or U24800 (N_24800,N_24553,N_24661);
or U24801 (N_24801,N_24628,N_24507);
and U24802 (N_24802,N_24736,N_24504);
nor U24803 (N_24803,N_24636,N_24673);
and U24804 (N_24804,N_24712,N_24546);
nor U24805 (N_24805,N_24677,N_24676);
nor U24806 (N_24806,N_24526,N_24648);
or U24807 (N_24807,N_24739,N_24700);
or U24808 (N_24808,N_24564,N_24655);
nand U24809 (N_24809,N_24626,N_24562);
or U24810 (N_24810,N_24535,N_24686);
and U24811 (N_24811,N_24706,N_24684);
or U24812 (N_24812,N_24653,N_24543);
xor U24813 (N_24813,N_24714,N_24587);
nor U24814 (N_24814,N_24590,N_24724);
or U24815 (N_24815,N_24577,N_24703);
or U24816 (N_24816,N_24701,N_24533);
or U24817 (N_24817,N_24607,N_24617);
and U24818 (N_24818,N_24603,N_24711);
or U24819 (N_24819,N_24726,N_24680);
or U24820 (N_24820,N_24583,N_24665);
xor U24821 (N_24821,N_24563,N_24681);
nand U24822 (N_24822,N_24619,N_24537);
nor U24823 (N_24823,N_24514,N_24594);
xor U24824 (N_24824,N_24666,N_24544);
xor U24825 (N_24825,N_24643,N_24588);
and U24826 (N_24826,N_24519,N_24505);
nand U24827 (N_24827,N_24521,N_24574);
or U24828 (N_24828,N_24709,N_24683);
nor U24829 (N_24829,N_24613,N_24503);
and U24830 (N_24830,N_24557,N_24707);
or U24831 (N_24831,N_24675,N_24671);
nor U24832 (N_24832,N_24742,N_24639);
nor U24833 (N_24833,N_24723,N_24589);
xor U24834 (N_24834,N_24623,N_24692);
nor U24835 (N_24835,N_24638,N_24644);
nor U24836 (N_24836,N_24620,N_24747);
nor U24837 (N_24837,N_24601,N_24559);
and U24838 (N_24838,N_24524,N_24710);
and U24839 (N_24839,N_24693,N_24576);
nor U24840 (N_24840,N_24560,N_24689);
or U24841 (N_24841,N_24745,N_24651);
nor U24842 (N_24842,N_24691,N_24593);
or U24843 (N_24843,N_24621,N_24578);
nor U24844 (N_24844,N_24547,N_24630);
xor U24845 (N_24845,N_24586,N_24730);
xnor U24846 (N_24846,N_24571,N_24502);
or U24847 (N_24847,N_24552,N_24749);
xor U24848 (N_24848,N_24664,N_24695);
or U24849 (N_24849,N_24678,N_24743);
nor U24850 (N_24850,N_24510,N_24517);
nand U24851 (N_24851,N_24518,N_24658);
xnor U24852 (N_24852,N_24744,N_24500);
and U24853 (N_24853,N_24629,N_24735);
nand U24854 (N_24854,N_24721,N_24705);
and U24855 (N_24855,N_24645,N_24605);
and U24856 (N_24856,N_24508,N_24556);
xor U24857 (N_24857,N_24532,N_24542);
xnor U24858 (N_24858,N_24716,N_24717);
nor U24859 (N_24859,N_24540,N_24668);
and U24860 (N_24860,N_24550,N_24649);
xnor U24861 (N_24861,N_24699,N_24733);
nor U24862 (N_24862,N_24568,N_24702);
and U24863 (N_24863,N_24646,N_24715);
and U24864 (N_24864,N_24554,N_24582);
nand U24865 (N_24865,N_24525,N_24608);
or U24866 (N_24866,N_24509,N_24738);
nor U24867 (N_24867,N_24569,N_24551);
and U24868 (N_24868,N_24625,N_24520);
nor U24869 (N_24869,N_24506,N_24545);
or U24870 (N_24870,N_24667,N_24694);
xnor U24871 (N_24871,N_24635,N_24536);
or U24872 (N_24872,N_24728,N_24734);
and U24873 (N_24873,N_24523,N_24652);
xnor U24874 (N_24874,N_24549,N_24642);
and U24875 (N_24875,N_24605,N_24652);
or U24876 (N_24876,N_24589,N_24560);
nor U24877 (N_24877,N_24529,N_24538);
nor U24878 (N_24878,N_24636,N_24747);
xnor U24879 (N_24879,N_24671,N_24509);
xor U24880 (N_24880,N_24577,N_24660);
or U24881 (N_24881,N_24622,N_24698);
and U24882 (N_24882,N_24723,N_24702);
nand U24883 (N_24883,N_24613,N_24650);
or U24884 (N_24884,N_24719,N_24737);
nor U24885 (N_24885,N_24647,N_24623);
xnor U24886 (N_24886,N_24638,N_24735);
or U24887 (N_24887,N_24687,N_24599);
or U24888 (N_24888,N_24697,N_24704);
nand U24889 (N_24889,N_24574,N_24513);
and U24890 (N_24890,N_24610,N_24575);
xnor U24891 (N_24891,N_24627,N_24668);
and U24892 (N_24892,N_24651,N_24559);
nor U24893 (N_24893,N_24512,N_24529);
nand U24894 (N_24894,N_24596,N_24628);
xor U24895 (N_24895,N_24718,N_24745);
and U24896 (N_24896,N_24685,N_24655);
nand U24897 (N_24897,N_24732,N_24544);
nor U24898 (N_24898,N_24574,N_24673);
or U24899 (N_24899,N_24610,N_24691);
nand U24900 (N_24900,N_24708,N_24603);
and U24901 (N_24901,N_24566,N_24704);
nor U24902 (N_24902,N_24573,N_24678);
nand U24903 (N_24903,N_24604,N_24545);
xnor U24904 (N_24904,N_24591,N_24533);
xnor U24905 (N_24905,N_24567,N_24726);
nand U24906 (N_24906,N_24621,N_24548);
nor U24907 (N_24907,N_24706,N_24643);
nand U24908 (N_24908,N_24528,N_24523);
nand U24909 (N_24909,N_24728,N_24640);
nor U24910 (N_24910,N_24586,N_24722);
nand U24911 (N_24911,N_24536,N_24653);
xor U24912 (N_24912,N_24716,N_24673);
and U24913 (N_24913,N_24745,N_24542);
or U24914 (N_24914,N_24504,N_24737);
and U24915 (N_24915,N_24526,N_24524);
xor U24916 (N_24916,N_24672,N_24561);
xor U24917 (N_24917,N_24617,N_24686);
xnor U24918 (N_24918,N_24679,N_24534);
xnor U24919 (N_24919,N_24655,N_24662);
xor U24920 (N_24920,N_24592,N_24536);
or U24921 (N_24921,N_24741,N_24564);
xor U24922 (N_24922,N_24737,N_24573);
nor U24923 (N_24923,N_24544,N_24686);
xnor U24924 (N_24924,N_24602,N_24533);
xnor U24925 (N_24925,N_24652,N_24700);
nor U24926 (N_24926,N_24683,N_24608);
and U24927 (N_24927,N_24605,N_24523);
nand U24928 (N_24928,N_24720,N_24600);
and U24929 (N_24929,N_24687,N_24626);
or U24930 (N_24930,N_24604,N_24530);
nor U24931 (N_24931,N_24599,N_24538);
nand U24932 (N_24932,N_24586,N_24601);
xnor U24933 (N_24933,N_24598,N_24536);
xnor U24934 (N_24934,N_24541,N_24667);
nand U24935 (N_24935,N_24656,N_24572);
or U24936 (N_24936,N_24639,N_24735);
or U24937 (N_24937,N_24547,N_24603);
xnor U24938 (N_24938,N_24504,N_24592);
nand U24939 (N_24939,N_24658,N_24712);
or U24940 (N_24940,N_24743,N_24653);
nor U24941 (N_24941,N_24729,N_24622);
xnor U24942 (N_24942,N_24505,N_24722);
nor U24943 (N_24943,N_24725,N_24575);
nor U24944 (N_24944,N_24701,N_24585);
xnor U24945 (N_24945,N_24647,N_24574);
xor U24946 (N_24946,N_24592,N_24593);
nand U24947 (N_24947,N_24553,N_24584);
and U24948 (N_24948,N_24658,N_24537);
xnor U24949 (N_24949,N_24747,N_24524);
xor U24950 (N_24950,N_24572,N_24676);
nor U24951 (N_24951,N_24690,N_24737);
and U24952 (N_24952,N_24596,N_24690);
and U24953 (N_24953,N_24719,N_24748);
nor U24954 (N_24954,N_24722,N_24576);
nand U24955 (N_24955,N_24722,N_24623);
xnor U24956 (N_24956,N_24732,N_24510);
or U24957 (N_24957,N_24574,N_24639);
nand U24958 (N_24958,N_24658,N_24630);
xnor U24959 (N_24959,N_24600,N_24693);
nand U24960 (N_24960,N_24653,N_24562);
nand U24961 (N_24961,N_24511,N_24544);
xor U24962 (N_24962,N_24521,N_24555);
and U24963 (N_24963,N_24689,N_24525);
or U24964 (N_24964,N_24537,N_24535);
or U24965 (N_24965,N_24622,N_24509);
nand U24966 (N_24966,N_24565,N_24713);
nor U24967 (N_24967,N_24522,N_24516);
nor U24968 (N_24968,N_24710,N_24726);
nand U24969 (N_24969,N_24557,N_24720);
or U24970 (N_24970,N_24730,N_24699);
xnor U24971 (N_24971,N_24524,N_24677);
nor U24972 (N_24972,N_24728,N_24585);
nand U24973 (N_24973,N_24538,N_24534);
and U24974 (N_24974,N_24705,N_24748);
nand U24975 (N_24975,N_24692,N_24748);
nand U24976 (N_24976,N_24526,N_24624);
and U24977 (N_24977,N_24619,N_24594);
nor U24978 (N_24978,N_24546,N_24682);
xnor U24979 (N_24979,N_24711,N_24745);
nor U24980 (N_24980,N_24614,N_24714);
or U24981 (N_24981,N_24607,N_24637);
or U24982 (N_24982,N_24710,N_24540);
nor U24983 (N_24983,N_24662,N_24632);
nand U24984 (N_24984,N_24716,N_24628);
and U24985 (N_24985,N_24727,N_24746);
xnor U24986 (N_24986,N_24742,N_24608);
or U24987 (N_24987,N_24649,N_24524);
nor U24988 (N_24988,N_24687,N_24556);
nand U24989 (N_24989,N_24561,N_24515);
xor U24990 (N_24990,N_24550,N_24581);
nand U24991 (N_24991,N_24683,N_24747);
or U24992 (N_24992,N_24624,N_24583);
nand U24993 (N_24993,N_24583,N_24718);
and U24994 (N_24994,N_24694,N_24740);
xnor U24995 (N_24995,N_24687,N_24584);
and U24996 (N_24996,N_24706,N_24529);
xor U24997 (N_24997,N_24645,N_24631);
nor U24998 (N_24998,N_24732,N_24637);
or U24999 (N_24999,N_24637,N_24547);
and UO_0 (O_0,N_24932,N_24925);
xor UO_1 (O_1,N_24804,N_24820);
and UO_2 (O_2,N_24852,N_24967);
and UO_3 (O_3,N_24878,N_24853);
or UO_4 (O_4,N_24965,N_24920);
xor UO_5 (O_5,N_24944,N_24949);
nand UO_6 (O_6,N_24809,N_24791);
xnor UO_7 (O_7,N_24936,N_24973);
nand UO_8 (O_8,N_24824,N_24797);
or UO_9 (O_9,N_24900,N_24847);
and UO_10 (O_10,N_24902,N_24773);
nand UO_11 (O_11,N_24998,N_24868);
and UO_12 (O_12,N_24871,N_24813);
or UO_13 (O_13,N_24891,N_24884);
or UO_14 (O_14,N_24986,N_24802);
nand UO_15 (O_15,N_24778,N_24882);
xnor UO_16 (O_16,N_24893,N_24975);
xnor UO_17 (O_17,N_24811,N_24751);
nor UO_18 (O_18,N_24772,N_24816);
nand UO_19 (O_19,N_24786,N_24908);
nand UO_20 (O_20,N_24832,N_24762);
or UO_21 (O_21,N_24960,N_24768);
and UO_22 (O_22,N_24927,N_24942);
and UO_23 (O_23,N_24827,N_24947);
and UO_24 (O_24,N_24770,N_24775);
xnor UO_25 (O_25,N_24880,N_24952);
nor UO_26 (O_26,N_24769,N_24765);
xor UO_27 (O_27,N_24752,N_24866);
nand UO_28 (O_28,N_24817,N_24859);
or UO_29 (O_29,N_24924,N_24989);
and UO_30 (O_30,N_24844,N_24777);
nor UO_31 (O_31,N_24899,N_24858);
or UO_32 (O_32,N_24764,N_24997);
and UO_33 (O_33,N_24890,N_24888);
xor UO_34 (O_34,N_24874,N_24800);
xor UO_35 (O_35,N_24935,N_24896);
nor UO_36 (O_36,N_24782,N_24787);
and UO_37 (O_37,N_24914,N_24962);
xor UO_38 (O_38,N_24870,N_24990);
nor UO_39 (O_39,N_24779,N_24867);
xnor UO_40 (O_40,N_24894,N_24943);
xor UO_41 (O_41,N_24819,N_24869);
nor UO_42 (O_42,N_24934,N_24938);
and UO_43 (O_43,N_24876,N_24849);
and UO_44 (O_44,N_24812,N_24839);
nor UO_45 (O_45,N_24833,N_24982);
or UO_46 (O_46,N_24864,N_24991);
or UO_47 (O_47,N_24756,N_24966);
and UO_48 (O_48,N_24848,N_24750);
and UO_49 (O_49,N_24984,N_24837);
nand UO_50 (O_50,N_24886,N_24857);
nor UO_51 (O_51,N_24854,N_24873);
nand UO_52 (O_52,N_24976,N_24805);
nand UO_53 (O_53,N_24789,N_24985);
xor UO_54 (O_54,N_24807,N_24838);
xnor UO_55 (O_55,N_24830,N_24753);
nor UO_56 (O_56,N_24948,N_24972);
nand UO_57 (O_57,N_24915,N_24788);
nand UO_58 (O_58,N_24834,N_24983);
xnor UO_59 (O_59,N_24970,N_24950);
nor UO_60 (O_60,N_24956,N_24821);
nor UO_61 (O_61,N_24763,N_24955);
nand UO_62 (O_62,N_24904,N_24856);
or UO_63 (O_63,N_24988,N_24885);
or UO_64 (O_64,N_24771,N_24954);
nand UO_65 (O_65,N_24922,N_24783);
and UO_66 (O_66,N_24977,N_24980);
nand UO_67 (O_67,N_24994,N_24959);
nand UO_68 (O_68,N_24795,N_24911);
and UO_69 (O_69,N_24861,N_24946);
xnor UO_70 (O_70,N_24918,N_24917);
and UO_71 (O_71,N_24754,N_24969);
nand UO_72 (O_72,N_24840,N_24968);
nand UO_73 (O_73,N_24790,N_24855);
nor UO_74 (O_74,N_24843,N_24826);
and UO_75 (O_75,N_24822,N_24964);
nor UO_76 (O_76,N_24889,N_24803);
xnor UO_77 (O_77,N_24905,N_24850);
xor UO_78 (O_78,N_24923,N_24971);
xor UO_79 (O_79,N_24883,N_24860);
and UO_80 (O_80,N_24825,N_24958);
and UO_81 (O_81,N_24758,N_24760);
and UO_82 (O_82,N_24828,N_24841);
or UO_83 (O_83,N_24879,N_24921);
xnor UO_84 (O_84,N_24862,N_24875);
and UO_85 (O_85,N_24910,N_24836);
nand UO_86 (O_86,N_24774,N_24814);
or UO_87 (O_87,N_24810,N_24755);
xor UO_88 (O_88,N_24993,N_24793);
nand UO_89 (O_89,N_24895,N_24981);
nand UO_90 (O_90,N_24806,N_24846);
nor UO_91 (O_91,N_24759,N_24792);
xor UO_92 (O_92,N_24999,N_24992);
or UO_93 (O_93,N_24877,N_24937);
nand UO_94 (O_94,N_24851,N_24930);
xnor UO_95 (O_95,N_24766,N_24987);
xor UO_96 (O_96,N_24951,N_24978);
nand UO_97 (O_97,N_24957,N_24767);
nor UO_98 (O_98,N_24801,N_24865);
nand UO_99 (O_99,N_24916,N_24898);
xnor UO_100 (O_100,N_24794,N_24829);
and UO_101 (O_101,N_24796,N_24798);
nor UO_102 (O_102,N_24933,N_24963);
nor UO_103 (O_103,N_24939,N_24897);
nor UO_104 (O_104,N_24784,N_24941);
and UO_105 (O_105,N_24776,N_24929);
xnor UO_106 (O_106,N_24799,N_24995);
xor UO_107 (O_107,N_24909,N_24996);
and UO_108 (O_108,N_24974,N_24780);
xnor UO_109 (O_109,N_24919,N_24757);
and UO_110 (O_110,N_24785,N_24815);
or UO_111 (O_111,N_24931,N_24901);
nor UO_112 (O_112,N_24881,N_24903);
and UO_113 (O_113,N_24872,N_24906);
nor UO_114 (O_114,N_24913,N_24863);
or UO_115 (O_115,N_24940,N_24845);
xnor UO_116 (O_116,N_24961,N_24912);
or UO_117 (O_117,N_24887,N_24979);
nand UO_118 (O_118,N_24892,N_24928);
nand UO_119 (O_119,N_24831,N_24926);
nor UO_120 (O_120,N_24953,N_24781);
nor UO_121 (O_121,N_24907,N_24761);
and UO_122 (O_122,N_24808,N_24835);
and UO_123 (O_123,N_24818,N_24842);
nand UO_124 (O_124,N_24823,N_24945);
and UO_125 (O_125,N_24827,N_24961);
and UO_126 (O_126,N_24899,N_24907);
nor UO_127 (O_127,N_24786,N_24949);
nor UO_128 (O_128,N_24967,N_24954);
or UO_129 (O_129,N_24996,N_24847);
nor UO_130 (O_130,N_24908,N_24988);
and UO_131 (O_131,N_24855,N_24930);
and UO_132 (O_132,N_24985,N_24996);
xnor UO_133 (O_133,N_24960,N_24796);
and UO_134 (O_134,N_24957,N_24874);
or UO_135 (O_135,N_24840,N_24853);
nor UO_136 (O_136,N_24995,N_24769);
xnor UO_137 (O_137,N_24792,N_24768);
or UO_138 (O_138,N_24842,N_24953);
xnor UO_139 (O_139,N_24774,N_24787);
nand UO_140 (O_140,N_24833,N_24775);
nand UO_141 (O_141,N_24770,N_24927);
nor UO_142 (O_142,N_24883,N_24799);
or UO_143 (O_143,N_24851,N_24946);
nand UO_144 (O_144,N_24969,N_24840);
and UO_145 (O_145,N_24954,N_24834);
xnor UO_146 (O_146,N_24949,N_24953);
or UO_147 (O_147,N_24816,N_24932);
and UO_148 (O_148,N_24888,N_24893);
nor UO_149 (O_149,N_24788,N_24805);
xnor UO_150 (O_150,N_24828,N_24980);
nand UO_151 (O_151,N_24973,N_24759);
and UO_152 (O_152,N_24991,N_24875);
and UO_153 (O_153,N_24811,N_24827);
and UO_154 (O_154,N_24980,N_24885);
nand UO_155 (O_155,N_24959,N_24793);
and UO_156 (O_156,N_24980,N_24894);
nor UO_157 (O_157,N_24948,N_24785);
nand UO_158 (O_158,N_24997,N_24923);
nand UO_159 (O_159,N_24790,N_24842);
nor UO_160 (O_160,N_24812,N_24981);
or UO_161 (O_161,N_24944,N_24797);
or UO_162 (O_162,N_24973,N_24908);
or UO_163 (O_163,N_24804,N_24982);
nand UO_164 (O_164,N_24981,N_24780);
nand UO_165 (O_165,N_24899,N_24924);
and UO_166 (O_166,N_24890,N_24901);
and UO_167 (O_167,N_24826,N_24812);
xnor UO_168 (O_168,N_24787,N_24984);
xnor UO_169 (O_169,N_24825,N_24848);
xnor UO_170 (O_170,N_24960,N_24836);
nand UO_171 (O_171,N_24958,N_24815);
or UO_172 (O_172,N_24916,N_24946);
nand UO_173 (O_173,N_24821,N_24816);
nand UO_174 (O_174,N_24910,N_24827);
xnor UO_175 (O_175,N_24991,N_24886);
nand UO_176 (O_176,N_24895,N_24868);
xnor UO_177 (O_177,N_24874,N_24790);
nand UO_178 (O_178,N_24895,N_24921);
and UO_179 (O_179,N_24752,N_24898);
nand UO_180 (O_180,N_24867,N_24856);
nand UO_181 (O_181,N_24819,N_24996);
nand UO_182 (O_182,N_24860,N_24786);
nor UO_183 (O_183,N_24796,N_24762);
and UO_184 (O_184,N_24790,N_24814);
nor UO_185 (O_185,N_24887,N_24995);
or UO_186 (O_186,N_24815,N_24910);
nor UO_187 (O_187,N_24877,N_24751);
nand UO_188 (O_188,N_24921,N_24943);
or UO_189 (O_189,N_24827,N_24838);
nor UO_190 (O_190,N_24825,N_24750);
or UO_191 (O_191,N_24893,N_24914);
xnor UO_192 (O_192,N_24951,N_24893);
xor UO_193 (O_193,N_24937,N_24840);
or UO_194 (O_194,N_24805,N_24965);
or UO_195 (O_195,N_24909,N_24831);
nand UO_196 (O_196,N_24970,N_24926);
and UO_197 (O_197,N_24907,N_24969);
or UO_198 (O_198,N_24904,N_24818);
nor UO_199 (O_199,N_24769,N_24844);
nor UO_200 (O_200,N_24973,N_24765);
and UO_201 (O_201,N_24909,N_24966);
and UO_202 (O_202,N_24864,N_24994);
nor UO_203 (O_203,N_24828,N_24873);
nor UO_204 (O_204,N_24836,N_24848);
xor UO_205 (O_205,N_24825,N_24912);
nand UO_206 (O_206,N_24911,N_24907);
and UO_207 (O_207,N_24767,N_24833);
nor UO_208 (O_208,N_24958,N_24942);
nor UO_209 (O_209,N_24818,N_24822);
xor UO_210 (O_210,N_24795,N_24942);
nand UO_211 (O_211,N_24996,N_24769);
and UO_212 (O_212,N_24831,N_24821);
nand UO_213 (O_213,N_24943,N_24779);
nand UO_214 (O_214,N_24759,N_24929);
or UO_215 (O_215,N_24870,N_24787);
xnor UO_216 (O_216,N_24784,N_24792);
and UO_217 (O_217,N_24782,N_24911);
or UO_218 (O_218,N_24971,N_24845);
xor UO_219 (O_219,N_24850,N_24897);
or UO_220 (O_220,N_24994,N_24989);
or UO_221 (O_221,N_24989,N_24891);
xnor UO_222 (O_222,N_24987,N_24891);
nor UO_223 (O_223,N_24870,N_24833);
xor UO_224 (O_224,N_24962,N_24933);
nand UO_225 (O_225,N_24992,N_24785);
or UO_226 (O_226,N_24793,N_24961);
nand UO_227 (O_227,N_24774,N_24919);
xnor UO_228 (O_228,N_24939,N_24943);
and UO_229 (O_229,N_24811,N_24867);
or UO_230 (O_230,N_24827,N_24850);
or UO_231 (O_231,N_24787,N_24840);
and UO_232 (O_232,N_24777,N_24867);
or UO_233 (O_233,N_24751,N_24795);
or UO_234 (O_234,N_24795,N_24897);
nor UO_235 (O_235,N_24894,N_24889);
or UO_236 (O_236,N_24925,N_24919);
xor UO_237 (O_237,N_24942,N_24882);
xor UO_238 (O_238,N_24785,N_24855);
and UO_239 (O_239,N_24772,N_24757);
nand UO_240 (O_240,N_24900,N_24790);
nor UO_241 (O_241,N_24775,N_24856);
or UO_242 (O_242,N_24841,N_24929);
nand UO_243 (O_243,N_24876,N_24967);
nand UO_244 (O_244,N_24841,N_24806);
xnor UO_245 (O_245,N_24944,N_24882);
and UO_246 (O_246,N_24818,N_24765);
nor UO_247 (O_247,N_24843,N_24979);
nand UO_248 (O_248,N_24869,N_24886);
xor UO_249 (O_249,N_24813,N_24912);
or UO_250 (O_250,N_24772,N_24774);
or UO_251 (O_251,N_24917,N_24778);
or UO_252 (O_252,N_24788,N_24913);
or UO_253 (O_253,N_24946,N_24932);
nor UO_254 (O_254,N_24840,N_24946);
xnor UO_255 (O_255,N_24945,N_24850);
or UO_256 (O_256,N_24888,N_24999);
and UO_257 (O_257,N_24937,N_24897);
or UO_258 (O_258,N_24900,N_24810);
or UO_259 (O_259,N_24764,N_24843);
and UO_260 (O_260,N_24865,N_24821);
nor UO_261 (O_261,N_24878,N_24986);
and UO_262 (O_262,N_24966,N_24777);
or UO_263 (O_263,N_24793,N_24764);
xnor UO_264 (O_264,N_24791,N_24917);
xor UO_265 (O_265,N_24895,N_24944);
or UO_266 (O_266,N_24921,N_24986);
and UO_267 (O_267,N_24954,N_24837);
nor UO_268 (O_268,N_24960,N_24757);
or UO_269 (O_269,N_24842,N_24805);
xor UO_270 (O_270,N_24823,N_24903);
nand UO_271 (O_271,N_24842,N_24889);
or UO_272 (O_272,N_24834,N_24780);
xor UO_273 (O_273,N_24967,N_24794);
nand UO_274 (O_274,N_24897,N_24751);
xnor UO_275 (O_275,N_24760,N_24849);
and UO_276 (O_276,N_24827,N_24801);
nor UO_277 (O_277,N_24872,N_24908);
nor UO_278 (O_278,N_24934,N_24881);
and UO_279 (O_279,N_24762,N_24989);
xnor UO_280 (O_280,N_24795,N_24991);
xor UO_281 (O_281,N_24939,N_24989);
and UO_282 (O_282,N_24862,N_24949);
and UO_283 (O_283,N_24841,N_24940);
nor UO_284 (O_284,N_24955,N_24789);
xor UO_285 (O_285,N_24908,N_24865);
xor UO_286 (O_286,N_24822,N_24886);
and UO_287 (O_287,N_24984,N_24768);
or UO_288 (O_288,N_24971,N_24918);
xor UO_289 (O_289,N_24878,N_24807);
nand UO_290 (O_290,N_24978,N_24783);
and UO_291 (O_291,N_24903,N_24802);
and UO_292 (O_292,N_24820,N_24905);
xor UO_293 (O_293,N_24891,N_24759);
or UO_294 (O_294,N_24977,N_24895);
nor UO_295 (O_295,N_24806,N_24783);
or UO_296 (O_296,N_24865,N_24783);
or UO_297 (O_297,N_24897,N_24770);
nand UO_298 (O_298,N_24770,N_24979);
xnor UO_299 (O_299,N_24839,N_24978);
nand UO_300 (O_300,N_24943,N_24973);
xnor UO_301 (O_301,N_24817,N_24920);
nand UO_302 (O_302,N_24795,N_24868);
xnor UO_303 (O_303,N_24866,N_24944);
nand UO_304 (O_304,N_24814,N_24925);
nor UO_305 (O_305,N_24877,N_24846);
xnor UO_306 (O_306,N_24937,N_24976);
and UO_307 (O_307,N_24808,N_24757);
nand UO_308 (O_308,N_24842,N_24782);
and UO_309 (O_309,N_24850,N_24977);
or UO_310 (O_310,N_24972,N_24946);
xor UO_311 (O_311,N_24820,N_24848);
xnor UO_312 (O_312,N_24800,N_24780);
and UO_313 (O_313,N_24846,N_24954);
nand UO_314 (O_314,N_24986,N_24903);
and UO_315 (O_315,N_24912,N_24932);
or UO_316 (O_316,N_24828,N_24769);
or UO_317 (O_317,N_24869,N_24772);
or UO_318 (O_318,N_24975,N_24964);
xnor UO_319 (O_319,N_24989,N_24895);
or UO_320 (O_320,N_24782,N_24795);
nor UO_321 (O_321,N_24835,N_24960);
nand UO_322 (O_322,N_24983,N_24902);
nand UO_323 (O_323,N_24963,N_24800);
or UO_324 (O_324,N_24851,N_24839);
and UO_325 (O_325,N_24782,N_24975);
nor UO_326 (O_326,N_24816,N_24768);
nor UO_327 (O_327,N_24788,N_24916);
nand UO_328 (O_328,N_24802,N_24807);
xnor UO_329 (O_329,N_24915,N_24929);
nand UO_330 (O_330,N_24959,N_24865);
or UO_331 (O_331,N_24787,N_24877);
or UO_332 (O_332,N_24956,N_24861);
and UO_333 (O_333,N_24789,N_24932);
nand UO_334 (O_334,N_24876,N_24786);
nand UO_335 (O_335,N_24868,N_24780);
or UO_336 (O_336,N_24949,N_24952);
xor UO_337 (O_337,N_24811,N_24993);
nand UO_338 (O_338,N_24938,N_24915);
nor UO_339 (O_339,N_24758,N_24963);
or UO_340 (O_340,N_24873,N_24846);
nand UO_341 (O_341,N_24831,N_24753);
nor UO_342 (O_342,N_24799,N_24786);
nor UO_343 (O_343,N_24920,N_24795);
xor UO_344 (O_344,N_24947,N_24885);
and UO_345 (O_345,N_24818,N_24887);
xor UO_346 (O_346,N_24837,N_24760);
or UO_347 (O_347,N_24937,N_24799);
nand UO_348 (O_348,N_24975,N_24909);
or UO_349 (O_349,N_24834,N_24888);
and UO_350 (O_350,N_24873,N_24997);
or UO_351 (O_351,N_24897,N_24780);
or UO_352 (O_352,N_24815,N_24813);
or UO_353 (O_353,N_24911,N_24928);
nor UO_354 (O_354,N_24862,N_24793);
nor UO_355 (O_355,N_24947,N_24785);
nand UO_356 (O_356,N_24846,N_24874);
nand UO_357 (O_357,N_24776,N_24979);
and UO_358 (O_358,N_24774,N_24756);
and UO_359 (O_359,N_24848,N_24958);
nand UO_360 (O_360,N_24847,N_24860);
nor UO_361 (O_361,N_24919,N_24857);
and UO_362 (O_362,N_24848,N_24894);
or UO_363 (O_363,N_24816,N_24910);
xor UO_364 (O_364,N_24968,N_24995);
and UO_365 (O_365,N_24944,N_24999);
nand UO_366 (O_366,N_24874,N_24865);
xnor UO_367 (O_367,N_24824,N_24930);
xor UO_368 (O_368,N_24994,N_24865);
nand UO_369 (O_369,N_24856,N_24942);
xor UO_370 (O_370,N_24951,N_24804);
nor UO_371 (O_371,N_24949,N_24913);
or UO_372 (O_372,N_24985,N_24983);
or UO_373 (O_373,N_24783,N_24917);
and UO_374 (O_374,N_24794,N_24998);
xor UO_375 (O_375,N_24801,N_24955);
xor UO_376 (O_376,N_24815,N_24916);
nor UO_377 (O_377,N_24926,N_24863);
nand UO_378 (O_378,N_24839,N_24909);
or UO_379 (O_379,N_24904,N_24868);
or UO_380 (O_380,N_24755,N_24863);
nand UO_381 (O_381,N_24916,N_24972);
nand UO_382 (O_382,N_24838,N_24996);
xnor UO_383 (O_383,N_24999,N_24956);
nor UO_384 (O_384,N_24897,N_24926);
or UO_385 (O_385,N_24940,N_24878);
or UO_386 (O_386,N_24998,N_24763);
and UO_387 (O_387,N_24767,N_24801);
and UO_388 (O_388,N_24802,N_24815);
nand UO_389 (O_389,N_24978,N_24860);
or UO_390 (O_390,N_24793,N_24922);
xnor UO_391 (O_391,N_24990,N_24882);
and UO_392 (O_392,N_24873,N_24970);
xnor UO_393 (O_393,N_24983,N_24818);
xor UO_394 (O_394,N_24838,N_24947);
and UO_395 (O_395,N_24872,N_24928);
nor UO_396 (O_396,N_24765,N_24913);
nand UO_397 (O_397,N_24936,N_24865);
nand UO_398 (O_398,N_24764,N_24928);
and UO_399 (O_399,N_24926,N_24795);
or UO_400 (O_400,N_24992,N_24964);
xor UO_401 (O_401,N_24782,N_24941);
nand UO_402 (O_402,N_24808,N_24899);
nand UO_403 (O_403,N_24949,N_24864);
or UO_404 (O_404,N_24987,N_24820);
xor UO_405 (O_405,N_24769,N_24890);
nor UO_406 (O_406,N_24882,N_24796);
xnor UO_407 (O_407,N_24788,N_24989);
xnor UO_408 (O_408,N_24801,N_24916);
nand UO_409 (O_409,N_24787,N_24966);
nor UO_410 (O_410,N_24921,N_24893);
and UO_411 (O_411,N_24750,N_24822);
and UO_412 (O_412,N_24909,N_24986);
nand UO_413 (O_413,N_24877,N_24894);
xor UO_414 (O_414,N_24757,N_24859);
xor UO_415 (O_415,N_24895,N_24983);
nand UO_416 (O_416,N_24955,N_24791);
nand UO_417 (O_417,N_24997,N_24918);
nor UO_418 (O_418,N_24996,N_24775);
nand UO_419 (O_419,N_24778,N_24844);
nor UO_420 (O_420,N_24944,N_24833);
xnor UO_421 (O_421,N_24971,N_24913);
nand UO_422 (O_422,N_24759,N_24854);
nand UO_423 (O_423,N_24989,N_24790);
or UO_424 (O_424,N_24976,N_24992);
xnor UO_425 (O_425,N_24839,N_24966);
nor UO_426 (O_426,N_24948,N_24982);
nand UO_427 (O_427,N_24819,N_24858);
xor UO_428 (O_428,N_24896,N_24977);
nand UO_429 (O_429,N_24838,N_24813);
nor UO_430 (O_430,N_24894,N_24797);
or UO_431 (O_431,N_24926,N_24825);
nor UO_432 (O_432,N_24814,N_24891);
nor UO_433 (O_433,N_24818,N_24918);
nor UO_434 (O_434,N_24905,N_24846);
xor UO_435 (O_435,N_24805,N_24874);
nand UO_436 (O_436,N_24865,N_24931);
xor UO_437 (O_437,N_24930,N_24960);
and UO_438 (O_438,N_24978,N_24811);
nand UO_439 (O_439,N_24942,N_24793);
xor UO_440 (O_440,N_24758,N_24813);
xnor UO_441 (O_441,N_24989,N_24995);
nand UO_442 (O_442,N_24787,N_24906);
nor UO_443 (O_443,N_24926,N_24946);
or UO_444 (O_444,N_24901,N_24828);
or UO_445 (O_445,N_24810,N_24793);
xnor UO_446 (O_446,N_24772,N_24781);
nor UO_447 (O_447,N_24766,N_24888);
and UO_448 (O_448,N_24875,N_24922);
or UO_449 (O_449,N_24863,N_24892);
nor UO_450 (O_450,N_24880,N_24879);
and UO_451 (O_451,N_24775,N_24899);
or UO_452 (O_452,N_24849,N_24784);
or UO_453 (O_453,N_24889,N_24920);
or UO_454 (O_454,N_24779,N_24798);
nor UO_455 (O_455,N_24809,N_24885);
xnor UO_456 (O_456,N_24830,N_24897);
or UO_457 (O_457,N_24774,N_24998);
xor UO_458 (O_458,N_24832,N_24994);
nor UO_459 (O_459,N_24926,N_24835);
xor UO_460 (O_460,N_24981,N_24772);
xnor UO_461 (O_461,N_24996,N_24846);
and UO_462 (O_462,N_24857,N_24848);
or UO_463 (O_463,N_24783,N_24782);
and UO_464 (O_464,N_24937,N_24841);
or UO_465 (O_465,N_24900,N_24938);
xor UO_466 (O_466,N_24857,N_24834);
nand UO_467 (O_467,N_24768,N_24821);
and UO_468 (O_468,N_24814,N_24788);
or UO_469 (O_469,N_24993,N_24851);
nand UO_470 (O_470,N_24846,N_24965);
and UO_471 (O_471,N_24842,N_24970);
or UO_472 (O_472,N_24957,N_24932);
nand UO_473 (O_473,N_24991,N_24915);
nor UO_474 (O_474,N_24972,N_24974);
nand UO_475 (O_475,N_24874,N_24854);
nor UO_476 (O_476,N_24925,N_24807);
xnor UO_477 (O_477,N_24820,N_24894);
nand UO_478 (O_478,N_24779,N_24751);
and UO_479 (O_479,N_24834,N_24837);
xor UO_480 (O_480,N_24940,N_24870);
or UO_481 (O_481,N_24766,N_24803);
or UO_482 (O_482,N_24953,N_24965);
and UO_483 (O_483,N_24890,N_24873);
nor UO_484 (O_484,N_24909,N_24834);
or UO_485 (O_485,N_24918,N_24871);
or UO_486 (O_486,N_24837,N_24945);
xnor UO_487 (O_487,N_24867,N_24953);
or UO_488 (O_488,N_24879,N_24751);
or UO_489 (O_489,N_24750,N_24836);
nor UO_490 (O_490,N_24847,N_24921);
xnor UO_491 (O_491,N_24926,N_24857);
or UO_492 (O_492,N_24884,N_24940);
or UO_493 (O_493,N_24997,N_24935);
nand UO_494 (O_494,N_24855,N_24951);
or UO_495 (O_495,N_24890,N_24852);
or UO_496 (O_496,N_24856,N_24758);
nor UO_497 (O_497,N_24911,N_24789);
nand UO_498 (O_498,N_24946,N_24793);
and UO_499 (O_499,N_24867,N_24986);
xor UO_500 (O_500,N_24862,N_24896);
nand UO_501 (O_501,N_24780,N_24881);
and UO_502 (O_502,N_24790,N_24999);
xor UO_503 (O_503,N_24754,N_24920);
nor UO_504 (O_504,N_24878,N_24906);
nor UO_505 (O_505,N_24774,N_24878);
and UO_506 (O_506,N_24975,N_24822);
nor UO_507 (O_507,N_24753,N_24993);
nor UO_508 (O_508,N_24997,N_24880);
nor UO_509 (O_509,N_24997,N_24924);
xnor UO_510 (O_510,N_24880,N_24761);
or UO_511 (O_511,N_24782,N_24895);
nor UO_512 (O_512,N_24942,N_24912);
xor UO_513 (O_513,N_24927,N_24841);
or UO_514 (O_514,N_24870,N_24754);
nand UO_515 (O_515,N_24784,N_24871);
nor UO_516 (O_516,N_24873,N_24809);
or UO_517 (O_517,N_24941,N_24920);
and UO_518 (O_518,N_24831,N_24920);
xnor UO_519 (O_519,N_24932,N_24759);
nand UO_520 (O_520,N_24810,N_24841);
nand UO_521 (O_521,N_24836,N_24788);
and UO_522 (O_522,N_24913,N_24894);
xor UO_523 (O_523,N_24763,N_24794);
and UO_524 (O_524,N_24901,N_24929);
or UO_525 (O_525,N_24759,N_24864);
nand UO_526 (O_526,N_24776,N_24955);
nand UO_527 (O_527,N_24751,N_24807);
xnor UO_528 (O_528,N_24915,N_24981);
xnor UO_529 (O_529,N_24772,N_24753);
nand UO_530 (O_530,N_24819,N_24870);
xnor UO_531 (O_531,N_24838,N_24904);
nor UO_532 (O_532,N_24860,N_24946);
and UO_533 (O_533,N_24898,N_24826);
nand UO_534 (O_534,N_24873,N_24845);
or UO_535 (O_535,N_24825,N_24832);
or UO_536 (O_536,N_24885,N_24859);
nand UO_537 (O_537,N_24829,N_24944);
or UO_538 (O_538,N_24801,N_24971);
and UO_539 (O_539,N_24870,N_24804);
or UO_540 (O_540,N_24826,N_24856);
or UO_541 (O_541,N_24857,N_24891);
or UO_542 (O_542,N_24960,N_24771);
or UO_543 (O_543,N_24757,N_24876);
xor UO_544 (O_544,N_24907,N_24926);
or UO_545 (O_545,N_24839,N_24753);
nor UO_546 (O_546,N_24850,N_24820);
xnor UO_547 (O_547,N_24880,N_24802);
or UO_548 (O_548,N_24872,N_24770);
nor UO_549 (O_549,N_24788,N_24828);
or UO_550 (O_550,N_24800,N_24902);
xor UO_551 (O_551,N_24951,N_24871);
nand UO_552 (O_552,N_24973,N_24920);
xnor UO_553 (O_553,N_24874,N_24987);
or UO_554 (O_554,N_24751,N_24885);
xor UO_555 (O_555,N_24962,N_24870);
or UO_556 (O_556,N_24758,N_24961);
nand UO_557 (O_557,N_24821,N_24967);
or UO_558 (O_558,N_24917,N_24774);
and UO_559 (O_559,N_24848,N_24930);
xnor UO_560 (O_560,N_24778,N_24879);
nor UO_561 (O_561,N_24893,N_24756);
and UO_562 (O_562,N_24847,N_24948);
xnor UO_563 (O_563,N_24779,N_24912);
or UO_564 (O_564,N_24897,N_24966);
xnor UO_565 (O_565,N_24785,N_24834);
and UO_566 (O_566,N_24809,N_24784);
nand UO_567 (O_567,N_24874,N_24822);
or UO_568 (O_568,N_24924,N_24750);
and UO_569 (O_569,N_24797,N_24800);
nor UO_570 (O_570,N_24975,N_24830);
and UO_571 (O_571,N_24993,N_24779);
or UO_572 (O_572,N_24768,N_24934);
and UO_573 (O_573,N_24899,N_24854);
or UO_574 (O_574,N_24769,N_24841);
and UO_575 (O_575,N_24869,N_24827);
and UO_576 (O_576,N_24759,N_24779);
nor UO_577 (O_577,N_24907,N_24773);
xor UO_578 (O_578,N_24941,N_24851);
and UO_579 (O_579,N_24756,N_24805);
and UO_580 (O_580,N_24926,N_24951);
nor UO_581 (O_581,N_24860,N_24814);
nor UO_582 (O_582,N_24950,N_24855);
xor UO_583 (O_583,N_24759,N_24974);
nand UO_584 (O_584,N_24796,N_24877);
or UO_585 (O_585,N_24872,N_24847);
and UO_586 (O_586,N_24937,N_24852);
and UO_587 (O_587,N_24819,N_24973);
and UO_588 (O_588,N_24789,N_24809);
xor UO_589 (O_589,N_24886,N_24849);
and UO_590 (O_590,N_24922,N_24784);
or UO_591 (O_591,N_24971,N_24897);
nor UO_592 (O_592,N_24975,N_24947);
nand UO_593 (O_593,N_24826,N_24910);
nand UO_594 (O_594,N_24861,N_24976);
and UO_595 (O_595,N_24930,N_24926);
or UO_596 (O_596,N_24779,N_24755);
and UO_597 (O_597,N_24917,N_24824);
xor UO_598 (O_598,N_24797,N_24829);
or UO_599 (O_599,N_24813,N_24916);
or UO_600 (O_600,N_24790,N_24782);
and UO_601 (O_601,N_24883,N_24809);
or UO_602 (O_602,N_24931,N_24934);
and UO_603 (O_603,N_24772,N_24918);
or UO_604 (O_604,N_24826,N_24835);
xor UO_605 (O_605,N_24765,N_24808);
and UO_606 (O_606,N_24795,N_24876);
xnor UO_607 (O_607,N_24892,N_24896);
or UO_608 (O_608,N_24778,N_24966);
xnor UO_609 (O_609,N_24866,N_24766);
or UO_610 (O_610,N_24919,N_24943);
nand UO_611 (O_611,N_24794,N_24965);
nand UO_612 (O_612,N_24958,N_24750);
and UO_613 (O_613,N_24912,N_24835);
nand UO_614 (O_614,N_24921,N_24873);
or UO_615 (O_615,N_24956,N_24878);
nor UO_616 (O_616,N_24994,N_24777);
xnor UO_617 (O_617,N_24989,N_24855);
and UO_618 (O_618,N_24858,N_24762);
nand UO_619 (O_619,N_24907,N_24769);
nand UO_620 (O_620,N_24906,N_24898);
nor UO_621 (O_621,N_24989,N_24796);
nand UO_622 (O_622,N_24946,N_24939);
and UO_623 (O_623,N_24933,N_24991);
xnor UO_624 (O_624,N_24785,N_24821);
or UO_625 (O_625,N_24946,N_24841);
xor UO_626 (O_626,N_24975,N_24844);
nor UO_627 (O_627,N_24940,N_24757);
and UO_628 (O_628,N_24838,N_24992);
or UO_629 (O_629,N_24942,N_24791);
and UO_630 (O_630,N_24809,N_24825);
nor UO_631 (O_631,N_24956,N_24883);
xnor UO_632 (O_632,N_24808,N_24797);
nor UO_633 (O_633,N_24770,N_24817);
xnor UO_634 (O_634,N_24823,N_24842);
and UO_635 (O_635,N_24886,N_24862);
nor UO_636 (O_636,N_24754,N_24760);
and UO_637 (O_637,N_24768,N_24886);
and UO_638 (O_638,N_24845,N_24934);
and UO_639 (O_639,N_24840,N_24765);
xnor UO_640 (O_640,N_24785,N_24872);
nor UO_641 (O_641,N_24969,N_24994);
xor UO_642 (O_642,N_24958,N_24949);
nor UO_643 (O_643,N_24857,N_24913);
nand UO_644 (O_644,N_24823,N_24864);
and UO_645 (O_645,N_24966,N_24983);
or UO_646 (O_646,N_24811,N_24984);
nor UO_647 (O_647,N_24964,N_24901);
nand UO_648 (O_648,N_24989,N_24845);
xor UO_649 (O_649,N_24826,N_24940);
nor UO_650 (O_650,N_24935,N_24903);
xor UO_651 (O_651,N_24851,N_24925);
nand UO_652 (O_652,N_24932,N_24811);
and UO_653 (O_653,N_24771,N_24765);
nand UO_654 (O_654,N_24886,N_24913);
nor UO_655 (O_655,N_24926,N_24778);
nor UO_656 (O_656,N_24786,N_24882);
and UO_657 (O_657,N_24943,N_24928);
xor UO_658 (O_658,N_24943,N_24822);
nand UO_659 (O_659,N_24965,N_24968);
nand UO_660 (O_660,N_24838,N_24896);
or UO_661 (O_661,N_24796,N_24990);
nor UO_662 (O_662,N_24752,N_24829);
xnor UO_663 (O_663,N_24751,N_24870);
and UO_664 (O_664,N_24901,N_24882);
nand UO_665 (O_665,N_24934,N_24769);
nand UO_666 (O_666,N_24764,N_24868);
or UO_667 (O_667,N_24825,N_24831);
nand UO_668 (O_668,N_24818,N_24825);
or UO_669 (O_669,N_24910,N_24783);
nor UO_670 (O_670,N_24870,N_24768);
and UO_671 (O_671,N_24926,N_24802);
or UO_672 (O_672,N_24790,N_24829);
xor UO_673 (O_673,N_24849,N_24811);
xor UO_674 (O_674,N_24782,N_24820);
and UO_675 (O_675,N_24972,N_24862);
xnor UO_676 (O_676,N_24803,N_24804);
or UO_677 (O_677,N_24894,N_24873);
nor UO_678 (O_678,N_24789,N_24813);
or UO_679 (O_679,N_24826,N_24779);
nor UO_680 (O_680,N_24936,N_24760);
xnor UO_681 (O_681,N_24825,N_24960);
and UO_682 (O_682,N_24893,N_24760);
nand UO_683 (O_683,N_24888,N_24949);
or UO_684 (O_684,N_24840,N_24885);
or UO_685 (O_685,N_24991,N_24796);
and UO_686 (O_686,N_24856,N_24899);
or UO_687 (O_687,N_24976,N_24972);
and UO_688 (O_688,N_24906,N_24770);
nor UO_689 (O_689,N_24912,N_24832);
xnor UO_690 (O_690,N_24820,N_24919);
or UO_691 (O_691,N_24875,N_24859);
and UO_692 (O_692,N_24834,N_24878);
or UO_693 (O_693,N_24833,N_24826);
or UO_694 (O_694,N_24839,N_24816);
nor UO_695 (O_695,N_24914,N_24840);
xor UO_696 (O_696,N_24768,N_24784);
and UO_697 (O_697,N_24823,N_24934);
nand UO_698 (O_698,N_24943,N_24877);
nor UO_699 (O_699,N_24756,N_24970);
nor UO_700 (O_700,N_24900,N_24795);
or UO_701 (O_701,N_24970,N_24752);
xnor UO_702 (O_702,N_24941,N_24945);
nand UO_703 (O_703,N_24891,N_24859);
or UO_704 (O_704,N_24869,N_24769);
nor UO_705 (O_705,N_24819,N_24786);
and UO_706 (O_706,N_24826,N_24752);
nor UO_707 (O_707,N_24848,N_24751);
and UO_708 (O_708,N_24948,N_24998);
and UO_709 (O_709,N_24821,N_24867);
nand UO_710 (O_710,N_24753,N_24968);
xnor UO_711 (O_711,N_24964,N_24793);
nor UO_712 (O_712,N_24952,N_24885);
and UO_713 (O_713,N_24765,N_24780);
xor UO_714 (O_714,N_24854,N_24791);
nor UO_715 (O_715,N_24828,N_24879);
and UO_716 (O_716,N_24775,N_24861);
xor UO_717 (O_717,N_24894,N_24964);
nand UO_718 (O_718,N_24764,N_24874);
and UO_719 (O_719,N_24830,N_24866);
xor UO_720 (O_720,N_24794,N_24768);
nand UO_721 (O_721,N_24778,N_24837);
and UO_722 (O_722,N_24970,N_24808);
or UO_723 (O_723,N_24816,N_24825);
and UO_724 (O_724,N_24907,N_24890);
or UO_725 (O_725,N_24794,N_24922);
or UO_726 (O_726,N_24819,N_24958);
or UO_727 (O_727,N_24888,N_24860);
and UO_728 (O_728,N_24829,N_24804);
or UO_729 (O_729,N_24863,N_24954);
nor UO_730 (O_730,N_24848,N_24790);
nand UO_731 (O_731,N_24845,N_24948);
and UO_732 (O_732,N_24896,N_24842);
and UO_733 (O_733,N_24774,N_24871);
nand UO_734 (O_734,N_24873,N_24892);
or UO_735 (O_735,N_24794,N_24828);
nor UO_736 (O_736,N_24998,N_24921);
and UO_737 (O_737,N_24912,N_24879);
nand UO_738 (O_738,N_24971,N_24822);
or UO_739 (O_739,N_24865,N_24983);
xor UO_740 (O_740,N_24825,N_24962);
nor UO_741 (O_741,N_24941,N_24967);
or UO_742 (O_742,N_24922,N_24838);
or UO_743 (O_743,N_24813,N_24956);
or UO_744 (O_744,N_24928,N_24758);
nand UO_745 (O_745,N_24914,N_24970);
xnor UO_746 (O_746,N_24779,N_24908);
nor UO_747 (O_747,N_24963,N_24782);
nand UO_748 (O_748,N_24907,N_24780);
or UO_749 (O_749,N_24849,N_24769);
and UO_750 (O_750,N_24923,N_24875);
nand UO_751 (O_751,N_24853,N_24891);
nand UO_752 (O_752,N_24950,N_24783);
nor UO_753 (O_753,N_24924,N_24786);
or UO_754 (O_754,N_24891,N_24795);
nor UO_755 (O_755,N_24947,N_24867);
nor UO_756 (O_756,N_24819,N_24989);
nand UO_757 (O_757,N_24971,N_24963);
nor UO_758 (O_758,N_24933,N_24806);
nor UO_759 (O_759,N_24788,N_24999);
nand UO_760 (O_760,N_24772,N_24851);
nor UO_761 (O_761,N_24886,N_24961);
and UO_762 (O_762,N_24810,N_24786);
nor UO_763 (O_763,N_24836,N_24802);
xnor UO_764 (O_764,N_24946,N_24890);
or UO_765 (O_765,N_24850,N_24813);
nor UO_766 (O_766,N_24984,N_24940);
or UO_767 (O_767,N_24829,N_24895);
nand UO_768 (O_768,N_24861,N_24964);
and UO_769 (O_769,N_24832,N_24999);
nor UO_770 (O_770,N_24766,N_24862);
nand UO_771 (O_771,N_24954,N_24756);
and UO_772 (O_772,N_24964,N_24909);
and UO_773 (O_773,N_24827,N_24763);
xor UO_774 (O_774,N_24832,N_24834);
or UO_775 (O_775,N_24992,N_24839);
nand UO_776 (O_776,N_24995,N_24793);
nand UO_777 (O_777,N_24989,N_24799);
or UO_778 (O_778,N_24892,N_24903);
and UO_779 (O_779,N_24751,N_24774);
or UO_780 (O_780,N_24871,N_24938);
and UO_781 (O_781,N_24842,N_24924);
and UO_782 (O_782,N_24845,N_24936);
nor UO_783 (O_783,N_24765,N_24767);
or UO_784 (O_784,N_24761,N_24752);
and UO_785 (O_785,N_24991,N_24938);
xnor UO_786 (O_786,N_24776,N_24905);
or UO_787 (O_787,N_24809,N_24971);
nor UO_788 (O_788,N_24868,N_24805);
nor UO_789 (O_789,N_24958,N_24809);
nand UO_790 (O_790,N_24788,N_24854);
xnor UO_791 (O_791,N_24952,N_24883);
or UO_792 (O_792,N_24822,N_24907);
and UO_793 (O_793,N_24783,N_24914);
nand UO_794 (O_794,N_24857,N_24770);
xor UO_795 (O_795,N_24883,N_24837);
and UO_796 (O_796,N_24919,N_24806);
nand UO_797 (O_797,N_24764,N_24953);
and UO_798 (O_798,N_24928,N_24932);
nand UO_799 (O_799,N_24934,N_24996);
or UO_800 (O_800,N_24912,N_24828);
nor UO_801 (O_801,N_24865,N_24805);
nor UO_802 (O_802,N_24946,N_24889);
nor UO_803 (O_803,N_24786,N_24870);
xnor UO_804 (O_804,N_24787,N_24975);
and UO_805 (O_805,N_24871,N_24988);
or UO_806 (O_806,N_24920,N_24833);
nor UO_807 (O_807,N_24903,N_24948);
nor UO_808 (O_808,N_24875,N_24828);
nor UO_809 (O_809,N_24866,N_24913);
nand UO_810 (O_810,N_24882,N_24803);
nand UO_811 (O_811,N_24848,N_24910);
or UO_812 (O_812,N_24788,N_24997);
nor UO_813 (O_813,N_24932,N_24877);
nor UO_814 (O_814,N_24763,N_24906);
nand UO_815 (O_815,N_24901,N_24773);
xnor UO_816 (O_816,N_24802,N_24773);
or UO_817 (O_817,N_24987,N_24864);
nand UO_818 (O_818,N_24957,N_24863);
and UO_819 (O_819,N_24884,N_24803);
nand UO_820 (O_820,N_24915,N_24815);
nand UO_821 (O_821,N_24956,N_24902);
nand UO_822 (O_822,N_24776,N_24833);
nand UO_823 (O_823,N_24976,N_24780);
or UO_824 (O_824,N_24857,N_24880);
nand UO_825 (O_825,N_24963,N_24944);
nor UO_826 (O_826,N_24891,N_24964);
or UO_827 (O_827,N_24963,N_24861);
xor UO_828 (O_828,N_24858,N_24796);
nor UO_829 (O_829,N_24875,N_24829);
or UO_830 (O_830,N_24839,N_24896);
and UO_831 (O_831,N_24858,N_24788);
nand UO_832 (O_832,N_24965,N_24770);
xor UO_833 (O_833,N_24790,N_24985);
xor UO_834 (O_834,N_24993,N_24904);
nor UO_835 (O_835,N_24834,N_24798);
xnor UO_836 (O_836,N_24820,N_24967);
or UO_837 (O_837,N_24906,N_24831);
xnor UO_838 (O_838,N_24759,N_24872);
or UO_839 (O_839,N_24914,N_24824);
nor UO_840 (O_840,N_24902,N_24957);
or UO_841 (O_841,N_24977,N_24778);
or UO_842 (O_842,N_24992,N_24807);
or UO_843 (O_843,N_24957,N_24979);
xor UO_844 (O_844,N_24870,N_24830);
and UO_845 (O_845,N_24905,N_24982);
xor UO_846 (O_846,N_24871,N_24818);
and UO_847 (O_847,N_24846,N_24925);
nor UO_848 (O_848,N_24780,N_24969);
xnor UO_849 (O_849,N_24909,N_24811);
xor UO_850 (O_850,N_24863,N_24932);
or UO_851 (O_851,N_24882,N_24902);
nand UO_852 (O_852,N_24986,N_24779);
xnor UO_853 (O_853,N_24959,N_24935);
and UO_854 (O_854,N_24896,N_24899);
nand UO_855 (O_855,N_24950,N_24778);
nand UO_856 (O_856,N_24970,N_24902);
xor UO_857 (O_857,N_24752,N_24991);
and UO_858 (O_858,N_24751,N_24862);
nand UO_859 (O_859,N_24824,N_24763);
nor UO_860 (O_860,N_24863,N_24852);
or UO_861 (O_861,N_24845,N_24756);
xnor UO_862 (O_862,N_24923,N_24788);
and UO_863 (O_863,N_24868,N_24818);
and UO_864 (O_864,N_24973,N_24807);
nand UO_865 (O_865,N_24915,N_24887);
nand UO_866 (O_866,N_24873,N_24954);
xor UO_867 (O_867,N_24864,N_24985);
xnor UO_868 (O_868,N_24768,N_24887);
xnor UO_869 (O_869,N_24898,N_24831);
and UO_870 (O_870,N_24993,N_24886);
or UO_871 (O_871,N_24901,N_24794);
nor UO_872 (O_872,N_24988,N_24990);
xor UO_873 (O_873,N_24924,N_24757);
or UO_874 (O_874,N_24967,N_24965);
or UO_875 (O_875,N_24971,N_24944);
nand UO_876 (O_876,N_24917,N_24984);
nand UO_877 (O_877,N_24912,N_24949);
nand UO_878 (O_878,N_24794,N_24788);
nand UO_879 (O_879,N_24792,N_24977);
nor UO_880 (O_880,N_24932,N_24929);
xor UO_881 (O_881,N_24936,N_24905);
nor UO_882 (O_882,N_24883,N_24986);
nor UO_883 (O_883,N_24951,N_24806);
nand UO_884 (O_884,N_24982,N_24814);
nor UO_885 (O_885,N_24961,N_24869);
nor UO_886 (O_886,N_24874,N_24870);
nor UO_887 (O_887,N_24758,N_24932);
nor UO_888 (O_888,N_24915,N_24931);
nand UO_889 (O_889,N_24866,N_24983);
nor UO_890 (O_890,N_24770,N_24957);
or UO_891 (O_891,N_24794,N_24872);
nor UO_892 (O_892,N_24989,N_24798);
xor UO_893 (O_893,N_24882,N_24756);
and UO_894 (O_894,N_24899,N_24913);
xnor UO_895 (O_895,N_24754,N_24860);
or UO_896 (O_896,N_24812,N_24978);
nor UO_897 (O_897,N_24974,N_24850);
and UO_898 (O_898,N_24890,N_24941);
or UO_899 (O_899,N_24917,N_24799);
and UO_900 (O_900,N_24927,N_24771);
nand UO_901 (O_901,N_24954,N_24824);
and UO_902 (O_902,N_24858,N_24822);
and UO_903 (O_903,N_24795,N_24821);
nor UO_904 (O_904,N_24885,N_24770);
nor UO_905 (O_905,N_24917,N_24941);
and UO_906 (O_906,N_24780,N_24763);
or UO_907 (O_907,N_24758,N_24967);
or UO_908 (O_908,N_24933,N_24944);
nor UO_909 (O_909,N_24912,N_24973);
xnor UO_910 (O_910,N_24817,N_24977);
nor UO_911 (O_911,N_24851,N_24867);
or UO_912 (O_912,N_24773,N_24873);
xor UO_913 (O_913,N_24904,N_24972);
nor UO_914 (O_914,N_24905,N_24972);
and UO_915 (O_915,N_24933,N_24973);
nand UO_916 (O_916,N_24889,N_24931);
and UO_917 (O_917,N_24874,N_24993);
nor UO_918 (O_918,N_24827,N_24996);
xor UO_919 (O_919,N_24982,N_24751);
xnor UO_920 (O_920,N_24890,N_24845);
xor UO_921 (O_921,N_24804,N_24931);
and UO_922 (O_922,N_24782,N_24873);
or UO_923 (O_923,N_24825,N_24851);
and UO_924 (O_924,N_24955,N_24813);
or UO_925 (O_925,N_24803,N_24822);
xor UO_926 (O_926,N_24919,N_24819);
nand UO_927 (O_927,N_24798,N_24873);
nor UO_928 (O_928,N_24817,N_24892);
or UO_929 (O_929,N_24991,N_24974);
xnor UO_930 (O_930,N_24861,N_24962);
or UO_931 (O_931,N_24961,N_24934);
nand UO_932 (O_932,N_24758,N_24891);
or UO_933 (O_933,N_24805,N_24962);
and UO_934 (O_934,N_24918,N_24942);
nor UO_935 (O_935,N_24922,N_24969);
and UO_936 (O_936,N_24939,N_24822);
or UO_937 (O_937,N_24805,N_24763);
nand UO_938 (O_938,N_24828,N_24948);
xnor UO_939 (O_939,N_24955,N_24949);
or UO_940 (O_940,N_24952,N_24831);
nor UO_941 (O_941,N_24896,N_24825);
nand UO_942 (O_942,N_24827,N_24784);
or UO_943 (O_943,N_24825,N_24863);
and UO_944 (O_944,N_24960,N_24914);
xnor UO_945 (O_945,N_24897,N_24967);
and UO_946 (O_946,N_24853,N_24896);
nand UO_947 (O_947,N_24932,N_24992);
nor UO_948 (O_948,N_24870,N_24955);
xnor UO_949 (O_949,N_24950,N_24888);
nand UO_950 (O_950,N_24903,N_24801);
nand UO_951 (O_951,N_24910,N_24882);
nor UO_952 (O_952,N_24891,N_24804);
nor UO_953 (O_953,N_24765,N_24996);
nor UO_954 (O_954,N_24870,N_24973);
xor UO_955 (O_955,N_24939,N_24986);
xnor UO_956 (O_956,N_24911,N_24837);
nand UO_957 (O_957,N_24868,N_24808);
nor UO_958 (O_958,N_24843,N_24751);
nor UO_959 (O_959,N_24963,N_24865);
or UO_960 (O_960,N_24803,N_24970);
nor UO_961 (O_961,N_24901,N_24767);
or UO_962 (O_962,N_24764,N_24958);
or UO_963 (O_963,N_24781,N_24969);
nand UO_964 (O_964,N_24943,N_24826);
xor UO_965 (O_965,N_24757,N_24918);
or UO_966 (O_966,N_24900,N_24774);
nand UO_967 (O_967,N_24754,N_24885);
nor UO_968 (O_968,N_24966,N_24763);
nand UO_969 (O_969,N_24931,N_24778);
or UO_970 (O_970,N_24787,N_24851);
nand UO_971 (O_971,N_24972,N_24831);
xnor UO_972 (O_972,N_24782,N_24986);
and UO_973 (O_973,N_24762,N_24783);
nand UO_974 (O_974,N_24909,N_24989);
nor UO_975 (O_975,N_24944,N_24862);
or UO_976 (O_976,N_24781,N_24843);
or UO_977 (O_977,N_24880,N_24848);
and UO_978 (O_978,N_24925,N_24861);
xnor UO_979 (O_979,N_24889,N_24892);
and UO_980 (O_980,N_24907,N_24981);
nor UO_981 (O_981,N_24895,N_24896);
nor UO_982 (O_982,N_24776,N_24761);
xor UO_983 (O_983,N_24998,N_24907);
xor UO_984 (O_984,N_24984,N_24827);
nor UO_985 (O_985,N_24993,N_24816);
nor UO_986 (O_986,N_24772,N_24974);
nand UO_987 (O_987,N_24769,N_24814);
and UO_988 (O_988,N_24860,N_24846);
nor UO_989 (O_989,N_24761,N_24816);
nand UO_990 (O_990,N_24942,N_24877);
and UO_991 (O_991,N_24853,N_24967);
xnor UO_992 (O_992,N_24956,N_24918);
or UO_993 (O_993,N_24809,N_24804);
nand UO_994 (O_994,N_24872,N_24867);
or UO_995 (O_995,N_24768,N_24836);
nand UO_996 (O_996,N_24779,N_24968);
nand UO_997 (O_997,N_24898,N_24800);
or UO_998 (O_998,N_24873,N_24772);
and UO_999 (O_999,N_24771,N_24980);
or UO_1000 (O_1000,N_24845,N_24815);
nor UO_1001 (O_1001,N_24981,N_24900);
xnor UO_1002 (O_1002,N_24786,N_24967);
nand UO_1003 (O_1003,N_24850,N_24991);
nand UO_1004 (O_1004,N_24823,N_24781);
or UO_1005 (O_1005,N_24770,N_24773);
xor UO_1006 (O_1006,N_24937,N_24971);
xnor UO_1007 (O_1007,N_24874,N_24774);
xor UO_1008 (O_1008,N_24895,N_24912);
nand UO_1009 (O_1009,N_24817,N_24889);
and UO_1010 (O_1010,N_24914,N_24940);
nand UO_1011 (O_1011,N_24984,N_24948);
xor UO_1012 (O_1012,N_24750,N_24834);
nor UO_1013 (O_1013,N_24753,N_24939);
or UO_1014 (O_1014,N_24836,N_24776);
or UO_1015 (O_1015,N_24782,N_24893);
xor UO_1016 (O_1016,N_24976,N_24924);
xnor UO_1017 (O_1017,N_24840,N_24836);
xnor UO_1018 (O_1018,N_24965,N_24933);
xnor UO_1019 (O_1019,N_24935,N_24886);
nor UO_1020 (O_1020,N_24883,N_24816);
and UO_1021 (O_1021,N_24759,N_24836);
and UO_1022 (O_1022,N_24966,N_24996);
and UO_1023 (O_1023,N_24908,N_24920);
or UO_1024 (O_1024,N_24890,N_24917);
nand UO_1025 (O_1025,N_24990,N_24798);
and UO_1026 (O_1026,N_24806,N_24786);
xor UO_1027 (O_1027,N_24894,N_24842);
nor UO_1028 (O_1028,N_24870,N_24956);
or UO_1029 (O_1029,N_24922,N_24981);
nand UO_1030 (O_1030,N_24892,N_24822);
and UO_1031 (O_1031,N_24750,N_24866);
and UO_1032 (O_1032,N_24773,N_24913);
nand UO_1033 (O_1033,N_24790,N_24885);
nor UO_1034 (O_1034,N_24833,N_24785);
xnor UO_1035 (O_1035,N_24919,N_24956);
and UO_1036 (O_1036,N_24935,N_24847);
nor UO_1037 (O_1037,N_24852,N_24825);
xnor UO_1038 (O_1038,N_24767,N_24795);
nand UO_1039 (O_1039,N_24802,N_24941);
nand UO_1040 (O_1040,N_24855,N_24822);
xnor UO_1041 (O_1041,N_24882,N_24955);
or UO_1042 (O_1042,N_24982,N_24856);
nor UO_1043 (O_1043,N_24885,N_24976);
xnor UO_1044 (O_1044,N_24825,N_24998);
and UO_1045 (O_1045,N_24961,N_24936);
and UO_1046 (O_1046,N_24807,N_24914);
xor UO_1047 (O_1047,N_24907,N_24851);
nor UO_1048 (O_1048,N_24940,N_24758);
xnor UO_1049 (O_1049,N_24841,N_24958);
nor UO_1050 (O_1050,N_24782,N_24850);
or UO_1051 (O_1051,N_24768,N_24847);
and UO_1052 (O_1052,N_24946,N_24772);
xnor UO_1053 (O_1053,N_24923,N_24766);
nor UO_1054 (O_1054,N_24779,N_24906);
xnor UO_1055 (O_1055,N_24800,N_24908);
nor UO_1056 (O_1056,N_24957,N_24916);
nand UO_1057 (O_1057,N_24976,N_24785);
xor UO_1058 (O_1058,N_24839,N_24772);
and UO_1059 (O_1059,N_24763,N_24956);
nand UO_1060 (O_1060,N_24975,N_24862);
or UO_1061 (O_1061,N_24994,N_24782);
xnor UO_1062 (O_1062,N_24755,N_24801);
xnor UO_1063 (O_1063,N_24896,N_24918);
nor UO_1064 (O_1064,N_24822,N_24832);
nand UO_1065 (O_1065,N_24977,N_24970);
xor UO_1066 (O_1066,N_24755,N_24915);
nand UO_1067 (O_1067,N_24750,N_24880);
nor UO_1068 (O_1068,N_24972,N_24754);
and UO_1069 (O_1069,N_24903,N_24858);
nor UO_1070 (O_1070,N_24892,N_24757);
nand UO_1071 (O_1071,N_24946,N_24895);
or UO_1072 (O_1072,N_24909,N_24875);
nand UO_1073 (O_1073,N_24805,N_24859);
or UO_1074 (O_1074,N_24779,N_24849);
nand UO_1075 (O_1075,N_24859,N_24967);
and UO_1076 (O_1076,N_24868,N_24902);
nor UO_1077 (O_1077,N_24830,N_24867);
or UO_1078 (O_1078,N_24798,N_24837);
nor UO_1079 (O_1079,N_24901,N_24827);
nand UO_1080 (O_1080,N_24930,N_24853);
nor UO_1081 (O_1081,N_24943,N_24860);
nand UO_1082 (O_1082,N_24917,N_24867);
nand UO_1083 (O_1083,N_24796,N_24931);
nand UO_1084 (O_1084,N_24945,N_24750);
or UO_1085 (O_1085,N_24984,N_24849);
xor UO_1086 (O_1086,N_24950,N_24949);
or UO_1087 (O_1087,N_24916,N_24866);
nor UO_1088 (O_1088,N_24843,N_24849);
nand UO_1089 (O_1089,N_24938,N_24898);
and UO_1090 (O_1090,N_24918,N_24911);
nand UO_1091 (O_1091,N_24979,N_24774);
nand UO_1092 (O_1092,N_24759,N_24987);
nor UO_1093 (O_1093,N_24813,N_24764);
or UO_1094 (O_1094,N_24752,N_24836);
and UO_1095 (O_1095,N_24788,N_24906);
or UO_1096 (O_1096,N_24960,N_24979);
nor UO_1097 (O_1097,N_24978,N_24989);
nand UO_1098 (O_1098,N_24861,N_24774);
xnor UO_1099 (O_1099,N_24915,N_24837);
or UO_1100 (O_1100,N_24919,N_24799);
xor UO_1101 (O_1101,N_24910,N_24924);
nor UO_1102 (O_1102,N_24769,N_24779);
and UO_1103 (O_1103,N_24886,N_24810);
and UO_1104 (O_1104,N_24933,N_24865);
or UO_1105 (O_1105,N_24802,N_24991);
nor UO_1106 (O_1106,N_24961,N_24752);
nand UO_1107 (O_1107,N_24918,N_24760);
and UO_1108 (O_1108,N_24845,N_24816);
and UO_1109 (O_1109,N_24804,N_24868);
xnor UO_1110 (O_1110,N_24893,N_24764);
or UO_1111 (O_1111,N_24892,N_24891);
nor UO_1112 (O_1112,N_24916,N_24986);
nor UO_1113 (O_1113,N_24773,N_24992);
or UO_1114 (O_1114,N_24907,N_24764);
nand UO_1115 (O_1115,N_24791,N_24836);
nand UO_1116 (O_1116,N_24985,N_24850);
and UO_1117 (O_1117,N_24935,N_24840);
and UO_1118 (O_1118,N_24770,N_24977);
or UO_1119 (O_1119,N_24899,N_24932);
xor UO_1120 (O_1120,N_24993,N_24873);
nand UO_1121 (O_1121,N_24776,N_24923);
xnor UO_1122 (O_1122,N_24751,N_24887);
nand UO_1123 (O_1123,N_24902,N_24853);
or UO_1124 (O_1124,N_24917,N_24926);
nor UO_1125 (O_1125,N_24922,N_24933);
and UO_1126 (O_1126,N_24796,N_24830);
nand UO_1127 (O_1127,N_24899,N_24815);
nand UO_1128 (O_1128,N_24751,N_24932);
nor UO_1129 (O_1129,N_24818,N_24947);
nor UO_1130 (O_1130,N_24993,N_24883);
or UO_1131 (O_1131,N_24898,N_24950);
or UO_1132 (O_1132,N_24761,N_24847);
nor UO_1133 (O_1133,N_24929,N_24956);
or UO_1134 (O_1134,N_24998,N_24775);
or UO_1135 (O_1135,N_24913,N_24947);
xnor UO_1136 (O_1136,N_24914,N_24957);
xor UO_1137 (O_1137,N_24978,N_24750);
or UO_1138 (O_1138,N_24901,N_24914);
or UO_1139 (O_1139,N_24967,N_24791);
and UO_1140 (O_1140,N_24846,N_24974);
nor UO_1141 (O_1141,N_24965,N_24945);
and UO_1142 (O_1142,N_24823,N_24996);
nor UO_1143 (O_1143,N_24755,N_24999);
and UO_1144 (O_1144,N_24751,N_24907);
nor UO_1145 (O_1145,N_24994,N_24892);
xnor UO_1146 (O_1146,N_24996,N_24859);
or UO_1147 (O_1147,N_24800,N_24809);
nand UO_1148 (O_1148,N_24833,N_24784);
nor UO_1149 (O_1149,N_24858,N_24874);
or UO_1150 (O_1150,N_24986,N_24825);
nand UO_1151 (O_1151,N_24847,N_24863);
and UO_1152 (O_1152,N_24874,N_24835);
nor UO_1153 (O_1153,N_24787,N_24885);
nand UO_1154 (O_1154,N_24986,N_24948);
nand UO_1155 (O_1155,N_24938,N_24760);
or UO_1156 (O_1156,N_24991,N_24977);
xor UO_1157 (O_1157,N_24831,N_24886);
nor UO_1158 (O_1158,N_24943,N_24771);
xor UO_1159 (O_1159,N_24787,N_24940);
and UO_1160 (O_1160,N_24992,N_24869);
and UO_1161 (O_1161,N_24988,N_24902);
nor UO_1162 (O_1162,N_24956,N_24934);
nor UO_1163 (O_1163,N_24797,N_24878);
xnor UO_1164 (O_1164,N_24769,N_24940);
nor UO_1165 (O_1165,N_24959,N_24901);
and UO_1166 (O_1166,N_24921,N_24825);
xor UO_1167 (O_1167,N_24841,N_24973);
or UO_1168 (O_1168,N_24885,N_24915);
or UO_1169 (O_1169,N_24930,N_24785);
xor UO_1170 (O_1170,N_24789,N_24953);
xnor UO_1171 (O_1171,N_24914,N_24769);
xnor UO_1172 (O_1172,N_24841,N_24819);
nor UO_1173 (O_1173,N_24908,N_24841);
nor UO_1174 (O_1174,N_24919,N_24814);
or UO_1175 (O_1175,N_24978,N_24819);
and UO_1176 (O_1176,N_24843,N_24820);
nand UO_1177 (O_1177,N_24964,N_24960);
nand UO_1178 (O_1178,N_24998,N_24816);
and UO_1179 (O_1179,N_24956,N_24921);
xor UO_1180 (O_1180,N_24852,N_24980);
xnor UO_1181 (O_1181,N_24865,N_24766);
nor UO_1182 (O_1182,N_24787,N_24862);
nand UO_1183 (O_1183,N_24877,N_24767);
nor UO_1184 (O_1184,N_24985,N_24883);
nand UO_1185 (O_1185,N_24953,N_24880);
and UO_1186 (O_1186,N_24948,N_24825);
and UO_1187 (O_1187,N_24813,N_24981);
and UO_1188 (O_1188,N_24871,N_24763);
nor UO_1189 (O_1189,N_24873,N_24753);
nand UO_1190 (O_1190,N_24812,N_24787);
or UO_1191 (O_1191,N_24862,N_24833);
xnor UO_1192 (O_1192,N_24881,N_24947);
nand UO_1193 (O_1193,N_24931,N_24844);
xnor UO_1194 (O_1194,N_24900,N_24750);
nor UO_1195 (O_1195,N_24771,N_24847);
nand UO_1196 (O_1196,N_24894,N_24849);
xnor UO_1197 (O_1197,N_24846,N_24927);
nor UO_1198 (O_1198,N_24899,N_24976);
nand UO_1199 (O_1199,N_24756,N_24994);
xor UO_1200 (O_1200,N_24871,N_24750);
xnor UO_1201 (O_1201,N_24788,N_24900);
nor UO_1202 (O_1202,N_24994,N_24761);
nand UO_1203 (O_1203,N_24764,N_24993);
xor UO_1204 (O_1204,N_24849,N_24906);
nor UO_1205 (O_1205,N_24929,N_24860);
and UO_1206 (O_1206,N_24831,N_24976);
nand UO_1207 (O_1207,N_24869,N_24875);
xnor UO_1208 (O_1208,N_24994,N_24839);
nor UO_1209 (O_1209,N_24940,N_24920);
nand UO_1210 (O_1210,N_24917,N_24768);
xnor UO_1211 (O_1211,N_24764,N_24802);
or UO_1212 (O_1212,N_24975,N_24828);
and UO_1213 (O_1213,N_24855,N_24889);
xor UO_1214 (O_1214,N_24863,N_24962);
nor UO_1215 (O_1215,N_24850,N_24756);
or UO_1216 (O_1216,N_24809,N_24867);
nand UO_1217 (O_1217,N_24916,N_24830);
and UO_1218 (O_1218,N_24775,N_24928);
xnor UO_1219 (O_1219,N_24850,N_24859);
nor UO_1220 (O_1220,N_24788,N_24948);
xnor UO_1221 (O_1221,N_24978,N_24901);
and UO_1222 (O_1222,N_24872,N_24831);
nor UO_1223 (O_1223,N_24991,N_24896);
xor UO_1224 (O_1224,N_24777,N_24845);
nand UO_1225 (O_1225,N_24936,N_24810);
xor UO_1226 (O_1226,N_24832,N_24989);
xor UO_1227 (O_1227,N_24965,N_24804);
nand UO_1228 (O_1228,N_24785,N_24964);
and UO_1229 (O_1229,N_24919,N_24978);
nor UO_1230 (O_1230,N_24834,N_24814);
xor UO_1231 (O_1231,N_24933,N_24750);
and UO_1232 (O_1232,N_24993,N_24977);
xnor UO_1233 (O_1233,N_24926,N_24881);
nor UO_1234 (O_1234,N_24802,N_24761);
and UO_1235 (O_1235,N_24895,N_24992);
xnor UO_1236 (O_1236,N_24802,N_24918);
or UO_1237 (O_1237,N_24915,N_24833);
nand UO_1238 (O_1238,N_24938,N_24911);
nand UO_1239 (O_1239,N_24837,N_24803);
nand UO_1240 (O_1240,N_24842,N_24996);
xor UO_1241 (O_1241,N_24937,N_24869);
nand UO_1242 (O_1242,N_24975,N_24940);
and UO_1243 (O_1243,N_24818,N_24877);
nor UO_1244 (O_1244,N_24783,N_24819);
nor UO_1245 (O_1245,N_24882,N_24929);
and UO_1246 (O_1246,N_24784,N_24860);
or UO_1247 (O_1247,N_24852,N_24873);
nand UO_1248 (O_1248,N_24755,N_24788);
nor UO_1249 (O_1249,N_24934,N_24852);
nor UO_1250 (O_1250,N_24765,N_24752);
xnor UO_1251 (O_1251,N_24783,N_24849);
xor UO_1252 (O_1252,N_24841,N_24822);
nor UO_1253 (O_1253,N_24847,N_24915);
and UO_1254 (O_1254,N_24775,N_24909);
nand UO_1255 (O_1255,N_24868,N_24939);
nor UO_1256 (O_1256,N_24952,N_24948);
nor UO_1257 (O_1257,N_24886,N_24772);
or UO_1258 (O_1258,N_24905,N_24882);
or UO_1259 (O_1259,N_24780,N_24874);
nor UO_1260 (O_1260,N_24842,N_24929);
and UO_1261 (O_1261,N_24957,N_24865);
xnor UO_1262 (O_1262,N_24969,N_24766);
nor UO_1263 (O_1263,N_24868,N_24879);
nor UO_1264 (O_1264,N_24804,N_24937);
or UO_1265 (O_1265,N_24883,N_24872);
and UO_1266 (O_1266,N_24838,N_24831);
nand UO_1267 (O_1267,N_24772,N_24909);
xnor UO_1268 (O_1268,N_24910,N_24942);
and UO_1269 (O_1269,N_24829,N_24825);
nand UO_1270 (O_1270,N_24909,N_24899);
or UO_1271 (O_1271,N_24921,N_24820);
and UO_1272 (O_1272,N_24861,N_24785);
nor UO_1273 (O_1273,N_24854,N_24848);
or UO_1274 (O_1274,N_24953,N_24864);
and UO_1275 (O_1275,N_24809,N_24783);
nor UO_1276 (O_1276,N_24981,N_24916);
and UO_1277 (O_1277,N_24755,N_24826);
or UO_1278 (O_1278,N_24863,N_24868);
xor UO_1279 (O_1279,N_24879,N_24884);
nor UO_1280 (O_1280,N_24872,N_24931);
and UO_1281 (O_1281,N_24832,N_24772);
and UO_1282 (O_1282,N_24978,N_24791);
nand UO_1283 (O_1283,N_24955,N_24887);
or UO_1284 (O_1284,N_24892,N_24777);
nor UO_1285 (O_1285,N_24990,N_24959);
nand UO_1286 (O_1286,N_24777,N_24768);
nand UO_1287 (O_1287,N_24802,N_24760);
and UO_1288 (O_1288,N_24899,N_24964);
or UO_1289 (O_1289,N_24870,N_24908);
xor UO_1290 (O_1290,N_24876,N_24960);
nor UO_1291 (O_1291,N_24903,N_24844);
or UO_1292 (O_1292,N_24895,N_24776);
or UO_1293 (O_1293,N_24970,N_24889);
nor UO_1294 (O_1294,N_24819,N_24871);
and UO_1295 (O_1295,N_24934,N_24882);
or UO_1296 (O_1296,N_24920,N_24914);
and UO_1297 (O_1297,N_24831,N_24871);
or UO_1298 (O_1298,N_24840,N_24846);
nand UO_1299 (O_1299,N_24770,N_24837);
and UO_1300 (O_1300,N_24823,N_24861);
and UO_1301 (O_1301,N_24890,N_24850);
xor UO_1302 (O_1302,N_24756,N_24757);
nor UO_1303 (O_1303,N_24949,N_24930);
nor UO_1304 (O_1304,N_24881,N_24761);
or UO_1305 (O_1305,N_24755,N_24781);
or UO_1306 (O_1306,N_24789,N_24913);
xnor UO_1307 (O_1307,N_24914,N_24844);
xnor UO_1308 (O_1308,N_24927,N_24833);
nand UO_1309 (O_1309,N_24975,N_24866);
or UO_1310 (O_1310,N_24969,N_24796);
and UO_1311 (O_1311,N_24792,N_24807);
or UO_1312 (O_1312,N_24971,N_24881);
nand UO_1313 (O_1313,N_24791,N_24933);
and UO_1314 (O_1314,N_24959,N_24874);
nor UO_1315 (O_1315,N_24808,N_24813);
nor UO_1316 (O_1316,N_24780,N_24750);
or UO_1317 (O_1317,N_24840,N_24963);
xnor UO_1318 (O_1318,N_24966,N_24848);
xnor UO_1319 (O_1319,N_24998,N_24991);
nand UO_1320 (O_1320,N_24972,N_24987);
nor UO_1321 (O_1321,N_24802,N_24843);
nand UO_1322 (O_1322,N_24876,N_24890);
nand UO_1323 (O_1323,N_24952,N_24961);
and UO_1324 (O_1324,N_24891,N_24933);
nand UO_1325 (O_1325,N_24851,N_24945);
or UO_1326 (O_1326,N_24890,N_24889);
and UO_1327 (O_1327,N_24969,N_24946);
xnor UO_1328 (O_1328,N_24954,N_24930);
nand UO_1329 (O_1329,N_24782,N_24811);
nand UO_1330 (O_1330,N_24949,N_24945);
nor UO_1331 (O_1331,N_24794,N_24824);
and UO_1332 (O_1332,N_24985,N_24877);
and UO_1333 (O_1333,N_24925,N_24751);
nand UO_1334 (O_1334,N_24760,N_24922);
nand UO_1335 (O_1335,N_24835,N_24915);
and UO_1336 (O_1336,N_24973,N_24947);
xnor UO_1337 (O_1337,N_24900,N_24863);
or UO_1338 (O_1338,N_24813,N_24931);
nand UO_1339 (O_1339,N_24853,N_24945);
nand UO_1340 (O_1340,N_24879,N_24945);
or UO_1341 (O_1341,N_24880,N_24772);
or UO_1342 (O_1342,N_24778,N_24959);
nand UO_1343 (O_1343,N_24890,N_24996);
nand UO_1344 (O_1344,N_24783,N_24990);
or UO_1345 (O_1345,N_24819,N_24905);
nand UO_1346 (O_1346,N_24839,N_24985);
nand UO_1347 (O_1347,N_24800,N_24750);
xnor UO_1348 (O_1348,N_24857,N_24779);
nand UO_1349 (O_1349,N_24975,N_24955);
xnor UO_1350 (O_1350,N_24800,N_24969);
xnor UO_1351 (O_1351,N_24831,N_24912);
and UO_1352 (O_1352,N_24909,N_24825);
or UO_1353 (O_1353,N_24795,N_24968);
or UO_1354 (O_1354,N_24824,N_24883);
and UO_1355 (O_1355,N_24897,N_24945);
or UO_1356 (O_1356,N_24789,N_24987);
and UO_1357 (O_1357,N_24999,N_24835);
and UO_1358 (O_1358,N_24996,N_24872);
and UO_1359 (O_1359,N_24817,N_24876);
nor UO_1360 (O_1360,N_24893,N_24908);
or UO_1361 (O_1361,N_24900,N_24818);
xor UO_1362 (O_1362,N_24846,N_24928);
nand UO_1363 (O_1363,N_24985,N_24974);
xnor UO_1364 (O_1364,N_24902,N_24848);
nor UO_1365 (O_1365,N_24844,N_24798);
nand UO_1366 (O_1366,N_24842,N_24897);
and UO_1367 (O_1367,N_24919,N_24896);
or UO_1368 (O_1368,N_24919,N_24831);
and UO_1369 (O_1369,N_24961,N_24943);
nor UO_1370 (O_1370,N_24951,N_24773);
nor UO_1371 (O_1371,N_24773,N_24849);
and UO_1372 (O_1372,N_24786,N_24835);
and UO_1373 (O_1373,N_24784,N_24985);
nand UO_1374 (O_1374,N_24833,N_24981);
and UO_1375 (O_1375,N_24796,N_24860);
nand UO_1376 (O_1376,N_24960,N_24898);
nand UO_1377 (O_1377,N_24829,N_24980);
and UO_1378 (O_1378,N_24771,N_24898);
and UO_1379 (O_1379,N_24914,N_24927);
xnor UO_1380 (O_1380,N_24898,N_24931);
nand UO_1381 (O_1381,N_24752,N_24782);
xnor UO_1382 (O_1382,N_24800,N_24970);
and UO_1383 (O_1383,N_24914,N_24755);
and UO_1384 (O_1384,N_24993,N_24755);
nor UO_1385 (O_1385,N_24968,N_24762);
or UO_1386 (O_1386,N_24985,N_24868);
xnor UO_1387 (O_1387,N_24912,N_24960);
nor UO_1388 (O_1388,N_24826,N_24969);
nor UO_1389 (O_1389,N_24950,N_24866);
nor UO_1390 (O_1390,N_24821,N_24843);
xor UO_1391 (O_1391,N_24786,N_24764);
or UO_1392 (O_1392,N_24975,N_24774);
nand UO_1393 (O_1393,N_24940,N_24753);
nand UO_1394 (O_1394,N_24830,N_24864);
or UO_1395 (O_1395,N_24791,N_24772);
nor UO_1396 (O_1396,N_24847,N_24905);
nor UO_1397 (O_1397,N_24891,N_24793);
xor UO_1398 (O_1398,N_24769,N_24789);
nand UO_1399 (O_1399,N_24815,N_24914);
and UO_1400 (O_1400,N_24768,N_24889);
or UO_1401 (O_1401,N_24812,N_24786);
or UO_1402 (O_1402,N_24762,N_24859);
or UO_1403 (O_1403,N_24929,N_24838);
or UO_1404 (O_1404,N_24815,N_24809);
nor UO_1405 (O_1405,N_24982,N_24871);
xnor UO_1406 (O_1406,N_24864,N_24952);
or UO_1407 (O_1407,N_24979,N_24759);
nor UO_1408 (O_1408,N_24775,N_24937);
or UO_1409 (O_1409,N_24772,N_24806);
nand UO_1410 (O_1410,N_24978,N_24944);
or UO_1411 (O_1411,N_24842,N_24762);
xnor UO_1412 (O_1412,N_24875,N_24999);
or UO_1413 (O_1413,N_24843,N_24977);
nor UO_1414 (O_1414,N_24836,N_24850);
or UO_1415 (O_1415,N_24872,N_24783);
xnor UO_1416 (O_1416,N_24941,N_24882);
xor UO_1417 (O_1417,N_24777,N_24828);
nand UO_1418 (O_1418,N_24993,N_24919);
nor UO_1419 (O_1419,N_24956,N_24769);
nor UO_1420 (O_1420,N_24908,N_24949);
nand UO_1421 (O_1421,N_24883,N_24827);
and UO_1422 (O_1422,N_24829,N_24853);
nand UO_1423 (O_1423,N_24887,N_24983);
nand UO_1424 (O_1424,N_24798,N_24861);
xor UO_1425 (O_1425,N_24787,N_24793);
or UO_1426 (O_1426,N_24901,N_24787);
nand UO_1427 (O_1427,N_24999,N_24985);
nand UO_1428 (O_1428,N_24879,N_24762);
nand UO_1429 (O_1429,N_24968,N_24956);
and UO_1430 (O_1430,N_24922,N_24765);
nor UO_1431 (O_1431,N_24806,N_24985);
xor UO_1432 (O_1432,N_24760,N_24993);
nand UO_1433 (O_1433,N_24907,N_24755);
xor UO_1434 (O_1434,N_24866,N_24838);
or UO_1435 (O_1435,N_24975,N_24762);
or UO_1436 (O_1436,N_24942,N_24919);
xor UO_1437 (O_1437,N_24838,N_24975);
nor UO_1438 (O_1438,N_24851,N_24813);
or UO_1439 (O_1439,N_24895,N_24821);
or UO_1440 (O_1440,N_24922,N_24751);
and UO_1441 (O_1441,N_24989,N_24984);
xor UO_1442 (O_1442,N_24883,N_24751);
xnor UO_1443 (O_1443,N_24891,N_24825);
xor UO_1444 (O_1444,N_24967,N_24875);
nor UO_1445 (O_1445,N_24828,N_24925);
xnor UO_1446 (O_1446,N_24949,N_24841);
nand UO_1447 (O_1447,N_24802,N_24881);
and UO_1448 (O_1448,N_24978,N_24980);
nand UO_1449 (O_1449,N_24921,N_24848);
xor UO_1450 (O_1450,N_24801,N_24850);
nand UO_1451 (O_1451,N_24950,N_24759);
and UO_1452 (O_1452,N_24978,N_24908);
xnor UO_1453 (O_1453,N_24949,N_24789);
nand UO_1454 (O_1454,N_24894,N_24994);
and UO_1455 (O_1455,N_24759,N_24914);
nor UO_1456 (O_1456,N_24844,N_24908);
and UO_1457 (O_1457,N_24990,N_24964);
nand UO_1458 (O_1458,N_24947,N_24884);
or UO_1459 (O_1459,N_24753,N_24750);
or UO_1460 (O_1460,N_24875,N_24903);
or UO_1461 (O_1461,N_24828,N_24884);
xor UO_1462 (O_1462,N_24795,N_24886);
nor UO_1463 (O_1463,N_24817,N_24803);
and UO_1464 (O_1464,N_24801,N_24979);
nand UO_1465 (O_1465,N_24814,N_24955);
xnor UO_1466 (O_1466,N_24984,N_24826);
and UO_1467 (O_1467,N_24776,N_24933);
nand UO_1468 (O_1468,N_24842,N_24802);
nand UO_1469 (O_1469,N_24956,N_24805);
xor UO_1470 (O_1470,N_24825,N_24950);
or UO_1471 (O_1471,N_24815,N_24893);
xor UO_1472 (O_1472,N_24872,N_24897);
xnor UO_1473 (O_1473,N_24754,N_24821);
or UO_1474 (O_1474,N_24803,N_24890);
or UO_1475 (O_1475,N_24929,N_24765);
nand UO_1476 (O_1476,N_24977,N_24759);
xnor UO_1477 (O_1477,N_24821,N_24930);
xnor UO_1478 (O_1478,N_24941,N_24932);
or UO_1479 (O_1479,N_24791,N_24997);
nand UO_1480 (O_1480,N_24918,N_24943);
xnor UO_1481 (O_1481,N_24788,N_24833);
or UO_1482 (O_1482,N_24917,N_24860);
xor UO_1483 (O_1483,N_24952,N_24974);
and UO_1484 (O_1484,N_24883,N_24802);
or UO_1485 (O_1485,N_24958,N_24940);
and UO_1486 (O_1486,N_24756,N_24855);
nand UO_1487 (O_1487,N_24881,N_24827);
xnor UO_1488 (O_1488,N_24771,N_24891);
xor UO_1489 (O_1489,N_24903,N_24857);
xnor UO_1490 (O_1490,N_24780,N_24802);
nor UO_1491 (O_1491,N_24965,N_24853);
xor UO_1492 (O_1492,N_24780,N_24987);
nor UO_1493 (O_1493,N_24860,N_24902);
nor UO_1494 (O_1494,N_24863,N_24943);
xor UO_1495 (O_1495,N_24981,N_24776);
nor UO_1496 (O_1496,N_24870,N_24992);
nor UO_1497 (O_1497,N_24984,N_24851);
nor UO_1498 (O_1498,N_24836,N_24824);
xor UO_1499 (O_1499,N_24784,N_24791);
nand UO_1500 (O_1500,N_24785,N_24799);
or UO_1501 (O_1501,N_24978,N_24975);
nand UO_1502 (O_1502,N_24864,N_24812);
nand UO_1503 (O_1503,N_24952,N_24918);
and UO_1504 (O_1504,N_24981,N_24837);
or UO_1505 (O_1505,N_24812,N_24763);
nand UO_1506 (O_1506,N_24820,N_24769);
nor UO_1507 (O_1507,N_24968,N_24944);
xnor UO_1508 (O_1508,N_24949,N_24812);
and UO_1509 (O_1509,N_24771,N_24912);
xor UO_1510 (O_1510,N_24757,N_24991);
or UO_1511 (O_1511,N_24983,N_24842);
xnor UO_1512 (O_1512,N_24787,N_24769);
nand UO_1513 (O_1513,N_24917,N_24952);
nand UO_1514 (O_1514,N_24827,N_24921);
or UO_1515 (O_1515,N_24932,N_24873);
and UO_1516 (O_1516,N_24839,N_24857);
and UO_1517 (O_1517,N_24943,N_24804);
and UO_1518 (O_1518,N_24985,N_24990);
nand UO_1519 (O_1519,N_24991,N_24922);
xnor UO_1520 (O_1520,N_24849,N_24788);
nor UO_1521 (O_1521,N_24781,N_24945);
nand UO_1522 (O_1522,N_24992,N_24897);
or UO_1523 (O_1523,N_24772,N_24915);
xnor UO_1524 (O_1524,N_24962,N_24758);
nand UO_1525 (O_1525,N_24809,N_24813);
nor UO_1526 (O_1526,N_24783,N_24961);
nand UO_1527 (O_1527,N_24892,N_24993);
and UO_1528 (O_1528,N_24815,N_24867);
nand UO_1529 (O_1529,N_24838,N_24861);
xnor UO_1530 (O_1530,N_24782,N_24923);
xnor UO_1531 (O_1531,N_24949,N_24785);
and UO_1532 (O_1532,N_24941,N_24962);
nand UO_1533 (O_1533,N_24964,N_24839);
nor UO_1534 (O_1534,N_24835,N_24763);
and UO_1535 (O_1535,N_24750,N_24901);
or UO_1536 (O_1536,N_24808,N_24825);
nor UO_1537 (O_1537,N_24849,N_24943);
nand UO_1538 (O_1538,N_24821,N_24974);
nand UO_1539 (O_1539,N_24886,N_24827);
nor UO_1540 (O_1540,N_24962,N_24997);
nand UO_1541 (O_1541,N_24816,N_24822);
xor UO_1542 (O_1542,N_24794,N_24773);
nor UO_1543 (O_1543,N_24788,N_24774);
nor UO_1544 (O_1544,N_24901,N_24871);
xnor UO_1545 (O_1545,N_24818,N_24830);
nand UO_1546 (O_1546,N_24969,N_24967);
and UO_1547 (O_1547,N_24777,N_24850);
nand UO_1548 (O_1548,N_24779,N_24750);
nand UO_1549 (O_1549,N_24756,N_24761);
nand UO_1550 (O_1550,N_24801,N_24901);
or UO_1551 (O_1551,N_24998,N_24812);
xor UO_1552 (O_1552,N_24993,N_24996);
xnor UO_1553 (O_1553,N_24852,N_24810);
nand UO_1554 (O_1554,N_24942,N_24939);
nor UO_1555 (O_1555,N_24816,N_24927);
nand UO_1556 (O_1556,N_24879,N_24814);
nand UO_1557 (O_1557,N_24973,N_24771);
xnor UO_1558 (O_1558,N_24912,N_24958);
nor UO_1559 (O_1559,N_24827,N_24995);
xor UO_1560 (O_1560,N_24880,N_24820);
nor UO_1561 (O_1561,N_24941,N_24885);
and UO_1562 (O_1562,N_24768,N_24857);
or UO_1563 (O_1563,N_24996,N_24897);
and UO_1564 (O_1564,N_24846,N_24753);
nor UO_1565 (O_1565,N_24929,N_24974);
nor UO_1566 (O_1566,N_24829,N_24989);
xor UO_1567 (O_1567,N_24965,N_24891);
nor UO_1568 (O_1568,N_24791,N_24777);
nand UO_1569 (O_1569,N_24892,N_24972);
xor UO_1570 (O_1570,N_24763,N_24898);
and UO_1571 (O_1571,N_24901,N_24970);
and UO_1572 (O_1572,N_24948,N_24923);
or UO_1573 (O_1573,N_24882,N_24865);
xnor UO_1574 (O_1574,N_24902,N_24908);
nor UO_1575 (O_1575,N_24907,N_24777);
nor UO_1576 (O_1576,N_24978,N_24947);
nand UO_1577 (O_1577,N_24980,N_24979);
xnor UO_1578 (O_1578,N_24945,N_24762);
nand UO_1579 (O_1579,N_24987,N_24975);
or UO_1580 (O_1580,N_24861,N_24845);
nor UO_1581 (O_1581,N_24938,N_24947);
xor UO_1582 (O_1582,N_24783,N_24877);
xnor UO_1583 (O_1583,N_24891,N_24774);
xnor UO_1584 (O_1584,N_24828,N_24856);
nand UO_1585 (O_1585,N_24855,N_24788);
and UO_1586 (O_1586,N_24835,N_24897);
xnor UO_1587 (O_1587,N_24957,N_24817);
and UO_1588 (O_1588,N_24988,N_24806);
xor UO_1589 (O_1589,N_24924,N_24772);
nand UO_1590 (O_1590,N_24987,N_24844);
xnor UO_1591 (O_1591,N_24809,N_24931);
xor UO_1592 (O_1592,N_24857,N_24900);
nor UO_1593 (O_1593,N_24865,N_24820);
xor UO_1594 (O_1594,N_24805,N_24808);
nor UO_1595 (O_1595,N_24886,N_24764);
and UO_1596 (O_1596,N_24876,N_24974);
nor UO_1597 (O_1597,N_24889,N_24805);
xnor UO_1598 (O_1598,N_24982,N_24900);
xor UO_1599 (O_1599,N_24870,N_24834);
and UO_1600 (O_1600,N_24982,N_24825);
or UO_1601 (O_1601,N_24838,N_24973);
nor UO_1602 (O_1602,N_24754,N_24841);
and UO_1603 (O_1603,N_24815,N_24998);
nand UO_1604 (O_1604,N_24792,N_24925);
and UO_1605 (O_1605,N_24944,N_24800);
xnor UO_1606 (O_1606,N_24868,N_24867);
xnor UO_1607 (O_1607,N_24785,N_24756);
nor UO_1608 (O_1608,N_24962,N_24836);
xnor UO_1609 (O_1609,N_24769,N_24878);
and UO_1610 (O_1610,N_24980,N_24773);
and UO_1611 (O_1611,N_24761,N_24778);
nor UO_1612 (O_1612,N_24792,N_24758);
nand UO_1613 (O_1613,N_24781,N_24761);
or UO_1614 (O_1614,N_24954,N_24976);
or UO_1615 (O_1615,N_24941,N_24849);
or UO_1616 (O_1616,N_24779,N_24815);
xnor UO_1617 (O_1617,N_24808,N_24886);
nor UO_1618 (O_1618,N_24860,N_24918);
xor UO_1619 (O_1619,N_24812,N_24772);
or UO_1620 (O_1620,N_24801,N_24870);
nand UO_1621 (O_1621,N_24769,N_24854);
and UO_1622 (O_1622,N_24876,N_24972);
nor UO_1623 (O_1623,N_24984,N_24891);
nor UO_1624 (O_1624,N_24830,N_24931);
or UO_1625 (O_1625,N_24829,N_24778);
xor UO_1626 (O_1626,N_24955,N_24822);
and UO_1627 (O_1627,N_24755,N_24888);
and UO_1628 (O_1628,N_24992,N_24924);
nand UO_1629 (O_1629,N_24760,N_24861);
or UO_1630 (O_1630,N_24824,N_24873);
nand UO_1631 (O_1631,N_24764,N_24903);
and UO_1632 (O_1632,N_24770,N_24810);
nand UO_1633 (O_1633,N_24933,N_24881);
or UO_1634 (O_1634,N_24978,N_24937);
and UO_1635 (O_1635,N_24859,N_24876);
and UO_1636 (O_1636,N_24816,N_24769);
nand UO_1637 (O_1637,N_24831,N_24984);
or UO_1638 (O_1638,N_24799,N_24872);
xnor UO_1639 (O_1639,N_24833,N_24860);
nor UO_1640 (O_1640,N_24930,N_24773);
nand UO_1641 (O_1641,N_24776,N_24816);
or UO_1642 (O_1642,N_24913,N_24946);
nand UO_1643 (O_1643,N_24871,N_24913);
and UO_1644 (O_1644,N_24808,N_24961);
and UO_1645 (O_1645,N_24870,N_24817);
nand UO_1646 (O_1646,N_24846,N_24921);
nand UO_1647 (O_1647,N_24974,N_24751);
nand UO_1648 (O_1648,N_24814,N_24985);
nand UO_1649 (O_1649,N_24910,N_24756);
xnor UO_1650 (O_1650,N_24751,N_24924);
nand UO_1651 (O_1651,N_24936,N_24843);
nand UO_1652 (O_1652,N_24914,N_24886);
xor UO_1653 (O_1653,N_24994,N_24996);
and UO_1654 (O_1654,N_24785,N_24839);
or UO_1655 (O_1655,N_24776,N_24909);
nand UO_1656 (O_1656,N_24862,N_24907);
nand UO_1657 (O_1657,N_24778,N_24890);
or UO_1658 (O_1658,N_24905,N_24852);
nor UO_1659 (O_1659,N_24927,N_24806);
or UO_1660 (O_1660,N_24913,N_24988);
nand UO_1661 (O_1661,N_24831,N_24922);
and UO_1662 (O_1662,N_24834,N_24815);
nand UO_1663 (O_1663,N_24783,N_24913);
nor UO_1664 (O_1664,N_24757,N_24761);
nand UO_1665 (O_1665,N_24989,N_24999);
xnor UO_1666 (O_1666,N_24908,N_24952);
nand UO_1667 (O_1667,N_24869,N_24882);
or UO_1668 (O_1668,N_24884,N_24793);
xor UO_1669 (O_1669,N_24979,N_24981);
and UO_1670 (O_1670,N_24958,N_24770);
or UO_1671 (O_1671,N_24868,N_24840);
xnor UO_1672 (O_1672,N_24750,N_24832);
xnor UO_1673 (O_1673,N_24856,N_24894);
nor UO_1674 (O_1674,N_24829,N_24943);
and UO_1675 (O_1675,N_24931,N_24842);
nor UO_1676 (O_1676,N_24889,N_24834);
xor UO_1677 (O_1677,N_24862,N_24904);
nor UO_1678 (O_1678,N_24917,N_24813);
nand UO_1679 (O_1679,N_24858,N_24816);
and UO_1680 (O_1680,N_24936,N_24891);
nand UO_1681 (O_1681,N_24948,N_24758);
or UO_1682 (O_1682,N_24915,N_24830);
nor UO_1683 (O_1683,N_24877,N_24840);
or UO_1684 (O_1684,N_24997,N_24986);
xnor UO_1685 (O_1685,N_24988,N_24939);
xor UO_1686 (O_1686,N_24784,N_24776);
or UO_1687 (O_1687,N_24866,N_24986);
and UO_1688 (O_1688,N_24931,N_24761);
nor UO_1689 (O_1689,N_24908,N_24898);
or UO_1690 (O_1690,N_24848,N_24889);
xnor UO_1691 (O_1691,N_24951,N_24980);
or UO_1692 (O_1692,N_24797,N_24759);
xnor UO_1693 (O_1693,N_24992,N_24753);
or UO_1694 (O_1694,N_24758,N_24816);
xor UO_1695 (O_1695,N_24816,N_24923);
nand UO_1696 (O_1696,N_24895,N_24780);
xnor UO_1697 (O_1697,N_24835,N_24914);
and UO_1698 (O_1698,N_24885,N_24899);
and UO_1699 (O_1699,N_24829,N_24784);
xor UO_1700 (O_1700,N_24824,N_24922);
or UO_1701 (O_1701,N_24964,N_24777);
nand UO_1702 (O_1702,N_24992,N_24984);
nand UO_1703 (O_1703,N_24889,N_24856);
nor UO_1704 (O_1704,N_24910,N_24859);
nor UO_1705 (O_1705,N_24850,N_24789);
nand UO_1706 (O_1706,N_24961,N_24992);
xnor UO_1707 (O_1707,N_24782,N_24877);
nand UO_1708 (O_1708,N_24799,N_24800);
xnor UO_1709 (O_1709,N_24877,N_24832);
nor UO_1710 (O_1710,N_24842,N_24974);
nand UO_1711 (O_1711,N_24945,N_24890);
or UO_1712 (O_1712,N_24962,N_24996);
and UO_1713 (O_1713,N_24785,N_24881);
nor UO_1714 (O_1714,N_24998,N_24857);
nor UO_1715 (O_1715,N_24911,N_24886);
nand UO_1716 (O_1716,N_24812,N_24879);
nand UO_1717 (O_1717,N_24870,N_24757);
or UO_1718 (O_1718,N_24907,N_24895);
xor UO_1719 (O_1719,N_24791,N_24869);
xnor UO_1720 (O_1720,N_24861,N_24935);
nor UO_1721 (O_1721,N_24852,N_24981);
nor UO_1722 (O_1722,N_24844,N_24921);
nand UO_1723 (O_1723,N_24856,N_24906);
and UO_1724 (O_1724,N_24872,N_24781);
xor UO_1725 (O_1725,N_24962,N_24824);
nor UO_1726 (O_1726,N_24956,N_24764);
nand UO_1727 (O_1727,N_24848,N_24980);
nor UO_1728 (O_1728,N_24999,N_24907);
and UO_1729 (O_1729,N_24862,N_24919);
or UO_1730 (O_1730,N_24941,N_24848);
nor UO_1731 (O_1731,N_24927,N_24891);
and UO_1732 (O_1732,N_24989,N_24951);
xor UO_1733 (O_1733,N_24807,N_24805);
and UO_1734 (O_1734,N_24797,N_24845);
nor UO_1735 (O_1735,N_24804,N_24985);
xnor UO_1736 (O_1736,N_24885,N_24866);
xor UO_1737 (O_1737,N_24880,N_24909);
and UO_1738 (O_1738,N_24759,N_24982);
xnor UO_1739 (O_1739,N_24909,N_24888);
and UO_1740 (O_1740,N_24801,N_24790);
xnor UO_1741 (O_1741,N_24796,N_24805);
nor UO_1742 (O_1742,N_24915,N_24782);
nor UO_1743 (O_1743,N_24916,N_24769);
nor UO_1744 (O_1744,N_24965,N_24904);
and UO_1745 (O_1745,N_24751,N_24988);
xor UO_1746 (O_1746,N_24817,N_24925);
nor UO_1747 (O_1747,N_24836,N_24989);
xor UO_1748 (O_1748,N_24968,N_24755);
or UO_1749 (O_1749,N_24995,N_24756);
or UO_1750 (O_1750,N_24914,N_24830);
nand UO_1751 (O_1751,N_24780,N_24990);
nand UO_1752 (O_1752,N_24923,N_24935);
nor UO_1753 (O_1753,N_24977,N_24862);
nor UO_1754 (O_1754,N_24766,N_24991);
xnor UO_1755 (O_1755,N_24811,N_24774);
xnor UO_1756 (O_1756,N_24932,N_24779);
nand UO_1757 (O_1757,N_24964,N_24874);
and UO_1758 (O_1758,N_24900,N_24755);
nor UO_1759 (O_1759,N_24826,N_24777);
and UO_1760 (O_1760,N_24978,N_24916);
nand UO_1761 (O_1761,N_24850,N_24791);
nor UO_1762 (O_1762,N_24853,N_24765);
and UO_1763 (O_1763,N_24958,N_24752);
xor UO_1764 (O_1764,N_24752,N_24798);
or UO_1765 (O_1765,N_24922,N_24921);
xnor UO_1766 (O_1766,N_24969,N_24786);
xnor UO_1767 (O_1767,N_24937,N_24807);
nand UO_1768 (O_1768,N_24854,N_24939);
xor UO_1769 (O_1769,N_24949,N_24951);
or UO_1770 (O_1770,N_24762,N_24985);
nand UO_1771 (O_1771,N_24948,N_24956);
or UO_1772 (O_1772,N_24786,N_24895);
nor UO_1773 (O_1773,N_24954,N_24859);
and UO_1774 (O_1774,N_24898,N_24874);
nand UO_1775 (O_1775,N_24865,N_24831);
and UO_1776 (O_1776,N_24811,N_24990);
nand UO_1777 (O_1777,N_24938,N_24974);
nor UO_1778 (O_1778,N_24809,N_24806);
nand UO_1779 (O_1779,N_24752,N_24920);
nor UO_1780 (O_1780,N_24937,N_24808);
and UO_1781 (O_1781,N_24757,N_24863);
nand UO_1782 (O_1782,N_24907,N_24758);
and UO_1783 (O_1783,N_24852,N_24876);
xnor UO_1784 (O_1784,N_24913,N_24768);
and UO_1785 (O_1785,N_24819,N_24920);
xnor UO_1786 (O_1786,N_24878,N_24855);
and UO_1787 (O_1787,N_24957,N_24880);
nor UO_1788 (O_1788,N_24936,N_24912);
xor UO_1789 (O_1789,N_24845,N_24985);
and UO_1790 (O_1790,N_24905,N_24947);
and UO_1791 (O_1791,N_24809,N_24801);
nor UO_1792 (O_1792,N_24939,N_24979);
xor UO_1793 (O_1793,N_24930,N_24932);
nand UO_1794 (O_1794,N_24765,N_24862);
and UO_1795 (O_1795,N_24896,N_24982);
xor UO_1796 (O_1796,N_24864,N_24888);
nand UO_1797 (O_1797,N_24947,N_24782);
or UO_1798 (O_1798,N_24960,N_24770);
and UO_1799 (O_1799,N_24897,N_24762);
or UO_1800 (O_1800,N_24797,N_24914);
xor UO_1801 (O_1801,N_24795,N_24939);
or UO_1802 (O_1802,N_24771,N_24845);
nand UO_1803 (O_1803,N_24975,N_24983);
xnor UO_1804 (O_1804,N_24917,N_24929);
nand UO_1805 (O_1805,N_24857,N_24879);
nor UO_1806 (O_1806,N_24979,N_24938);
or UO_1807 (O_1807,N_24912,N_24858);
and UO_1808 (O_1808,N_24934,N_24797);
or UO_1809 (O_1809,N_24816,N_24990);
nand UO_1810 (O_1810,N_24835,N_24965);
nand UO_1811 (O_1811,N_24884,N_24848);
nor UO_1812 (O_1812,N_24966,N_24803);
or UO_1813 (O_1813,N_24923,N_24938);
xor UO_1814 (O_1814,N_24840,N_24849);
nand UO_1815 (O_1815,N_24930,N_24933);
or UO_1816 (O_1816,N_24809,N_24901);
nor UO_1817 (O_1817,N_24834,N_24923);
or UO_1818 (O_1818,N_24924,N_24935);
xor UO_1819 (O_1819,N_24887,N_24926);
xor UO_1820 (O_1820,N_24813,N_24870);
or UO_1821 (O_1821,N_24953,N_24947);
and UO_1822 (O_1822,N_24913,N_24973);
nor UO_1823 (O_1823,N_24799,N_24894);
nand UO_1824 (O_1824,N_24770,N_24790);
and UO_1825 (O_1825,N_24969,N_24954);
nand UO_1826 (O_1826,N_24908,N_24875);
and UO_1827 (O_1827,N_24864,N_24905);
and UO_1828 (O_1828,N_24909,N_24802);
nand UO_1829 (O_1829,N_24965,N_24912);
nand UO_1830 (O_1830,N_24866,N_24946);
xor UO_1831 (O_1831,N_24988,N_24935);
nand UO_1832 (O_1832,N_24897,N_24807);
and UO_1833 (O_1833,N_24777,N_24773);
nand UO_1834 (O_1834,N_24818,N_24783);
and UO_1835 (O_1835,N_24978,N_24847);
or UO_1836 (O_1836,N_24997,N_24767);
xor UO_1837 (O_1837,N_24760,N_24854);
nand UO_1838 (O_1838,N_24987,N_24949);
xor UO_1839 (O_1839,N_24850,N_24774);
nand UO_1840 (O_1840,N_24802,N_24798);
and UO_1841 (O_1841,N_24790,N_24780);
xnor UO_1842 (O_1842,N_24988,N_24844);
or UO_1843 (O_1843,N_24800,N_24850);
and UO_1844 (O_1844,N_24750,N_24792);
or UO_1845 (O_1845,N_24816,N_24787);
xnor UO_1846 (O_1846,N_24886,N_24866);
xor UO_1847 (O_1847,N_24840,N_24809);
nand UO_1848 (O_1848,N_24899,N_24850);
xnor UO_1849 (O_1849,N_24758,N_24903);
nor UO_1850 (O_1850,N_24883,N_24937);
nor UO_1851 (O_1851,N_24783,N_24768);
nand UO_1852 (O_1852,N_24841,N_24799);
and UO_1853 (O_1853,N_24806,N_24958);
xor UO_1854 (O_1854,N_24819,N_24953);
and UO_1855 (O_1855,N_24967,N_24900);
xnor UO_1856 (O_1856,N_24977,N_24783);
or UO_1857 (O_1857,N_24993,N_24906);
or UO_1858 (O_1858,N_24807,N_24835);
and UO_1859 (O_1859,N_24895,N_24758);
and UO_1860 (O_1860,N_24878,N_24799);
nand UO_1861 (O_1861,N_24979,N_24864);
xor UO_1862 (O_1862,N_24890,N_24982);
nand UO_1863 (O_1863,N_24893,N_24854);
or UO_1864 (O_1864,N_24923,N_24940);
nor UO_1865 (O_1865,N_24890,N_24785);
and UO_1866 (O_1866,N_24781,N_24987);
or UO_1867 (O_1867,N_24985,N_24984);
nand UO_1868 (O_1868,N_24888,N_24762);
nand UO_1869 (O_1869,N_24982,N_24958);
nor UO_1870 (O_1870,N_24843,N_24942);
nand UO_1871 (O_1871,N_24954,N_24915);
nor UO_1872 (O_1872,N_24848,N_24830);
nand UO_1873 (O_1873,N_24807,N_24781);
and UO_1874 (O_1874,N_24893,N_24998);
nand UO_1875 (O_1875,N_24845,N_24878);
or UO_1876 (O_1876,N_24784,N_24813);
xor UO_1877 (O_1877,N_24836,N_24999);
or UO_1878 (O_1878,N_24779,N_24937);
nand UO_1879 (O_1879,N_24923,N_24882);
xor UO_1880 (O_1880,N_24916,N_24947);
xnor UO_1881 (O_1881,N_24876,N_24780);
or UO_1882 (O_1882,N_24916,N_24959);
or UO_1883 (O_1883,N_24816,N_24911);
nand UO_1884 (O_1884,N_24933,N_24918);
nor UO_1885 (O_1885,N_24765,N_24969);
xnor UO_1886 (O_1886,N_24770,N_24860);
and UO_1887 (O_1887,N_24975,N_24899);
nand UO_1888 (O_1888,N_24906,N_24893);
and UO_1889 (O_1889,N_24968,N_24786);
xnor UO_1890 (O_1890,N_24815,N_24773);
nand UO_1891 (O_1891,N_24758,N_24784);
or UO_1892 (O_1892,N_24832,N_24860);
xor UO_1893 (O_1893,N_24990,N_24897);
nor UO_1894 (O_1894,N_24958,N_24844);
or UO_1895 (O_1895,N_24938,N_24956);
xor UO_1896 (O_1896,N_24823,N_24995);
and UO_1897 (O_1897,N_24762,N_24873);
nand UO_1898 (O_1898,N_24935,N_24758);
xor UO_1899 (O_1899,N_24867,N_24913);
nand UO_1900 (O_1900,N_24886,N_24899);
and UO_1901 (O_1901,N_24904,N_24881);
xor UO_1902 (O_1902,N_24912,N_24896);
nand UO_1903 (O_1903,N_24789,N_24980);
or UO_1904 (O_1904,N_24966,N_24926);
xnor UO_1905 (O_1905,N_24912,N_24778);
nor UO_1906 (O_1906,N_24759,N_24801);
or UO_1907 (O_1907,N_24766,N_24916);
nand UO_1908 (O_1908,N_24853,N_24839);
nand UO_1909 (O_1909,N_24901,N_24876);
and UO_1910 (O_1910,N_24946,N_24944);
nand UO_1911 (O_1911,N_24918,N_24759);
or UO_1912 (O_1912,N_24982,N_24926);
nor UO_1913 (O_1913,N_24824,N_24760);
or UO_1914 (O_1914,N_24863,N_24866);
nand UO_1915 (O_1915,N_24942,N_24923);
or UO_1916 (O_1916,N_24876,N_24956);
and UO_1917 (O_1917,N_24991,N_24964);
nand UO_1918 (O_1918,N_24787,N_24923);
nor UO_1919 (O_1919,N_24803,N_24825);
xnor UO_1920 (O_1920,N_24818,N_24908);
and UO_1921 (O_1921,N_24906,N_24977);
nand UO_1922 (O_1922,N_24931,N_24773);
nor UO_1923 (O_1923,N_24811,N_24883);
xnor UO_1924 (O_1924,N_24853,N_24985);
nor UO_1925 (O_1925,N_24970,N_24787);
nor UO_1926 (O_1926,N_24882,N_24962);
nand UO_1927 (O_1927,N_24979,N_24755);
and UO_1928 (O_1928,N_24754,N_24807);
nor UO_1929 (O_1929,N_24788,N_24968);
xor UO_1930 (O_1930,N_24957,N_24846);
or UO_1931 (O_1931,N_24840,N_24976);
nor UO_1932 (O_1932,N_24770,N_24822);
nand UO_1933 (O_1933,N_24883,N_24828);
and UO_1934 (O_1934,N_24902,N_24776);
nor UO_1935 (O_1935,N_24902,N_24903);
and UO_1936 (O_1936,N_24937,N_24870);
nand UO_1937 (O_1937,N_24848,N_24948);
nand UO_1938 (O_1938,N_24899,N_24783);
or UO_1939 (O_1939,N_24799,N_24820);
xnor UO_1940 (O_1940,N_24989,N_24936);
or UO_1941 (O_1941,N_24850,N_24980);
or UO_1942 (O_1942,N_24797,N_24788);
nor UO_1943 (O_1943,N_24833,N_24852);
and UO_1944 (O_1944,N_24994,N_24910);
and UO_1945 (O_1945,N_24990,N_24792);
nor UO_1946 (O_1946,N_24817,N_24998);
nor UO_1947 (O_1947,N_24849,N_24980);
nand UO_1948 (O_1948,N_24891,N_24798);
or UO_1949 (O_1949,N_24763,N_24987);
nor UO_1950 (O_1950,N_24800,N_24830);
nor UO_1951 (O_1951,N_24751,N_24826);
or UO_1952 (O_1952,N_24985,N_24857);
or UO_1953 (O_1953,N_24942,N_24861);
nor UO_1954 (O_1954,N_24797,N_24867);
nand UO_1955 (O_1955,N_24795,N_24877);
nor UO_1956 (O_1956,N_24833,N_24758);
or UO_1957 (O_1957,N_24992,N_24916);
xor UO_1958 (O_1958,N_24906,N_24999);
nand UO_1959 (O_1959,N_24803,N_24978);
or UO_1960 (O_1960,N_24844,N_24820);
or UO_1961 (O_1961,N_24922,N_24802);
xor UO_1962 (O_1962,N_24751,N_24841);
nand UO_1963 (O_1963,N_24819,N_24854);
nand UO_1964 (O_1964,N_24807,N_24971);
nor UO_1965 (O_1965,N_24906,N_24806);
xnor UO_1966 (O_1966,N_24935,N_24830);
nand UO_1967 (O_1967,N_24885,N_24975);
nor UO_1968 (O_1968,N_24911,N_24759);
or UO_1969 (O_1969,N_24763,N_24952);
nor UO_1970 (O_1970,N_24835,N_24996);
nand UO_1971 (O_1971,N_24887,N_24828);
and UO_1972 (O_1972,N_24884,N_24982);
nand UO_1973 (O_1973,N_24881,N_24959);
and UO_1974 (O_1974,N_24888,N_24758);
or UO_1975 (O_1975,N_24838,N_24820);
nor UO_1976 (O_1976,N_24779,N_24766);
and UO_1977 (O_1977,N_24766,N_24947);
and UO_1978 (O_1978,N_24966,N_24838);
xor UO_1979 (O_1979,N_24854,N_24919);
nor UO_1980 (O_1980,N_24950,N_24980);
nor UO_1981 (O_1981,N_24949,N_24802);
or UO_1982 (O_1982,N_24950,N_24787);
nor UO_1983 (O_1983,N_24861,N_24884);
xor UO_1984 (O_1984,N_24921,N_24930);
and UO_1985 (O_1985,N_24882,N_24918);
or UO_1986 (O_1986,N_24893,N_24793);
and UO_1987 (O_1987,N_24799,N_24752);
nor UO_1988 (O_1988,N_24904,N_24827);
nand UO_1989 (O_1989,N_24761,N_24887);
xnor UO_1990 (O_1990,N_24968,N_24982);
xnor UO_1991 (O_1991,N_24866,N_24881);
nor UO_1992 (O_1992,N_24781,N_24909);
nand UO_1993 (O_1993,N_24848,N_24985);
nand UO_1994 (O_1994,N_24788,N_24947);
nand UO_1995 (O_1995,N_24904,N_24817);
or UO_1996 (O_1996,N_24942,N_24970);
nand UO_1997 (O_1997,N_24958,N_24837);
nand UO_1998 (O_1998,N_24848,N_24779);
nand UO_1999 (O_1999,N_24964,N_24870);
nand UO_2000 (O_2000,N_24873,N_24768);
xor UO_2001 (O_2001,N_24786,N_24964);
and UO_2002 (O_2002,N_24922,N_24819);
xnor UO_2003 (O_2003,N_24770,N_24911);
xor UO_2004 (O_2004,N_24896,N_24852);
nand UO_2005 (O_2005,N_24916,N_24927);
xor UO_2006 (O_2006,N_24892,N_24956);
nor UO_2007 (O_2007,N_24997,N_24801);
and UO_2008 (O_2008,N_24844,N_24923);
xnor UO_2009 (O_2009,N_24876,N_24924);
xnor UO_2010 (O_2010,N_24915,N_24895);
nor UO_2011 (O_2011,N_24822,N_24900);
xnor UO_2012 (O_2012,N_24833,N_24922);
and UO_2013 (O_2013,N_24851,N_24765);
nand UO_2014 (O_2014,N_24827,N_24780);
or UO_2015 (O_2015,N_24968,N_24988);
or UO_2016 (O_2016,N_24770,N_24999);
or UO_2017 (O_2017,N_24763,N_24876);
or UO_2018 (O_2018,N_24921,N_24767);
or UO_2019 (O_2019,N_24838,N_24799);
nor UO_2020 (O_2020,N_24943,N_24972);
or UO_2021 (O_2021,N_24893,N_24938);
xor UO_2022 (O_2022,N_24863,N_24867);
xor UO_2023 (O_2023,N_24890,N_24953);
nand UO_2024 (O_2024,N_24931,N_24794);
nand UO_2025 (O_2025,N_24834,N_24838);
and UO_2026 (O_2026,N_24973,N_24883);
nor UO_2027 (O_2027,N_24882,N_24790);
xor UO_2028 (O_2028,N_24927,N_24962);
or UO_2029 (O_2029,N_24852,N_24752);
and UO_2030 (O_2030,N_24881,N_24853);
and UO_2031 (O_2031,N_24797,N_24896);
or UO_2032 (O_2032,N_24832,N_24783);
and UO_2033 (O_2033,N_24912,N_24986);
or UO_2034 (O_2034,N_24897,N_24806);
and UO_2035 (O_2035,N_24940,N_24842);
nor UO_2036 (O_2036,N_24829,N_24838);
and UO_2037 (O_2037,N_24812,N_24962);
nor UO_2038 (O_2038,N_24988,N_24899);
nand UO_2039 (O_2039,N_24941,N_24776);
nor UO_2040 (O_2040,N_24761,N_24750);
xor UO_2041 (O_2041,N_24816,N_24801);
or UO_2042 (O_2042,N_24850,N_24970);
and UO_2043 (O_2043,N_24804,N_24928);
nor UO_2044 (O_2044,N_24916,N_24764);
or UO_2045 (O_2045,N_24975,N_24965);
nand UO_2046 (O_2046,N_24919,N_24755);
and UO_2047 (O_2047,N_24856,N_24804);
and UO_2048 (O_2048,N_24951,N_24946);
or UO_2049 (O_2049,N_24957,N_24908);
or UO_2050 (O_2050,N_24927,N_24787);
nand UO_2051 (O_2051,N_24868,N_24757);
and UO_2052 (O_2052,N_24953,N_24849);
nand UO_2053 (O_2053,N_24981,N_24763);
or UO_2054 (O_2054,N_24979,N_24943);
and UO_2055 (O_2055,N_24795,N_24829);
nor UO_2056 (O_2056,N_24996,N_24865);
nand UO_2057 (O_2057,N_24890,N_24821);
or UO_2058 (O_2058,N_24761,N_24937);
and UO_2059 (O_2059,N_24798,N_24975);
or UO_2060 (O_2060,N_24966,N_24794);
nand UO_2061 (O_2061,N_24791,N_24895);
xor UO_2062 (O_2062,N_24896,N_24784);
nor UO_2063 (O_2063,N_24857,N_24932);
nand UO_2064 (O_2064,N_24983,N_24822);
or UO_2065 (O_2065,N_24812,N_24835);
and UO_2066 (O_2066,N_24995,N_24977);
or UO_2067 (O_2067,N_24822,N_24780);
xnor UO_2068 (O_2068,N_24918,N_24905);
and UO_2069 (O_2069,N_24813,N_24841);
xnor UO_2070 (O_2070,N_24906,N_24775);
nand UO_2071 (O_2071,N_24755,N_24855);
xnor UO_2072 (O_2072,N_24941,N_24840);
or UO_2073 (O_2073,N_24988,N_24989);
nor UO_2074 (O_2074,N_24867,N_24765);
nand UO_2075 (O_2075,N_24891,N_24912);
xor UO_2076 (O_2076,N_24824,N_24855);
nor UO_2077 (O_2077,N_24782,N_24786);
or UO_2078 (O_2078,N_24984,N_24928);
or UO_2079 (O_2079,N_24941,N_24950);
nor UO_2080 (O_2080,N_24998,N_24761);
and UO_2081 (O_2081,N_24876,N_24941);
nand UO_2082 (O_2082,N_24968,N_24950);
nor UO_2083 (O_2083,N_24905,N_24805);
or UO_2084 (O_2084,N_24773,N_24843);
nor UO_2085 (O_2085,N_24772,N_24961);
and UO_2086 (O_2086,N_24872,N_24991);
nor UO_2087 (O_2087,N_24895,N_24985);
nor UO_2088 (O_2088,N_24876,N_24777);
and UO_2089 (O_2089,N_24930,N_24945);
or UO_2090 (O_2090,N_24917,N_24966);
xnor UO_2091 (O_2091,N_24763,N_24957);
or UO_2092 (O_2092,N_24965,N_24899);
and UO_2093 (O_2093,N_24750,N_24776);
or UO_2094 (O_2094,N_24999,N_24958);
or UO_2095 (O_2095,N_24771,N_24998);
xnor UO_2096 (O_2096,N_24998,N_24757);
and UO_2097 (O_2097,N_24851,N_24809);
xor UO_2098 (O_2098,N_24767,N_24965);
xor UO_2099 (O_2099,N_24922,N_24804);
or UO_2100 (O_2100,N_24989,N_24934);
and UO_2101 (O_2101,N_24991,N_24784);
and UO_2102 (O_2102,N_24836,N_24822);
xor UO_2103 (O_2103,N_24806,N_24921);
nor UO_2104 (O_2104,N_24987,N_24984);
nand UO_2105 (O_2105,N_24804,N_24921);
nor UO_2106 (O_2106,N_24876,N_24933);
and UO_2107 (O_2107,N_24794,N_24910);
nand UO_2108 (O_2108,N_24916,N_24989);
nor UO_2109 (O_2109,N_24870,N_24781);
xnor UO_2110 (O_2110,N_24862,N_24817);
nor UO_2111 (O_2111,N_24928,N_24969);
nor UO_2112 (O_2112,N_24759,N_24857);
and UO_2113 (O_2113,N_24775,N_24876);
or UO_2114 (O_2114,N_24819,N_24817);
xnor UO_2115 (O_2115,N_24940,N_24752);
and UO_2116 (O_2116,N_24965,N_24856);
or UO_2117 (O_2117,N_24963,N_24883);
xor UO_2118 (O_2118,N_24780,N_24795);
and UO_2119 (O_2119,N_24886,N_24879);
xor UO_2120 (O_2120,N_24932,N_24869);
nor UO_2121 (O_2121,N_24982,N_24840);
nor UO_2122 (O_2122,N_24945,N_24827);
nor UO_2123 (O_2123,N_24890,N_24751);
and UO_2124 (O_2124,N_24837,N_24774);
xnor UO_2125 (O_2125,N_24904,N_24788);
xor UO_2126 (O_2126,N_24766,N_24761);
xnor UO_2127 (O_2127,N_24921,N_24807);
nand UO_2128 (O_2128,N_24776,N_24828);
nor UO_2129 (O_2129,N_24941,N_24852);
nor UO_2130 (O_2130,N_24758,N_24964);
xor UO_2131 (O_2131,N_24983,N_24799);
or UO_2132 (O_2132,N_24827,N_24808);
nor UO_2133 (O_2133,N_24891,N_24903);
or UO_2134 (O_2134,N_24845,N_24876);
nor UO_2135 (O_2135,N_24839,N_24907);
or UO_2136 (O_2136,N_24804,N_24994);
nand UO_2137 (O_2137,N_24991,N_24798);
nand UO_2138 (O_2138,N_24973,N_24809);
and UO_2139 (O_2139,N_24929,N_24822);
and UO_2140 (O_2140,N_24829,N_24927);
and UO_2141 (O_2141,N_24799,N_24831);
nor UO_2142 (O_2142,N_24807,N_24822);
nor UO_2143 (O_2143,N_24793,N_24812);
xor UO_2144 (O_2144,N_24999,N_24838);
xnor UO_2145 (O_2145,N_24926,N_24820);
and UO_2146 (O_2146,N_24972,N_24941);
and UO_2147 (O_2147,N_24822,N_24924);
nand UO_2148 (O_2148,N_24938,N_24825);
or UO_2149 (O_2149,N_24875,N_24946);
nor UO_2150 (O_2150,N_24884,N_24906);
nor UO_2151 (O_2151,N_24829,N_24845);
xnor UO_2152 (O_2152,N_24936,N_24761);
or UO_2153 (O_2153,N_24868,N_24900);
nor UO_2154 (O_2154,N_24904,N_24910);
nand UO_2155 (O_2155,N_24935,N_24890);
and UO_2156 (O_2156,N_24867,N_24942);
or UO_2157 (O_2157,N_24999,N_24961);
xor UO_2158 (O_2158,N_24980,N_24762);
nor UO_2159 (O_2159,N_24904,N_24989);
or UO_2160 (O_2160,N_24904,N_24836);
nand UO_2161 (O_2161,N_24903,N_24907);
and UO_2162 (O_2162,N_24963,N_24918);
or UO_2163 (O_2163,N_24798,N_24908);
xnor UO_2164 (O_2164,N_24762,N_24994);
nor UO_2165 (O_2165,N_24902,N_24913);
nand UO_2166 (O_2166,N_24970,N_24763);
nand UO_2167 (O_2167,N_24820,N_24808);
and UO_2168 (O_2168,N_24780,N_24841);
or UO_2169 (O_2169,N_24811,N_24897);
nor UO_2170 (O_2170,N_24886,N_24865);
nor UO_2171 (O_2171,N_24832,N_24763);
or UO_2172 (O_2172,N_24933,N_24906);
nand UO_2173 (O_2173,N_24754,N_24790);
xnor UO_2174 (O_2174,N_24999,N_24909);
or UO_2175 (O_2175,N_24911,N_24979);
nand UO_2176 (O_2176,N_24870,N_24812);
and UO_2177 (O_2177,N_24891,N_24937);
nand UO_2178 (O_2178,N_24878,N_24870);
nor UO_2179 (O_2179,N_24881,N_24835);
nor UO_2180 (O_2180,N_24867,N_24814);
or UO_2181 (O_2181,N_24885,N_24924);
nand UO_2182 (O_2182,N_24852,N_24894);
xor UO_2183 (O_2183,N_24896,N_24904);
nand UO_2184 (O_2184,N_24903,N_24834);
nand UO_2185 (O_2185,N_24783,N_24904);
and UO_2186 (O_2186,N_24960,N_24862);
xor UO_2187 (O_2187,N_24796,N_24889);
xor UO_2188 (O_2188,N_24881,N_24980);
nor UO_2189 (O_2189,N_24843,N_24870);
or UO_2190 (O_2190,N_24928,N_24773);
xnor UO_2191 (O_2191,N_24868,N_24771);
xor UO_2192 (O_2192,N_24868,N_24979);
xor UO_2193 (O_2193,N_24775,N_24973);
nor UO_2194 (O_2194,N_24915,N_24761);
xnor UO_2195 (O_2195,N_24948,N_24853);
or UO_2196 (O_2196,N_24957,N_24821);
nand UO_2197 (O_2197,N_24877,N_24810);
or UO_2198 (O_2198,N_24817,N_24927);
nor UO_2199 (O_2199,N_24939,N_24761);
nor UO_2200 (O_2200,N_24807,N_24779);
xnor UO_2201 (O_2201,N_24974,N_24968);
or UO_2202 (O_2202,N_24849,N_24889);
nand UO_2203 (O_2203,N_24761,N_24753);
and UO_2204 (O_2204,N_24949,N_24889);
nand UO_2205 (O_2205,N_24791,N_24940);
and UO_2206 (O_2206,N_24827,N_24817);
xor UO_2207 (O_2207,N_24818,N_24845);
or UO_2208 (O_2208,N_24925,N_24898);
nand UO_2209 (O_2209,N_24879,N_24889);
or UO_2210 (O_2210,N_24772,N_24833);
xor UO_2211 (O_2211,N_24953,N_24998);
xor UO_2212 (O_2212,N_24765,N_24892);
xor UO_2213 (O_2213,N_24971,N_24953);
nor UO_2214 (O_2214,N_24976,N_24999);
or UO_2215 (O_2215,N_24996,N_24755);
and UO_2216 (O_2216,N_24997,N_24836);
or UO_2217 (O_2217,N_24876,N_24944);
nor UO_2218 (O_2218,N_24767,N_24780);
or UO_2219 (O_2219,N_24891,N_24968);
nor UO_2220 (O_2220,N_24788,N_24785);
and UO_2221 (O_2221,N_24987,N_24842);
or UO_2222 (O_2222,N_24957,N_24844);
or UO_2223 (O_2223,N_24898,N_24923);
and UO_2224 (O_2224,N_24860,N_24842);
and UO_2225 (O_2225,N_24995,N_24767);
or UO_2226 (O_2226,N_24783,N_24788);
nor UO_2227 (O_2227,N_24751,N_24985);
nor UO_2228 (O_2228,N_24892,N_24798);
or UO_2229 (O_2229,N_24802,N_24946);
xor UO_2230 (O_2230,N_24920,N_24780);
and UO_2231 (O_2231,N_24895,N_24831);
xor UO_2232 (O_2232,N_24774,N_24802);
or UO_2233 (O_2233,N_24953,N_24814);
nor UO_2234 (O_2234,N_24800,N_24837);
xor UO_2235 (O_2235,N_24788,N_24767);
xnor UO_2236 (O_2236,N_24906,N_24794);
nor UO_2237 (O_2237,N_24895,N_24838);
nand UO_2238 (O_2238,N_24977,N_24890);
or UO_2239 (O_2239,N_24991,N_24844);
or UO_2240 (O_2240,N_24785,N_24985);
nor UO_2241 (O_2241,N_24844,N_24762);
or UO_2242 (O_2242,N_24868,N_24936);
and UO_2243 (O_2243,N_24871,N_24992);
nor UO_2244 (O_2244,N_24958,N_24789);
and UO_2245 (O_2245,N_24893,N_24892);
and UO_2246 (O_2246,N_24841,N_24794);
xnor UO_2247 (O_2247,N_24820,N_24793);
xor UO_2248 (O_2248,N_24854,N_24976);
xnor UO_2249 (O_2249,N_24918,N_24962);
nor UO_2250 (O_2250,N_24752,N_24962);
or UO_2251 (O_2251,N_24922,N_24890);
or UO_2252 (O_2252,N_24912,N_24974);
or UO_2253 (O_2253,N_24998,N_24930);
or UO_2254 (O_2254,N_24849,N_24815);
or UO_2255 (O_2255,N_24817,N_24938);
xnor UO_2256 (O_2256,N_24861,N_24941);
nand UO_2257 (O_2257,N_24914,N_24898);
nand UO_2258 (O_2258,N_24899,N_24872);
nor UO_2259 (O_2259,N_24861,N_24924);
and UO_2260 (O_2260,N_24979,N_24790);
nand UO_2261 (O_2261,N_24936,N_24778);
or UO_2262 (O_2262,N_24925,N_24955);
and UO_2263 (O_2263,N_24778,N_24896);
and UO_2264 (O_2264,N_24947,N_24795);
nor UO_2265 (O_2265,N_24969,N_24771);
nand UO_2266 (O_2266,N_24888,N_24781);
or UO_2267 (O_2267,N_24933,N_24926);
nor UO_2268 (O_2268,N_24756,N_24849);
nor UO_2269 (O_2269,N_24951,N_24785);
nor UO_2270 (O_2270,N_24806,N_24926);
nor UO_2271 (O_2271,N_24815,N_24837);
or UO_2272 (O_2272,N_24999,N_24903);
and UO_2273 (O_2273,N_24958,N_24974);
nor UO_2274 (O_2274,N_24784,N_24840);
or UO_2275 (O_2275,N_24776,N_24848);
nand UO_2276 (O_2276,N_24901,N_24776);
nor UO_2277 (O_2277,N_24916,N_24941);
nand UO_2278 (O_2278,N_24978,N_24885);
nor UO_2279 (O_2279,N_24968,N_24883);
or UO_2280 (O_2280,N_24963,N_24945);
nand UO_2281 (O_2281,N_24959,N_24987);
or UO_2282 (O_2282,N_24956,N_24781);
nand UO_2283 (O_2283,N_24876,N_24803);
xnor UO_2284 (O_2284,N_24968,N_24767);
nor UO_2285 (O_2285,N_24783,N_24770);
nor UO_2286 (O_2286,N_24807,N_24791);
nor UO_2287 (O_2287,N_24789,N_24753);
xor UO_2288 (O_2288,N_24977,N_24750);
nor UO_2289 (O_2289,N_24898,N_24798);
or UO_2290 (O_2290,N_24878,N_24902);
nand UO_2291 (O_2291,N_24948,N_24819);
or UO_2292 (O_2292,N_24943,N_24756);
or UO_2293 (O_2293,N_24851,N_24986);
nor UO_2294 (O_2294,N_24871,N_24916);
and UO_2295 (O_2295,N_24926,N_24937);
nand UO_2296 (O_2296,N_24794,N_24844);
and UO_2297 (O_2297,N_24875,N_24936);
and UO_2298 (O_2298,N_24787,N_24855);
nand UO_2299 (O_2299,N_24867,N_24776);
nor UO_2300 (O_2300,N_24819,N_24935);
nor UO_2301 (O_2301,N_24800,N_24775);
or UO_2302 (O_2302,N_24904,N_24909);
nand UO_2303 (O_2303,N_24791,N_24986);
nor UO_2304 (O_2304,N_24871,N_24954);
nand UO_2305 (O_2305,N_24847,N_24995);
nor UO_2306 (O_2306,N_24864,N_24820);
xor UO_2307 (O_2307,N_24961,N_24922);
nand UO_2308 (O_2308,N_24990,N_24924);
nand UO_2309 (O_2309,N_24852,N_24794);
or UO_2310 (O_2310,N_24782,N_24806);
nor UO_2311 (O_2311,N_24986,N_24902);
and UO_2312 (O_2312,N_24794,N_24808);
nand UO_2313 (O_2313,N_24943,N_24865);
or UO_2314 (O_2314,N_24820,N_24851);
xor UO_2315 (O_2315,N_24974,N_24987);
nand UO_2316 (O_2316,N_24889,N_24787);
xor UO_2317 (O_2317,N_24806,N_24789);
and UO_2318 (O_2318,N_24877,N_24866);
nand UO_2319 (O_2319,N_24823,N_24771);
xnor UO_2320 (O_2320,N_24828,N_24861);
or UO_2321 (O_2321,N_24955,N_24754);
and UO_2322 (O_2322,N_24948,N_24909);
xor UO_2323 (O_2323,N_24810,N_24781);
and UO_2324 (O_2324,N_24769,N_24898);
nand UO_2325 (O_2325,N_24879,N_24775);
or UO_2326 (O_2326,N_24866,N_24937);
xnor UO_2327 (O_2327,N_24959,N_24822);
and UO_2328 (O_2328,N_24843,N_24933);
nand UO_2329 (O_2329,N_24949,N_24956);
or UO_2330 (O_2330,N_24859,N_24766);
or UO_2331 (O_2331,N_24972,N_24914);
or UO_2332 (O_2332,N_24930,N_24754);
nand UO_2333 (O_2333,N_24772,N_24956);
xor UO_2334 (O_2334,N_24870,N_24960);
or UO_2335 (O_2335,N_24803,N_24880);
and UO_2336 (O_2336,N_24991,N_24763);
nor UO_2337 (O_2337,N_24887,N_24928);
xnor UO_2338 (O_2338,N_24901,N_24879);
and UO_2339 (O_2339,N_24934,N_24783);
nor UO_2340 (O_2340,N_24888,N_24933);
nand UO_2341 (O_2341,N_24909,N_24836);
and UO_2342 (O_2342,N_24788,N_24862);
and UO_2343 (O_2343,N_24830,N_24874);
or UO_2344 (O_2344,N_24804,N_24945);
nand UO_2345 (O_2345,N_24930,N_24910);
and UO_2346 (O_2346,N_24772,N_24925);
nor UO_2347 (O_2347,N_24989,N_24778);
nor UO_2348 (O_2348,N_24810,N_24899);
and UO_2349 (O_2349,N_24814,N_24904);
or UO_2350 (O_2350,N_24827,N_24865);
and UO_2351 (O_2351,N_24996,N_24826);
or UO_2352 (O_2352,N_24792,N_24770);
and UO_2353 (O_2353,N_24826,N_24924);
nor UO_2354 (O_2354,N_24862,N_24995);
or UO_2355 (O_2355,N_24759,N_24852);
xnor UO_2356 (O_2356,N_24763,N_24945);
and UO_2357 (O_2357,N_24780,N_24938);
nand UO_2358 (O_2358,N_24791,N_24770);
nand UO_2359 (O_2359,N_24930,N_24823);
and UO_2360 (O_2360,N_24938,N_24964);
nor UO_2361 (O_2361,N_24912,N_24786);
and UO_2362 (O_2362,N_24816,N_24891);
nor UO_2363 (O_2363,N_24806,N_24805);
xor UO_2364 (O_2364,N_24972,N_24804);
and UO_2365 (O_2365,N_24875,N_24755);
and UO_2366 (O_2366,N_24838,N_24903);
xnor UO_2367 (O_2367,N_24943,N_24993);
xor UO_2368 (O_2368,N_24777,N_24952);
or UO_2369 (O_2369,N_24964,N_24798);
or UO_2370 (O_2370,N_24979,N_24802);
and UO_2371 (O_2371,N_24875,N_24797);
nand UO_2372 (O_2372,N_24873,N_24979);
or UO_2373 (O_2373,N_24886,N_24859);
xnor UO_2374 (O_2374,N_24792,N_24956);
or UO_2375 (O_2375,N_24946,N_24892);
or UO_2376 (O_2376,N_24957,N_24927);
and UO_2377 (O_2377,N_24933,N_24992);
xor UO_2378 (O_2378,N_24782,N_24978);
or UO_2379 (O_2379,N_24971,N_24999);
or UO_2380 (O_2380,N_24834,N_24768);
and UO_2381 (O_2381,N_24959,N_24985);
nand UO_2382 (O_2382,N_24855,N_24767);
nand UO_2383 (O_2383,N_24884,N_24753);
or UO_2384 (O_2384,N_24846,N_24933);
xnor UO_2385 (O_2385,N_24848,N_24773);
nor UO_2386 (O_2386,N_24937,N_24872);
nand UO_2387 (O_2387,N_24895,N_24919);
nand UO_2388 (O_2388,N_24949,N_24876);
xor UO_2389 (O_2389,N_24962,N_24772);
and UO_2390 (O_2390,N_24979,N_24860);
xor UO_2391 (O_2391,N_24872,N_24973);
or UO_2392 (O_2392,N_24845,N_24848);
nand UO_2393 (O_2393,N_24828,N_24878);
or UO_2394 (O_2394,N_24956,N_24996);
nor UO_2395 (O_2395,N_24910,N_24938);
nand UO_2396 (O_2396,N_24911,N_24910);
nand UO_2397 (O_2397,N_24755,N_24912);
or UO_2398 (O_2398,N_24764,N_24820);
or UO_2399 (O_2399,N_24925,N_24806);
xnor UO_2400 (O_2400,N_24815,N_24909);
or UO_2401 (O_2401,N_24947,N_24833);
xnor UO_2402 (O_2402,N_24955,N_24979);
nand UO_2403 (O_2403,N_24967,N_24882);
and UO_2404 (O_2404,N_24932,N_24783);
nand UO_2405 (O_2405,N_24849,N_24823);
or UO_2406 (O_2406,N_24920,N_24969);
and UO_2407 (O_2407,N_24800,N_24918);
nor UO_2408 (O_2408,N_24879,N_24806);
and UO_2409 (O_2409,N_24998,N_24984);
xor UO_2410 (O_2410,N_24774,N_24993);
or UO_2411 (O_2411,N_24872,N_24981);
nor UO_2412 (O_2412,N_24866,N_24932);
xor UO_2413 (O_2413,N_24963,N_24863);
nor UO_2414 (O_2414,N_24931,N_24793);
nand UO_2415 (O_2415,N_24866,N_24973);
nor UO_2416 (O_2416,N_24933,N_24912);
and UO_2417 (O_2417,N_24800,N_24783);
nand UO_2418 (O_2418,N_24786,N_24953);
or UO_2419 (O_2419,N_24982,N_24850);
or UO_2420 (O_2420,N_24951,N_24986);
and UO_2421 (O_2421,N_24831,N_24994);
nand UO_2422 (O_2422,N_24895,N_24754);
and UO_2423 (O_2423,N_24805,N_24945);
xor UO_2424 (O_2424,N_24987,N_24997);
nand UO_2425 (O_2425,N_24912,N_24994);
or UO_2426 (O_2426,N_24917,N_24985);
or UO_2427 (O_2427,N_24897,N_24905);
xor UO_2428 (O_2428,N_24813,N_24898);
xor UO_2429 (O_2429,N_24847,N_24759);
or UO_2430 (O_2430,N_24817,N_24987);
or UO_2431 (O_2431,N_24833,N_24808);
nor UO_2432 (O_2432,N_24816,N_24836);
nor UO_2433 (O_2433,N_24964,N_24864);
or UO_2434 (O_2434,N_24856,N_24873);
nor UO_2435 (O_2435,N_24872,N_24846);
or UO_2436 (O_2436,N_24904,N_24786);
or UO_2437 (O_2437,N_24847,N_24974);
or UO_2438 (O_2438,N_24825,N_24991);
xnor UO_2439 (O_2439,N_24755,N_24881);
or UO_2440 (O_2440,N_24938,N_24921);
and UO_2441 (O_2441,N_24792,N_24951);
and UO_2442 (O_2442,N_24998,N_24784);
nand UO_2443 (O_2443,N_24999,N_24878);
nand UO_2444 (O_2444,N_24923,N_24870);
or UO_2445 (O_2445,N_24882,N_24785);
nand UO_2446 (O_2446,N_24955,N_24844);
xor UO_2447 (O_2447,N_24843,N_24975);
and UO_2448 (O_2448,N_24975,N_24856);
or UO_2449 (O_2449,N_24880,N_24931);
or UO_2450 (O_2450,N_24801,N_24785);
xnor UO_2451 (O_2451,N_24863,N_24876);
and UO_2452 (O_2452,N_24892,N_24929);
nor UO_2453 (O_2453,N_24945,N_24980);
and UO_2454 (O_2454,N_24940,N_24768);
and UO_2455 (O_2455,N_24875,N_24811);
nor UO_2456 (O_2456,N_24751,N_24825);
and UO_2457 (O_2457,N_24919,N_24750);
nand UO_2458 (O_2458,N_24774,N_24926);
xnor UO_2459 (O_2459,N_24856,N_24794);
or UO_2460 (O_2460,N_24923,N_24761);
nor UO_2461 (O_2461,N_24997,N_24978);
nand UO_2462 (O_2462,N_24960,N_24966);
and UO_2463 (O_2463,N_24903,N_24806);
and UO_2464 (O_2464,N_24788,N_24929);
nand UO_2465 (O_2465,N_24961,N_24920);
or UO_2466 (O_2466,N_24762,N_24949);
and UO_2467 (O_2467,N_24977,N_24840);
or UO_2468 (O_2468,N_24826,N_24775);
and UO_2469 (O_2469,N_24989,N_24834);
or UO_2470 (O_2470,N_24799,N_24847);
or UO_2471 (O_2471,N_24880,N_24797);
xnor UO_2472 (O_2472,N_24947,N_24794);
xor UO_2473 (O_2473,N_24770,N_24836);
nand UO_2474 (O_2474,N_24781,N_24750);
nor UO_2475 (O_2475,N_24853,N_24892);
nor UO_2476 (O_2476,N_24964,N_24892);
nor UO_2477 (O_2477,N_24987,N_24963);
xnor UO_2478 (O_2478,N_24934,N_24983);
nor UO_2479 (O_2479,N_24784,N_24832);
nand UO_2480 (O_2480,N_24812,N_24895);
and UO_2481 (O_2481,N_24797,N_24963);
and UO_2482 (O_2482,N_24797,N_24781);
xnor UO_2483 (O_2483,N_24923,N_24860);
and UO_2484 (O_2484,N_24888,N_24899);
and UO_2485 (O_2485,N_24928,N_24906);
nand UO_2486 (O_2486,N_24813,N_24896);
and UO_2487 (O_2487,N_24755,N_24798);
nand UO_2488 (O_2488,N_24842,N_24959);
nor UO_2489 (O_2489,N_24836,N_24755);
nand UO_2490 (O_2490,N_24992,N_24962);
xnor UO_2491 (O_2491,N_24789,N_24868);
or UO_2492 (O_2492,N_24786,N_24855);
xor UO_2493 (O_2493,N_24897,N_24827);
and UO_2494 (O_2494,N_24955,N_24890);
and UO_2495 (O_2495,N_24773,N_24942);
or UO_2496 (O_2496,N_24898,N_24808);
or UO_2497 (O_2497,N_24979,N_24948);
or UO_2498 (O_2498,N_24930,N_24961);
and UO_2499 (O_2499,N_24852,N_24943);
nor UO_2500 (O_2500,N_24847,N_24827);
or UO_2501 (O_2501,N_24775,N_24959);
nor UO_2502 (O_2502,N_24950,N_24983);
nor UO_2503 (O_2503,N_24986,N_24960);
and UO_2504 (O_2504,N_24840,N_24916);
nand UO_2505 (O_2505,N_24897,N_24838);
or UO_2506 (O_2506,N_24959,N_24836);
nor UO_2507 (O_2507,N_24912,N_24882);
or UO_2508 (O_2508,N_24798,N_24931);
or UO_2509 (O_2509,N_24866,N_24957);
nand UO_2510 (O_2510,N_24887,N_24849);
nor UO_2511 (O_2511,N_24915,N_24783);
nand UO_2512 (O_2512,N_24963,N_24873);
xor UO_2513 (O_2513,N_24969,N_24913);
nor UO_2514 (O_2514,N_24814,N_24993);
or UO_2515 (O_2515,N_24849,N_24913);
or UO_2516 (O_2516,N_24887,N_24793);
nand UO_2517 (O_2517,N_24830,N_24850);
and UO_2518 (O_2518,N_24861,N_24810);
nor UO_2519 (O_2519,N_24875,N_24787);
or UO_2520 (O_2520,N_24863,N_24798);
nand UO_2521 (O_2521,N_24927,N_24834);
or UO_2522 (O_2522,N_24790,N_24797);
nand UO_2523 (O_2523,N_24862,N_24807);
xor UO_2524 (O_2524,N_24917,N_24826);
nor UO_2525 (O_2525,N_24993,N_24877);
or UO_2526 (O_2526,N_24771,N_24904);
xnor UO_2527 (O_2527,N_24920,N_24993);
or UO_2528 (O_2528,N_24965,N_24931);
xor UO_2529 (O_2529,N_24752,N_24760);
nor UO_2530 (O_2530,N_24953,N_24930);
and UO_2531 (O_2531,N_24993,N_24875);
or UO_2532 (O_2532,N_24959,N_24814);
nand UO_2533 (O_2533,N_24881,N_24969);
and UO_2534 (O_2534,N_24755,N_24828);
or UO_2535 (O_2535,N_24834,N_24987);
or UO_2536 (O_2536,N_24799,N_24909);
or UO_2537 (O_2537,N_24946,N_24931);
nor UO_2538 (O_2538,N_24825,N_24939);
nand UO_2539 (O_2539,N_24955,N_24946);
nand UO_2540 (O_2540,N_24869,N_24855);
or UO_2541 (O_2541,N_24939,N_24809);
or UO_2542 (O_2542,N_24902,N_24818);
nor UO_2543 (O_2543,N_24794,N_24934);
or UO_2544 (O_2544,N_24983,N_24955);
and UO_2545 (O_2545,N_24818,N_24827);
xor UO_2546 (O_2546,N_24894,N_24844);
and UO_2547 (O_2547,N_24992,N_24791);
and UO_2548 (O_2548,N_24858,N_24902);
or UO_2549 (O_2549,N_24755,N_24753);
xnor UO_2550 (O_2550,N_24809,N_24835);
and UO_2551 (O_2551,N_24857,N_24833);
or UO_2552 (O_2552,N_24871,N_24760);
nand UO_2553 (O_2553,N_24849,N_24810);
nand UO_2554 (O_2554,N_24915,N_24890);
nand UO_2555 (O_2555,N_24866,N_24936);
xnor UO_2556 (O_2556,N_24753,N_24932);
nand UO_2557 (O_2557,N_24950,N_24957);
or UO_2558 (O_2558,N_24953,N_24802);
or UO_2559 (O_2559,N_24790,N_24808);
nand UO_2560 (O_2560,N_24855,N_24867);
and UO_2561 (O_2561,N_24802,N_24784);
nor UO_2562 (O_2562,N_24848,N_24856);
or UO_2563 (O_2563,N_24983,N_24785);
nor UO_2564 (O_2564,N_24928,N_24874);
and UO_2565 (O_2565,N_24799,N_24775);
and UO_2566 (O_2566,N_24839,N_24770);
and UO_2567 (O_2567,N_24874,N_24963);
and UO_2568 (O_2568,N_24994,N_24854);
and UO_2569 (O_2569,N_24928,N_24790);
or UO_2570 (O_2570,N_24841,N_24816);
xor UO_2571 (O_2571,N_24853,N_24883);
and UO_2572 (O_2572,N_24896,N_24792);
or UO_2573 (O_2573,N_24870,N_24941);
or UO_2574 (O_2574,N_24841,N_24891);
and UO_2575 (O_2575,N_24938,N_24803);
or UO_2576 (O_2576,N_24767,N_24865);
or UO_2577 (O_2577,N_24895,N_24958);
xor UO_2578 (O_2578,N_24920,N_24948);
nor UO_2579 (O_2579,N_24798,N_24922);
nand UO_2580 (O_2580,N_24855,N_24863);
nor UO_2581 (O_2581,N_24766,N_24805);
xnor UO_2582 (O_2582,N_24862,N_24764);
xor UO_2583 (O_2583,N_24809,N_24849);
nand UO_2584 (O_2584,N_24945,N_24795);
nor UO_2585 (O_2585,N_24918,N_24866);
nand UO_2586 (O_2586,N_24845,N_24947);
nor UO_2587 (O_2587,N_24810,N_24759);
xnor UO_2588 (O_2588,N_24764,N_24895);
or UO_2589 (O_2589,N_24861,N_24836);
xor UO_2590 (O_2590,N_24945,N_24880);
xnor UO_2591 (O_2591,N_24915,N_24891);
or UO_2592 (O_2592,N_24979,N_24791);
nor UO_2593 (O_2593,N_24756,N_24751);
or UO_2594 (O_2594,N_24847,N_24926);
or UO_2595 (O_2595,N_24869,N_24814);
xnor UO_2596 (O_2596,N_24838,N_24786);
xnor UO_2597 (O_2597,N_24886,N_24934);
nor UO_2598 (O_2598,N_24926,N_24848);
nand UO_2599 (O_2599,N_24872,N_24881);
or UO_2600 (O_2600,N_24757,N_24978);
or UO_2601 (O_2601,N_24966,N_24841);
xnor UO_2602 (O_2602,N_24803,N_24928);
nand UO_2603 (O_2603,N_24915,N_24992);
nor UO_2604 (O_2604,N_24894,N_24997);
nand UO_2605 (O_2605,N_24870,N_24902);
or UO_2606 (O_2606,N_24826,N_24816);
xor UO_2607 (O_2607,N_24979,N_24852);
nor UO_2608 (O_2608,N_24894,N_24953);
xnor UO_2609 (O_2609,N_24975,N_24842);
and UO_2610 (O_2610,N_24917,N_24983);
or UO_2611 (O_2611,N_24889,N_24965);
nand UO_2612 (O_2612,N_24891,N_24924);
nand UO_2613 (O_2613,N_24953,N_24886);
or UO_2614 (O_2614,N_24771,N_24872);
and UO_2615 (O_2615,N_24773,N_24949);
nor UO_2616 (O_2616,N_24870,N_24802);
and UO_2617 (O_2617,N_24830,N_24969);
and UO_2618 (O_2618,N_24771,N_24910);
and UO_2619 (O_2619,N_24839,N_24838);
nor UO_2620 (O_2620,N_24756,N_24955);
or UO_2621 (O_2621,N_24970,N_24941);
nor UO_2622 (O_2622,N_24759,N_24849);
nand UO_2623 (O_2623,N_24943,N_24835);
and UO_2624 (O_2624,N_24862,N_24767);
or UO_2625 (O_2625,N_24974,N_24792);
nor UO_2626 (O_2626,N_24894,N_24990);
or UO_2627 (O_2627,N_24857,N_24856);
nor UO_2628 (O_2628,N_24840,N_24949);
xor UO_2629 (O_2629,N_24787,N_24944);
nand UO_2630 (O_2630,N_24945,N_24973);
xnor UO_2631 (O_2631,N_24948,N_24805);
or UO_2632 (O_2632,N_24877,N_24915);
xor UO_2633 (O_2633,N_24852,N_24884);
xnor UO_2634 (O_2634,N_24795,N_24901);
nor UO_2635 (O_2635,N_24989,N_24795);
nand UO_2636 (O_2636,N_24775,N_24938);
nand UO_2637 (O_2637,N_24774,N_24996);
nand UO_2638 (O_2638,N_24927,N_24994);
and UO_2639 (O_2639,N_24867,N_24966);
xor UO_2640 (O_2640,N_24958,N_24899);
and UO_2641 (O_2641,N_24797,N_24982);
nor UO_2642 (O_2642,N_24752,N_24775);
nor UO_2643 (O_2643,N_24870,N_24891);
nand UO_2644 (O_2644,N_24898,N_24825);
nand UO_2645 (O_2645,N_24982,N_24784);
nor UO_2646 (O_2646,N_24826,N_24990);
xor UO_2647 (O_2647,N_24878,N_24806);
nand UO_2648 (O_2648,N_24755,N_24792);
xnor UO_2649 (O_2649,N_24810,N_24856);
nor UO_2650 (O_2650,N_24796,N_24930);
xor UO_2651 (O_2651,N_24816,N_24906);
or UO_2652 (O_2652,N_24869,N_24965);
xor UO_2653 (O_2653,N_24798,N_24801);
nand UO_2654 (O_2654,N_24984,N_24976);
xor UO_2655 (O_2655,N_24780,N_24873);
nor UO_2656 (O_2656,N_24946,N_24986);
xnor UO_2657 (O_2657,N_24760,N_24968);
or UO_2658 (O_2658,N_24868,N_24970);
nor UO_2659 (O_2659,N_24871,N_24889);
and UO_2660 (O_2660,N_24971,N_24837);
xnor UO_2661 (O_2661,N_24925,N_24770);
nor UO_2662 (O_2662,N_24877,N_24805);
or UO_2663 (O_2663,N_24863,N_24750);
xor UO_2664 (O_2664,N_24852,N_24917);
nand UO_2665 (O_2665,N_24906,N_24927);
nor UO_2666 (O_2666,N_24784,N_24808);
xor UO_2667 (O_2667,N_24847,N_24836);
xor UO_2668 (O_2668,N_24906,N_24817);
xnor UO_2669 (O_2669,N_24868,N_24842);
nand UO_2670 (O_2670,N_24785,N_24894);
xor UO_2671 (O_2671,N_24795,N_24997);
nand UO_2672 (O_2672,N_24867,N_24841);
nand UO_2673 (O_2673,N_24973,N_24887);
nand UO_2674 (O_2674,N_24998,N_24851);
or UO_2675 (O_2675,N_24910,N_24767);
or UO_2676 (O_2676,N_24890,N_24931);
and UO_2677 (O_2677,N_24979,N_24969);
nand UO_2678 (O_2678,N_24838,N_24790);
nor UO_2679 (O_2679,N_24925,N_24777);
nor UO_2680 (O_2680,N_24808,N_24875);
nor UO_2681 (O_2681,N_24856,N_24813);
nor UO_2682 (O_2682,N_24805,N_24904);
nand UO_2683 (O_2683,N_24821,N_24935);
and UO_2684 (O_2684,N_24983,N_24889);
xor UO_2685 (O_2685,N_24898,N_24868);
and UO_2686 (O_2686,N_24891,N_24916);
xnor UO_2687 (O_2687,N_24992,N_24949);
nor UO_2688 (O_2688,N_24886,N_24804);
nand UO_2689 (O_2689,N_24991,N_24824);
nand UO_2690 (O_2690,N_24959,N_24967);
nor UO_2691 (O_2691,N_24887,N_24984);
and UO_2692 (O_2692,N_24908,N_24772);
nor UO_2693 (O_2693,N_24868,N_24822);
or UO_2694 (O_2694,N_24837,N_24903);
and UO_2695 (O_2695,N_24781,N_24877);
xnor UO_2696 (O_2696,N_24929,N_24960);
nand UO_2697 (O_2697,N_24970,N_24875);
nand UO_2698 (O_2698,N_24928,N_24987);
nand UO_2699 (O_2699,N_24806,N_24922);
nor UO_2700 (O_2700,N_24808,N_24814);
or UO_2701 (O_2701,N_24803,N_24757);
or UO_2702 (O_2702,N_24970,N_24839);
and UO_2703 (O_2703,N_24945,N_24915);
nand UO_2704 (O_2704,N_24836,N_24832);
nand UO_2705 (O_2705,N_24975,N_24942);
nor UO_2706 (O_2706,N_24765,N_24941);
xnor UO_2707 (O_2707,N_24999,N_24786);
and UO_2708 (O_2708,N_24821,N_24802);
nor UO_2709 (O_2709,N_24885,N_24814);
nand UO_2710 (O_2710,N_24801,N_24839);
xor UO_2711 (O_2711,N_24850,N_24764);
or UO_2712 (O_2712,N_24841,N_24962);
nor UO_2713 (O_2713,N_24858,N_24922);
nor UO_2714 (O_2714,N_24800,N_24881);
or UO_2715 (O_2715,N_24840,N_24907);
nand UO_2716 (O_2716,N_24799,N_24769);
and UO_2717 (O_2717,N_24989,N_24957);
nor UO_2718 (O_2718,N_24964,N_24886);
nor UO_2719 (O_2719,N_24909,N_24970);
nor UO_2720 (O_2720,N_24848,N_24844);
xor UO_2721 (O_2721,N_24828,N_24812);
and UO_2722 (O_2722,N_24837,N_24953);
nor UO_2723 (O_2723,N_24872,N_24904);
and UO_2724 (O_2724,N_24934,N_24876);
nor UO_2725 (O_2725,N_24772,N_24970);
and UO_2726 (O_2726,N_24785,N_24775);
nor UO_2727 (O_2727,N_24861,N_24782);
or UO_2728 (O_2728,N_24854,N_24888);
nand UO_2729 (O_2729,N_24921,N_24776);
and UO_2730 (O_2730,N_24803,N_24939);
xnor UO_2731 (O_2731,N_24812,N_24970);
or UO_2732 (O_2732,N_24751,N_24768);
and UO_2733 (O_2733,N_24969,N_24900);
and UO_2734 (O_2734,N_24965,N_24766);
and UO_2735 (O_2735,N_24928,N_24798);
nand UO_2736 (O_2736,N_24997,N_24860);
nor UO_2737 (O_2737,N_24934,N_24907);
and UO_2738 (O_2738,N_24888,N_24756);
nor UO_2739 (O_2739,N_24773,N_24936);
nor UO_2740 (O_2740,N_24900,N_24838);
nand UO_2741 (O_2741,N_24879,N_24793);
xnor UO_2742 (O_2742,N_24800,N_24968);
or UO_2743 (O_2743,N_24836,N_24787);
nor UO_2744 (O_2744,N_24940,N_24817);
nor UO_2745 (O_2745,N_24997,N_24951);
nor UO_2746 (O_2746,N_24845,N_24984);
xor UO_2747 (O_2747,N_24875,N_24776);
nand UO_2748 (O_2748,N_24970,N_24782);
nor UO_2749 (O_2749,N_24875,N_24894);
nand UO_2750 (O_2750,N_24952,N_24786);
nand UO_2751 (O_2751,N_24879,N_24861);
xnor UO_2752 (O_2752,N_24927,N_24857);
xnor UO_2753 (O_2753,N_24792,N_24933);
nor UO_2754 (O_2754,N_24758,N_24881);
and UO_2755 (O_2755,N_24892,N_24895);
or UO_2756 (O_2756,N_24895,N_24877);
nor UO_2757 (O_2757,N_24930,N_24992);
nor UO_2758 (O_2758,N_24842,N_24851);
nor UO_2759 (O_2759,N_24955,N_24785);
or UO_2760 (O_2760,N_24769,N_24768);
nand UO_2761 (O_2761,N_24762,N_24869);
xor UO_2762 (O_2762,N_24843,N_24956);
nor UO_2763 (O_2763,N_24931,N_24768);
and UO_2764 (O_2764,N_24778,N_24865);
or UO_2765 (O_2765,N_24945,N_24787);
xor UO_2766 (O_2766,N_24882,N_24961);
xor UO_2767 (O_2767,N_24899,N_24929);
or UO_2768 (O_2768,N_24917,N_24944);
nor UO_2769 (O_2769,N_24850,N_24986);
xnor UO_2770 (O_2770,N_24967,N_24998);
nand UO_2771 (O_2771,N_24889,N_24979);
nand UO_2772 (O_2772,N_24923,N_24755);
nor UO_2773 (O_2773,N_24848,N_24989);
xor UO_2774 (O_2774,N_24911,N_24804);
and UO_2775 (O_2775,N_24949,N_24819);
or UO_2776 (O_2776,N_24794,N_24873);
and UO_2777 (O_2777,N_24899,N_24993);
and UO_2778 (O_2778,N_24967,N_24815);
or UO_2779 (O_2779,N_24940,N_24971);
nor UO_2780 (O_2780,N_24952,N_24792);
nand UO_2781 (O_2781,N_24923,N_24900);
xor UO_2782 (O_2782,N_24775,N_24883);
xor UO_2783 (O_2783,N_24759,N_24949);
and UO_2784 (O_2784,N_24998,N_24906);
or UO_2785 (O_2785,N_24948,N_24866);
nor UO_2786 (O_2786,N_24827,N_24781);
nor UO_2787 (O_2787,N_24896,N_24857);
and UO_2788 (O_2788,N_24968,N_24822);
xor UO_2789 (O_2789,N_24849,N_24767);
nand UO_2790 (O_2790,N_24865,N_24756);
and UO_2791 (O_2791,N_24811,N_24794);
or UO_2792 (O_2792,N_24768,N_24763);
xnor UO_2793 (O_2793,N_24973,N_24822);
xnor UO_2794 (O_2794,N_24806,N_24857);
nand UO_2795 (O_2795,N_24776,N_24861);
nand UO_2796 (O_2796,N_24995,N_24921);
nand UO_2797 (O_2797,N_24887,N_24814);
or UO_2798 (O_2798,N_24858,N_24831);
nor UO_2799 (O_2799,N_24981,N_24756);
and UO_2800 (O_2800,N_24792,N_24811);
nor UO_2801 (O_2801,N_24885,N_24895);
nor UO_2802 (O_2802,N_24815,N_24960);
nor UO_2803 (O_2803,N_24939,N_24991);
nor UO_2804 (O_2804,N_24811,N_24824);
or UO_2805 (O_2805,N_24774,N_24790);
and UO_2806 (O_2806,N_24977,N_24979);
and UO_2807 (O_2807,N_24785,N_24935);
xor UO_2808 (O_2808,N_24762,N_24867);
xnor UO_2809 (O_2809,N_24921,N_24980);
or UO_2810 (O_2810,N_24950,N_24792);
nor UO_2811 (O_2811,N_24824,N_24887);
nor UO_2812 (O_2812,N_24944,N_24867);
or UO_2813 (O_2813,N_24887,N_24898);
nand UO_2814 (O_2814,N_24778,N_24967);
nor UO_2815 (O_2815,N_24948,N_24932);
and UO_2816 (O_2816,N_24788,N_24811);
or UO_2817 (O_2817,N_24901,N_24971);
nor UO_2818 (O_2818,N_24942,N_24876);
nand UO_2819 (O_2819,N_24855,N_24813);
nor UO_2820 (O_2820,N_24855,N_24956);
or UO_2821 (O_2821,N_24809,N_24826);
and UO_2822 (O_2822,N_24947,N_24803);
or UO_2823 (O_2823,N_24769,N_24800);
nand UO_2824 (O_2824,N_24977,N_24994);
or UO_2825 (O_2825,N_24799,N_24835);
nor UO_2826 (O_2826,N_24840,N_24780);
and UO_2827 (O_2827,N_24912,N_24875);
or UO_2828 (O_2828,N_24871,N_24952);
or UO_2829 (O_2829,N_24879,N_24891);
xnor UO_2830 (O_2830,N_24791,N_24983);
xor UO_2831 (O_2831,N_24877,N_24853);
and UO_2832 (O_2832,N_24871,N_24980);
xor UO_2833 (O_2833,N_24800,N_24826);
or UO_2834 (O_2834,N_24926,N_24781);
xnor UO_2835 (O_2835,N_24778,N_24839);
nor UO_2836 (O_2836,N_24894,N_24838);
or UO_2837 (O_2837,N_24769,N_24874);
and UO_2838 (O_2838,N_24963,N_24848);
or UO_2839 (O_2839,N_24893,N_24903);
or UO_2840 (O_2840,N_24838,N_24772);
or UO_2841 (O_2841,N_24790,N_24870);
or UO_2842 (O_2842,N_24953,N_24818);
nor UO_2843 (O_2843,N_24770,N_24944);
nand UO_2844 (O_2844,N_24960,N_24957);
and UO_2845 (O_2845,N_24904,N_24975);
nand UO_2846 (O_2846,N_24975,N_24771);
nand UO_2847 (O_2847,N_24967,N_24928);
xnor UO_2848 (O_2848,N_24777,N_24861);
xor UO_2849 (O_2849,N_24999,N_24914);
or UO_2850 (O_2850,N_24944,N_24985);
or UO_2851 (O_2851,N_24821,N_24864);
nor UO_2852 (O_2852,N_24849,N_24842);
xnor UO_2853 (O_2853,N_24841,N_24934);
or UO_2854 (O_2854,N_24994,N_24770);
and UO_2855 (O_2855,N_24760,N_24859);
and UO_2856 (O_2856,N_24838,N_24824);
and UO_2857 (O_2857,N_24764,N_24944);
nor UO_2858 (O_2858,N_24843,N_24750);
nand UO_2859 (O_2859,N_24879,N_24819);
and UO_2860 (O_2860,N_24925,N_24943);
nor UO_2861 (O_2861,N_24931,N_24845);
xor UO_2862 (O_2862,N_24967,N_24914);
nor UO_2863 (O_2863,N_24845,N_24928);
or UO_2864 (O_2864,N_24981,N_24788);
xor UO_2865 (O_2865,N_24967,N_24896);
or UO_2866 (O_2866,N_24886,N_24954);
xor UO_2867 (O_2867,N_24943,N_24866);
and UO_2868 (O_2868,N_24754,N_24944);
nor UO_2869 (O_2869,N_24802,N_24861);
and UO_2870 (O_2870,N_24770,N_24827);
or UO_2871 (O_2871,N_24998,N_24772);
and UO_2872 (O_2872,N_24946,N_24899);
nor UO_2873 (O_2873,N_24827,N_24934);
xnor UO_2874 (O_2874,N_24958,N_24954);
or UO_2875 (O_2875,N_24951,N_24868);
nor UO_2876 (O_2876,N_24859,N_24862);
nor UO_2877 (O_2877,N_24899,N_24875);
nor UO_2878 (O_2878,N_24811,N_24900);
nand UO_2879 (O_2879,N_24771,N_24876);
nor UO_2880 (O_2880,N_24888,N_24885);
nor UO_2881 (O_2881,N_24854,N_24983);
and UO_2882 (O_2882,N_24806,N_24932);
nor UO_2883 (O_2883,N_24861,N_24874);
xor UO_2884 (O_2884,N_24877,N_24794);
and UO_2885 (O_2885,N_24810,N_24876);
or UO_2886 (O_2886,N_24974,N_24827);
nand UO_2887 (O_2887,N_24940,N_24938);
nor UO_2888 (O_2888,N_24949,N_24980);
xnor UO_2889 (O_2889,N_24997,N_24888);
nor UO_2890 (O_2890,N_24882,N_24827);
xor UO_2891 (O_2891,N_24939,N_24815);
nor UO_2892 (O_2892,N_24837,N_24934);
nor UO_2893 (O_2893,N_24959,N_24774);
or UO_2894 (O_2894,N_24896,N_24755);
or UO_2895 (O_2895,N_24971,N_24750);
and UO_2896 (O_2896,N_24957,N_24901);
nor UO_2897 (O_2897,N_24969,N_24837);
and UO_2898 (O_2898,N_24992,N_24858);
nand UO_2899 (O_2899,N_24860,N_24769);
nor UO_2900 (O_2900,N_24984,N_24909);
and UO_2901 (O_2901,N_24790,N_24932);
or UO_2902 (O_2902,N_24979,N_24815);
and UO_2903 (O_2903,N_24922,N_24929);
xnor UO_2904 (O_2904,N_24899,N_24893);
nor UO_2905 (O_2905,N_24896,N_24952);
nor UO_2906 (O_2906,N_24760,N_24950);
xnor UO_2907 (O_2907,N_24973,N_24901);
nand UO_2908 (O_2908,N_24948,N_24863);
nand UO_2909 (O_2909,N_24892,N_24856);
xnor UO_2910 (O_2910,N_24847,N_24786);
nand UO_2911 (O_2911,N_24966,N_24820);
or UO_2912 (O_2912,N_24992,N_24786);
and UO_2913 (O_2913,N_24912,N_24940);
or UO_2914 (O_2914,N_24890,N_24967);
nand UO_2915 (O_2915,N_24997,N_24932);
nand UO_2916 (O_2916,N_24918,N_24954);
or UO_2917 (O_2917,N_24904,N_24760);
and UO_2918 (O_2918,N_24990,N_24932);
nand UO_2919 (O_2919,N_24976,N_24752);
xor UO_2920 (O_2920,N_24751,N_24902);
nand UO_2921 (O_2921,N_24802,N_24947);
xnor UO_2922 (O_2922,N_24892,N_24980);
nand UO_2923 (O_2923,N_24903,N_24812);
nand UO_2924 (O_2924,N_24754,N_24995);
nand UO_2925 (O_2925,N_24801,N_24776);
xnor UO_2926 (O_2926,N_24763,N_24976);
and UO_2927 (O_2927,N_24769,N_24753);
and UO_2928 (O_2928,N_24783,N_24867);
or UO_2929 (O_2929,N_24866,N_24751);
nor UO_2930 (O_2930,N_24973,N_24889);
and UO_2931 (O_2931,N_24994,N_24791);
xor UO_2932 (O_2932,N_24858,N_24820);
xnor UO_2933 (O_2933,N_24864,N_24896);
nor UO_2934 (O_2934,N_24870,N_24914);
nand UO_2935 (O_2935,N_24832,N_24925);
nand UO_2936 (O_2936,N_24919,N_24852);
nand UO_2937 (O_2937,N_24853,N_24784);
xor UO_2938 (O_2938,N_24971,N_24993);
and UO_2939 (O_2939,N_24791,N_24939);
nor UO_2940 (O_2940,N_24757,N_24931);
xnor UO_2941 (O_2941,N_24777,N_24936);
or UO_2942 (O_2942,N_24828,N_24815);
or UO_2943 (O_2943,N_24959,N_24790);
nand UO_2944 (O_2944,N_24821,N_24989);
or UO_2945 (O_2945,N_24936,N_24895);
nor UO_2946 (O_2946,N_24990,N_24962);
or UO_2947 (O_2947,N_24862,N_24848);
xnor UO_2948 (O_2948,N_24960,N_24845);
nor UO_2949 (O_2949,N_24970,N_24786);
or UO_2950 (O_2950,N_24787,N_24953);
nor UO_2951 (O_2951,N_24976,N_24815);
and UO_2952 (O_2952,N_24785,N_24957);
or UO_2953 (O_2953,N_24975,N_24903);
or UO_2954 (O_2954,N_24773,N_24863);
nor UO_2955 (O_2955,N_24981,N_24796);
nor UO_2956 (O_2956,N_24879,N_24997);
xnor UO_2957 (O_2957,N_24962,N_24928);
nor UO_2958 (O_2958,N_24770,N_24913);
or UO_2959 (O_2959,N_24822,N_24815);
and UO_2960 (O_2960,N_24769,N_24751);
xnor UO_2961 (O_2961,N_24913,N_24776);
or UO_2962 (O_2962,N_24758,N_24936);
or UO_2963 (O_2963,N_24926,N_24956);
xor UO_2964 (O_2964,N_24797,N_24989);
nand UO_2965 (O_2965,N_24773,N_24821);
and UO_2966 (O_2966,N_24830,N_24807);
and UO_2967 (O_2967,N_24783,N_24869);
xnor UO_2968 (O_2968,N_24910,N_24863);
nand UO_2969 (O_2969,N_24858,N_24887);
nor UO_2970 (O_2970,N_24911,N_24913);
xor UO_2971 (O_2971,N_24765,N_24953);
nor UO_2972 (O_2972,N_24895,N_24963);
nand UO_2973 (O_2973,N_24796,N_24982);
nand UO_2974 (O_2974,N_24895,N_24924);
nor UO_2975 (O_2975,N_24841,N_24989);
nor UO_2976 (O_2976,N_24755,N_24995);
nand UO_2977 (O_2977,N_24786,N_24945);
xnor UO_2978 (O_2978,N_24879,N_24972);
nand UO_2979 (O_2979,N_24961,N_24797);
xor UO_2980 (O_2980,N_24897,N_24817);
nand UO_2981 (O_2981,N_24956,N_24993);
and UO_2982 (O_2982,N_24805,N_24782);
and UO_2983 (O_2983,N_24801,N_24872);
nand UO_2984 (O_2984,N_24949,N_24895);
and UO_2985 (O_2985,N_24836,N_24996);
and UO_2986 (O_2986,N_24890,N_24822);
xnor UO_2987 (O_2987,N_24983,N_24764);
nand UO_2988 (O_2988,N_24890,N_24862);
or UO_2989 (O_2989,N_24969,N_24784);
xnor UO_2990 (O_2990,N_24791,N_24906);
or UO_2991 (O_2991,N_24914,N_24924);
or UO_2992 (O_2992,N_24954,N_24801);
or UO_2993 (O_2993,N_24895,N_24911);
xor UO_2994 (O_2994,N_24901,N_24850);
or UO_2995 (O_2995,N_24857,N_24841);
nand UO_2996 (O_2996,N_24953,N_24753);
nor UO_2997 (O_2997,N_24848,N_24823);
nand UO_2998 (O_2998,N_24775,N_24760);
nor UO_2999 (O_2999,N_24886,N_24999);
endmodule