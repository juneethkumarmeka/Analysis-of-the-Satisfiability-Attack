module basic_1000_10000_1500_2_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5001,N_5002,N_5003,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5013,N_5014,N_5021,N_5023,N_5024,N_5025,N_5028,N_5030,N_5032,N_5033,N_5034,N_5035,N_5037,N_5038,N_5039,N_5044,N_5045,N_5047,N_5050,N_5053,N_5055,N_5056,N_5057,N_5060,N_5061,N_5065,N_5070,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5080,N_5081,N_5083,N_5088,N_5089,N_5091,N_5093,N_5096,N_5097,N_5099,N_5100,N_5102,N_5104,N_5105,N_5106,N_5107,N_5109,N_5111,N_5115,N_5116,N_5117,N_5118,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5130,N_5132,N_5136,N_5137,N_5138,N_5139,N_5140,N_5142,N_5145,N_5146,N_5151,N_5154,N_5155,N_5157,N_5158,N_5163,N_5164,N_5166,N_5167,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5180,N_5181,N_5183,N_5184,N_5186,N_5187,N_5188,N_5189,N_5190,N_5193,N_5194,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5209,N_5210,N_5211,N_5213,N_5215,N_5216,N_5217,N_5220,N_5222,N_5223,N_5228,N_5231,N_5232,N_5233,N_5234,N_5236,N_5237,N_5243,N_5244,N_5245,N_5249,N_5251,N_5253,N_5255,N_5258,N_5259,N_5262,N_5263,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5275,N_5276,N_5278,N_5279,N_5280,N_5283,N_5284,N_5286,N_5287,N_5288,N_5291,N_5292,N_5294,N_5295,N_5296,N_5300,N_5301,N_5304,N_5305,N_5306,N_5307,N_5310,N_5311,N_5313,N_5314,N_5317,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5330,N_5331,N_5333,N_5334,N_5335,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5344,N_5346,N_5347,N_5348,N_5349,N_5351,N_5352,N_5353,N_5354,N_5355,N_5358,N_5359,N_5360,N_5361,N_5363,N_5364,N_5365,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5376,N_5377,N_5378,N_5380,N_5382,N_5383,N_5385,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5398,N_5401,N_5402,N_5403,N_5404,N_5406,N_5408,N_5409,N_5410,N_5411,N_5413,N_5414,N_5416,N_5418,N_5419,N_5425,N_5426,N_5427,N_5430,N_5431,N_5433,N_5435,N_5437,N_5438,N_5439,N_5441,N_5445,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5456,N_5457,N_5460,N_5461,N_5462,N_5464,N_5465,N_5467,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5477,N_5478,N_5481,N_5482,N_5483,N_5484,N_5487,N_5488,N_5490,N_5493,N_5494,N_5495,N_5497,N_5498,N_5500,N_5501,N_5502,N_5503,N_5504,N_5507,N_5509,N_5510,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5522,N_5524,N_5526,N_5527,N_5533,N_5534,N_5535,N_5536,N_5538,N_5540,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5552,N_5554,N_5557,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5573,N_5575,N_5576,N_5578,N_5579,N_5582,N_5583,N_5584,N_5588,N_5589,N_5590,N_5592,N_5593,N_5598,N_5599,N_5601,N_5603,N_5604,N_5605,N_5606,N_5608,N_5610,N_5611,N_5613,N_5614,N_5619,N_5620,N_5622,N_5624,N_5626,N_5627,N_5628,N_5629,N_5631,N_5633,N_5635,N_5636,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5650,N_5652,N_5653,N_5655,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5665,N_5668,N_5670,N_5671,N_5672,N_5674,N_5676,N_5677,N_5678,N_5680,N_5682,N_5684,N_5685,N_5686,N_5687,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5699,N_5701,N_5702,N_5703,N_5705,N_5706,N_5708,N_5709,N_5715,N_5717,N_5719,N_5721,N_5722,N_5723,N_5724,N_5725,N_5728,N_5729,N_5730,N_5732,N_5733,N_5734,N_5738,N_5739,N_5740,N_5742,N_5743,N_5745,N_5746,N_5747,N_5748,N_5749,N_5754,N_5755,N_5757,N_5758,N_5759,N_5762,N_5763,N_5768,N_5769,N_5770,N_5772,N_5779,N_5780,N_5782,N_5783,N_5785,N_5788,N_5790,N_5791,N_5793,N_5799,N_5805,N_5806,N_5807,N_5808,N_5809,N_5811,N_5812,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5821,N_5823,N_5824,N_5825,N_5826,N_5828,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5837,N_5838,N_5840,N_5841,N_5843,N_5844,N_5845,N_5846,N_5851,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5864,N_5867,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5886,N_5888,N_5890,N_5891,N_5892,N_5893,N_5896,N_5897,N_5898,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5909,N_5910,N_5912,N_5914,N_5915,N_5917,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5930,N_5931,N_5935,N_5936,N_5937,N_5943,N_5944,N_5945,N_5947,N_5948,N_5950,N_5952,N_5953,N_5954,N_5955,N_5956,N_5958,N_5959,N_5960,N_5961,N_5962,N_5966,N_5968,N_5969,N_5971,N_5972,N_5976,N_5977,N_5978,N_5979,N_5980,N_5983,N_5984,N_5987,N_5990,N_5991,N_5992,N_5994,N_5996,N_5999,N_6002,N_6003,N_6004,N_6005,N_6006,N_6009,N_6011,N_6014,N_6015,N_6018,N_6019,N_6021,N_6022,N_6023,N_6025,N_6027,N_6029,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6040,N_6042,N_6044,N_6047,N_6048,N_6049,N_6050,N_6052,N_6054,N_6056,N_6057,N_6061,N_6062,N_6063,N_6064,N_6066,N_6070,N_6071,N_6073,N_6077,N_6078,N_6079,N_6081,N_6083,N_6084,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6093,N_6094,N_6095,N_6098,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6110,N_6113,N_6115,N_6116,N_6117,N_6120,N_6121,N_6122,N_6124,N_6125,N_6126,N_6128,N_6129,N_6130,N_6131,N_6132,N_6135,N_6138,N_6139,N_6143,N_6144,N_6147,N_6148,N_6150,N_6151,N_6152,N_6153,N_6156,N_6157,N_6162,N_6165,N_6166,N_6168,N_6169,N_6170,N_6171,N_6173,N_6174,N_6175,N_6176,N_6178,N_6183,N_6184,N_6186,N_6187,N_6188,N_6189,N_6190,N_6193,N_6194,N_6196,N_6201,N_6204,N_6205,N_6206,N_6207,N_6208,N_6210,N_6211,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6220,N_6221,N_6223,N_6227,N_6228,N_6234,N_6237,N_6242,N_6243,N_6244,N_6246,N_6247,N_6252,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6262,N_6266,N_6267,N_6268,N_6271,N_6272,N_6274,N_6275,N_6280,N_6281,N_6283,N_6284,N_6285,N_6288,N_6289,N_6290,N_6291,N_6293,N_6294,N_6296,N_6297,N_6300,N_6301,N_6302,N_6305,N_6306,N_6308,N_6309,N_6311,N_6312,N_6314,N_6315,N_6322,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6331,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6342,N_6344,N_6346,N_6347,N_6348,N_6349,N_6350,N_6352,N_6353,N_6354,N_6355,N_6357,N_6359,N_6360,N_6361,N_6366,N_6368,N_6371,N_6372,N_6374,N_6375,N_6376,N_6379,N_6382,N_6386,N_6388,N_6389,N_6390,N_6392,N_6395,N_6396,N_6397,N_6398,N_6399,N_6401,N_6404,N_6406,N_6407,N_6408,N_6410,N_6413,N_6414,N_6415,N_6416,N_6419,N_6421,N_6422,N_6423,N_6424,N_6425,N_6429,N_6430,N_6431,N_6434,N_6439,N_6440,N_6442,N_6443,N_6444,N_6445,N_6446,N_6448,N_6449,N_6450,N_6451,N_6452,N_6454,N_6456,N_6457,N_6458,N_6459,N_6462,N_6464,N_6465,N_6466,N_6467,N_6468,N_6472,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6483,N_6484,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6496,N_6497,N_6498,N_6503,N_6504,N_6505,N_6508,N_6509,N_6510,N_6513,N_6514,N_6518,N_6520,N_6523,N_6524,N_6526,N_6528,N_6529,N_6530,N_6531,N_6532,N_6534,N_6535,N_6536,N_6538,N_6539,N_6540,N_6541,N_6542,N_6545,N_6546,N_6547,N_6548,N_6551,N_6552,N_6553,N_6554,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6571,N_6573,N_6576,N_6577,N_6579,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6588,N_6590,N_6595,N_6597,N_6600,N_6601,N_6602,N_6604,N_6606,N_6608,N_6609,N_6614,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6630,N_6631,N_6633,N_6635,N_6636,N_6637,N_6640,N_6641,N_6643,N_6644,N_6645,N_6646,N_6650,N_6654,N_6655,N_6656,N_6657,N_6658,N_6660,N_6661,N_6667,N_6668,N_6670,N_6671,N_6673,N_6675,N_6679,N_6681,N_6682,N_6685,N_6686,N_6687,N_6689,N_6690,N_6694,N_6695,N_6696,N_6699,N_6700,N_6703,N_6704,N_6708,N_6709,N_6710,N_6714,N_6716,N_6719,N_6721,N_6722,N_6727,N_6728,N_6729,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6739,N_6740,N_6741,N_6742,N_6743,N_6745,N_6747,N_6749,N_6750,N_6752,N_6753,N_6754,N_6755,N_6759,N_6760,N_6762,N_6763,N_6764,N_6765,N_6767,N_6768,N_6769,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6778,N_6780,N_6781,N_6783,N_6784,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6793,N_6794,N_6797,N_6799,N_6801,N_6802,N_6803,N_6804,N_6805,N_6807,N_6811,N_6812,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6825,N_6826,N_6828,N_6829,N_6832,N_6833,N_6835,N_6836,N_6837,N_6838,N_6839,N_6842,N_6843,N_6844,N_6845,N_6848,N_6851,N_6852,N_6854,N_6855,N_6857,N_6858,N_6859,N_6863,N_6865,N_6867,N_6868,N_6869,N_6870,N_6871,N_6874,N_6877,N_6878,N_6879,N_6880,N_6882,N_6884,N_6885,N_6886,N_6889,N_6891,N_6893,N_6894,N_6897,N_6898,N_6900,N_6901,N_6903,N_6907,N_6908,N_6909,N_6912,N_6913,N_6917,N_6919,N_6921,N_6922,N_6924,N_6925,N_6926,N_6928,N_6930,N_6931,N_6932,N_6933,N_6935,N_6936,N_6938,N_6939,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6948,N_6950,N_6951,N_6952,N_6954,N_6955,N_6956,N_6957,N_6959,N_6961,N_6962,N_6963,N_6965,N_6966,N_6967,N_6968,N_6972,N_6976,N_6978,N_6981,N_6982,N_6983,N_6984,N_6986,N_6987,N_6989,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7004,N_7006,N_7008,N_7009,N_7011,N_7015,N_7016,N_7022,N_7023,N_7026,N_7027,N_7028,N_7030,N_7031,N_7034,N_7035,N_7037,N_7039,N_7041,N_7043,N_7046,N_7047,N_7049,N_7051,N_7052,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7063,N_7066,N_7068,N_7069,N_7071,N_7072,N_7073,N_7075,N_7077,N_7078,N_7080,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7089,N_7090,N_7091,N_7093,N_7094,N_7095,N_7097,N_7098,N_7100,N_7101,N_7102,N_7103,N_7106,N_7107,N_7108,N_7110,N_7111,N_7114,N_7115,N_7117,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7130,N_7131,N_7136,N_7137,N_7139,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7150,N_7155,N_7156,N_7159,N_7160,N_7161,N_7164,N_7165,N_7168,N_7172,N_7173,N_7176,N_7177,N_7180,N_7181,N_7183,N_7184,N_7185,N_7188,N_7189,N_7190,N_7191,N_7194,N_7195,N_7196,N_7198,N_7200,N_7202,N_7204,N_7205,N_7206,N_7207,N_7208,N_7210,N_7215,N_7216,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7233,N_7234,N_7236,N_7237,N_7238,N_7240,N_7241,N_7243,N_7245,N_7246,N_7247,N_7248,N_7254,N_7257,N_7258,N_7259,N_7261,N_7262,N_7264,N_7267,N_7268,N_7270,N_7271,N_7274,N_7275,N_7276,N_7277,N_7278,N_7280,N_7281,N_7284,N_7285,N_7286,N_7287,N_7288,N_7291,N_7293,N_7294,N_7297,N_7298,N_7299,N_7300,N_7304,N_7307,N_7308,N_7309,N_7310,N_7311,N_7313,N_7314,N_7317,N_7318,N_7319,N_7320,N_7321,N_7323,N_7325,N_7326,N_7327,N_7329,N_7330,N_7331,N_7335,N_7336,N_7337,N_7339,N_7340,N_7341,N_7342,N_7343,N_7345,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7357,N_7358,N_7359,N_7361,N_7362,N_7363,N_7366,N_7367,N_7369,N_7373,N_7374,N_7375,N_7376,N_7380,N_7381,N_7382,N_7384,N_7385,N_7386,N_7388,N_7390,N_7392,N_7393,N_7396,N_7398,N_7399,N_7400,N_7401,N_7404,N_7406,N_7408,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7422,N_7423,N_7425,N_7427,N_7428,N_7430,N_7431,N_7432,N_7433,N_7435,N_7436,N_7437,N_7438,N_7440,N_7442,N_7444,N_7445,N_7446,N_7448,N_7451,N_7452,N_7453,N_7454,N_7455,N_7458,N_7459,N_7460,N_7461,N_7462,N_7465,N_7468,N_7470,N_7471,N_7473,N_7475,N_7477,N_7479,N_7480,N_7481,N_7483,N_7485,N_7487,N_7488,N_7490,N_7492,N_7493,N_7496,N_7497,N_7500,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7513,N_7517,N_7518,N_7519,N_7520,N_7523,N_7524,N_7526,N_7528,N_7529,N_7531,N_7533,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7547,N_7548,N_7551,N_7552,N_7553,N_7559,N_7563,N_7564,N_7565,N_7567,N_7569,N_7570,N_7573,N_7574,N_7575,N_7576,N_7577,N_7580,N_7581,N_7582,N_7583,N_7586,N_7587,N_7588,N_7589,N_7590,N_7593,N_7595,N_7598,N_7599,N_7600,N_7602,N_7603,N_7604,N_7606,N_7607,N_7608,N_7609,N_7611,N_7612,N_7613,N_7615,N_7616,N_7617,N_7618,N_7620,N_7624,N_7626,N_7628,N_7631,N_7633,N_7635,N_7639,N_7640,N_7642,N_7643,N_7646,N_7649,N_7650,N_7652,N_7654,N_7655,N_7657,N_7659,N_7660,N_7661,N_7662,N_7664,N_7666,N_7668,N_7669,N_7670,N_7671,N_7672,N_7674,N_7680,N_7682,N_7684,N_7685,N_7688,N_7689,N_7691,N_7692,N_7693,N_7696,N_7700,N_7704,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7715,N_7716,N_7717,N_7720,N_7721,N_7722,N_7723,N_7724,N_7727,N_7729,N_7734,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7745,N_7748,N_7749,N_7751,N_7753,N_7754,N_7758,N_7759,N_7762,N_7763,N_7764,N_7765,N_7766,N_7768,N_7770,N_7771,N_7774,N_7775,N_7776,N_7778,N_7779,N_7780,N_7784,N_7792,N_7794,N_7796,N_7800,N_7802,N_7803,N_7804,N_7807,N_7810,N_7812,N_7813,N_7816,N_7820,N_7821,N_7823,N_7826,N_7827,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7838,N_7839,N_7842,N_7843,N_7844,N_7846,N_7849,N_7850,N_7851,N_7853,N_7854,N_7855,N_7857,N_7858,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7869,N_7870,N_7872,N_7873,N_7874,N_7875,N_7878,N_7881,N_7883,N_7884,N_7886,N_7887,N_7888,N_7890,N_7891,N_7892,N_7895,N_7897,N_7899,N_7901,N_7902,N_7903,N_7905,N_7906,N_7907,N_7908,N_7911,N_7912,N_7914,N_7917,N_7921,N_7922,N_7925,N_7930,N_7933,N_7934,N_7935,N_7937,N_7939,N_7940,N_7941,N_7945,N_7952,N_7953,N_7956,N_7957,N_7958,N_7959,N_7961,N_7963,N_7964,N_7965,N_7966,N_7967,N_7970,N_7971,N_7973,N_7974,N_7976,N_7977,N_7979,N_7980,N_7983,N_7985,N_7986,N_7989,N_7990,N_7991,N_7992,N_7993,N_7999,N_8001,N_8002,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8020,N_8023,N_8024,N_8025,N_8028,N_8029,N_8030,N_8031,N_8034,N_8037,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8046,N_8048,N_8049,N_8050,N_8054,N_8058,N_8060,N_8061,N_8062,N_8063,N_8065,N_8066,N_8067,N_8068,N_8070,N_8071,N_8072,N_8075,N_8076,N_8077,N_8082,N_8083,N_8085,N_8089,N_8090,N_8093,N_8094,N_8096,N_8097,N_8098,N_8099,N_8101,N_8102,N_8103,N_8104,N_8106,N_8107,N_8108,N_8109,N_8110,N_8112,N_8113,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8124,N_8126,N_8127,N_8130,N_8131,N_8132,N_8134,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8143,N_8145,N_8146,N_8147,N_8148,N_8149,N_8151,N_8157,N_8158,N_8160,N_8161,N_8163,N_8164,N_8165,N_8166,N_8167,N_8169,N_8170,N_8173,N_8174,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8185,N_8189,N_8190,N_8192,N_8195,N_8196,N_8197,N_8199,N_8201,N_8203,N_8204,N_8205,N_8206,N_8209,N_8211,N_8212,N_8215,N_8216,N_8217,N_8219,N_8220,N_8223,N_8225,N_8228,N_8229,N_8230,N_8231,N_8232,N_8234,N_8235,N_8236,N_8237,N_8238,N_8242,N_8243,N_8244,N_8248,N_8249,N_8253,N_8254,N_8258,N_8259,N_8260,N_8261,N_8263,N_8264,N_8267,N_8269,N_8270,N_8271,N_8273,N_8274,N_8278,N_8280,N_8282,N_8284,N_8286,N_8288,N_8290,N_8293,N_8295,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8307,N_8308,N_8310,N_8312,N_8313,N_8314,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8324,N_8325,N_8330,N_8333,N_8334,N_8336,N_8337,N_8339,N_8340,N_8341,N_8344,N_8348,N_8351,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8367,N_8371,N_8372,N_8376,N_8378,N_8379,N_8380,N_8382,N_8383,N_8386,N_8387,N_8388,N_8390,N_8391,N_8392,N_8393,N_8397,N_8398,N_8399,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8410,N_8411,N_8412,N_8413,N_8415,N_8416,N_8417,N_8418,N_8421,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8435,N_8436,N_8437,N_8438,N_8440,N_8444,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8455,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8467,N_8469,N_8470,N_8472,N_8475,N_8477,N_8478,N_8480,N_8481,N_8482,N_8483,N_8486,N_8487,N_8488,N_8491,N_8492,N_8493,N_8495,N_8496,N_8497,N_8498,N_8500,N_8501,N_8502,N_8506,N_8507,N_8508,N_8509,N_8511,N_8513,N_8514,N_8515,N_8517,N_8518,N_8520,N_8521,N_8523,N_8525,N_8526,N_8529,N_8530,N_8531,N_8532,N_8540,N_8542,N_8543,N_8544,N_8546,N_8547,N_8549,N_8551,N_8552,N_8554,N_8557,N_8558,N_8560,N_8563,N_8566,N_8567,N_8572,N_8573,N_8574,N_8577,N_8580,N_8583,N_8585,N_8586,N_8587,N_8588,N_8589,N_8591,N_8594,N_8596,N_8597,N_8598,N_8600,N_8601,N_8603,N_8604,N_8605,N_8608,N_8609,N_8610,N_8612,N_8613,N_8615,N_8616,N_8617,N_8620,N_8621,N_8622,N_8623,N_8624,N_8626,N_8627,N_8628,N_8630,N_8631,N_8632,N_8633,N_8634,N_8637,N_8638,N_8639,N_8640,N_8644,N_8648,N_8649,N_8650,N_8651,N_8652,N_8654,N_8658,N_8659,N_8660,N_8663,N_8664,N_8665,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8678,N_8681,N_8682,N_8683,N_8685,N_8686,N_8687,N_8688,N_8689,N_8692,N_8693,N_8694,N_8695,N_8697,N_8700,N_8701,N_8703,N_8704,N_8705,N_8707,N_8709,N_8710,N_8711,N_8712,N_8713,N_8716,N_8717,N_8718,N_8721,N_8723,N_8726,N_8728,N_8729,N_8731,N_8732,N_8733,N_8735,N_8737,N_8739,N_8741,N_8742,N_8744,N_8745,N_8746,N_8747,N_8748,N_8750,N_8751,N_8753,N_8756,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8766,N_8768,N_8772,N_8773,N_8774,N_8775,N_8777,N_8778,N_8779,N_8781,N_8783,N_8784,N_8786,N_8787,N_8788,N_8794,N_8795,N_8796,N_8797,N_8799,N_8801,N_8803,N_8804,N_8805,N_8806,N_8810,N_8814,N_8815,N_8816,N_8818,N_8821,N_8822,N_8825,N_8826,N_8827,N_8831,N_8832,N_8835,N_8836,N_8837,N_8838,N_8840,N_8841,N_8842,N_8843,N_8845,N_8849,N_8851,N_8852,N_8853,N_8855,N_8856,N_8857,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8868,N_8869,N_8870,N_8872,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8889,N_8890,N_8892,N_8893,N_8895,N_8896,N_8898,N_8902,N_8903,N_8906,N_8909,N_8911,N_8913,N_8915,N_8918,N_8919,N_8920,N_8922,N_8924,N_8925,N_8926,N_8930,N_8931,N_8933,N_8934,N_8935,N_8939,N_8941,N_8942,N_8943,N_8944,N_8946,N_8949,N_8952,N_8954,N_8955,N_8957,N_8958,N_8960,N_8961,N_8964,N_8965,N_8969,N_8971,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8991,N_8992,N_8996,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9005,N_9006,N_9007,N_9008,N_9010,N_9013,N_9014,N_9015,N_9017,N_9018,N_9021,N_9022,N_9024,N_9025,N_9026,N_9027,N_9029,N_9030,N_9031,N_9033,N_9036,N_9038,N_9043,N_9044,N_9045,N_9046,N_9047,N_9049,N_9050,N_9053,N_9054,N_9055,N_9057,N_9058,N_9059,N_9060,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9080,N_9081,N_9082,N_9083,N_9084,N_9086,N_9087,N_9088,N_9089,N_9091,N_9092,N_9096,N_9099,N_9101,N_9103,N_9106,N_9108,N_9111,N_9112,N_9113,N_9114,N_9115,N_9117,N_9118,N_9119,N_9121,N_9123,N_9124,N_9125,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9137,N_9139,N_9140,N_9141,N_9142,N_9144,N_9145,N_9146,N_9150,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9160,N_9161,N_9162,N_9163,N_9165,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9174,N_9176,N_9178,N_9182,N_9186,N_9187,N_9189,N_9191,N_9192,N_9194,N_9195,N_9202,N_9203,N_9205,N_9210,N_9211,N_9212,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9221,N_9223,N_9225,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9237,N_9238,N_9239,N_9242,N_9244,N_9245,N_9248,N_9249,N_9252,N_9253,N_9254,N_9255,N_9257,N_9259,N_9260,N_9262,N_9266,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9291,N_9292,N_9293,N_9297,N_9298,N_9300,N_9301,N_9304,N_9306,N_9307,N_9309,N_9310,N_9311,N_9312,N_9314,N_9315,N_9316,N_9317,N_9320,N_9321,N_9322,N_9323,N_9325,N_9331,N_9332,N_9333,N_9336,N_9338,N_9339,N_9341,N_9342,N_9344,N_9346,N_9347,N_9348,N_9349,N_9352,N_9353,N_9354,N_9355,N_9357,N_9358,N_9359,N_9360,N_9362,N_9363,N_9364,N_9366,N_9367,N_9368,N_9369,N_9370,N_9373,N_9374,N_9376,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9387,N_9389,N_9391,N_9394,N_9395,N_9396,N_9398,N_9399,N_9402,N_9403,N_9405,N_9409,N_9410,N_9412,N_9413,N_9415,N_9417,N_9419,N_9420,N_9421,N_9422,N_9423,N_9425,N_9426,N_9428,N_9429,N_9430,N_9433,N_9434,N_9435,N_9436,N_9438,N_9439,N_9440,N_9442,N_9443,N_9444,N_9446,N_9448,N_9451,N_9452,N_9456,N_9457,N_9460,N_9461,N_9463,N_9464,N_9466,N_9467,N_9468,N_9469,N_9475,N_9477,N_9478,N_9480,N_9481,N_9484,N_9487,N_9488,N_9489,N_9490,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9503,N_9504,N_9505,N_9508,N_9509,N_9512,N_9513,N_9515,N_9516,N_9517,N_9519,N_9523,N_9525,N_9526,N_9527,N_9529,N_9532,N_9534,N_9535,N_9537,N_9538,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9553,N_9556,N_9557,N_9558,N_9560,N_9562,N_9564,N_9566,N_9567,N_9569,N_9570,N_9576,N_9577,N_9579,N_9580,N_9583,N_9584,N_9586,N_9588,N_9589,N_9590,N_9592,N_9595,N_9596,N_9597,N_9598,N_9601,N_9602,N_9603,N_9605,N_9606,N_9607,N_9608,N_9610,N_9611,N_9612,N_9613,N_9615,N_9616,N_9617,N_9619,N_9621,N_9623,N_9624,N_9626,N_9628,N_9631,N_9632,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9646,N_9648,N_9649,N_9650,N_9654,N_9655,N_9656,N_9657,N_9659,N_9663,N_9665,N_9667,N_9670,N_9672,N_9676,N_9677,N_9678,N_9679,N_9681,N_9683,N_9684,N_9685,N_9686,N_9687,N_9691,N_9692,N_9693,N_9695,N_9700,N_9701,N_9702,N_9705,N_9708,N_9710,N_9712,N_9717,N_9718,N_9719,N_9722,N_9723,N_9727,N_9729,N_9730,N_9731,N_9732,N_9737,N_9738,N_9741,N_9743,N_9748,N_9749,N_9750,N_9751,N_9753,N_9754,N_9755,N_9757,N_9758,N_9761,N_9762,N_9764,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9774,N_9775,N_9783,N_9784,N_9786,N_9787,N_9790,N_9791,N_9792,N_9793,N_9795,N_9797,N_9798,N_9801,N_9803,N_9805,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9816,N_9817,N_9818,N_9821,N_9824,N_9825,N_9827,N_9828,N_9829,N_9832,N_9834,N_9835,N_9836,N_9837,N_9838,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9859,N_9860,N_9862,N_9863,N_9864,N_9867,N_9868,N_9871,N_9872,N_9875,N_9876,N_9877,N_9878,N_9881,N_9885,N_9887,N_9889,N_9890,N_9891,N_9892,N_9894,N_9895,N_9897,N_9898,N_9900,N_9901,N_9902,N_9907,N_9908,N_9909,N_9910,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9919,N_9924,N_9926,N_9931,N_9933,N_9934,N_9935,N_9936,N_9938,N_9940,N_9941,N_9942,N_9943,N_9945,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9955,N_9957,N_9958,N_9959,N_9962,N_9966,N_9967,N_9973,N_9974,N_9975,N_9977,N_9978,N_9979,N_9980,N_9981,N_9984,N_9986,N_9987,N_9991,N_9992,N_9995,N_9996,N_9998,N_9999;
and U0 (N_0,In_500,In_974);
or U1 (N_1,In_618,In_227);
nor U2 (N_2,In_557,In_178);
xnor U3 (N_3,In_341,In_738);
nand U4 (N_4,In_773,In_816);
nor U5 (N_5,In_718,In_496);
nand U6 (N_6,In_774,In_754);
or U7 (N_7,In_20,In_890);
or U8 (N_8,In_471,In_592);
and U9 (N_9,In_111,In_719);
xnor U10 (N_10,In_884,In_89);
and U11 (N_11,In_934,In_583);
or U12 (N_12,In_770,In_271);
and U13 (N_13,In_748,In_840);
nor U14 (N_14,In_595,In_625);
or U15 (N_15,In_425,In_80);
nand U16 (N_16,In_538,In_165);
nand U17 (N_17,In_732,In_485);
or U18 (N_18,In_530,In_250);
nand U19 (N_19,In_503,In_932);
nand U20 (N_20,In_358,In_286);
or U21 (N_21,In_217,In_906);
nor U22 (N_22,In_190,In_104);
nor U23 (N_23,In_326,In_237);
nand U24 (N_24,In_376,In_836);
or U25 (N_25,In_465,In_173);
nor U26 (N_26,In_815,In_486);
or U27 (N_27,In_631,In_479);
or U28 (N_28,In_148,In_25);
nand U29 (N_29,In_848,In_222);
and U30 (N_30,In_612,In_208);
nor U31 (N_31,In_454,In_438);
nor U32 (N_32,In_593,In_751);
nor U33 (N_33,In_188,In_877);
and U34 (N_34,In_299,In_501);
or U35 (N_35,In_517,In_586);
nand U36 (N_36,In_229,In_123);
nor U37 (N_37,In_135,In_643);
and U38 (N_38,In_895,In_183);
and U39 (N_39,In_636,In_931);
or U40 (N_40,In_985,In_708);
or U41 (N_41,In_675,In_524);
nand U42 (N_42,In_131,In_457);
nor U43 (N_43,In_713,In_555);
and U44 (N_44,In_377,In_186);
xnor U45 (N_45,In_975,In_633);
nor U46 (N_46,In_180,In_16);
nand U47 (N_47,In_752,In_772);
nand U48 (N_48,In_126,In_319);
and U49 (N_49,In_615,In_847);
nor U50 (N_50,In_144,In_857);
or U51 (N_51,In_936,In_296);
and U52 (N_52,In_494,In_887);
or U53 (N_53,In_771,In_150);
nor U54 (N_54,In_843,In_921);
and U55 (N_55,In_100,In_32);
and U56 (N_56,In_819,In_584);
and U57 (N_57,In_176,In_458);
or U58 (N_58,In_408,In_291);
and U59 (N_59,In_775,In_629);
nand U60 (N_60,In_546,In_415);
nand U61 (N_61,In_858,In_410);
and U62 (N_62,In_572,In_269);
nand U63 (N_63,In_39,In_516);
and U64 (N_64,In_670,In_422);
nand U65 (N_65,In_317,In_842);
and U66 (N_66,In_927,In_396);
nand U67 (N_67,In_810,In_78);
and U68 (N_68,In_203,In_363);
nor U69 (N_69,In_303,In_833);
or U70 (N_70,In_147,In_107);
and U71 (N_71,In_321,In_912);
or U72 (N_72,In_266,In_556);
and U73 (N_73,In_63,In_276);
or U74 (N_74,In_917,In_978);
nand U75 (N_75,In_506,In_994);
or U76 (N_76,In_431,In_657);
and U77 (N_77,In_864,In_987);
nand U78 (N_78,In_66,In_806);
nand U79 (N_79,In_798,In_54);
and U80 (N_80,In_329,In_582);
or U81 (N_81,In_862,In_692);
and U82 (N_82,In_813,In_574);
or U83 (N_83,In_273,In_22);
and U84 (N_84,In_98,In_310);
and U85 (N_85,In_225,In_268);
nand U86 (N_86,In_280,In_43);
nor U87 (N_87,In_255,In_325);
nand U88 (N_88,In_720,In_620);
nand U89 (N_89,In_980,In_818);
or U90 (N_90,In_929,In_984);
and U91 (N_91,In_497,In_627);
nand U92 (N_92,In_866,In_328);
and U93 (N_93,In_499,In_821);
nand U94 (N_94,In_743,In_294);
nor U95 (N_95,In_982,In_248);
and U96 (N_96,In_852,In_99);
nor U97 (N_97,In_507,In_102);
nor U98 (N_98,In_172,In_502);
or U99 (N_99,In_232,In_382);
nor U100 (N_100,In_215,In_849);
and U101 (N_101,In_691,In_312);
nand U102 (N_102,In_826,In_683);
or U103 (N_103,In_746,In_449);
and U104 (N_104,In_401,In_558);
nand U105 (N_105,In_324,In_529);
nand U106 (N_106,In_990,In_734);
nor U107 (N_107,In_292,In_809);
nor U108 (N_108,In_421,In_570);
and U109 (N_109,In_699,In_249);
nor U110 (N_110,In_967,In_694);
nor U111 (N_111,In_483,In_820);
nor U112 (N_112,In_939,In_76);
nor U113 (N_113,In_999,In_366);
nor U114 (N_114,In_976,In_653);
and U115 (N_115,In_903,In_715);
or U116 (N_116,In_608,In_542);
or U117 (N_117,In_690,In_997);
nor U118 (N_118,In_776,In_265);
nand U119 (N_119,In_70,In_744);
and U120 (N_120,In_941,In_461);
and U121 (N_121,In_834,In_17);
nand U122 (N_122,In_198,In_588);
nor U123 (N_123,In_88,In_441);
nand U124 (N_124,In_474,In_221);
nor U125 (N_125,In_938,In_49);
and U126 (N_126,In_606,In_737);
nand U127 (N_127,In_220,In_343);
nor U128 (N_128,In_455,In_837);
nand U129 (N_129,In_440,In_405);
nor U130 (N_130,In_196,In_12);
nand U131 (N_131,In_892,In_124);
nand U132 (N_132,In_65,In_492);
or U133 (N_133,In_381,In_640);
nor U134 (N_134,In_874,In_412);
nand U135 (N_135,In_308,In_762);
nand U136 (N_136,In_240,In_136);
nor U137 (N_137,In_375,In_62);
or U138 (N_138,In_672,In_965);
nor U139 (N_139,In_780,In_48);
and U140 (N_140,In_913,In_119);
or U141 (N_141,In_52,In_498);
xor U142 (N_142,In_56,In_693);
or U143 (N_143,In_716,In_753);
and U144 (N_144,In_860,In_665);
or U145 (N_145,In_658,In_908);
and U146 (N_146,In_493,In_400);
and U147 (N_147,In_561,In_766);
or U148 (N_148,In_814,In_649);
nor U149 (N_149,In_623,In_345);
or U150 (N_150,In_962,In_210);
nor U151 (N_151,In_742,In_6);
nand U152 (N_152,In_365,In_706);
nor U153 (N_153,In_897,In_241);
or U154 (N_154,In_611,In_85);
nor U155 (N_155,In_21,In_424);
nor U156 (N_156,In_477,In_96);
and U157 (N_157,In_263,In_224);
nand U158 (N_158,In_423,In_669);
nor U159 (N_159,In_270,In_945);
or U160 (N_160,In_130,In_831);
nor U161 (N_161,In_384,In_302);
nor U162 (N_162,In_537,In_77);
nor U163 (N_163,In_703,In_86);
nand U164 (N_164,In_246,In_407);
or U165 (N_165,In_368,In_369);
nand U166 (N_166,In_552,In_433);
or U167 (N_167,In_207,In_597);
and U168 (N_168,In_782,In_630);
and U169 (N_169,In_191,In_406);
and U170 (N_170,In_152,In_184);
nand U171 (N_171,In_947,In_937);
nand U172 (N_172,In_617,In_998);
nor U173 (N_173,In_888,In_260);
or U174 (N_174,In_889,In_698);
nand U175 (N_175,In_609,In_958);
and U176 (N_176,In_125,In_656);
or U177 (N_177,In_374,In_568);
nand U178 (N_178,In_654,In_614);
and U179 (N_179,In_995,In_515);
or U180 (N_180,In_581,In_540);
and U181 (N_181,In_404,In_37);
and U182 (N_182,In_74,In_340);
nor U183 (N_183,In_613,In_3);
and U184 (N_184,In_437,In_855);
nor U185 (N_185,In_961,In_214);
and U186 (N_186,In_704,In_488);
nand U187 (N_187,In_940,In_262);
or U188 (N_188,In_372,In_952);
nand U189 (N_189,In_277,In_791);
or U190 (N_190,In_235,In_315);
nand U191 (N_191,In_311,In_784);
nand U192 (N_192,In_149,In_680);
or U193 (N_193,In_469,In_946);
nand U194 (N_194,In_101,In_769);
nand U195 (N_195,In_92,In_579);
or U196 (N_196,In_659,In_896);
and U197 (N_197,In_571,In_259);
nand U198 (N_198,In_907,In_764);
xor U199 (N_199,In_676,In_953);
or U200 (N_200,In_812,In_380);
nor U201 (N_201,In_881,In_914);
nand U202 (N_202,In_31,In_272);
or U203 (N_203,In_899,In_389);
or U204 (N_204,In_370,In_918);
nor U205 (N_205,In_520,In_484);
and U206 (N_206,In_601,In_393);
nor U207 (N_207,In_662,In_242);
nand U208 (N_208,In_120,In_607);
and U209 (N_209,In_795,In_414);
or U210 (N_210,In_105,In_632);
or U211 (N_211,In_674,In_443);
and U212 (N_212,In_979,In_828);
and U213 (N_213,In_970,In_373);
and U214 (N_214,In_724,In_922);
nor U215 (N_215,In_853,In_948);
and U216 (N_216,In_830,In_371);
xor U217 (N_217,In_599,In_863);
nand U218 (N_218,In_468,In_902);
nor U219 (N_219,In_205,In_297);
nor U220 (N_220,In_236,In_445);
or U221 (N_221,In_228,In_60);
or U222 (N_222,In_452,In_949);
nor U223 (N_223,In_304,In_256);
nor U224 (N_224,In_508,In_278);
nand U225 (N_225,In_346,In_456);
and U226 (N_226,In_434,In_331);
or U227 (N_227,In_564,In_915);
or U228 (N_228,In_40,In_977);
and U229 (N_229,In_689,In_113);
nor U230 (N_230,In_44,In_344);
nand U231 (N_231,In_53,In_58);
and U232 (N_232,In_824,In_963);
nor U233 (N_233,In_285,In_578);
and U234 (N_234,In_886,In_204);
and U235 (N_235,In_306,In_551);
nor U236 (N_236,In_827,In_712);
and U237 (N_237,In_986,In_905);
nor U238 (N_238,In_67,In_846);
or U239 (N_239,In_154,In_330);
and U240 (N_240,In_335,In_731);
xor U241 (N_241,In_347,In_314);
nand U242 (N_242,In_298,In_115);
or U243 (N_243,In_153,In_167);
or U244 (N_244,In_349,In_655);
nand U245 (N_245,In_252,In_851);
and U246 (N_246,In_75,In_893);
and U247 (N_247,In_996,In_287);
or U248 (N_248,In_175,In_528);
nor U249 (N_249,In_158,In_24);
nor U250 (N_250,In_829,In_935);
or U251 (N_251,In_900,In_333);
nand U252 (N_252,In_856,In_671);
nor U253 (N_253,In_554,In_591);
nand U254 (N_254,In_293,In_57);
and U255 (N_255,In_223,In_413);
nand U256 (N_256,In_361,In_687);
nor U257 (N_257,In_392,In_789);
or U258 (N_258,In_476,In_177);
nor U259 (N_259,In_402,In_450);
nor U260 (N_260,In_391,In_518);
nand U261 (N_261,In_122,In_234);
or U262 (N_262,In_710,In_957);
nand U263 (N_263,In_390,In_467);
and U264 (N_264,In_805,In_462);
nand U265 (N_265,In_489,In_447);
and U266 (N_266,In_761,In_850);
or U267 (N_267,In_735,In_417);
and U268 (N_268,In_811,In_141);
or U269 (N_269,In_94,In_109);
and U270 (N_270,In_543,In_127);
nor U271 (N_271,In_663,In_162);
and U272 (N_272,In_602,In_245);
nand U273 (N_273,In_928,In_202);
and U274 (N_274,In_28,In_8);
and U275 (N_275,In_721,In_960);
nand U276 (N_276,In_650,In_164);
nand U277 (N_277,In_71,In_7);
nor U278 (N_278,In_352,In_861);
nor U279 (N_279,In_134,In_868);
and U280 (N_280,In_81,In_835);
and U281 (N_281,In_169,In_30);
and U282 (N_282,In_128,In_825);
or U283 (N_283,In_702,In_667);
or U284 (N_284,In_394,In_759);
nor U285 (N_285,In_334,In_736);
nor U286 (N_286,In_513,In_527);
nand U287 (N_287,In_420,In_803);
nand U288 (N_288,In_727,In_93);
and U289 (N_289,In_968,In_45);
or U290 (N_290,In_364,In_729);
nand U291 (N_291,In_487,In_589);
nor U292 (N_292,In_714,In_788);
and U293 (N_293,In_399,In_356);
and U294 (N_294,In_726,In_218);
xor U295 (N_295,In_114,In_637);
nor U296 (N_296,In_750,In_757);
or U297 (N_297,In_981,In_639);
nand U298 (N_298,In_573,In_925);
and U299 (N_299,In_47,In_875);
or U300 (N_300,In_274,In_84);
or U301 (N_301,In_873,In_403);
nand U302 (N_302,In_845,In_920);
nand U303 (N_303,In_876,In_351);
nor U304 (N_304,In_563,In_869);
and U305 (N_305,In_504,In_569);
and U306 (N_306,In_944,In_785);
and U307 (N_307,In_163,In_604);
or U308 (N_308,In_741,In_59);
and U309 (N_309,In_289,In_865);
nor U310 (N_310,In_9,In_709);
nor U311 (N_311,In_992,In_733);
nor U312 (N_312,In_779,In_257);
or U313 (N_313,In_323,In_185);
and U314 (N_314,In_90,In_679);
nand U315 (N_315,In_661,In_332);
nor U316 (N_316,In_478,In_435);
or U317 (N_317,In_264,In_839);
and U318 (N_318,In_547,In_802);
and U319 (N_319,In_969,In_495);
nor U320 (N_320,In_796,In_82);
nor U321 (N_321,In_660,In_348);
nor U322 (N_322,In_580,In_27);
nor U323 (N_323,In_682,In_747);
or U324 (N_324,In_490,In_778);
nand U325 (N_325,In_418,In_168);
nand U326 (N_326,In_686,In_97);
nand U327 (N_327,In_281,In_531);
nand U328 (N_328,In_439,In_666);
nand U329 (N_329,In_238,In_605);
or U330 (N_330,In_339,In_73);
nand U331 (N_331,In_510,In_219);
and U332 (N_332,In_678,In_916);
nor U333 (N_333,In_521,In_132);
nand U334 (N_334,In_541,In_787);
or U335 (N_335,In_910,In_777);
nor U336 (N_336,In_956,In_472);
or U337 (N_337,In_626,In_247);
nor U338 (N_338,In_398,In_179);
nor U339 (N_339,In_919,In_426);
and U340 (N_340,In_146,In_129);
nor U341 (N_341,In_35,In_951);
or U342 (N_342,In_212,In_475);
nor U343 (N_343,In_275,In_797);
nand U344 (N_344,In_891,In_705);
or U345 (N_345,In_139,In_522);
and U346 (N_346,In_505,In_594);
or U347 (N_347,In_972,In_231);
and U348 (N_348,In_117,In_526);
and U349 (N_349,In_318,In_0);
and U350 (N_350,In_768,In_717);
nor U351 (N_351,In_622,In_879);
or U352 (N_352,In_790,In_195);
or U353 (N_353,In_781,In_901);
nor U354 (N_354,In_353,In_587);
or U355 (N_355,In_695,In_133);
nor U356 (N_356,In_585,In_383);
or U357 (N_357,In_544,In_320);
and U358 (N_358,In_519,In_282);
or U359 (N_359,In_385,In_959);
and U360 (N_360,In_964,In_201);
and U361 (N_361,In_145,In_924);
nand U362 (N_362,In_397,In_577);
and U363 (N_363,In_446,In_942);
or U364 (N_364,In_598,In_971);
nand U365 (N_365,In_182,In_562);
and U366 (N_366,In_432,In_616);
or U367 (N_367,In_4,In_156);
or U368 (N_368,In_251,In_233);
and U369 (N_369,In_711,In_668);
nor U370 (N_370,In_295,In_10);
nand U371 (N_371,In_696,In_428);
nor U372 (N_372,In_808,In_646);
or U373 (N_373,In_955,In_95);
and U374 (N_374,In_41,In_549);
and U375 (N_375,In_26,In_46);
and U376 (N_376,In_641,In_429);
and U377 (N_377,In_253,In_697);
nand U378 (N_378,In_822,In_159);
nand U379 (N_379,In_336,In_444);
nor U380 (N_380,In_64,In_137);
or U381 (N_381,In_239,In_230);
and U382 (N_382,In_898,In_756);
or U383 (N_383,In_823,In_322);
or U384 (N_384,In_871,In_38);
or U385 (N_385,In_430,In_973);
nor U386 (N_386,In_170,In_923);
and U387 (N_387,In_553,In_142);
or U388 (N_388,In_279,In_290);
and U389 (N_389,In_387,In_792);
and U390 (N_390,In_15,In_909);
and U391 (N_391,In_647,In_832);
and U392 (N_392,In_739,In_118);
xor U393 (N_393,In_13,In_560);
nand U394 (N_394,In_301,In_197);
xnor U395 (N_395,In_327,In_859);
or U396 (N_396,In_254,In_23);
nand U397 (N_397,In_470,In_395);
or U398 (N_398,In_379,In_596);
nand U399 (N_399,In_50,In_313);
nor U400 (N_400,In_480,In_192);
and U401 (N_401,In_993,In_817);
or U402 (N_402,In_619,In_463);
nor U403 (N_403,In_590,In_29);
nor U404 (N_404,In_106,In_989);
nand U405 (N_405,In_841,In_83);
or U406 (N_406,In_894,In_648);
nor U407 (N_407,In_532,In_652);
and U408 (N_408,In_359,In_638);
nand U409 (N_409,In_350,In_566);
or U410 (N_410,In_645,In_760);
or U411 (N_411,In_800,In_700);
or U412 (N_412,In_804,In_793);
nor U413 (N_413,In_309,In_110);
nand U414 (N_414,In_688,In_966);
and U415 (N_415,In_155,In_464);
and U416 (N_416,In_261,In_283);
or U417 (N_417,In_491,In_885);
and U418 (N_418,In_36,In_878);
nand U419 (N_419,In_765,In_5);
nor U420 (N_420,In_536,In_116);
xor U421 (N_421,In_193,In_157);
nand U422 (N_422,In_416,In_872);
and U423 (N_423,In_386,In_69);
and U424 (N_424,In_466,In_728);
and U425 (N_425,In_883,In_342);
nor U426 (N_426,In_644,In_535);
or U427 (N_427,In_11,In_621);
nand U428 (N_428,In_151,In_539);
nor U429 (N_429,In_783,In_799);
nor U430 (N_430,In_870,In_844);
or U431 (N_431,In_243,In_904);
xnor U432 (N_432,In_473,In_211);
and U433 (N_433,In_482,In_305);
and U434 (N_434,In_161,In_533);
nand U435 (N_435,In_174,In_300);
and U436 (N_436,In_226,In_87);
nand U437 (N_437,In_681,In_725);
or U438 (N_438,In_801,In_481);
nand U439 (N_439,In_258,In_189);
nor U440 (N_440,In_51,In_701);
or U441 (N_441,In_545,In_61);
nor U442 (N_442,In_360,In_288);
and U443 (N_443,In_453,In_103);
or U444 (N_444,In_685,In_565);
or U445 (N_445,In_33,In_509);
nand U446 (N_446,In_388,In_988);
nor U447 (N_447,In_677,In_459);
nor U448 (N_448,In_112,In_880);
or U449 (N_449,In_603,In_930);
and U450 (N_450,In_807,In_673);
nand U451 (N_451,In_138,In_284);
nand U452 (N_452,In_514,In_200);
nor U453 (N_453,In_635,In_18);
nand U454 (N_454,In_436,In_550);
and U455 (N_455,In_943,In_451);
nand U456 (N_456,In_378,In_749);
and U457 (N_457,In_79,In_991);
or U458 (N_458,In_427,In_723);
or U459 (N_459,In_357,In_338);
nand U460 (N_460,In_181,In_911);
and U461 (N_461,In_367,In_448);
or U462 (N_462,In_337,In_19);
nand U463 (N_463,In_316,In_722);
nand U464 (N_464,In_307,In_624);
nand U465 (N_465,In_460,In_525);
nor U466 (N_466,In_854,In_763);
or U467 (N_467,In_42,In_419);
or U468 (N_468,In_642,In_206);
nand U469 (N_469,In_511,In_409);
nor U470 (N_470,In_664,In_160);
nand U471 (N_471,In_55,In_355);
nand U472 (N_472,In_882,In_121);
and U473 (N_473,In_213,In_767);
or U474 (N_474,In_628,In_548);
and U475 (N_475,In_267,In_72);
nor U476 (N_476,In_143,In_730);
and U477 (N_477,In_108,In_216);
nand U478 (N_478,In_34,In_14);
and U479 (N_479,In_244,In_534);
and U480 (N_480,In_171,In_794);
nand U481 (N_481,In_194,In_755);
nor U482 (N_482,In_933,In_684);
and U483 (N_483,In_576,In_166);
nand U484 (N_484,In_634,In_926);
nand U485 (N_485,In_950,In_651);
or U486 (N_486,In_786,In_2);
or U487 (N_487,In_199,In_600);
and U488 (N_488,In_140,In_707);
nor U489 (N_489,In_362,In_740);
or U490 (N_490,In_575,In_411);
or U491 (N_491,In_745,In_1);
nand U492 (N_492,In_187,In_91);
or U493 (N_493,In_983,In_209);
nand U494 (N_494,In_354,In_567);
and U495 (N_495,In_523,In_867);
and U496 (N_496,In_442,In_512);
and U497 (N_497,In_954,In_68);
and U498 (N_498,In_610,In_559);
and U499 (N_499,In_838,In_758);
nand U500 (N_500,In_793,In_859);
and U501 (N_501,In_528,In_205);
nand U502 (N_502,In_826,In_6);
nand U503 (N_503,In_485,In_981);
or U504 (N_504,In_905,In_677);
and U505 (N_505,In_206,In_342);
nand U506 (N_506,In_752,In_510);
nand U507 (N_507,In_676,In_140);
nor U508 (N_508,In_996,In_804);
and U509 (N_509,In_63,In_759);
and U510 (N_510,In_506,In_353);
and U511 (N_511,In_655,In_192);
or U512 (N_512,In_547,In_341);
or U513 (N_513,In_267,In_261);
nand U514 (N_514,In_131,In_594);
nand U515 (N_515,In_184,In_676);
xor U516 (N_516,In_99,In_438);
and U517 (N_517,In_726,In_377);
nand U518 (N_518,In_905,In_742);
or U519 (N_519,In_366,In_983);
or U520 (N_520,In_931,In_94);
xor U521 (N_521,In_722,In_677);
and U522 (N_522,In_989,In_908);
nand U523 (N_523,In_495,In_305);
and U524 (N_524,In_426,In_149);
or U525 (N_525,In_580,In_917);
and U526 (N_526,In_71,In_345);
nor U527 (N_527,In_631,In_638);
and U528 (N_528,In_651,In_805);
or U529 (N_529,In_458,In_691);
nand U530 (N_530,In_485,In_589);
nand U531 (N_531,In_369,In_265);
nand U532 (N_532,In_326,In_655);
nand U533 (N_533,In_903,In_448);
or U534 (N_534,In_212,In_954);
nor U535 (N_535,In_71,In_532);
or U536 (N_536,In_506,In_867);
nor U537 (N_537,In_985,In_346);
nor U538 (N_538,In_938,In_753);
and U539 (N_539,In_520,In_181);
xnor U540 (N_540,In_649,In_947);
or U541 (N_541,In_243,In_702);
and U542 (N_542,In_163,In_715);
nand U543 (N_543,In_835,In_544);
nand U544 (N_544,In_827,In_730);
nand U545 (N_545,In_511,In_919);
or U546 (N_546,In_905,In_942);
nor U547 (N_547,In_28,In_648);
and U548 (N_548,In_27,In_622);
nand U549 (N_549,In_654,In_490);
nand U550 (N_550,In_133,In_983);
nand U551 (N_551,In_334,In_9);
xnor U552 (N_552,In_544,In_311);
or U553 (N_553,In_779,In_263);
nand U554 (N_554,In_838,In_862);
or U555 (N_555,In_678,In_479);
and U556 (N_556,In_448,In_71);
and U557 (N_557,In_768,In_813);
and U558 (N_558,In_480,In_698);
or U559 (N_559,In_388,In_156);
or U560 (N_560,In_338,In_668);
and U561 (N_561,In_501,In_27);
and U562 (N_562,In_733,In_109);
nand U563 (N_563,In_307,In_604);
and U564 (N_564,In_0,In_227);
or U565 (N_565,In_649,In_691);
nor U566 (N_566,In_886,In_282);
nand U567 (N_567,In_175,In_974);
and U568 (N_568,In_457,In_259);
nand U569 (N_569,In_559,In_869);
nand U570 (N_570,In_224,In_322);
or U571 (N_571,In_716,In_338);
nor U572 (N_572,In_158,In_610);
or U573 (N_573,In_816,In_692);
and U574 (N_574,In_788,In_398);
and U575 (N_575,In_223,In_163);
nand U576 (N_576,In_480,In_618);
nor U577 (N_577,In_277,In_113);
and U578 (N_578,In_50,In_546);
or U579 (N_579,In_738,In_109);
nor U580 (N_580,In_672,In_786);
xnor U581 (N_581,In_408,In_839);
nor U582 (N_582,In_748,In_46);
nand U583 (N_583,In_231,In_389);
and U584 (N_584,In_650,In_803);
and U585 (N_585,In_599,In_694);
and U586 (N_586,In_498,In_579);
and U587 (N_587,In_613,In_492);
or U588 (N_588,In_848,In_635);
nand U589 (N_589,In_528,In_124);
nand U590 (N_590,In_682,In_720);
and U591 (N_591,In_595,In_735);
nor U592 (N_592,In_628,In_678);
nor U593 (N_593,In_811,In_264);
and U594 (N_594,In_48,In_912);
or U595 (N_595,In_743,In_583);
nand U596 (N_596,In_16,In_768);
and U597 (N_597,In_988,In_571);
and U598 (N_598,In_417,In_934);
nor U599 (N_599,In_496,In_49);
nand U600 (N_600,In_539,In_135);
or U601 (N_601,In_781,In_356);
and U602 (N_602,In_916,In_302);
nor U603 (N_603,In_619,In_566);
nand U604 (N_604,In_907,In_371);
and U605 (N_605,In_19,In_830);
or U606 (N_606,In_336,In_163);
or U607 (N_607,In_787,In_466);
or U608 (N_608,In_179,In_594);
and U609 (N_609,In_46,In_267);
nor U610 (N_610,In_943,In_768);
nand U611 (N_611,In_572,In_660);
nand U612 (N_612,In_944,In_766);
nand U613 (N_613,In_346,In_351);
nand U614 (N_614,In_622,In_42);
and U615 (N_615,In_403,In_561);
and U616 (N_616,In_397,In_947);
nor U617 (N_617,In_459,In_977);
nand U618 (N_618,In_856,In_664);
nand U619 (N_619,In_595,In_416);
nor U620 (N_620,In_32,In_942);
or U621 (N_621,In_853,In_870);
and U622 (N_622,In_550,In_685);
nor U623 (N_623,In_834,In_903);
nor U624 (N_624,In_139,In_453);
or U625 (N_625,In_751,In_353);
and U626 (N_626,In_137,In_978);
xor U627 (N_627,In_925,In_933);
or U628 (N_628,In_524,In_411);
nor U629 (N_629,In_803,In_233);
nand U630 (N_630,In_254,In_156);
nand U631 (N_631,In_727,In_799);
nor U632 (N_632,In_907,In_464);
and U633 (N_633,In_982,In_959);
nor U634 (N_634,In_666,In_521);
and U635 (N_635,In_795,In_484);
nand U636 (N_636,In_98,In_926);
or U637 (N_637,In_425,In_263);
xnor U638 (N_638,In_682,In_223);
nand U639 (N_639,In_394,In_216);
and U640 (N_640,In_673,In_116);
and U641 (N_641,In_58,In_986);
or U642 (N_642,In_193,In_865);
or U643 (N_643,In_83,In_486);
xnor U644 (N_644,In_895,In_673);
nand U645 (N_645,In_889,In_409);
or U646 (N_646,In_608,In_136);
nor U647 (N_647,In_398,In_741);
and U648 (N_648,In_44,In_666);
nand U649 (N_649,In_276,In_583);
nor U650 (N_650,In_193,In_6);
nor U651 (N_651,In_838,In_885);
or U652 (N_652,In_893,In_70);
and U653 (N_653,In_580,In_86);
nand U654 (N_654,In_684,In_850);
nor U655 (N_655,In_498,In_957);
nor U656 (N_656,In_587,In_529);
nand U657 (N_657,In_763,In_321);
or U658 (N_658,In_653,In_850);
nand U659 (N_659,In_813,In_60);
nor U660 (N_660,In_124,In_894);
and U661 (N_661,In_529,In_192);
or U662 (N_662,In_123,In_588);
and U663 (N_663,In_462,In_597);
and U664 (N_664,In_496,In_365);
nor U665 (N_665,In_832,In_967);
and U666 (N_666,In_163,In_951);
nor U667 (N_667,In_824,In_36);
nand U668 (N_668,In_639,In_968);
or U669 (N_669,In_282,In_182);
nor U670 (N_670,In_875,In_244);
and U671 (N_671,In_764,In_265);
nor U672 (N_672,In_358,In_965);
nor U673 (N_673,In_448,In_845);
or U674 (N_674,In_66,In_626);
and U675 (N_675,In_471,In_318);
nor U676 (N_676,In_608,In_318);
or U677 (N_677,In_176,In_213);
or U678 (N_678,In_998,In_281);
nor U679 (N_679,In_886,In_682);
nor U680 (N_680,In_45,In_937);
nor U681 (N_681,In_389,In_619);
nand U682 (N_682,In_32,In_76);
or U683 (N_683,In_558,In_687);
or U684 (N_684,In_772,In_31);
xnor U685 (N_685,In_115,In_5);
nor U686 (N_686,In_346,In_46);
and U687 (N_687,In_228,In_325);
nor U688 (N_688,In_536,In_865);
and U689 (N_689,In_536,In_602);
and U690 (N_690,In_793,In_78);
nor U691 (N_691,In_594,In_946);
or U692 (N_692,In_514,In_292);
and U693 (N_693,In_18,In_412);
xor U694 (N_694,In_441,In_305);
and U695 (N_695,In_15,In_18);
and U696 (N_696,In_575,In_588);
nand U697 (N_697,In_983,In_895);
or U698 (N_698,In_980,In_759);
or U699 (N_699,In_879,In_830);
or U700 (N_700,In_183,In_648);
nor U701 (N_701,In_938,In_512);
nand U702 (N_702,In_182,In_478);
and U703 (N_703,In_869,In_244);
xnor U704 (N_704,In_586,In_744);
and U705 (N_705,In_530,In_531);
nor U706 (N_706,In_636,In_635);
nor U707 (N_707,In_635,In_460);
nor U708 (N_708,In_487,In_988);
nand U709 (N_709,In_342,In_638);
nand U710 (N_710,In_550,In_889);
and U711 (N_711,In_729,In_966);
or U712 (N_712,In_852,In_579);
xnor U713 (N_713,In_581,In_590);
and U714 (N_714,In_979,In_506);
nor U715 (N_715,In_568,In_40);
and U716 (N_716,In_968,In_17);
nor U717 (N_717,In_423,In_535);
xnor U718 (N_718,In_518,In_617);
nor U719 (N_719,In_220,In_509);
nand U720 (N_720,In_305,In_74);
or U721 (N_721,In_927,In_520);
nor U722 (N_722,In_147,In_711);
or U723 (N_723,In_143,In_856);
or U724 (N_724,In_946,In_509);
nor U725 (N_725,In_31,In_418);
nor U726 (N_726,In_95,In_143);
or U727 (N_727,In_93,In_884);
nor U728 (N_728,In_840,In_560);
nor U729 (N_729,In_347,In_788);
nor U730 (N_730,In_948,In_304);
nand U731 (N_731,In_230,In_894);
or U732 (N_732,In_27,In_136);
and U733 (N_733,In_311,In_887);
or U734 (N_734,In_161,In_87);
and U735 (N_735,In_286,In_582);
nand U736 (N_736,In_613,In_995);
or U737 (N_737,In_428,In_609);
nand U738 (N_738,In_708,In_253);
nand U739 (N_739,In_895,In_692);
nand U740 (N_740,In_256,In_66);
and U741 (N_741,In_462,In_585);
and U742 (N_742,In_110,In_520);
nand U743 (N_743,In_374,In_234);
or U744 (N_744,In_676,In_803);
and U745 (N_745,In_399,In_72);
nor U746 (N_746,In_153,In_915);
nor U747 (N_747,In_159,In_503);
or U748 (N_748,In_274,In_82);
and U749 (N_749,In_611,In_110);
nor U750 (N_750,In_221,In_920);
or U751 (N_751,In_555,In_185);
or U752 (N_752,In_37,In_712);
nor U753 (N_753,In_206,In_820);
nand U754 (N_754,In_120,In_725);
and U755 (N_755,In_302,In_604);
nor U756 (N_756,In_585,In_324);
and U757 (N_757,In_712,In_316);
nand U758 (N_758,In_560,In_994);
or U759 (N_759,In_118,In_741);
nand U760 (N_760,In_607,In_681);
nor U761 (N_761,In_688,In_942);
nor U762 (N_762,In_12,In_995);
nand U763 (N_763,In_121,In_459);
nor U764 (N_764,In_131,In_103);
nor U765 (N_765,In_187,In_490);
or U766 (N_766,In_597,In_897);
nand U767 (N_767,In_967,In_32);
and U768 (N_768,In_596,In_370);
nor U769 (N_769,In_61,In_645);
xor U770 (N_770,In_81,In_749);
nand U771 (N_771,In_370,In_266);
xnor U772 (N_772,In_599,In_662);
nand U773 (N_773,In_798,In_81);
nor U774 (N_774,In_988,In_647);
nor U775 (N_775,In_665,In_551);
or U776 (N_776,In_525,In_465);
nor U777 (N_777,In_901,In_915);
or U778 (N_778,In_761,In_233);
or U779 (N_779,In_945,In_337);
nor U780 (N_780,In_144,In_971);
nand U781 (N_781,In_371,In_757);
nor U782 (N_782,In_64,In_54);
or U783 (N_783,In_134,In_991);
or U784 (N_784,In_353,In_725);
and U785 (N_785,In_86,In_466);
and U786 (N_786,In_670,In_331);
and U787 (N_787,In_489,In_955);
and U788 (N_788,In_975,In_352);
xnor U789 (N_789,In_936,In_148);
nand U790 (N_790,In_818,In_647);
or U791 (N_791,In_455,In_592);
or U792 (N_792,In_633,In_907);
nor U793 (N_793,In_848,In_846);
and U794 (N_794,In_910,In_369);
or U795 (N_795,In_860,In_598);
nor U796 (N_796,In_545,In_902);
and U797 (N_797,In_358,In_125);
nor U798 (N_798,In_372,In_376);
nor U799 (N_799,In_772,In_196);
and U800 (N_800,In_98,In_399);
or U801 (N_801,In_961,In_154);
or U802 (N_802,In_340,In_406);
nor U803 (N_803,In_130,In_10);
and U804 (N_804,In_713,In_404);
and U805 (N_805,In_425,In_740);
and U806 (N_806,In_248,In_500);
xor U807 (N_807,In_960,In_733);
nor U808 (N_808,In_617,In_323);
and U809 (N_809,In_340,In_472);
or U810 (N_810,In_558,In_78);
nand U811 (N_811,In_380,In_806);
or U812 (N_812,In_684,In_121);
or U813 (N_813,In_648,In_397);
nand U814 (N_814,In_964,In_50);
nor U815 (N_815,In_635,In_242);
or U816 (N_816,In_326,In_136);
and U817 (N_817,In_686,In_294);
and U818 (N_818,In_823,In_724);
nand U819 (N_819,In_165,In_326);
nand U820 (N_820,In_973,In_366);
or U821 (N_821,In_449,In_325);
nand U822 (N_822,In_479,In_564);
or U823 (N_823,In_225,In_704);
nor U824 (N_824,In_817,In_415);
nand U825 (N_825,In_331,In_557);
and U826 (N_826,In_638,In_540);
nor U827 (N_827,In_897,In_541);
and U828 (N_828,In_407,In_876);
and U829 (N_829,In_445,In_774);
and U830 (N_830,In_355,In_671);
nand U831 (N_831,In_536,In_231);
or U832 (N_832,In_464,In_938);
or U833 (N_833,In_805,In_330);
or U834 (N_834,In_441,In_932);
and U835 (N_835,In_143,In_179);
or U836 (N_836,In_887,In_623);
or U837 (N_837,In_527,In_233);
nand U838 (N_838,In_291,In_541);
nand U839 (N_839,In_777,In_575);
or U840 (N_840,In_711,In_328);
xnor U841 (N_841,In_545,In_386);
or U842 (N_842,In_557,In_815);
nand U843 (N_843,In_282,In_512);
nor U844 (N_844,In_143,In_686);
and U845 (N_845,In_335,In_405);
and U846 (N_846,In_225,In_150);
or U847 (N_847,In_387,In_313);
nand U848 (N_848,In_242,In_670);
nor U849 (N_849,In_37,In_216);
xnor U850 (N_850,In_515,In_790);
nor U851 (N_851,In_359,In_558);
and U852 (N_852,In_771,In_471);
or U853 (N_853,In_287,In_807);
nand U854 (N_854,In_616,In_77);
and U855 (N_855,In_104,In_244);
nor U856 (N_856,In_733,In_916);
nor U857 (N_857,In_154,In_432);
and U858 (N_858,In_694,In_475);
xor U859 (N_859,In_241,In_894);
or U860 (N_860,In_620,In_722);
nor U861 (N_861,In_681,In_701);
and U862 (N_862,In_148,In_792);
nand U863 (N_863,In_808,In_604);
and U864 (N_864,In_754,In_434);
nand U865 (N_865,In_225,In_455);
nand U866 (N_866,In_228,In_935);
nor U867 (N_867,In_789,In_837);
or U868 (N_868,In_813,In_252);
or U869 (N_869,In_594,In_690);
nand U870 (N_870,In_262,In_562);
and U871 (N_871,In_881,In_70);
or U872 (N_872,In_615,In_478);
xor U873 (N_873,In_276,In_281);
and U874 (N_874,In_78,In_200);
nand U875 (N_875,In_33,In_303);
and U876 (N_876,In_48,In_948);
and U877 (N_877,In_356,In_984);
and U878 (N_878,In_61,In_662);
nand U879 (N_879,In_221,In_574);
or U880 (N_880,In_854,In_972);
and U881 (N_881,In_288,In_603);
and U882 (N_882,In_103,In_645);
nor U883 (N_883,In_416,In_526);
nor U884 (N_884,In_897,In_544);
nor U885 (N_885,In_623,In_897);
and U886 (N_886,In_965,In_906);
nand U887 (N_887,In_416,In_292);
nor U888 (N_888,In_829,In_204);
nor U889 (N_889,In_846,In_684);
or U890 (N_890,In_60,In_176);
nor U891 (N_891,In_716,In_217);
nor U892 (N_892,In_583,In_335);
nand U893 (N_893,In_12,In_987);
and U894 (N_894,In_82,In_949);
nor U895 (N_895,In_176,In_460);
nor U896 (N_896,In_59,In_433);
and U897 (N_897,In_998,In_429);
nand U898 (N_898,In_88,In_365);
or U899 (N_899,In_458,In_133);
or U900 (N_900,In_714,In_455);
or U901 (N_901,In_19,In_77);
and U902 (N_902,In_896,In_450);
and U903 (N_903,In_680,In_354);
nor U904 (N_904,In_617,In_597);
and U905 (N_905,In_625,In_150);
nor U906 (N_906,In_171,In_498);
and U907 (N_907,In_715,In_609);
nand U908 (N_908,In_212,In_833);
or U909 (N_909,In_237,In_735);
nor U910 (N_910,In_887,In_61);
or U911 (N_911,In_793,In_988);
nor U912 (N_912,In_449,In_113);
nor U913 (N_913,In_220,In_919);
and U914 (N_914,In_245,In_443);
or U915 (N_915,In_431,In_591);
and U916 (N_916,In_524,In_837);
and U917 (N_917,In_816,In_817);
nor U918 (N_918,In_338,In_779);
nor U919 (N_919,In_777,In_352);
and U920 (N_920,In_546,In_660);
or U921 (N_921,In_795,In_793);
nand U922 (N_922,In_860,In_699);
or U923 (N_923,In_612,In_856);
nor U924 (N_924,In_485,In_301);
nand U925 (N_925,In_66,In_278);
nand U926 (N_926,In_459,In_938);
and U927 (N_927,In_766,In_940);
nor U928 (N_928,In_716,In_333);
or U929 (N_929,In_131,In_487);
and U930 (N_930,In_519,In_53);
nand U931 (N_931,In_289,In_203);
nor U932 (N_932,In_718,In_98);
nand U933 (N_933,In_751,In_303);
nand U934 (N_934,In_17,In_430);
nor U935 (N_935,In_310,In_883);
or U936 (N_936,In_204,In_883);
and U937 (N_937,In_90,In_752);
nand U938 (N_938,In_742,In_577);
or U939 (N_939,In_766,In_895);
nor U940 (N_940,In_603,In_329);
or U941 (N_941,In_123,In_372);
or U942 (N_942,In_617,In_681);
nor U943 (N_943,In_715,In_381);
and U944 (N_944,In_423,In_856);
nand U945 (N_945,In_117,In_223);
nor U946 (N_946,In_667,In_981);
and U947 (N_947,In_728,In_664);
nor U948 (N_948,In_797,In_525);
and U949 (N_949,In_569,In_713);
nor U950 (N_950,In_740,In_732);
and U951 (N_951,In_45,In_913);
or U952 (N_952,In_762,In_103);
nor U953 (N_953,In_250,In_361);
or U954 (N_954,In_731,In_659);
nor U955 (N_955,In_325,In_184);
nand U956 (N_956,In_728,In_690);
nor U957 (N_957,In_138,In_687);
or U958 (N_958,In_789,In_757);
nor U959 (N_959,In_349,In_445);
and U960 (N_960,In_796,In_888);
nand U961 (N_961,In_777,In_213);
or U962 (N_962,In_117,In_266);
nand U963 (N_963,In_102,In_594);
or U964 (N_964,In_189,In_648);
and U965 (N_965,In_789,In_459);
nand U966 (N_966,In_160,In_538);
nand U967 (N_967,In_861,In_887);
nand U968 (N_968,In_755,In_540);
nor U969 (N_969,In_894,In_482);
nor U970 (N_970,In_650,In_741);
and U971 (N_971,In_339,In_618);
nand U972 (N_972,In_681,In_498);
nor U973 (N_973,In_910,In_646);
or U974 (N_974,In_934,In_939);
and U975 (N_975,In_550,In_933);
nand U976 (N_976,In_626,In_421);
or U977 (N_977,In_705,In_947);
and U978 (N_978,In_988,In_47);
and U979 (N_979,In_922,In_248);
or U980 (N_980,In_376,In_893);
and U981 (N_981,In_171,In_86);
nand U982 (N_982,In_150,In_213);
or U983 (N_983,In_599,In_867);
and U984 (N_984,In_810,In_569);
nand U985 (N_985,In_328,In_889);
xor U986 (N_986,In_304,In_19);
and U987 (N_987,In_11,In_205);
nand U988 (N_988,In_817,In_745);
nand U989 (N_989,In_451,In_759);
or U990 (N_990,In_244,In_12);
nor U991 (N_991,In_537,In_123);
and U992 (N_992,In_118,In_3);
or U993 (N_993,In_965,In_512);
or U994 (N_994,In_572,In_679);
nand U995 (N_995,In_78,In_40);
and U996 (N_996,In_475,In_883);
or U997 (N_997,In_748,In_684);
and U998 (N_998,In_979,In_167);
nor U999 (N_999,In_395,In_602);
or U1000 (N_1000,In_587,In_854);
nand U1001 (N_1001,In_42,In_394);
nand U1002 (N_1002,In_747,In_698);
xnor U1003 (N_1003,In_670,In_49);
nand U1004 (N_1004,In_541,In_222);
nand U1005 (N_1005,In_653,In_848);
or U1006 (N_1006,In_499,In_450);
xnor U1007 (N_1007,In_266,In_288);
or U1008 (N_1008,In_200,In_787);
nand U1009 (N_1009,In_664,In_297);
and U1010 (N_1010,In_890,In_634);
nand U1011 (N_1011,In_792,In_227);
and U1012 (N_1012,In_978,In_679);
nor U1013 (N_1013,In_159,In_761);
or U1014 (N_1014,In_520,In_15);
nor U1015 (N_1015,In_965,In_501);
nand U1016 (N_1016,In_971,In_454);
or U1017 (N_1017,In_719,In_911);
nor U1018 (N_1018,In_842,In_587);
and U1019 (N_1019,In_27,In_321);
and U1020 (N_1020,In_498,In_265);
or U1021 (N_1021,In_287,In_340);
nor U1022 (N_1022,In_675,In_323);
or U1023 (N_1023,In_436,In_503);
or U1024 (N_1024,In_137,In_452);
and U1025 (N_1025,In_999,In_513);
nor U1026 (N_1026,In_343,In_462);
nand U1027 (N_1027,In_637,In_303);
nand U1028 (N_1028,In_37,In_501);
nand U1029 (N_1029,In_861,In_45);
or U1030 (N_1030,In_138,In_148);
and U1031 (N_1031,In_206,In_712);
nor U1032 (N_1032,In_748,In_599);
nand U1033 (N_1033,In_987,In_453);
or U1034 (N_1034,In_862,In_61);
nor U1035 (N_1035,In_733,In_362);
nor U1036 (N_1036,In_396,In_176);
nor U1037 (N_1037,In_461,In_76);
nand U1038 (N_1038,In_769,In_888);
nand U1039 (N_1039,In_283,In_22);
and U1040 (N_1040,In_169,In_765);
nor U1041 (N_1041,In_495,In_856);
or U1042 (N_1042,In_83,In_982);
nor U1043 (N_1043,In_46,In_545);
nor U1044 (N_1044,In_510,In_693);
xor U1045 (N_1045,In_58,In_754);
or U1046 (N_1046,In_405,In_824);
and U1047 (N_1047,In_38,In_593);
and U1048 (N_1048,In_654,In_145);
nor U1049 (N_1049,In_831,In_633);
nor U1050 (N_1050,In_327,In_101);
nor U1051 (N_1051,In_280,In_306);
and U1052 (N_1052,In_68,In_965);
and U1053 (N_1053,In_635,In_850);
or U1054 (N_1054,In_113,In_887);
or U1055 (N_1055,In_906,In_376);
and U1056 (N_1056,In_696,In_734);
nand U1057 (N_1057,In_537,In_885);
and U1058 (N_1058,In_50,In_117);
nor U1059 (N_1059,In_68,In_278);
and U1060 (N_1060,In_209,In_515);
nor U1061 (N_1061,In_115,In_80);
nand U1062 (N_1062,In_149,In_369);
and U1063 (N_1063,In_808,In_629);
and U1064 (N_1064,In_784,In_251);
or U1065 (N_1065,In_796,In_34);
or U1066 (N_1066,In_229,In_539);
nor U1067 (N_1067,In_467,In_654);
nand U1068 (N_1068,In_535,In_814);
and U1069 (N_1069,In_606,In_180);
nor U1070 (N_1070,In_96,In_797);
or U1071 (N_1071,In_281,In_852);
or U1072 (N_1072,In_477,In_217);
nor U1073 (N_1073,In_862,In_480);
or U1074 (N_1074,In_234,In_798);
and U1075 (N_1075,In_695,In_991);
nand U1076 (N_1076,In_737,In_95);
nand U1077 (N_1077,In_514,In_57);
nor U1078 (N_1078,In_583,In_926);
nand U1079 (N_1079,In_742,In_303);
and U1080 (N_1080,In_599,In_13);
nor U1081 (N_1081,In_926,In_138);
nor U1082 (N_1082,In_564,In_617);
nor U1083 (N_1083,In_730,In_19);
or U1084 (N_1084,In_273,In_392);
nand U1085 (N_1085,In_272,In_564);
or U1086 (N_1086,In_90,In_602);
and U1087 (N_1087,In_349,In_901);
and U1088 (N_1088,In_75,In_121);
nand U1089 (N_1089,In_631,In_484);
nand U1090 (N_1090,In_479,In_77);
and U1091 (N_1091,In_39,In_274);
or U1092 (N_1092,In_332,In_555);
or U1093 (N_1093,In_925,In_820);
nor U1094 (N_1094,In_276,In_555);
and U1095 (N_1095,In_999,In_936);
or U1096 (N_1096,In_518,In_234);
and U1097 (N_1097,In_860,In_883);
and U1098 (N_1098,In_359,In_531);
nand U1099 (N_1099,In_333,In_2);
nor U1100 (N_1100,In_392,In_929);
nor U1101 (N_1101,In_293,In_368);
or U1102 (N_1102,In_989,In_582);
or U1103 (N_1103,In_882,In_11);
and U1104 (N_1104,In_830,In_17);
and U1105 (N_1105,In_97,In_171);
and U1106 (N_1106,In_643,In_779);
or U1107 (N_1107,In_968,In_654);
or U1108 (N_1108,In_261,In_151);
or U1109 (N_1109,In_754,In_724);
or U1110 (N_1110,In_422,In_16);
and U1111 (N_1111,In_788,In_583);
nor U1112 (N_1112,In_585,In_432);
xor U1113 (N_1113,In_661,In_901);
or U1114 (N_1114,In_947,In_545);
nor U1115 (N_1115,In_555,In_604);
nand U1116 (N_1116,In_533,In_900);
or U1117 (N_1117,In_291,In_100);
and U1118 (N_1118,In_625,In_19);
nand U1119 (N_1119,In_938,In_521);
and U1120 (N_1120,In_186,In_98);
and U1121 (N_1121,In_438,In_691);
nor U1122 (N_1122,In_981,In_350);
nand U1123 (N_1123,In_511,In_789);
nor U1124 (N_1124,In_539,In_749);
and U1125 (N_1125,In_610,In_382);
nand U1126 (N_1126,In_893,In_331);
nor U1127 (N_1127,In_426,In_599);
nor U1128 (N_1128,In_598,In_415);
nor U1129 (N_1129,In_755,In_508);
nor U1130 (N_1130,In_286,In_296);
nor U1131 (N_1131,In_109,In_770);
nor U1132 (N_1132,In_895,In_732);
nor U1133 (N_1133,In_549,In_362);
nand U1134 (N_1134,In_22,In_833);
nor U1135 (N_1135,In_730,In_951);
or U1136 (N_1136,In_863,In_50);
and U1137 (N_1137,In_200,In_222);
nor U1138 (N_1138,In_697,In_679);
nand U1139 (N_1139,In_762,In_918);
nand U1140 (N_1140,In_88,In_568);
nand U1141 (N_1141,In_65,In_814);
nor U1142 (N_1142,In_871,In_472);
and U1143 (N_1143,In_921,In_85);
nor U1144 (N_1144,In_705,In_796);
nor U1145 (N_1145,In_13,In_943);
and U1146 (N_1146,In_244,In_873);
and U1147 (N_1147,In_236,In_333);
and U1148 (N_1148,In_20,In_815);
and U1149 (N_1149,In_253,In_150);
or U1150 (N_1150,In_446,In_799);
or U1151 (N_1151,In_996,In_606);
nor U1152 (N_1152,In_783,In_793);
nand U1153 (N_1153,In_770,In_654);
and U1154 (N_1154,In_747,In_913);
or U1155 (N_1155,In_988,In_821);
or U1156 (N_1156,In_807,In_740);
nor U1157 (N_1157,In_614,In_124);
nand U1158 (N_1158,In_200,In_505);
and U1159 (N_1159,In_44,In_511);
or U1160 (N_1160,In_537,In_551);
nor U1161 (N_1161,In_264,In_620);
and U1162 (N_1162,In_669,In_644);
or U1163 (N_1163,In_646,In_629);
nor U1164 (N_1164,In_531,In_820);
and U1165 (N_1165,In_712,In_797);
nor U1166 (N_1166,In_538,In_993);
or U1167 (N_1167,In_56,In_149);
and U1168 (N_1168,In_202,In_268);
nor U1169 (N_1169,In_342,In_118);
or U1170 (N_1170,In_859,In_757);
and U1171 (N_1171,In_683,In_188);
or U1172 (N_1172,In_960,In_878);
xnor U1173 (N_1173,In_903,In_684);
nor U1174 (N_1174,In_273,In_0);
nor U1175 (N_1175,In_975,In_219);
or U1176 (N_1176,In_708,In_537);
or U1177 (N_1177,In_184,In_118);
nor U1178 (N_1178,In_177,In_685);
nor U1179 (N_1179,In_677,In_749);
and U1180 (N_1180,In_270,In_810);
and U1181 (N_1181,In_637,In_117);
and U1182 (N_1182,In_384,In_181);
nand U1183 (N_1183,In_393,In_659);
nor U1184 (N_1184,In_783,In_331);
and U1185 (N_1185,In_214,In_627);
and U1186 (N_1186,In_703,In_498);
nand U1187 (N_1187,In_858,In_327);
nor U1188 (N_1188,In_51,In_774);
and U1189 (N_1189,In_708,In_656);
or U1190 (N_1190,In_682,In_950);
nor U1191 (N_1191,In_149,In_876);
and U1192 (N_1192,In_584,In_152);
or U1193 (N_1193,In_56,In_67);
nand U1194 (N_1194,In_181,In_903);
and U1195 (N_1195,In_449,In_14);
and U1196 (N_1196,In_430,In_826);
and U1197 (N_1197,In_843,In_470);
and U1198 (N_1198,In_109,In_781);
nand U1199 (N_1199,In_824,In_678);
nand U1200 (N_1200,In_317,In_552);
or U1201 (N_1201,In_316,In_954);
or U1202 (N_1202,In_299,In_48);
or U1203 (N_1203,In_434,In_58);
or U1204 (N_1204,In_670,In_451);
nand U1205 (N_1205,In_527,In_2);
nor U1206 (N_1206,In_112,In_504);
nand U1207 (N_1207,In_191,In_902);
and U1208 (N_1208,In_682,In_68);
nor U1209 (N_1209,In_956,In_830);
nor U1210 (N_1210,In_747,In_78);
nand U1211 (N_1211,In_665,In_882);
nor U1212 (N_1212,In_108,In_976);
and U1213 (N_1213,In_258,In_111);
nand U1214 (N_1214,In_319,In_548);
nor U1215 (N_1215,In_17,In_770);
or U1216 (N_1216,In_836,In_639);
or U1217 (N_1217,In_188,In_290);
and U1218 (N_1218,In_230,In_457);
or U1219 (N_1219,In_235,In_958);
nand U1220 (N_1220,In_895,In_547);
xnor U1221 (N_1221,In_477,In_614);
nor U1222 (N_1222,In_615,In_473);
and U1223 (N_1223,In_613,In_214);
nor U1224 (N_1224,In_594,In_340);
nor U1225 (N_1225,In_753,In_493);
nor U1226 (N_1226,In_554,In_336);
nor U1227 (N_1227,In_778,In_908);
or U1228 (N_1228,In_188,In_810);
nand U1229 (N_1229,In_896,In_922);
nand U1230 (N_1230,In_582,In_90);
and U1231 (N_1231,In_531,In_120);
and U1232 (N_1232,In_532,In_214);
nor U1233 (N_1233,In_614,In_432);
or U1234 (N_1234,In_385,In_6);
or U1235 (N_1235,In_608,In_797);
or U1236 (N_1236,In_501,In_98);
or U1237 (N_1237,In_926,In_677);
nand U1238 (N_1238,In_272,In_729);
nor U1239 (N_1239,In_169,In_893);
nor U1240 (N_1240,In_971,In_739);
and U1241 (N_1241,In_362,In_618);
nand U1242 (N_1242,In_680,In_489);
nor U1243 (N_1243,In_895,In_14);
or U1244 (N_1244,In_617,In_698);
nand U1245 (N_1245,In_286,In_465);
nand U1246 (N_1246,In_748,In_159);
xnor U1247 (N_1247,In_430,In_405);
nor U1248 (N_1248,In_81,In_703);
or U1249 (N_1249,In_989,In_396);
or U1250 (N_1250,In_954,In_56);
nand U1251 (N_1251,In_547,In_244);
nor U1252 (N_1252,In_449,In_118);
or U1253 (N_1253,In_334,In_730);
nand U1254 (N_1254,In_423,In_947);
nand U1255 (N_1255,In_506,In_54);
nand U1256 (N_1256,In_786,In_402);
and U1257 (N_1257,In_537,In_457);
or U1258 (N_1258,In_973,In_558);
or U1259 (N_1259,In_817,In_786);
and U1260 (N_1260,In_108,In_689);
nand U1261 (N_1261,In_363,In_369);
nor U1262 (N_1262,In_167,In_947);
nand U1263 (N_1263,In_447,In_16);
or U1264 (N_1264,In_473,In_635);
or U1265 (N_1265,In_397,In_244);
nor U1266 (N_1266,In_450,In_890);
nor U1267 (N_1267,In_682,In_394);
and U1268 (N_1268,In_695,In_800);
nand U1269 (N_1269,In_840,In_28);
nor U1270 (N_1270,In_685,In_938);
nor U1271 (N_1271,In_659,In_792);
or U1272 (N_1272,In_604,In_400);
or U1273 (N_1273,In_694,In_491);
xnor U1274 (N_1274,In_788,In_231);
nor U1275 (N_1275,In_462,In_177);
or U1276 (N_1276,In_710,In_920);
nand U1277 (N_1277,In_746,In_783);
nor U1278 (N_1278,In_291,In_526);
nand U1279 (N_1279,In_328,In_998);
or U1280 (N_1280,In_262,In_621);
nor U1281 (N_1281,In_403,In_570);
or U1282 (N_1282,In_933,In_256);
nand U1283 (N_1283,In_70,In_336);
and U1284 (N_1284,In_739,In_132);
and U1285 (N_1285,In_72,In_679);
or U1286 (N_1286,In_716,In_719);
nand U1287 (N_1287,In_677,In_208);
xor U1288 (N_1288,In_168,In_829);
or U1289 (N_1289,In_810,In_843);
or U1290 (N_1290,In_56,In_193);
and U1291 (N_1291,In_309,In_385);
or U1292 (N_1292,In_505,In_725);
nand U1293 (N_1293,In_140,In_448);
nand U1294 (N_1294,In_670,In_639);
or U1295 (N_1295,In_231,In_158);
nand U1296 (N_1296,In_134,In_87);
nor U1297 (N_1297,In_243,In_816);
nor U1298 (N_1298,In_428,In_53);
and U1299 (N_1299,In_981,In_279);
and U1300 (N_1300,In_51,In_855);
and U1301 (N_1301,In_916,In_415);
nor U1302 (N_1302,In_900,In_73);
nand U1303 (N_1303,In_632,In_636);
and U1304 (N_1304,In_0,In_874);
nand U1305 (N_1305,In_698,In_347);
and U1306 (N_1306,In_912,In_837);
nand U1307 (N_1307,In_825,In_777);
nor U1308 (N_1308,In_922,In_234);
nor U1309 (N_1309,In_682,In_605);
and U1310 (N_1310,In_222,In_268);
and U1311 (N_1311,In_84,In_546);
nor U1312 (N_1312,In_263,In_497);
and U1313 (N_1313,In_883,In_988);
nor U1314 (N_1314,In_750,In_618);
and U1315 (N_1315,In_976,In_715);
xor U1316 (N_1316,In_853,In_781);
and U1317 (N_1317,In_410,In_185);
nor U1318 (N_1318,In_853,In_236);
nand U1319 (N_1319,In_428,In_784);
nand U1320 (N_1320,In_647,In_385);
and U1321 (N_1321,In_45,In_581);
and U1322 (N_1322,In_517,In_848);
nor U1323 (N_1323,In_635,In_833);
or U1324 (N_1324,In_825,In_233);
or U1325 (N_1325,In_598,In_591);
or U1326 (N_1326,In_263,In_797);
nor U1327 (N_1327,In_233,In_632);
or U1328 (N_1328,In_230,In_665);
nor U1329 (N_1329,In_753,In_589);
and U1330 (N_1330,In_794,In_80);
nor U1331 (N_1331,In_696,In_456);
nand U1332 (N_1332,In_983,In_36);
nor U1333 (N_1333,In_237,In_418);
nor U1334 (N_1334,In_64,In_468);
or U1335 (N_1335,In_416,In_290);
and U1336 (N_1336,In_251,In_603);
nor U1337 (N_1337,In_13,In_865);
nor U1338 (N_1338,In_699,In_700);
or U1339 (N_1339,In_361,In_446);
nand U1340 (N_1340,In_276,In_489);
or U1341 (N_1341,In_577,In_661);
nand U1342 (N_1342,In_959,In_581);
nand U1343 (N_1343,In_44,In_891);
nor U1344 (N_1344,In_305,In_153);
or U1345 (N_1345,In_873,In_611);
or U1346 (N_1346,In_862,In_125);
nand U1347 (N_1347,In_296,In_589);
nor U1348 (N_1348,In_160,In_595);
or U1349 (N_1349,In_385,In_79);
or U1350 (N_1350,In_401,In_673);
nand U1351 (N_1351,In_702,In_27);
nor U1352 (N_1352,In_68,In_868);
or U1353 (N_1353,In_222,In_859);
and U1354 (N_1354,In_677,In_299);
nand U1355 (N_1355,In_525,In_539);
or U1356 (N_1356,In_780,In_321);
nor U1357 (N_1357,In_281,In_364);
and U1358 (N_1358,In_323,In_454);
and U1359 (N_1359,In_129,In_151);
nor U1360 (N_1360,In_793,In_100);
or U1361 (N_1361,In_137,In_784);
nand U1362 (N_1362,In_710,In_748);
nand U1363 (N_1363,In_685,In_630);
or U1364 (N_1364,In_876,In_629);
xor U1365 (N_1365,In_236,In_346);
nor U1366 (N_1366,In_540,In_66);
nand U1367 (N_1367,In_630,In_407);
nand U1368 (N_1368,In_47,In_125);
nand U1369 (N_1369,In_254,In_408);
nand U1370 (N_1370,In_947,In_602);
and U1371 (N_1371,In_119,In_292);
nor U1372 (N_1372,In_53,In_729);
and U1373 (N_1373,In_608,In_540);
or U1374 (N_1374,In_638,In_740);
xnor U1375 (N_1375,In_398,In_183);
nor U1376 (N_1376,In_627,In_15);
or U1377 (N_1377,In_494,In_565);
nand U1378 (N_1378,In_907,In_421);
and U1379 (N_1379,In_504,In_815);
and U1380 (N_1380,In_769,In_943);
or U1381 (N_1381,In_951,In_910);
nand U1382 (N_1382,In_402,In_491);
or U1383 (N_1383,In_403,In_781);
nor U1384 (N_1384,In_975,In_349);
and U1385 (N_1385,In_763,In_995);
and U1386 (N_1386,In_453,In_821);
or U1387 (N_1387,In_325,In_80);
or U1388 (N_1388,In_765,In_970);
xnor U1389 (N_1389,In_972,In_491);
nand U1390 (N_1390,In_731,In_837);
nand U1391 (N_1391,In_87,In_753);
or U1392 (N_1392,In_931,In_176);
and U1393 (N_1393,In_869,In_906);
nor U1394 (N_1394,In_773,In_136);
nor U1395 (N_1395,In_39,In_500);
nor U1396 (N_1396,In_419,In_909);
nor U1397 (N_1397,In_621,In_827);
or U1398 (N_1398,In_961,In_926);
xnor U1399 (N_1399,In_495,In_559);
and U1400 (N_1400,In_220,In_93);
nand U1401 (N_1401,In_885,In_535);
nand U1402 (N_1402,In_190,In_685);
and U1403 (N_1403,In_681,In_539);
nor U1404 (N_1404,In_714,In_593);
or U1405 (N_1405,In_568,In_903);
or U1406 (N_1406,In_399,In_916);
xnor U1407 (N_1407,In_815,In_387);
or U1408 (N_1408,In_130,In_861);
or U1409 (N_1409,In_706,In_976);
nand U1410 (N_1410,In_304,In_356);
or U1411 (N_1411,In_956,In_918);
or U1412 (N_1412,In_59,In_592);
xor U1413 (N_1413,In_477,In_528);
nand U1414 (N_1414,In_375,In_286);
and U1415 (N_1415,In_809,In_380);
nor U1416 (N_1416,In_499,In_806);
and U1417 (N_1417,In_518,In_91);
nand U1418 (N_1418,In_515,In_573);
nor U1419 (N_1419,In_720,In_552);
and U1420 (N_1420,In_436,In_870);
nor U1421 (N_1421,In_176,In_91);
or U1422 (N_1422,In_964,In_757);
nand U1423 (N_1423,In_560,In_820);
or U1424 (N_1424,In_778,In_712);
nand U1425 (N_1425,In_581,In_94);
nand U1426 (N_1426,In_255,In_786);
nand U1427 (N_1427,In_32,In_164);
or U1428 (N_1428,In_833,In_320);
nor U1429 (N_1429,In_569,In_43);
nand U1430 (N_1430,In_502,In_854);
and U1431 (N_1431,In_640,In_638);
or U1432 (N_1432,In_729,In_387);
nand U1433 (N_1433,In_147,In_429);
and U1434 (N_1434,In_628,In_754);
or U1435 (N_1435,In_279,In_832);
nor U1436 (N_1436,In_937,In_831);
and U1437 (N_1437,In_885,In_739);
nor U1438 (N_1438,In_262,In_2);
or U1439 (N_1439,In_564,In_93);
nor U1440 (N_1440,In_335,In_76);
or U1441 (N_1441,In_426,In_670);
nand U1442 (N_1442,In_31,In_438);
xnor U1443 (N_1443,In_535,In_367);
nand U1444 (N_1444,In_177,In_179);
nand U1445 (N_1445,In_996,In_230);
or U1446 (N_1446,In_247,In_174);
or U1447 (N_1447,In_14,In_288);
or U1448 (N_1448,In_287,In_263);
and U1449 (N_1449,In_115,In_9);
and U1450 (N_1450,In_845,In_896);
xnor U1451 (N_1451,In_27,In_99);
nand U1452 (N_1452,In_69,In_699);
nor U1453 (N_1453,In_27,In_875);
nor U1454 (N_1454,In_403,In_267);
and U1455 (N_1455,In_361,In_980);
nand U1456 (N_1456,In_448,In_196);
and U1457 (N_1457,In_456,In_375);
or U1458 (N_1458,In_697,In_628);
xor U1459 (N_1459,In_353,In_262);
and U1460 (N_1460,In_714,In_115);
and U1461 (N_1461,In_440,In_182);
nor U1462 (N_1462,In_84,In_987);
or U1463 (N_1463,In_437,In_579);
nand U1464 (N_1464,In_341,In_757);
or U1465 (N_1465,In_771,In_775);
nand U1466 (N_1466,In_386,In_344);
and U1467 (N_1467,In_868,In_313);
nor U1468 (N_1468,In_872,In_342);
and U1469 (N_1469,In_959,In_6);
or U1470 (N_1470,In_929,In_228);
nor U1471 (N_1471,In_50,In_738);
or U1472 (N_1472,In_719,In_456);
and U1473 (N_1473,In_27,In_422);
nand U1474 (N_1474,In_161,In_712);
or U1475 (N_1475,In_676,In_701);
nor U1476 (N_1476,In_781,In_869);
nor U1477 (N_1477,In_19,In_953);
nor U1478 (N_1478,In_161,In_517);
xor U1479 (N_1479,In_462,In_843);
and U1480 (N_1480,In_159,In_381);
nand U1481 (N_1481,In_456,In_578);
or U1482 (N_1482,In_777,In_737);
nand U1483 (N_1483,In_342,In_849);
and U1484 (N_1484,In_432,In_816);
and U1485 (N_1485,In_802,In_855);
and U1486 (N_1486,In_378,In_54);
nor U1487 (N_1487,In_556,In_61);
nor U1488 (N_1488,In_865,In_527);
and U1489 (N_1489,In_805,In_125);
and U1490 (N_1490,In_539,In_240);
nand U1491 (N_1491,In_136,In_636);
nor U1492 (N_1492,In_479,In_265);
xor U1493 (N_1493,In_903,In_623);
or U1494 (N_1494,In_70,In_362);
nand U1495 (N_1495,In_27,In_578);
or U1496 (N_1496,In_288,In_750);
and U1497 (N_1497,In_364,In_579);
and U1498 (N_1498,In_51,In_262);
or U1499 (N_1499,In_908,In_94);
nand U1500 (N_1500,In_54,In_702);
nand U1501 (N_1501,In_141,In_626);
and U1502 (N_1502,In_312,In_206);
xor U1503 (N_1503,In_186,In_767);
or U1504 (N_1504,In_310,In_104);
nand U1505 (N_1505,In_569,In_668);
and U1506 (N_1506,In_826,In_213);
and U1507 (N_1507,In_164,In_626);
and U1508 (N_1508,In_333,In_959);
and U1509 (N_1509,In_9,In_381);
and U1510 (N_1510,In_39,In_671);
nor U1511 (N_1511,In_397,In_508);
nor U1512 (N_1512,In_641,In_517);
or U1513 (N_1513,In_362,In_669);
nor U1514 (N_1514,In_967,In_942);
nor U1515 (N_1515,In_495,In_764);
nor U1516 (N_1516,In_522,In_80);
nand U1517 (N_1517,In_799,In_506);
or U1518 (N_1518,In_812,In_156);
and U1519 (N_1519,In_842,In_998);
nor U1520 (N_1520,In_156,In_2);
nand U1521 (N_1521,In_474,In_983);
nor U1522 (N_1522,In_738,In_876);
or U1523 (N_1523,In_986,In_964);
or U1524 (N_1524,In_749,In_618);
and U1525 (N_1525,In_306,In_500);
and U1526 (N_1526,In_672,In_979);
nand U1527 (N_1527,In_154,In_923);
or U1528 (N_1528,In_191,In_282);
or U1529 (N_1529,In_317,In_226);
xnor U1530 (N_1530,In_666,In_590);
or U1531 (N_1531,In_402,In_211);
and U1532 (N_1532,In_389,In_149);
or U1533 (N_1533,In_986,In_308);
and U1534 (N_1534,In_557,In_577);
or U1535 (N_1535,In_443,In_195);
and U1536 (N_1536,In_431,In_190);
nand U1537 (N_1537,In_385,In_734);
and U1538 (N_1538,In_795,In_895);
nand U1539 (N_1539,In_806,In_966);
or U1540 (N_1540,In_305,In_406);
nand U1541 (N_1541,In_254,In_914);
or U1542 (N_1542,In_601,In_683);
and U1543 (N_1543,In_330,In_831);
or U1544 (N_1544,In_447,In_741);
nand U1545 (N_1545,In_870,In_827);
nand U1546 (N_1546,In_619,In_544);
or U1547 (N_1547,In_973,In_299);
nand U1548 (N_1548,In_640,In_552);
or U1549 (N_1549,In_976,In_594);
nor U1550 (N_1550,In_175,In_480);
and U1551 (N_1551,In_870,In_223);
xor U1552 (N_1552,In_659,In_595);
and U1553 (N_1553,In_330,In_997);
nor U1554 (N_1554,In_292,In_319);
nor U1555 (N_1555,In_284,In_454);
or U1556 (N_1556,In_627,In_174);
or U1557 (N_1557,In_495,In_292);
nor U1558 (N_1558,In_91,In_908);
nor U1559 (N_1559,In_48,In_435);
or U1560 (N_1560,In_762,In_879);
nor U1561 (N_1561,In_55,In_859);
or U1562 (N_1562,In_331,In_30);
nor U1563 (N_1563,In_751,In_48);
and U1564 (N_1564,In_51,In_428);
nor U1565 (N_1565,In_633,In_484);
and U1566 (N_1566,In_338,In_573);
nand U1567 (N_1567,In_483,In_919);
nor U1568 (N_1568,In_14,In_562);
nor U1569 (N_1569,In_735,In_803);
nand U1570 (N_1570,In_748,In_662);
nand U1571 (N_1571,In_50,In_100);
and U1572 (N_1572,In_163,In_272);
nand U1573 (N_1573,In_720,In_120);
nor U1574 (N_1574,In_588,In_949);
and U1575 (N_1575,In_277,In_909);
nor U1576 (N_1576,In_149,In_185);
nand U1577 (N_1577,In_698,In_96);
nor U1578 (N_1578,In_141,In_935);
nor U1579 (N_1579,In_685,In_5);
and U1580 (N_1580,In_364,In_93);
nor U1581 (N_1581,In_979,In_264);
nand U1582 (N_1582,In_829,In_433);
nor U1583 (N_1583,In_231,In_370);
nor U1584 (N_1584,In_511,In_257);
nand U1585 (N_1585,In_202,In_649);
or U1586 (N_1586,In_108,In_433);
and U1587 (N_1587,In_624,In_317);
nand U1588 (N_1588,In_990,In_628);
or U1589 (N_1589,In_955,In_28);
nor U1590 (N_1590,In_646,In_188);
and U1591 (N_1591,In_16,In_569);
nor U1592 (N_1592,In_557,In_834);
nor U1593 (N_1593,In_576,In_647);
nor U1594 (N_1594,In_258,In_64);
and U1595 (N_1595,In_532,In_28);
nand U1596 (N_1596,In_451,In_556);
nor U1597 (N_1597,In_896,In_646);
nor U1598 (N_1598,In_74,In_209);
or U1599 (N_1599,In_878,In_158);
and U1600 (N_1600,In_348,In_780);
nor U1601 (N_1601,In_385,In_207);
or U1602 (N_1602,In_865,In_219);
and U1603 (N_1603,In_743,In_651);
and U1604 (N_1604,In_417,In_278);
nor U1605 (N_1605,In_349,In_615);
and U1606 (N_1606,In_126,In_552);
nand U1607 (N_1607,In_900,In_523);
nor U1608 (N_1608,In_334,In_469);
or U1609 (N_1609,In_749,In_829);
and U1610 (N_1610,In_318,In_129);
nand U1611 (N_1611,In_465,In_73);
or U1612 (N_1612,In_35,In_352);
nand U1613 (N_1613,In_157,In_19);
nor U1614 (N_1614,In_325,In_566);
or U1615 (N_1615,In_359,In_475);
and U1616 (N_1616,In_697,In_605);
nor U1617 (N_1617,In_11,In_742);
nand U1618 (N_1618,In_858,In_990);
nand U1619 (N_1619,In_675,In_527);
and U1620 (N_1620,In_508,In_598);
nor U1621 (N_1621,In_780,In_541);
or U1622 (N_1622,In_717,In_71);
and U1623 (N_1623,In_180,In_521);
or U1624 (N_1624,In_744,In_736);
nand U1625 (N_1625,In_862,In_250);
and U1626 (N_1626,In_241,In_950);
nand U1627 (N_1627,In_858,In_802);
and U1628 (N_1628,In_408,In_537);
nor U1629 (N_1629,In_408,In_354);
and U1630 (N_1630,In_678,In_464);
or U1631 (N_1631,In_323,In_594);
and U1632 (N_1632,In_795,In_508);
and U1633 (N_1633,In_505,In_52);
or U1634 (N_1634,In_37,In_340);
xor U1635 (N_1635,In_183,In_652);
nand U1636 (N_1636,In_418,In_400);
or U1637 (N_1637,In_479,In_543);
or U1638 (N_1638,In_833,In_928);
or U1639 (N_1639,In_1,In_761);
xnor U1640 (N_1640,In_139,In_275);
nor U1641 (N_1641,In_621,In_293);
and U1642 (N_1642,In_681,In_691);
or U1643 (N_1643,In_696,In_164);
or U1644 (N_1644,In_433,In_617);
or U1645 (N_1645,In_771,In_577);
nand U1646 (N_1646,In_877,In_336);
or U1647 (N_1647,In_971,In_540);
and U1648 (N_1648,In_399,In_715);
or U1649 (N_1649,In_610,In_968);
nand U1650 (N_1650,In_718,In_380);
nor U1651 (N_1651,In_888,In_818);
nand U1652 (N_1652,In_486,In_662);
nor U1653 (N_1653,In_909,In_561);
nor U1654 (N_1654,In_469,In_635);
nand U1655 (N_1655,In_532,In_622);
or U1656 (N_1656,In_909,In_522);
and U1657 (N_1657,In_846,In_131);
and U1658 (N_1658,In_616,In_481);
nand U1659 (N_1659,In_771,In_207);
and U1660 (N_1660,In_162,In_826);
and U1661 (N_1661,In_246,In_872);
and U1662 (N_1662,In_630,In_581);
nand U1663 (N_1663,In_674,In_596);
and U1664 (N_1664,In_155,In_845);
or U1665 (N_1665,In_427,In_69);
and U1666 (N_1666,In_983,In_936);
or U1667 (N_1667,In_804,In_306);
and U1668 (N_1668,In_85,In_131);
nand U1669 (N_1669,In_836,In_257);
nor U1670 (N_1670,In_86,In_651);
nand U1671 (N_1671,In_825,In_796);
or U1672 (N_1672,In_788,In_635);
nand U1673 (N_1673,In_897,In_257);
nand U1674 (N_1674,In_341,In_160);
and U1675 (N_1675,In_984,In_20);
and U1676 (N_1676,In_906,In_497);
or U1677 (N_1677,In_989,In_728);
or U1678 (N_1678,In_519,In_769);
or U1679 (N_1679,In_944,In_209);
nand U1680 (N_1680,In_808,In_439);
or U1681 (N_1681,In_680,In_702);
nand U1682 (N_1682,In_436,In_116);
nor U1683 (N_1683,In_953,In_341);
or U1684 (N_1684,In_546,In_481);
or U1685 (N_1685,In_89,In_258);
and U1686 (N_1686,In_895,In_611);
or U1687 (N_1687,In_268,In_153);
nor U1688 (N_1688,In_976,In_457);
or U1689 (N_1689,In_590,In_801);
nand U1690 (N_1690,In_471,In_576);
nand U1691 (N_1691,In_510,In_884);
and U1692 (N_1692,In_930,In_20);
nor U1693 (N_1693,In_324,In_330);
or U1694 (N_1694,In_242,In_794);
and U1695 (N_1695,In_410,In_228);
and U1696 (N_1696,In_155,In_199);
or U1697 (N_1697,In_998,In_9);
nand U1698 (N_1698,In_227,In_327);
nor U1699 (N_1699,In_504,In_801);
and U1700 (N_1700,In_949,In_167);
and U1701 (N_1701,In_783,In_385);
xnor U1702 (N_1702,In_1,In_706);
nand U1703 (N_1703,In_76,In_657);
nor U1704 (N_1704,In_594,In_467);
nand U1705 (N_1705,In_654,In_442);
and U1706 (N_1706,In_207,In_327);
nand U1707 (N_1707,In_679,In_859);
nor U1708 (N_1708,In_190,In_146);
or U1709 (N_1709,In_245,In_424);
nand U1710 (N_1710,In_417,In_281);
nand U1711 (N_1711,In_453,In_773);
nand U1712 (N_1712,In_791,In_164);
xnor U1713 (N_1713,In_559,In_119);
nor U1714 (N_1714,In_213,In_198);
and U1715 (N_1715,In_769,In_348);
nand U1716 (N_1716,In_340,In_10);
or U1717 (N_1717,In_877,In_420);
nor U1718 (N_1718,In_929,In_796);
or U1719 (N_1719,In_280,In_79);
xnor U1720 (N_1720,In_587,In_294);
or U1721 (N_1721,In_390,In_582);
nand U1722 (N_1722,In_493,In_214);
or U1723 (N_1723,In_456,In_177);
nor U1724 (N_1724,In_990,In_293);
nand U1725 (N_1725,In_349,In_272);
and U1726 (N_1726,In_785,In_677);
and U1727 (N_1727,In_686,In_131);
and U1728 (N_1728,In_738,In_780);
or U1729 (N_1729,In_114,In_761);
nor U1730 (N_1730,In_828,In_380);
and U1731 (N_1731,In_653,In_887);
and U1732 (N_1732,In_466,In_998);
nand U1733 (N_1733,In_168,In_676);
nand U1734 (N_1734,In_314,In_144);
nand U1735 (N_1735,In_665,In_897);
or U1736 (N_1736,In_333,In_590);
or U1737 (N_1737,In_716,In_803);
nor U1738 (N_1738,In_339,In_807);
and U1739 (N_1739,In_392,In_52);
or U1740 (N_1740,In_806,In_929);
or U1741 (N_1741,In_810,In_288);
or U1742 (N_1742,In_384,In_545);
nand U1743 (N_1743,In_442,In_950);
or U1744 (N_1744,In_950,In_250);
or U1745 (N_1745,In_335,In_893);
nor U1746 (N_1746,In_555,In_799);
nor U1747 (N_1747,In_128,In_16);
and U1748 (N_1748,In_852,In_735);
nand U1749 (N_1749,In_646,In_571);
nand U1750 (N_1750,In_516,In_737);
nor U1751 (N_1751,In_895,In_568);
nand U1752 (N_1752,In_266,In_265);
and U1753 (N_1753,In_986,In_894);
or U1754 (N_1754,In_395,In_774);
or U1755 (N_1755,In_661,In_62);
nand U1756 (N_1756,In_130,In_647);
and U1757 (N_1757,In_643,In_434);
and U1758 (N_1758,In_422,In_766);
nand U1759 (N_1759,In_61,In_214);
or U1760 (N_1760,In_216,In_288);
or U1761 (N_1761,In_731,In_821);
nand U1762 (N_1762,In_460,In_213);
xor U1763 (N_1763,In_985,In_202);
or U1764 (N_1764,In_253,In_455);
nand U1765 (N_1765,In_946,In_869);
xnor U1766 (N_1766,In_1,In_727);
and U1767 (N_1767,In_420,In_777);
xnor U1768 (N_1768,In_812,In_246);
nand U1769 (N_1769,In_517,In_580);
and U1770 (N_1770,In_266,In_915);
and U1771 (N_1771,In_571,In_169);
or U1772 (N_1772,In_490,In_378);
or U1773 (N_1773,In_270,In_146);
and U1774 (N_1774,In_489,In_159);
nor U1775 (N_1775,In_883,In_196);
and U1776 (N_1776,In_147,In_735);
nor U1777 (N_1777,In_824,In_421);
and U1778 (N_1778,In_708,In_457);
and U1779 (N_1779,In_280,In_243);
or U1780 (N_1780,In_151,In_969);
nor U1781 (N_1781,In_353,In_835);
nor U1782 (N_1782,In_666,In_300);
xnor U1783 (N_1783,In_770,In_810);
nor U1784 (N_1784,In_940,In_188);
nand U1785 (N_1785,In_93,In_851);
and U1786 (N_1786,In_469,In_502);
or U1787 (N_1787,In_660,In_673);
nor U1788 (N_1788,In_23,In_628);
xnor U1789 (N_1789,In_115,In_930);
or U1790 (N_1790,In_348,In_928);
or U1791 (N_1791,In_517,In_888);
and U1792 (N_1792,In_214,In_57);
nor U1793 (N_1793,In_423,In_982);
or U1794 (N_1794,In_42,In_577);
nor U1795 (N_1795,In_725,In_283);
xnor U1796 (N_1796,In_212,In_763);
nor U1797 (N_1797,In_966,In_743);
xor U1798 (N_1798,In_810,In_925);
nand U1799 (N_1799,In_718,In_673);
or U1800 (N_1800,In_372,In_26);
nor U1801 (N_1801,In_729,In_4);
and U1802 (N_1802,In_77,In_510);
or U1803 (N_1803,In_371,In_750);
nand U1804 (N_1804,In_649,In_917);
or U1805 (N_1805,In_910,In_506);
and U1806 (N_1806,In_594,In_555);
or U1807 (N_1807,In_29,In_417);
and U1808 (N_1808,In_975,In_507);
nand U1809 (N_1809,In_317,In_858);
or U1810 (N_1810,In_858,In_881);
nor U1811 (N_1811,In_108,In_610);
nor U1812 (N_1812,In_110,In_566);
or U1813 (N_1813,In_723,In_476);
nor U1814 (N_1814,In_191,In_970);
or U1815 (N_1815,In_572,In_595);
or U1816 (N_1816,In_533,In_342);
nor U1817 (N_1817,In_211,In_873);
nor U1818 (N_1818,In_966,In_672);
and U1819 (N_1819,In_383,In_254);
nand U1820 (N_1820,In_322,In_978);
nor U1821 (N_1821,In_168,In_305);
xnor U1822 (N_1822,In_74,In_539);
xnor U1823 (N_1823,In_327,In_95);
or U1824 (N_1824,In_58,In_833);
or U1825 (N_1825,In_452,In_420);
or U1826 (N_1826,In_820,In_449);
or U1827 (N_1827,In_361,In_411);
or U1828 (N_1828,In_490,In_718);
and U1829 (N_1829,In_964,In_7);
and U1830 (N_1830,In_42,In_803);
and U1831 (N_1831,In_314,In_143);
nand U1832 (N_1832,In_585,In_87);
or U1833 (N_1833,In_728,In_923);
nor U1834 (N_1834,In_117,In_700);
and U1835 (N_1835,In_578,In_732);
or U1836 (N_1836,In_592,In_99);
nor U1837 (N_1837,In_617,In_527);
nand U1838 (N_1838,In_680,In_531);
and U1839 (N_1839,In_60,In_519);
and U1840 (N_1840,In_582,In_708);
nor U1841 (N_1841,In_551,In_827);
or U1842 (N_1842,In_342,In_130);
or U1843 (N_1843,In_983,In_240);
nor U1844 (N_1844,In_879,In_426);
or U1845 (N_1845,In_996,In_660);
nand U1846 (N_1846,In_763,In_225);
and U1847 (N_1847,In_483,In_684);
nand U1848 (N_1848,In_203,In_136);
nor U1849 (N_1849,In_920,In_402);
and U1850 (N_1850,In_233,In_19);
or U1851 (N_1851,In_980,In_522);
or U1852 (N_1852,In_31,In_550);
or U1853 (N_1853,In_348,In_379);
nand U1854 (N_1854,In_805,In_83);
or U1855 (N_1855,In_626,In_796);
or U1856 (N_1856,In_645,In_230);
nor U1857 (N_1857,In_94,In_441);
and U1858 (N_1858,In_365,In_676);
and U1859 (N_1859,In_340,In_67);
and U1860 (N_1860,In_519,In_174);
nor U1861 (N_1861,In_11,In_504);
and U1862 (N_1862,In_781,In_183);
or U1863 (N_1863,In_478,In_821);
xnor U1864 (N_1864,In_539,In_926);
and U1865 (N_1865,In_579,In_662);
and U1866 (N_1866,In_582,In_670);
nand U1867 (N_1867,In_778,In_78);
or U1868 (N_1868,In_17,In_61);
and U1869 (N_1869,In_977,In_371);
and U1870 (N_1870,In_802,In_715);
nor U1871 (N_1871,In_588,In_430);
nor U1872 (N_1872,In_369,In_377);
nor U1873 (N_1873,In_53,In_68);
and U1874 (N_1874,In_490,In_469);
or U1875 (N_1875,In_102,In_138);
or U1876 (N_1876,In_876,In_81);
and U1877 (N_1877,In_739,In_337);
nor U1878 (N_1878,In_859,In_855);
nand U1879 (N_1879,In_868,In_259);
and U1880 (N_1880,In_28,In_176);
nand U1881 (N_1881,In_691,In_849);
nor U1882 (N_1882,In_297,In_142);
nor U1883 (N_1883,In_993,In_730);
and U1884 (N_1884,In_678,In_102);
nor U1885 (N_1885,In_985,In_414);
nor U1886 (N_1886,In_999,In_453);
and U1887 (N_1887,In_961,In_577);
nor U1888 (N_1888,In_785,In_124);
nor U1889 (N_1889,In_910,In_463);
nor U1890 (N_1890,In_14,In_232);
xnor U1891 (N_1891,In_261,In_48);
nand U1892 (N_1892,In_63,In_576);
or U1893 (N_1893,In_244,In_551);
or U1894 (N_1894,In_433,In_485);
or U1895 (N_1895,In_251,In_128);
or U1896 (N_1896,In_574,In_134);
nand U1897 (N_1897,In_228,In_432);
nand U1898 (N_1898,In_923,In_352);
and U1899 (N_1899,In_66,In_287);
nor U1900 (N_1900,In_943,In_65);
and U1901 (N_1901,In_717,In_729);
and U1902 (N_1902,In_923,In_975);
nand U1903 (N_1903,In_974,In_221);
and U1904 (N_1904,In_357,In_200);
and U1905 (N_1905,In_539,In_191);
nand U1906 (N_1906,In_532,In_80);
and U1907 (N_1907,In_290,In_621);
nor U1908 (N_1908,In_897,In_179);
xnor U1909 (N_1909,In_727,In_692);
nor U1910 (N_1910,In_907,In_865);
or U1911 (N_1911,In_705,In_471);
nor U1912 (N_1912,In_694,In_940);
nor U1913 (N_1913,In_95,In_968);
or U1914 (N_1914,In_632,In_918);
nand U1915 (N_1915,In_622,In_271);
nor U1916 (N_1916,In_793,In_447);
or U1917 (N_1917,In_579,In_167);
and U1918 (N_1918,In_741,In_72);
nand U1919 (N_1919,In_794,In_962);
nor U1920 (N_1920,In_131,In_144);
nor U1921 (N_1921,In_275,In_94);
or U1922 (N_1922,In_691,In_997);
and U1923 (N_1923,In_986,In_833);
or U1924 (N_1924,In_550,In_311);
nor U1925 (N_1925,In_712,In_168);
and U1926 (N_1926,In_827,In_181);
nand U1927 (N_1927,In_149,In_23);
nand U1928 (N_1928,In_220,In_201);
nand U1929 (N_1929,In_86,In_330);
or U1930 (N_1930,In_592,In_237);
nand U1931 (N_1931,In_70,In_6);
and U1932 (N_1932,In_287,In_780);
or U1933 (N_1933,In_420,In_947);
and U1934 (N_1934,In_82,In_189);
or U1935 (N_1935,In_104,In_124);
or U1936 (N_1936,In_382,In_689);
and U1937 (N_1937,In_45,In_750);
nand U1938 (N_1938,In_996,In_37);
and U1939 (N_1939,In_156,In_844);
xor U1940 (N_1940,In_678,In_496);
nand U1941 (N_1941,In_870,In_938);
or U1942 (N_1942,In_762,In_458);
and U1943 (N_1943,In_486,In_209);
nor U1944 (N_1944,In_555,In_652);
or U1945 (N_1945,In_982,In_516);
nand U1946 (N_1946,In_242,In_145);
and U1947 (N_1947,In_757,In_304);
or U1948 (N_1948,In_312,In_592);
nor U1949 (N_1949,In_593,In_982);
and U1950 (N_1950,In_874,In_604);
nor U1951 (N_1951,In_637,In_245);
or U1952 (N_1952,In_75,In_802);
nand U1953 (N_1953,In_260,In_612);
or U1954 (N_1954,In_719,In_264);
xnor U1955 (N_1955,In_596,In_390);
or U1956 (N_1956,In_703,In_220);
nor U1957 (N_1957,In_567,In_955);
and U1958 (N_1958,In_569,In_223);
nor U1959 (N_1959,In_172,In_800);
or U1960 (N_1960,In_788,In_412);
nand U1961 (N_1961,In_824,In_212);
and U1962 (N_1962,In_943,In_178);
nand U1963 (N_1963,In_130,In_959);
or U1964 (N_1964,In_465,In_202);
and U1965 (N_1965,In_312,In_129);
or U1966 (N_1966,In_204,In_290);
or U1967 (N_1967,In_114,In_421);
or U1968 (N_1968,In_915,In_164);
nor U1969 (N_1969,In_66,In_462);
or U1970 (N_1970,In_891,In_522);
nand U1971 (N_1971,In_402,In_858);
and U1972 (N_1972,In_979,In_483);
or U1973 (N_1973,In_817,In_114);
nand U1974 (N_1974,In_52,In_804);
or U1975 (N_1975,In_421,In_323);
or U1976 (N_1976,In_716,In_834);
or U1977 (N_1977,In_943,In_341);
and U1978 (N_1978,In_910,In_66);
and U1979 (N_1979,In_302,In_818);
nor U1980 (N_1980,In_305,In_946);
and U1981 (N_1981,In_597,In_598);
and U1982 (N_1982,In_672,In_201);
xnor U1983 (N_1983,In_512,In_316);
nor U1984 (N_1984,In_809,In_935);
nand U1985 (N_1985,In_128,In_847);
and U1986 (N_1986,In_284,In_533);
or U1987 (N_1987,In_872,In_47);
nor U1988 (N_1988,In_879,In_575);
nand U1989 (N_1989,In_104,In_416);
nand U1990 (N_1990,In_577,In_844);
and U1991 (N_1991,In_432,In_118);
and U1992 (N_1992,In_969,In_857);
and U1993 (N_1993,In_839,In_828);
and U1994 (N_1994,In_146,In_271);
nor U1995 (N_1995,In_261,In_186);
nand U1996 (N_1996,In_776,In_169);
nand U1997 (N_1997,In_103,In_530);
nor U1998 (N_1998,In_842,In_118);
nor U1999 (N_1999,In_404,In_540);
nor U2000 (N_2000,In_486,In_184);
nand U2001 (N_2001,In_691,In_830);
nand U2002 (N_2002,In_439,In_588);
and U2003 (N_2003,In_271,In_314);
nand U2004 (N_2004,In_603,In_336);
and U2005 (N_2005,In_481,In_426);
or U2006 (N_2006,In_583,In_575);
or U2007 (N_2007,In_610,In_420);
or U2008 (N_2008,In_597,In_239);
nor U2009 (N_2009,In_495,In_948);
nor U2010 (N_2010,In_624,In_241);
nor U2011 (N_2011,In_306,In_643);
or U2012 (N_2012,In_409,In_444);
or U2013 (N_2013,In_807,In_224);
and U2014 (N_2014,In_659,In_797);
nand U2015 (N_2015,In_321,In_390);
nor U2016 (N_2016,In_479,In_355);
nand U2017 (N_2017,In_707,In_338);
nand U2018 (N_2018,In_894,In_627);
nand U2019 (N_2019,In_862,In_346);
nor U2020 (N_2020,In_844,In_381);
and U2021 (N_2021,In_458,In_184);
or U2022 (N_2022,In_965,In_98);
nand U2023 (N_2023,In_676,In_698);
nor U2024 (N_2024,In_411,In_251);
nand U2025 (N_2025,In_3,In_544);
and U2026 (N_2026,In_352,In_680);
nor U2027 (N_2027,In_873,In_944);
nand U2028 (N_2028,In_83,In_188);
or U2029 (N_2029,In_761,In_983);
nand U2030 (N_2030,In_664,In_153);
or U2031 (N_2031,In_53,In_574);
nand U2032 (N_2032,In_425,In_840);
and U2033 (N_2033,In_54,In_726);
and U2034 (N_2034,In_480,In_123);
nor U2035 (N_2035,In_700,In_915);
nand U2036 (N_2036,In_104,In_509);
nor U2037 (N_2037,In_615,In_278);
nand U2038 (N_2038,In_75,In_196);
nand U2039 (N_2039,In_117,In_769);
and U2040 (N_2040,In_738,In_950);
nor U2041 (N_2041,In_184,In_589);
and U2042 (N_2042,In_805,In_243);
and U2043 (N_2043,In_620,In_596);
nor U2044 (N_2044,In_67,In_987);
nand U2045 (N_2045,In_731,In_931);
nor U2046 (N_2046,In_667,In_334);
nand U2047 (N_2047,In_702,In_624);
nand U2048 (N_2048,In_772,In_63);
and U2049 (N_2049,In_790,In_203);
and U2050 (N_2050,In_681,In_474);
nand U2051 (N_2051,In_478,In_570);
nor U2052 (N_2052,In_966,In_698);
nor U2053 (N_2053,In_25,In_809);
or U2054 (N_2054,In_768,In_737);
or U2055 (N_2055,In_744,In_262);
and U2056 (N_2056,In_436,In_119);
and U2057 (N_2057,In_657,In_731);
or U2058 (N_2058,In_128,In_12);
nand U2059 (N_2059,In_903,In_552);
and U2060 (N_2060,In_442,In_521);
nand U2061 (N_2061,In_351,In_909);
and U2062 (N_2062,In_509,In_279);
nand U2063 (N_2063,In_727,In_7);
and U2064 (N_2064,In_433,In_270);
or U2065 (N_2065,In_104,In_953);
nand U2066 (N_2066,In_465,In_64);
nor U2067 (N_2067,In_283,In_303);
or U2068 (N_2068,In_870,In_898);
nor U2069 (N_2069,In_163,In_739);
and U2070 (N_2070,In_921,In_168);
nand U2071 (N_2071,In_326,In_377);
or U2072 (N_2072,In_94,In_705);
nor U2073 (N_2073,In_883,In_90);
and U2074 (N_2074,In_746,In_807);
nor U2075 (N_2075,In_761,In_987);
or U2076 (N_2076,In_890,In_79);
nor U2077 (N_2077,In_668,In_69);
nor U2078 (N_2078,In_967,In_524);
and U2079 (N_2079,In_430,In_524);
nand U2080 (N_2080,In_703,In_778);
and U2081 (N_2081,In_513,In_217);
xnor U2082 (N_2082,In_269,In_173);
nor U2083 (N_2083,In_256,In_238);
nand U2084 (N_2084,In_672,In_814);
and U2085 (N_2085,In_205,In_120);
and U2086 (N_2086,In_434,In_77);
nand U2087 (N_2087,In_575,In_916);
or U2088 (N_2088,In_75,In_870);
nor U2089 (N_2089,In_740,In_829);
or U2090 (N_2090,In_572,In_990);
nor U2091 (N_2091,In_731,In_998);
nand U2092 (N_2092,In_908,In_267);
nand U2093 (N_2093,In_797,In_592);
and U2094 (N_2094,In_655,In_989);
and U2095 (N_2095,In_568,In_779);
or U2096 (N_2096,In_220,In_895);
or U2097 (N_2097,In_134,In_778);
nand U2098 (N_2098,In_199,In_993);
nor U2099 (N_2099,In_833,In_590);
or U2100 (N_2100,In_492,In_251);
nand U2101 (N_2101,In_528,In_620);
nand U2102 (N_2102,In_455,In_956);
and U2103 (N_2103,In_161,In_29);
nor U2104 (N_2104,In_437,In_644);
nand U2105 (N_2105,In_279,In_864);
nand U2106 (N_2106,In_20,In_516);
nand U2107 (N_2107,In_382,In_173);
and U2108 (N_2108,In_130,In_215);
or U2109 (N_2109,In_854,In_362);
and U2110 (N_2110,In_967,In_595);
nand U2111 (N_2111,In_198,In_94);
nand U2112 (N_2112,In_88,In_746);
nor U2113 (N_2113,In_842,In_812);
and U2114 (N_2114,In_526,In_566);
nor U2115 (N_2115,In_956,In_552);
nor U2116 (N_2116,In_217,In_972);
nor U2117 (N_2117,In_735,In_349);
and U2118 (N_2118,In_484,In_727);
or U2119 (N_2119,In_309,In_679);
nand U2120 (N_2120,In_442,In_360);
and U2121 (N_2121,In_315,In_307);
and U2122 (N_2122,In_224,In_965);
nor U2123 (N_2123,In_741,In_317);
nand U2124 (N_2124,In_472,In_338);
or U2125 (N_2125,In_142,In_412);
nor U2126 (N_2126,In_103,In_4);
nor U2127 (N_2127,In_370,In_537);
nor U2128 (N_2128,In_374,In_735);
and U2129 (N_2129,In_969,In_765);
or U2130 (N_2130,In_473,In_388);
nor U2131 (N_2131,In_827,In_373);
nor U2132 (N_2132,In_260,In_45);
nand U2133 (N_2133,In_139,In_872);
and U2134 (N_2134,In_374,In_584);
or U2135 (N_2135,In_698,In_400);
nand U2136 (N_2136,In_338,In_29);
nor U2137 (N_2137,In_752,In_788);
and U2138 (N_2138,In_156,In_584);
nand U2139 (N_2139,In_666,In_583);
or U2140 (N_2140,In_200,In_176);
or U2141 (N_2141,In_209,In_612);
or U2142 (N_2142,In_292,In_793);
or U2143 (N_2143,In_178,In_999);
and U2144 (N_2144,In_831,In_37);
or U2145 (N_2145,In_973,In_273);
nand U2146 (N_2146,In_71,In_634);
nor U2147 (N_2147,In_906,In_97);
and U2148 (N_2148,In_19,In_614);
or U2149 (N_2149,In_729,In_69);
nor U2150 (N_2150,In_900,In_833);
xor U2151 (N_2151,In_241,In_566);
nor U2152 (N_2152,In_530,In_821);
nand U2153 (N_2153,In_655,In_104);
and U2154 (N_2154,In_783,In_382);
and U2155 (N_2155,In_754,In_399);
nand U2156 (N_2156,In_509,In_725);
nor U2157 (N_2157,In_216,In_750);
nand U2158 (N_2158,In_656,In_794);
nor U2159 (N_2159,In_376,In_267);
nand U2160 (N_2160,In_177,In_444);
nand U2161 (N_2161,In_454,In_596);
and U2162 (N_2162,In_328,In_989);
and U2163 (N_2163,In_936,In_845);
or U2164 (N_2164,In_637,In_977);
nor U2165 (N_2165,In_378,In_2);
and U2166 (N_2166,In_86,In_681);
nand U2167 (N_2167,In_448,In_271);
and U2168 (N_2168,In_473,In_586);
and U2169 (N_2169,In_441,In_623);
and U2170 (N_2170,In_876,In_192);
nand U2171 (N_2171,In_790,In_29);
nand U2172 (N_2172,In_389,In_820);
or U2173 (N_2173,In_484,In_270);
or U2174 (N_2174,In_51,In_879);
nand U2175 (N_2175,In_150,In_583);
nand U2176 (N_2176,In_830,In_877);
nand U2177 (N_2177,In_305,In_335);
xnor U2178 (N_2178,In_586,In_903);
nor U2179 (N_2179,In_252,In_525);
nor U2180 (N_2180,In_853,In_958);
or U2181 (N_2181,In_207,In_519);
or U2182 (N_2182,In_645,In_132);
or U2183 (N_2183,In_605,In_17);
nor U2184 (N_2184,In_407,In_993);
nand U2185 (N_2185,In_737,In_764);
or U2186 (N_2186,In_231,In_881);
and U2187 (N_2187,In_794,In_145);
and U2188 (N_2188,In_432,In_375);
nand U2189 (N_2189,In_89,In_122);
nor U2190 (N_2190,In_734,In_27);
or U2191 (N_2191,In_140,In_144);
or U2192 (N_2192,In_12,In_564);
and U2193 (N_2193,In_451,In_469);
nand U2194 (N_2194,In_942,In_676);
nand U2195 (N_2195,In_50,In_699);
nor U2196 (N_2196,In_301,In_331);
or U2197 (N_2197,In_879,In_82);
nor U2198 (N_2198,In_830,In_709);
and U2199 (N_2199,In_728,In_401);
and U2200 (N_2200,In_438,In_849);
or U2201 (N_2201,In_634,In_842);
or U2202 (N_2202,In_706,In_470);
nor U2203 (N_2203,In_738,In_180);
and U2204 (N_2204,In_184,In_740);
or U2205 (N_2205,In_495,In_570);
nand U2206 (N_2206,In_694,In_221);
and U2207 (N_2207,In_589,In_367);
or U2208 (N_2208,In_696,In_193);
and U2209 (N_2209,In_999,In_935);
nand U2210 (N_2210,In_856,In_353);
nand U2211 (N_2211,In_259,In_427);
nor U2212 (N_2212,In_199,In_590);
or U2213 (N_2213,In_177,In_90);
nor U2214 (N_2214,In_399,In_126);
nand U2215 (N_2215,In_532,In_265);
nor U2216 (N_2216,In_332,In_546);
nand U2217 (N_2217,In_593,In_533);
nor U2218 (N_2218,In_934,In_347);
nand U2219 (N_2219,In_77,In_225);
and U2220 (N_2220,In_793,In_24);
nand U2221 (N_2221,In_590,In_491);
nand U2222 (N_2222,In_333,In_301);
nor U2223 (N_2223,In_129,In_805);
and U2224 (N_2224,In_128,In_724);
nand U2225 (N_2225,In_462,In_376);
or U2226 (N_2226,In_812,In_882);
nor U2227 (N_2227,In_881,In_295);
or U2228 (N_2228,In_834,In_843);
or U2229 (N_2229,In_847,In_428);
nand U2230 (N_2230,In_301,In_869);
and U2231 (N_2231,In_57,In_201);
and U2232 (N_2232,In_329,In_524);
and U2233 (N_2233,In_386,In_447);
nand U2234 (N_2234,In_412,In_423);
nand U2235 (N_2235,In_827,In_274);
nand U2236 (N_2236,In_310,In_502);
or U2237 (N_2237,In_530,In_792);
nor U2238 (N_2238,In_304,In_684);
and U2239 (N_2239,In_898,In_959);
nand U2240 (N_2240,In_779,In_337);
or U2241 (N_2241,In_62,In_751);
nor U2242 (N_2242,In_67,In_320);
nand U2243 (N_2243,In_728,In_128);
and U2244 (N_2244,In_251,In_352);
and U2245 (N_2245,In_10,In_33);
or U2246 (N_2246,In_725,In_68);
nand U2247 (N_2247,In_1,In_999);
or U2248 (N_2248,In_532,In_852);
nand U2249 (N_2249,In_281,In_89);
nand U2250 (N_2250,In_656,In_786);
and U2251 (N_2251,In_118,In_318);
or U2252 (N_2252,In_380,In_206);
and U2253 (N_2253,In_246,In_718);
and U2254 (N_2254,In_63,In_112);
nand U2255 (N_2255,In_413,In_93);
nor U2256 (N_2256,In_590,In_683);
nand U2257 (N_2257,In_766,In_615);
and U2258 (N_2258,In_739,In_858);
and U2259 (N_2259,In_919,In_42);
nor U2260 (N_2260,In_423,In_69);
and U2261 (N_2261,In_98,In_380);
nand U2262 (N_2262,In_651,In_533);
nor U2263 (N_2263,In_162,In_702);
nor U2264 (N_2264,In_763,In_848);
or U2265 (N_2265,In_703,In_796);
and U2266 (N_2266,In_489,In_690);
and U2267 (N_2267,In_490,In_493);
and U2268 (N_2268,In_55,In_669);
or U2269 (N_2269,In_897,In_554);
and U2270 (N_2270,In_825,In_498);
or U2271 (N_2271,In_786,In_639);
or U2272 (N_2272,In_176,In_690);
nand U2273 (N_2273,In_45,In_800);
and U2274 (N_2274,In_299,In_920);
nor U2275 (N_2275,In_788,In_792);
nand U2276 (N_2276,In_712,In_780);
and U2277 (N_2277,In_356,In_342);
or U2278 (N_2278,In_489,In_976);
nor U2279 (N_2279,In_664,In_238);
nor U2280 (N_2280,In_500,In_999);
or U2281 (N_2281,In_794,In_770);
and U2282 (N_2282,In_954,In_154);
and U2283 (N_2283,In_93,In_223);
or U2284 (N_2284,In_205,In_382);
and U2285 (N_2285,In_134,In_946);
nor U2286 (N_2286,In_200,In_558);
nand U2287 (N_2287,In_115,In_408);
nor U2288 (N_2288,In_261,In_481);
nor U2289 (N_2289,In_720,In_650);
nand U2290 (N_2290,In_252,In_993);
nor U2291 (N_2291,In_419,In_127);
and U2292 (N_2292,In_277,In_340);
or U2293 (N_2293,In_95,In_714);
or U2294 (N_2294,In_138,In_310);
nand U2295 (N_2295,In_249,In_217);
or U2296 (N_2296,In_132,In_830);
or U2297 (N_2297,In_901,In_670);
and U2298 (N_2298,In_488,In_580);
or U2299 (N_2299,In_912,In_409);
and U2300 (N_2300,In_861,In_403);
and U2301 (N_2301,In_743,In_868);
nand U2302 (N_2302,In_785,In_650);
xnor U2303 (N_2303,In_428,In_608);
or U2304 (N_2304,In_177,In_562);
or U2305 (N_2305,In_891,In_719);
nand U2306 (N_2306,In_395,In_883);
nor U2307 (N_2307,In_333,In_84);
nand U2308 (N_2308,In_702,In_852);
nand U2309 (N_2309,In_98,In_175);
and U2310 (N_2310,In_226,In_441);
xor U2311 (N_2311,In_29,In_691);
or U2312 (N_2312,In_523,In_875);
nand U2313 (N_2313,In_670,In_53);
nor U2314 (N_2314,In_493,In_416);
nand U2315 (N_2315,In_979,In_537);
nor U2316 (N_2316,In_934,In_316);
nand U2317 (N_2317,In_325,In_979);
xor U2318 (N_2318,In_858,In_517);
or U2319 (N_2319,In_869,In_674);
nand U2320 (N_2320,In_152,In_385);
or U2321 (N_2321,In_501,In_273);
and U2322 (N_2322,In_50,In_560);
or U2323 (N_2323,In_280,In_356);
xor U2324 (N_2324,In_552,In_245);
or U2325 (N_2325,In_631,In_397);
xor U2326 (N_2326,In_69,In_631);
or U2327 (N_2327,In_354,In_889);
nor U2328 (N_2328,In_491,In_29);
nor U2329 (N_2329,In_16,In_808);
or U2330 (N_2330,In_647,In_333);
nor U2331 (N_2331,In_508,In_175);
nand U2332 (N_2332,In_541,In_274);
or U2333 (N_2333,In_775,In_220);
nand U2334 (N_2334,In_648,In_295);
nand U2335 (N_2335,In_859,In_114);
and U2336 (N_2336,In_942,In_291);
and U2337 (N_2337,In_621,In_187);
nor U2338 (N_2338,In_279,In_562);
nand U2339 (N_2339,In_42,In_333);
or U2340 (N_2340,In_878,In_701);
nor U2341 (N_2341,In_347,In_122);
xnor U2342 (N_2342,In_100,In_110);
nor U2343 (N_2343,In_943,In_277);
and U2344 (N_2344,In_920,In_532);
nor U2345 (N_2345,In_273,In_372);
and U2346 (N_2346,In_638,In_105);
nor U2347 (N_2347,In_501,In_933);
and U2348 (N_2348,In_700,In_742);
xor U2349 (N_2349,In_863,In_350);
or U2350 (N_2350,In_166,In_737);
and U2351 (N_2351,In_542,In_944);
and U2352 (N_2352,In_699,In_613);
nand U2353 (N_2353,In_716,In_981);
nor U2354 (N_2354,In_653,In_600);
xor U2355 (N_2355,In_382,In_172);
and U2356 (N_2356,In_497,In_644);
nor U2357 (N_2357,In_458,In_916);
nand U2358 (N_2358,In_231,In_654);
and U2359 (N_2359,In_20,In_401);
nand U2360 (N_2360,In_843,In_872);
nor U2361 (N_2361,In_113,In_984);
nor U2362 (N_2362,In_529,In_507);
or U2363 (N_2363,In_79,In_136);
or U2364 (N_2364,In_771,In_815);
nand U2365 (N_2365,In_364,In_29);
or U2366 (N_2366,In_902,In_776);
nand U2367 (N_2367,In_415,In_565);
xnor U2368 (N_2368,In_473,In_607);
and U2369 (N_2369,In_918,In_949);
nor U2370 (N_2370,In_274,In_491);
nand U2371 (N_2371,In_169,In_331);
and U2372 (N_2372,In_575,In_977);
and U2373 (N_2373,In_723,In_872);
and U2374 (N_2374,In_143,In_806);
nand U2375 (N_2375,In_0,In_424);
nor U2376 (N_2376,In_395,In_641);
xor U2377 (N_2377,In_328,In_931);
nor U2378 (N_2378,In_751,In_476);
and U2379 (N_2379,In_564,In_258);
and U2380 (N_2380,In_160,In_113);
nor U2381 (N_2381,In_102,In_32);
nor U2382 (N_2382,In_539,In_78);
and U2383 (N_2383,In_25,In_734);
and U2384 (N_2384,In_531,In_836);
nor U2385 (N_2385,In_736,In_597);
nand U2386 (N_2386,In_278,In_337);
nand U2387 (N_2387,In_951,In_693);
nor U2388 (N_2388,In_496,In_628);
nor U2389 (N_2389,In_603,In_137);
and U2390 (N_2390,In_358,In_266);
nor U2391 (N_2391,In_438,In_24);
xnor U2392 (N_2392,In_505,In_575);
nand U2393 (N_2393,In_482,In_445);
nor U2394 (N_2394,In_17,In_751);
or U2395 (N_2395,In_966,In_136);
or U2396 (N_2396,In_663,In_806);
nand U2397 (N_2397,In_130,In_388);
or U2398 (N_2398,In_529,In_673);
nand U2399 (N_2399,In_933,In_937);
nor U2400 (N_2400,In_866,In_403);
nand U2401 (N_2401,In_293,In_440);
or U2402 (N_2402,In_149,In_256);
nor U2403 (N_2403,In_12,In_705);
nor U2404 (N_2404,In_625,In_259);
xnor U2405 (N_2405,In_799,In_468);
nor U2406 (N_2406,In_171,In_926);
and U2407 (N_2407,In_490,In_981);
nand U2408 (N_2408,In_581,In_960);
and U2409 (N_2409,In_158,In_283);
and U2410 (N_2410,In_356,In_739);
or U2411 (N_2411,In_884,In_602);
nand U2412 (N_2412,In_686,In_923);
nand U2413 (N_2413,In_588,In_395);
and U2414 (N_2414,In_748,In_706);
nand U2415 (N_2415,In_626,In_542);
and U2416 (N_2416,In_170,In_99);
or U2417 (N_2417,In_289,In_902);
nor U2418 (N_2418,In_596,In_469);
nor U2419 (N_2419,In_516,In_823);
xnor U2420 (N_2420,In_224,In_203);
nand U2421 (N_2421,In_880,In_838);
or U2422 (N_2422,In_549,In_212);
and U2423 (N_2423,In_298,In_749);
nand U2424 (N_2424,In_892,In_392);
or U2425 (N_2425,In_416,In_267);
nand U2426 (N_2426,In_500,In_867);
nor U2427 (N_2427,In_672,In_585);
nor U2428 (N_2428,In_22,In_935);
nand U2429 (N_2429,In_937,In_310);
and U2430 (N_2430,In_591,In_620);
nor U2431 (N_2431,In_182,In_177);
nand U2432 (N_2432,In_58,In_144);
nand U2433 (N_2433,In_147,In_367);
nand U2434 (N_2434,In_253,In_339);
and U2435 (N_2435,In_929,In_952);
nand U2436 (N_2436,In_621,In_730);
or U2437 (N_2437,In_614,In_75);
nor U2438 (N_2438,In_334,In_945);
nor U2439 (N_2439,In_716,In_14);
or U2440 (N_2440,In_806,In_191);
xor U2441 (N_2441,In_235,In_622);
or U2442 (N_2442,In_697,In_775);
nor U2443 (N_2443,In_257,In_415);
and U2444 (N_2444,In_531,In_998);
nand U2445 (N_2445,In_883,In_837);
nand U2446 (N_2446,In_947,In_291);
or U2447 (N_2447,In_205,In_694);
or U2448 (N_2448,In_743,In_93);
or U2449 (N_2449,In_949,In_838);
nand U2450 (N_2450,In_111,In_759);
nand U2451 (N_2451,In_495,In_11);
and U2452 (N_2452,In_381,In_68);
nor U2453 (N_2453,In_873,In_187);
nand U2454 (N_2454,In_59,In_837);
and U2455 (N_2455,In_402,In_117);
or U2456 (N_2456,In_966,In_932);
and U2457 (N_2457,In_129,In_665);
and U2458 (N_2458,In_394,In_276);
nand U2459 (N_2459,In_750,In_785);
or U2460 (N_2460,In_791,In_77);
and U2461 (N_2461,In_481,In_108);
nor U2462 (N_2462,In_979,In_499);
nor U2463 (N_2463,In_257,In_337);
nand U2464 (N_2464,In_672,In_174);
or U2465 (N_2465,In_545,In_852);
or U2466 (N_2466,In_836,In_529);
or U2467 (N_2467,In_416,In_742);
and U2468 (N_2468,In_363,In_9);
and U2469 (N_2469,In_37,In_478);
and U2470 (N_2470,In_912,In_663);
xnor U2471 (N_2471,In_997,In_567);
nor U2472 (N_2472,In_847,In_999);
and U2473 (N_2473,In_998,In_545);
or U2474 (N_2474,In_408,In_746);
nand U2475 (N_2475,In_336,In_659);
or U2476 (N_2476,In_658,In_814);
and U2477 (N_2477,In_171,In_861);
nand U2478 (N_2478,In_822,In_545);
or U2479 (N_2479,In_500,In_707);
nand U2480 (N_2480,In_586,In_712);
or U2481 (N_2481,In_798,In_20);
and U2482 (N_2482,In_477,In_1);
and U2483 (N_2483,In_898,In_490);
and U2484 (N_2484,In_120,In_695);
or U2485 (N_2485,In_980,In_826);
nand U2486 (N_2486,In_528,In_172);
nand U2487 (N_2487,In_273,In_711);
and U2488 (N_2488,In_533,In_346);
nand U2489 (N_2489,In_389,In_69);
or U2490 (N_2490,In_357,In_310);
nand U2491 (N_2491,In_163,In_68);
nand U2492 (N_2492,In_766,In_492);
nor U2493 (N_2493,In_936,In_826);
and U2494 (N_2494,In_186,In_554);
and U2495 (N_2495,In_560,In_960);
nor U2496 (N_2496,In_290,In_521);
nor U2497 (N_2497,In_90,In_373);
nor U2498 (N_2498,In_545,In_926);
and U2499 (N_2499,In_946,In_791);
nor U2500 (N_2500,In_637,In_925);
and U2501 (N_2501,In_983,In_378);
or U2502 (N_2502,In_625,In_233);
nor U2503 (N_2503,In_290,In_225);
and U2504 (N_2504,In_572,In_675);
or U2505 (N_2505,In_405,In_86);
xnor U2506 (N_2506,In_642,In_507);
or U2507 (N_2507,In_544,In_885);
nor U2508 (N_2508,In_213,In_580);
nor U2509 (N_2509,In_653,In_903);
or U2510 (N_2510,In_100,In_670);
nand U2511 (N_2511,In_286,In_48);
and U2512 (N_2512,In_117,In_345);
and U2513 (N_2513,In_558,In_258);
nand U2514 (N_2514,In_668,In_989);
xnor U2515 (N_2515,In_794,In_816);
nand U2516 (N_2516,In_876,In_288);
or U2517 (N_2517,In_546,In_530);
or U2518 (N_2518,In_225,In_184);
nor U2519 (N_2519,In_619,In_161);
and U2520 (N_2520,In_79,In_967);
and U2521 (N_2521,In_573,In_718);
nand U2522 (N_2522,In_302,In_549);
nand U2523 (N_2523,In_257,In_522);
nand U2524 (N_2524,In_419,In_100);
or U2525 (N_2525,In_728,In_143);
and U2526 (N_2526,In_419,In_54);
and U2527 (N_2527,In_650,In_693);
or U2528 (N_2528,In_412,In_356);
nor U2529 (N_2529,In_604,In_716);
and U2530 (N_2530,In_988,In_11);
or U2531 (N_2531,In_731,In_146);
and U2532 (N_2532,In_190,In_983);
or U2533 (N_2533,In_164,In_903);
xnor U2534 (N_2534,In_957,In_829);
nand U2535 (N_2535,In_858,In_377);
nand U2536 (N_2536,In_21,In_199);
nand U2537 (N_2537,In_509,In_763);
or U2538 (N_2538,In_554,In_689);
nor U2539 (N_2539,In_765,In_930);
nor U2540 (N_2540,In_286,In_748);
nand U2541 (N_2541,In_679,In_393);
nand U2542 (N_2542,In_944,In_754);
nand U2543 (N_2543,In_654,In_98);
nor U2544 (N_2544,In_245,In_273);
or U2545 (N_2545,In_297,In_942);
nand U2546 (N_2546,In_511,In_945);
nor U2547 (N_2547,In_808,In_598);
nor U2548 (N_2548,In_899,In_933);
or U2549 (N_2549,In_540,In_563);
or U2550 (N_2550,In_986,In_395);
and U2551 (N_2551,In_527,In_416);
nor U2552 (N_2552,In_902,In_180);
or U2553 (N_2553,In_71,In_335);
and U2554 (N_2554,In_39,In_552);
nand U2555 (N_2555,In_938,In_937);
nor U2556 (N_2556,In_499,In_201);
nor U2557 (N_2557,In_875,In_952);
and U2558 (N_2558,In_889,In_104);
and U2559 (N_2559,In_988,In_10);
nor U2560 (N_2560,In_196,In_968);
xor U2561 (N_2561,In_778,In_523);
and U2562 (N_2562,In_951,In_632);
nor U2563 (N_2563,In_82,In_664);
nand U2564 (N_2564,In_71,In_963);
or U2565 (N_2565,In_112,In_740);
nor U2566 (N_2566,In_374,In_129);
xor U2567 (N_2567,In_225,In_471);
nor U2568 (N_2568,In_176,In_456);
nor U2569 (N_2569,In_524,In_314);
xnor U2570 (N_2570,In_886,In_454);
nor U2571 (N_2571,In_166,In_208);
or U2572 (N_2572,In_353,In_475);
and U2573 (N_2573,In_883,In_561);
nor U2574 (N_2574,In_868,In_230);
nor U2575 (N_2575,In_155,In_392);
nor U2576 (N_2576,In_275,In_699);
nand U2577 (N_2577,In_503,In_666);
nor U2578 (N_2578,In_68,In_811);
or U2579 (N_2579,In_259,In_80);
and U2580 (N_2580,In_504,In_926);
nor U2581 (N_2581,In_427,In_352);
nor U2582 (N_2582,In_819,In_531);
nor U2583 (N_2583,In_610,In_157);
nand U2584 (N_2584,In_538,In_282);
nand U2585 (N_2585,In_941,In_610);
or U2586 (N_2586,In_212,In_308);
nand U2587 (N_2587,In_632,In_116);
or U2588 (N_2588,In_714,In_191);
nand U2589 (N_2589,In_184,In_919);
nor U2590 (N_2590,In_0,In_255);
and U2591 (N_2591,In_927,In_246);
nor U2592 (N_2592,In_855,In_106);
or U2593 (N_2593,In_153,In_357);
and U2594 (N_2594,In_610,In_406);
or U2595 (N_2595,In_663,In_474);
nand U2596 (N_2596,In_377,In_518);
and U2597 (N_2597,In_439,In_268);
and U2598 (N_2598,In_116,In_286);
or U2599 (N_2599,In_429,In_873);
and U2600 (N_2600,In_265,In_557);
or U2601 (N_2601,In_161,In_974);
nand U2602 (N_2602,In_889,In_670);
or U2603 (N_2603,In_645,In_784);
or U2604 (N_2604,In_26,In_317);
nand U2605 (N_2605,In_930,In_149);
and U2606 (N_2606,In_547,In_22);
nand U2607 (N_2607,In_609,In_152);
or U2608 (N_2608,In_487,In_506);
and U2609 (N_2609,In_491,In_503);
nor U2610 (N_2610,In_499,In_241);
and U2611 (N_2611,In_606,In_479);
or U2612 (N_2612,In_454,In_373);
or U2613 (N_2613,In_391,In_44);
nor U2614 (N_2614,In_595,In_880);
nor U2615 (N_2615,In_742,In_672);
and U2616 (N_2616,In_927,In_386);
and U2617 (N_2617,In_129,In_473);
and U2618 (N_2618,In_304,In_720);
nor U2619 (N_2619,In_613,In_752);
xor U2620 (N_2620,In_416,In_552);
xnor U2621 (N_2621,In_876,In_898);
or U2622 (N_2622,In_977,In_543);
nand U2623 (N_2623,In_628,In_637);
nor U2624 (N_2624,In_366,In_687);
and U2625 (N_2625,In_914,In_266);
nor U2626 (N_2626,In_268,In_999);
nor U2627 (N_2627,In_752,In_198);
nand U2628 (N_2628,In_560,In_134);
or U2629 (N_2629,In_420,In_643);
or U2630 (N_2630,In_354,In_575);
nand U2631 (N_2631,In_847,In_524);
nor U2632 (N_2632,In_440,In_500);
nand U2633 (N_2633,In_683,In_351);
nor U2634 (N_2634,In_624,In_846);
nand U2635 (N_2635,In_41,In_453);
and U2636 (N_2636,In_198,In_536);
xor U2637 (N_2637,In_327,In_218);
or U2638 (N_2638,In_264,In_974);
nand U2639 (N_2639,In_887,In_788);
nand U2640 (N_2640,In_592,In_948);
nor U2641 (N_2641,In_583,In_641);
and U2642 (N_2642,In_78,In_858);
nand U2643 (N_2643,In_637,In_806);
nand U2644 (N_2644,In_950,In_85);
xnor U2645 (N_2645,In_51,In_44);
or U2646 (N_2646,In_554,In_938);
nor U2647 (N_2647,In_163,In_62);
nand U2648 (N_2648,In_798,In_479);
or U2649 (N_2649,In_157,In_397);
and U2650 (N_2650,In_557,In_221);
nand U2651 (N_2651,In_54,In_613);
nor U2652 (N_2652,In_334,In_61);
or U2653 (N_2653,In_770,In_649);
nor U2654 (N_2654,In_386,In_68);
or U2655 (N_2655,In_977,In_959);
nand U2656 (N_2656,In_695,In_718);
or U2657 (N_2657,In_414,In_364);
or U2658 (N_2658,In_561,In_530);
and U2659 (N_2659,In_761,In_232);
or U2660 (N_2660,In_906,In_159);
nor U2661 (N_2661,In_452,In_274);
or U2662 (N_2662,In_513,In_666);
nor U2663 (N_2663,In_759,In_153);
or U2664 (N_2664,In_259,In_294);
xor U2665 (N_2665,In_551,In_361);
and U2666 (N_2666,In_776,In_458);
nand U2667 (N_2667,In_101,In_860);
and U2668 (N_2668,In_437,In_445);
and U2669 (N_2669,In_949,In_719);
xor U2670 (N_2670,In_297,In_826);
and U2671 (N_2671,In_10,In_527);
nand U2672 (N_2672,In_315,In_18);
and U2673 (N_2673,In_568,In_574);
nand U2674 (N_2674,In_103,In_43);
nor U2675 (N_2675,In_623,In_424);
nand U2676 (N_2676,In_420,In_981);
nor U2677 (N_2677,In_37,In_995);
or U2678 (N_2678,In_496,In_726);
nor U2679 (N_2679,In_350,In_98);
and U2680 (N_2680,In_484,In_760);
nor U2681 (N_2681,In_135,In_273);
nand U2682 (N_2682,In_852,In_636);
nand U2683 (N_2683,In_938,In_284);
nand U2684 (N_2684,In_545,In_692);
nor U2685 (N_2685,In_404,In_251);
nor U2686 (N_2686,In_122,In_658);
or U2687 (N_2687,In_470,In_455);
xor U2688 (N_2688,In_161,In_438);
and U2689 (N_2689,In_426,In_209);
and U2690 (N_2690,In_708,In_203);
and U2691 (N_2691,In_754,In_397);
or U2692 (N_2692,In_571,In_701);
or U2693 (N_2693,In_55,In_723);
nor U2694 (N_2694,In_672,In_749);
or U2695 (N_2695,In_693,In_888);
nor U2696 (N_2696,In_666,In_177);
or U2697 (N_2697,In_781,In_333);
nor U2698 (N_2698,In_32,In_385);
and U2699 (N_2699,In_831,In_736);
nor U2700 (N_2700,In_539,In_548);
and U2701 (N_2701,In_762,In_993);
or U2702 (N_2702,In_594,In_422);
or U2703 (N_2703,In_972,In_317);
or U2704 (N_2704,In_90,In_936);
nand U2705 (N_2705,In_82,In_127);
nand U2706 (N_2706,In_423,In_308);
nand U2707 (N_2707,In_676,In_968);
nand U2708 (N_2708,In_582,In_952);
and U2709 (N_2709,In_72,In_872);
or U2710 (N_2710,In_457,In_942);
nand U2711 (N_2711,In_643,In_511);
nand U2712 (N_2712,In_322,In_231);
or U2713 (N_2713,In_487,In_184);
or U2714 (N_2714,In_424,In_293);
or U2715 (N_2715,In_967,In_135);
nand U2716 (N_2716,In_838,In_922);
nor U2717 (N_2717,In_330,In_479);
nor U2718 (N_2718,In_687,In_436);
or U2719 (N_2719,In_173,In_968);
xor U2720 (N_2720,In_275,In_249);
nor U2721 (N_2721,In_551,In_913);
nor U2722 (N_2722,In_883,In_110);
and U2723 (N_2723,In_239,In_246);
or U2724 (N_2724,In_196,In_428);
nor U2725 (N_2725,In_83,In_851);
nor U2726 (N_2726,In_531,In_927);
and U2727 (N_2727,In_311,In_740);
nand U2728 (N_2728,In_125,In_879);
nor U2729 (N_2729,In_688,In_173);
and U2730 (N_2730,In_482,In_867);
nor U2731 (N_2731,In_424,In_533);
or U2732 (N_2732,In_737,In_792);
and U2733 (N_2733,In_1,In_288);
nor U2734 (N_2734,In_561,In_794);
and U2735 (N_2735,In_39,In_418);
and U2736 (N_2736,In_673,In_76);
nor U2737 (N_2737,In_973,In_50);
or U2738 (N_2738,In_356,In_994);
and U2739 (N_2739,In_178,In_773);
nand U2740 (N_2740,In_811,In_121);
and U2741 (N_2741,In_561,In_593);
nand U2742 (N_2742,In_809,In_974);
or U2743 (N_2743,In_935,In_216);
or U2744 (N_2744,In_88,In_146);
nand U2745 (N_2745,In_33,In_989);
nor U2746 (N_2746,In_128,In_102);
and U2747 (N_2747,In_864,In_25);
nor U2748 (N_2748,In_503,In_223);
or U2749 (N_2749,In_903,In_344);
nor U2750 (N_2750,In_729,In_346);
nor U2751 (N_2751,In_430,In_424);
and U2752 (N_2752,In_833,In_805);
nor U2753 (N_2753,In_397,In_670);
or U2754 (N_2754,In_225,In_543);
nand U2755 (N_2755,In_476,In_528);
nor U2756 (N_2756,In_464,In_440);
nor U2757 (N_2757,In_477,In_265);
and U2758 (N_2758,In_555,In_175);
nor U2759 (N_2759,In_689,In_123);
nor U2760 (N_2760,In_691,In_303);
nand U2761 (N_2761,In_74,In_190);
nand U2762 (N_2762,In_241,In_550);
nor U2763 (N_2763,In_915,In_895);
nand U2764 (N_2764,In_789,In_827);
nand U2765 (N_2765,In_694,In_622);
nor U2766 (N_2766,In_287,In_365);
nand U2767 (N_2767,In_193,In_905);
nor U2768 (N_2768,In_389,In_506);
or U2769 (N_2769,In_777,In_537);
or U2770 (N_2770,In_50,In_353);
nor U2771 (N_2771,In_574,In_313);
or U2772 (N_2772,In_413,In_986);
nor U2773 (N_2773,In_378,In_986);
xnor U2774 (N_2774,In_731,In_157);
or U2775 (N_2775,In_829,In_230);
and U2776 (N_2776,In_530,In_579);
nor U2777 (N_2777,In_504,In_741);
and U2778 (N_2778,In_584,In_973);
nand U2779 (N_2779,In_734,In_707);
nor U2780 (N_2780,In_300,In_453);
and U2781 (N_2781,In_827,In_806);
nand U2782 (N_2782,In_84,In_26);
xnor U2783 (N_2783,In_300,In_898);
and U2784 (N_2784,In_584,In_946);
and U2785 (N_2785,In_900,In_494);
nor U2786 (N_2786,In_257,In_570);
and U2787 (N_2787,In_666,In_321);
nor U2788 (N_2788,In_637,In_185);
or U2789 (N_2789,In_224,In_475);
and U2790 (N_2790,In_355,In_68);
nor U2791 (N_2791,In_884,In_900);
nand U2792 (N_2792,In_146,In_806);
or U2793 (N_2793,In_781,In_538);
and U2794 (N_2794,In_187,In_411);
nor U2795 (N_2795,In_574,In_424);
nand U2796 (N_2796,In_109,In_894);
or U2797 (N_2797,In_561,In_862);
nor U2798 (N_2798,In_696,In_337);
nor U2799 (N_2799,In_446,In_964);
or U2800 (N_2800,In_903,In_642);
nor U2801 (N_2801,In_310,In_296);
nand U2802 (N_2802,In_219,In_447);
and U2803 (N_2803,In_284,In_571);
nand U2804 (N_2804,In_942,In_848);
nand U2805 (N_2805,In_974,In_227);
and U2806 (N_2806,In_24,In_510);
or U2807 (N_2807,In_271,In_643);
nor U2808 (N_2808,In_851,In_693);
and U2809 (N_2809,In_681,In_292);
nor U2810 (N_2810,In_306,In_219);
nand U2811 (N_2811,In_147,In_186);
or U2812 (N_2812,In_931,In_529);
or U2813 (N_2813,In_968,In_241);
nand U2814 (N_2814,In_101,In_797);
or U2815 (N_2815,In_743,In_169);
and U2816 (N_2816,In_119,In_93);
or U2817 (N_2817,In_112,In_194);
nand U2818 (N_2818,In_156,In_650);
and U2819 (N_2819,In_983,In_329);
nand U2820 (N_2820,In_888,In_662);
nand U2821 (N_2821,In_282,In_135);
or U2822 (N_2822,In_363,In_401);
and U2823 (N_2823,In_632,In_660);
and U2824 (N_2824,In_93,In_328);
or U2825 (N_2825,In_811,In_127);
nand U2826 (N_2826,In_695,In_571);
xor U2827 (N_2827,In_494,In_367);
or U2828 (N_2828,In_90,In_458);
nor U2829 (N_2829,In_212,In_290);
and U2830 (N_2830,In_633,In_752);
xor U2831 (N_2831,In_643,In_186);
or U2832 (N_2832,In_797,In_756);
nor U2833 (N_2833,In_858,In_597);
xor U2834 (N_2834,In_225,In_315);
and U2835 (N_2835,In_788,In_5);
nand U2836 (N_2836,In_814,In_397);
or U2837 (N_2837,In_100,In_401);
and U2838 (N_2838,In_956,In_484);
nor U2839 (N_2839,In_308,In_942);
nand U2840 (N_2840,In_159,In_420);
nand U2841 (N_2841,In_887,In_508);
xor U2842 (N_2842,In_753,In_245);
and U2843 (N_2843,In_275,In_302);
nor U2844 (N_2844,In_65,In_372);
nor U2845 (N_2845,In_481,In_787);
or U2846 (N_2846,In_933,In_137);
and U2847 (N_2847,In_770,In_858);
or U2848 (N_2848,In_467,In_274);
or U2849 (N_2849,In_278,In_351);
nor U2850 (N_2850,In_918,In_845);
nor U2851 (N_2851,In_614,In_122);
nand U2852 (N_2852,In_617,In_121);
and U2853 (N_2853,In_39,In_773);
nor U2854 (N_2854,In_778,In_527);
or U2855 (N_2855,In_734,In_555);
or U2856 (N_2856,In_685,In_340);
and U2857 (N_2857,In_5,In_555);
nor U2858 (N_2858,In_668,In_892);
or U2859 (N_2859,In_137,In_812);
nor U2860 (N_2860,In_819,In_500);
or U2861 (N_2861,In_378,In_972);
or U2862 (N_2862,In_764,In_711);
or U2863 (N_2863,In_569,In_472);
nand U2864 (N_2864,In_72,In_745);
or U2865 (N_2865,In_499,In_453);
nand U2866 (N_2866,In_230,In_495);
or U2867 (N_2867,In_314,In_522);
nor U2868 (N_2868,In_759,In_699);
or U2869 (N_2869,In_725,In_642);
nor U2870 (N_2870,In_548,In_480);
nor U2871 (N_2871,In_105,In_550);
nand U2872 (N_2872,In_726,In_450);
and U2873 (N_2873,In_574,In_280);
nand U2874 (N_2874,In_712,In_118);
nor U2875 (N_2875,In_617,In_471);
nor U2876 (N_2876,In_46,In_9);
nor U2877 (N_2877,In_214,In_670);
and U2878 (N_2878,In_903,In_934);
nor U2879 (N_2879,In_344,In_614);
nor U2880 (N_2880,In_911,In_356);
nand U2881 (N_2881,In_888,In_941);
or U2882 (N_2882,In_694,In_602);
nor U2883 (N_2883,In_543,In_601);
or U2884 (N_2884,In_73,In_36);
nor U2885 (N_2885,In_31,In_780);
or U2886 (N_2886,In_163,In_775);
nor U2887 (N_2887,In_548,In_88);
or U2888 (N_2888,In_120,In_502);
nand U2889 (N_2889,In_531,In_771);
or U2890 (N_2890,In_643,In_541);
or U2891 (N_2891,In_19,In_666);
and U2892 (N_2892,In_857,In_572);
and U2893 (N_2893,In_653,In_819);
or U2894 (N_2894,In_238,In_521);
nand U2895 (N_2895,In_51,In_978);
nand U2896 (N_2896,In_914,In_58);
and U2897 (N_2897,In_840,In_119);
nor U2898 (N_2898,In_341,In_864);
and U2899 (N_2899,In_181,In_33);
and U2900 (N_2900,In_936,In_842);
or U2901 (N_2901,In_170,In_195);
nor U2902 (N_2902,In_687,In_55);
or U2903 (N_2903,In_128,In_749);
nor U2904 (N_2904,In_893,In_596);
or U2905 (N_2905,In_56,In_990);
nand U2906 (N_2906,In_853,In_459);
nor U2907 (N_2907,In_824,In_581);
or U2908 (N_2908,In_515,In_80);
and U2909 (N_2909,In_474,In_170);
and U2910 (N_2910,In_269,In_919);
or U2911 (N_2911,In_891,In_183);
and U2912 (N_2912,In_601,In_348);
nand U2913 (N_2913,In_657,In_57);
nand U2914 (N_2914,In_375,In_719);
and U2915 (N_2915,In_874,In_151);
and U2916 (N_2916,In_857,In_852);
nor U2917 (N_2917,In_350,In_597);
and U2918 (N_2918,In_791,In_38);
nand U2919 (N_2919,In_652,In_354);
nand U2920 (N_2920,In_671,In_150);
or U2921 (N_2921,In_650,In_79);
or U2922 (N_2922,In_154,In_149);
or U2923 (N_2923,In_875,In_340);
or U2924 (N_2924,In_657,In_381);
nor U2925 (N_2925,In_921,In_422);
nor U2926 (N_2926,In_812,In_274);
nor U2927 (N_2927,In_540,In_195);
and U2928 (N_2928,In_402,In_693);
nand U2929 (N_2929,In_672,In_707);
and U2930 (N_2930,In_998,In_719);
nor U2931 (N_2931,In_405,In_714);
or U2932 (N_2932,In_771,In_889);
or U2933 (N_2933,In_203,In_898);
or U2934 (N_2934,In_228,In_135);
nand U2935 (N_2935,In_114,In_135);
xor U2936 (N_2936,In_414,In_407);
nor U2937 (N_2937,In_22,In_557);
nand U2938 (N_2938,In_204,In_32);
and U2939 (N_2939,In_546,In_854);
nor U2940 (N_2940,In_928,In_567);
nor U2941 (N_2941,In_709,In_208);
nor U2942 (N_2942,In_541,In_658);
nand U2943 (N_2943,In_146,In_301);
nand U2944 (N_2944,In_18,In_191);
or U2945 (N_2945,In_628,In_289);
nor U2946 (N_2946,In_59,In_489);
nor U2947 (N_2947,In_470,In_673);
or U2948 (N_2948,In_856,In_905);
nand U2949 (N_2949,In_392,In_594);
and U2950 (N_2950,In_875,In_747);
or U2951 (N_2951,In_215,In_884);
and U2952 (N_2952,In_796,In_880);
nor U2953 (N_2953,In_540,In_783);
nand U2954 (N_2954,In_675,In_60);
or U2955 (N_2955,In_868,In_880);
nand U2956 (N_2956,In_96,In_436);
and U2957 (N_2957,In_453,In_887);
and U2958 (N_2958,In_586,In_113);
or U2959 (N_2959,In_988,In_662);
and U2960 (N_2960,In_963,In_213);
or U2961 (N_2961,In_153,In_962);
nand U2962 (N_2962,In_547,In_790);
nand U2963 (N_2963,In_539,In_9);
nor U2964 (N_2964,In_174,In_302);
nor U2965 (N_2965,In_534,In_557);
or U2966 (N_2966,In_677,In_427);
or U2967 (N_2967,In_421,In_523);
nor U2968 (N_2968,In_337,In_366);
and U2969 (N_2969,In_128,In_752);
nand U2970 (N_2970,In_579,In_974);
or U2971 (N_2971,In_662,In_798);
nor U2972 (N_2972,In_866,In_806);
nand U2973 (N_2973,In_421,In_822);
nand U2974 (N_2974,In_46,In_651);
nor U2975 (N_2975,In_883,In_254);
nor U2976 (N_2976,In_292,In_842);
nand U2977 (N_2977,In_661,In_912);
and U2978 (N_2978,In_925,In_804);
or U2979 (N_2979,In_368,In_739);
nand U2980 (N_2980,In_437,In_433);
or U2981 (N_2981,In_31,In_500);
nand U2982 (N_2982,In_583,In_269);
or U2983 (N_2983,In_346,In_847);
nand U2984 (N_2984,In_947,In_191);
or U2985 (N_2985,In_305,In_705);
nand U2986 (N_2986,In_167,In_410);
xnor U2987 (N_2987,In_491,In_372);
nand U2988 (N_2988,In_962,In_278);
nand U2989 (N_2989,In_585,In_358);
or U2990 (N_2990,In_88,In_566);
and U2991 (N_2991,In_881,In_779);
xnor U2992 (N_2992,In_57,In_622);
nand U2993 (N_2993,In_178,In_295);
or U2994 (N_2994,In_275,In_218);
nand U2995 (N_2995,In_798,In_652);
or U2996 (N_2996,In_561,In_770);
and U2997 (N_2997,In_506,In_782);
nand U2998 (N_2998,In_242,In_432);
and U2999 (N_2999,In_445,In_553);
nor U3000 (N_3000,In_14,In_145);
and U3001 (N_3001,In_187,In_887);
nor U3002 (N_3002,In_90,In_584);
nor U3003 (N_3003,In_342,In_508);
and U3004 (N_3004,In_173,In_301);
and U3005 (N_3005,In_166,In_768);
nand U3006 (N_3006,In_851,In_199);
nor U3007 (N_3007,In_332,In_818);
and U3008 (N_3008,In_428,In_444);
and U3009 (N_3009,In_500,In_904);
nand U3010 (N_3010,In_973,In_479);
or U3011 (N_3011,In_922,In_154);
nand U3012 (N_3012,In_159,In_661);
nand U3013 (N_3013,In_601,In_811);
or U3014 (N_3014,In_563,In_370);
or U3015 (N_3015,In_457,In_177);
nand U3016 (N_3016,In_816,In_661);
and U3017 (N_3017,In_807,In_374);
nor U3018 (N_3018,In_890,In_278);
nand U3019 (N_3019,In_246,In_479);
and U3020 (N_3020,In_4,In_489);
nor U3021 (N_3021,In_418,In_925);
xor U3022 (N_3022,In_553,In_886);
and U3023 (N_3023,In_232,In_251);
nand U3024 (N_3024,In_551,In_212);
or U3025 (N_3025,In_1,In_431);
nand U3026 (N_3026,In_153,In_795);
nand U3027 (N_3027,In_528,In_80);
and U3028 (N_3028,In_85,In_614);
nand U3029 (N_3029,In_145,In_188);
nor U3030 (N_3030,In_926,In_36);
nand U3031 (N_3031,In_566,In_676);
nand U3032 (N_3032,In_584,In_199);
nor U3033 (N_3033,In_9,In_382);
xor U3034 (N_3034,In_656,In_923);
or U3035 (N_3035,In_412,In_88);
nor U3036 (N_3036,In_774,In_678);
nand U3037 (N_3037,In_389,In_458);
nor U3038 (N_3038,In_0,In_252);
nor U3039 (N_3039,In_47,In_282);
and U3040 (N_3040,In_542,In_869);
or U3041 (N_3041,In_862,In_761);
and U3042 (N_3042,In_259,In_897);
and U3043 (N_3043,In_492,In_851);
nand U3044 (N_3044,In_13,In_938);
or U3045 (N_3045,In_53,In_735);
nand U3046 (N_3046,In_367,In_565);
and U3047 (N_3047,In_749,In_253);
or U3048 (N_3048,In_509,In_598);
or U3049 (N_3049,In_51,In_580);
and U3050 (N_3050,In_455,In_308);
xnor U3051 (N_3051,In_999,In_559);
nand U3052 (N_3052,In_448,In_973);
and U3053 (N_3053,In_186,In_860);
xor U3054 (N_3054,In_790,In_62);
nand U3055 (N_3055,In_872,In_927);
or U3056 (N_3056,In_120,In_779);
nor U3057 (N_3057,In_930,In_881);
nand U3058 (N_3058,In_393,In_474);
or U3059 (N_3059,In_330,In_407);
and U3060 (N_3060,In_378,In_159);
or U3061 (N_3061,In_995,In_330);
or U3062 (N_3062,In_594,In_755);
nor U3063 (N_3063,In_716,In_844);
and U3064 (N_3064,In_2,In_587);
or U3065 (N_3065,In_117,In_950);
and U3066 (N_3066,In_630,In_822);
nor U3067 (N_3067,In_371,In_362);
nor U3068 (N_3068,In_76,In_637);
xor U3069 (N_3069,In_331,In_520);
and U3070 (N_3070,In_454,In_28);
nor U3071 (N_3071,In_379,In_372);
xnor U3072 (N_3072,In_631,In_944);
nor U3073 (N_3073,In_586,In_342);
or U3074 (N_3074,In_24,In_664);
or U3075 (N_3075,In_127,In_683);
nor U3076 (N_3076,In_830,In_988);
nor U3077 (N_3077,In_456,In_277);
nand U3078 (N_3078,In_629,In_376);
and U3079 (N_3079,In_207,In_791);
or U3080 (N_3080,In_309,In_811);
nor U3081 (N_3081,In_40,In_93);
nand U3082 (N_3082,In_587,In_872);
nand U3083 (N_3083,In_137,In_808);
nand U3084 (N_3084,In_862,In_893);
nand U3085 (N_3085,In_199,In_591);
nor U3086 (N_3086,In_871,In_9);
and U3087 (N_3087,In_115,In_675);
or U3088 (N_3088,In_703,In_412);
or U3089 (N_3089,In_30,In_966);
xor U3090 (N_3090,In_853,In_894);
and U3091 (N_3091,In_630,In_459);
nor U3092 (N_3092,In_861,In_7);
or U3093 (N_3093,In_604,In_344);
or U3094 (N_3094,In_81,In_420);
or U3095 (N_3095,In_870,In_577);
nand U3096 (N_3096,In_591,In_31);
or U3097 (N_3097,In_364,In_82);
or U3098 (N_3098,In_180,In_583);
nor U3099 (N_3099,In_532,In_538);
or U3100 (N_3100,In_438,In_986);
or U3101 (N_3101,In_612,In_285);
nand U3102 (N_3102,In_268,In_148);
and U3103 (N_3103,In_226,In_694);
nand U3104 (N_3104,In_799,In_336);
nand U3105 (N_3105,In_518,In_20);
and U3106 (N_3106,In_964,In_943);
or U3107 (N_3107,In_196,In_831);
and U3108 (N_3108,In_288,In_761);
nor U3109 (N_3109,In_814,In_736);
nor U3110 (N_3110,In_48,In_449);
and U3111 (N_3111,In_533,In_118);
nor U3112 (N_3112,In_597,In_105);
or U3113 (N_3113,In_388,In_373);
nor U3114 (N_3114,In_306,In_640);
nand U3115 (N_3115,In_956,In_732);
and U3116 (N_3116,In_612,In_659);
or U3117 (N_3117,In_847,In_738);
and U3118 (N_3118,In_400,In_832);
nand U3119 (N_3119,In_392,In_753);
nand U3120 (N_3120,In_46,In_228);
and U3121 (N_3121,In_327,In_894);
xnor U3122 (N_3122,In_685,In_233);
or U3123 (N_3123,In_661,In_350);
and U3124 (N_3124,In_324,In_921);
or U3125 (N_3125,In_425,In_645);
or U3126 (N_3126,In_182,In_342);
nand U3127 (N_3127,In_139,In_19);
and U3128 (N_3128,In_203,In_913);
or U3129 (N_3129,In_376,In_135);
nor U3130 (N_3130,In_229,In_256);
and U3131 (N_3131,In_693,In_922);
and U3132 (N_3132,In_978,In_508);
and U3133 (N_3133,In_781,In_861);
nor U3134 (N_3134,In_345,In_417);
nor U3135 (N_3135,In_361,In_571);
and U3136 (N_3136,In_295,In_649);
nor U3137 (N_3137,In_564,In_110);
or U3138 (N_3138,In_274,In_292);
and U3139 (N_3139,In_132,In_388);
nand U3140 (N_3140,In_671,In_716);
or U3141 (N_3141,In_972,In_330);
nand U3142 (N_3142,In_420,In_852);
nand U3143 (N_3143,In_483,In_724);
and U3144 (N_3144,In_878,In_495);
xnor U3145 (N_3145,In_854,In_479);
nor U3146 (N_3146,In_462,In_863);
or U3147 (N_3147,In_95,In_571);
and U3148 (N_3148,In_117,In_678);
or U3149 (N_3149,In_298,In_1);
nand U3150 (N_3150,In_838,In_958);
nor U3151 (N_3151,In_432,In_77);
or U3152 (N_3152,In_650,In_252);
nand U3153 (N_3153,In_965,In_395);
nor U3154 (N_3154,In_927,In_474);
nor U3155 (N_3155,In_939,In_601);
xnor U3156 (N_3156,In_65,In_784);
and U3157 (N_3157,In_700,In_969);
nand U3158 (N_3158,In_787,In_904);
or U3159 (N_3159,In_58,In_867);
or U3160 (N_3160,In_969,In_422);
nor U3161 (N_3161,In_143,In_386);
xor U3162 (N_3162,In_962,In_603);
and U3163 (N_3163,In_853,In_34);
and U3164 (N_3164,In_95,In_118);
and U3165 (N_3165,In_273,In_479);
nor U3166 (N_3166,In_718,In_581);
or U3167 (N_3167,In_811,In_674);
nor U3168 (N_3168,In_170,In_465);
nor U3169 (N_3169,In_241,In_962);
nor U3170 (N_3170,In_572,In_704);
or U3171 (N_3171,In_664,In_855);
nor U3172 (N_3172,In_167,In_547);
nor U3173 (N_3173,In_798,In_913);
and U3174 (N_3174,In_12,In_556);
nand U3175 (N_3175,In_805,In_372);
and U3176 (N_3176,In_950,In_34);
nand U3177 (N_3177,In_208,In_200);
and U3178 (N_3178,In_621,In_73);
or U3179 (N_3179,In_139,In_769);
nand U3180 (N_3180,In_845,In_818);
or U3181 (N_3181,In_135,In_943);
and U3182 (N_3182,In_653,In_863);
nor U3183 (N_3183,In_572,In_209);
and U3184 (N_3184,In_464,In_976);
or U3185 (N_3185,In_476,In_748);
and U3186 (N_3186,In_539,In_89);
and U3187 (N_3187,In_393,In_143);
nor U3188 (N_3188,In_757,In_336);
or U3189 (N_3189,In_873,In_913);
and U3190 (N_3190,In_363,In_848);
and U3191 (N_3191,In_220,In_866);
and U3192 (N_3192,In_656,In_810);
nor U3193 (N_3193,In_314,In_744);
nor U3194 (N_3194,In_812,In_979);
and U3195 (N_3195,In_265,In_526);
nor U3196 (N_3196,In_193,In_126);
nand U3197 (N_3197,In_944,In_340);
and U3198 (N_3198,In_252,In_320);
nand U3199 (N_3199,In_673,In_55);
or U3200 (N_3200,In_441,In_990);
or U3201 (N_3201,In_21,In_391);
or U3202 (N_3202,In_990,In_784);
nor U3203 (N_3203,In_970,In_992);
and U3204 (N_3204,In_640,In_367);
nor U3205 (N_3205,In_52,In_91);
and U3206 (N_3206,In_282,In_23);
and U3207 (N_3207,In_759,In_491);
or U3208 (N_3208,In_827,In_376);
nand U3209 (N_3209,In_479,In_920);
nand U3210 (N_3210,In_265,In_538);
nand U3211 (N_3211,In_618,In_247);
nor U3212 (N_3212,In_717,In_777);
nor U3213 (N_3213,In_923,In_616);
nand U3214 (N_3214,In_272,In_302);
nand U3215 (N_3215,In_604,In_799);
nand U3216 (N_3216,In_421,In_796);
or U3217 (N_3217,In_369,In_777);
nand U3218 (N_3218,In_659,In_780);
nand U3219 (N_3219,In_984,In_779);
nand U3220 (N_3220,In_41,In_830);
or U3221 (N_3221,In_696,In_622);
nand U3222 (N_3222,In_360,In_30);
nor U3223 (N_3223,In_313,In_407);
nand U3224 (N_3224,In_319,In_907);
nor U3225 (N_3225,In_658,In_156);
nor U3226 (N_3226,In_547,In_839);
or U3227 (N_3227,In_487,In_471);
xnor U3228 (N_3228,In_398,In_868);
nor U3229 (N_3229,In_454,In_673);
or U3230 (N_3230,In_414,In_14);
nand U3231 (N_3231,In_714,In_540);
and U3232 (N_3232,In_685,In_851);
and U3233 (N_3233,In_790,In_650);
nor U3234 (N_3234,In_151,In_933);
nand U3235 (N_3235,In_425,In_209);
nand U3236 (N_3236,In_189,In_463);
nor U3237 (N_3237,In_757,In_293);
and U3238 (N_3238,In_940,In_502);
nor U3239 (N_3239,In_665,In_834);
or U3240 (N_3240,In_814,In_136);
and U3241 (N_3241,In_95,In_804);
and U3242 (N_3242,In_754,In_783);
nand U3243 (N_3243,In_156,In_338);
or U3244 (N_3244,In_553,In_461);
or U3245 (N_3245,In_996,In_601);
xor U3246 (N_3246,In_112,In_975);
nor U3247 (N_3247,In_400,In_575);
nor U3248 (N_3248,In_323,In_641);
nand U3249 (N_3249,In_265,In_516);
nor U3250 (N_3250,In_73,In_953);
nor U3251 (N_3251,In_50,In_7);
nand U3252 (N_3252,In_629,In_62);
or U3253 (N_3253,In_211,In_742);
or U3254 (N_3254,In_792,In_80);
or U3255 (N_3255,In_84,In_863);
and U3256 (N_3256,In_84,In_101);
or U3257 (N_3257,In_102,In_308);
nand U3258 (N_3258,In_772,In_329);
nor U3259 (N_3259,In_5,In_751);
nor U3260 (N_3260,In_770,In_691);
and U3261 (N_3261,In_468,In_125);
and U3262 (N_3262,In_984,In_558);
nand U3263 (N_3263,In_144,In_595);
nand U3264 (N_3264,In_331,In_510);
nor U3265 (N_3265,In_981,In_610);
nor U3266 (N_3266,In_95,In_370);
nor U3267 (N_3267,In_359,In_645);
and U3268 (N_3268,In_392,In_686);
nor U3269 (N_3269,In_530,In_470);
and U3270 (N_3270,In_194,In_144);
or U3271 (N_3271,In_374,In_448);
nand U3272 (N_3272,In_545,In_44);
or U3273 (N_3273,In_74,In_830);
nor U3274 (N_3274,In_778,In_677);
or U3275 (N_3275,In_479,In_113);
or U3276 (N_3276,In_194,In_318);
nor U3277 (N_3277,In_526,In_814);
nand U3278 (N_3278,In_279,In_432);
or U3279 (N_3279,In_424,In_611);
or U3280 (N_3280,In_223,In_977);
nor U3281 (N_3281,In_21,In_548);
nand U3282 (N_3282,In_817,In_585);
xor U3283 (N_3283,In_134,In_287);
or U3284 (N_3284,In_327,In_965);
nor U3285 (N_3285,In_654,In_848);
or U3286 (N_3286,In_569,In_307);
or U3287 (N_3287,In_924,In_138);
or U3288 (N_3288,In_337,In_207);
or U3289 (N_3289,In_140,In_278);
and U3290 (N_3290,In_887,In_160);
nand U3291 (N_3291,In_941,In_968);
or U3292 (N_3292,In_967,In_185);
nor U3293 (N_3293,In_997,In_884);
or U3294 (N_3294,In_164,In_557);
nand U3295 (N_3295,In_213,In_41);
or U3296 (N_3296,In_600,In_838);
nand U3297 (N_3297,In_480,In_917);
and U3298 (N_3298,In_469,In_981);
and U3299 (N_3299,In_490,In_136);
or U3300 (N_3300,In_9,In_942);
or U3301 (N_3301,In_76,In_884);
nand U3302 (N_3302,In_226,In_208);
and U3303 (N_3303,In_466,In_168);
nor U3304 (N_3304,In_916,In_966);
nor U3305 (N_3305,In_128,In_551);
nor U3306 (N_3306,In_912,In_238);
nor U3307 (N_3307,In_730,In_219);
or U3308 (N_3308,In_578,In_976);
nand U3309 (N_3309,In_863,In_12);
and U3310 (N_3310,In_259,In_70);
and U3311 (N_3311,In_781,In_435);
nand U3312 (N_3312,In_157,In_457);
nor U3313 (N_3313,In_568,In_482);
nor U3314 (N_3314,In_14,In_573);
nand U3315 (N_3315,In_138,In_97);
and U3316 (N_3316,In_691,In_929);
or U3317 (N_3317,In_700,In_528);
nor U3318 (N_3318,In_151,In_514);
or U3319 (N_3319,In_852,In_487);
nor U3320 (N_3320,In_407,In_916);
or U3321 (N_3321,In_946,In_662);
and U3322 (N_3322,In_425,In_463);
or U3323 (N_3323,In_581,In_820);
nor U3324 (N_3324,In_327,In_166);
or U3325 (N_3325,In_444,In_871);
nor U3326 (N_3326,In_76,In_782);
nand U3327 (N_3327,In_434,In_365);
and U3328 (N_3328,In_79,In_767);
xor U3329 (N_3329,In_837,In_701);
and U3330 (N_3330,In_757,In_860);
nor U3331 (N_3331,In_600,In_271);
and U3332 (N_3332,In_959,In_761);
nand U3333 (N_3333,In_769,In_998);
nor U3334 (N_3334,In_497,In_53);
nand U3335 (N_3335,In_99,In_439);
nor U3336 (N_3336,In_865,In_10);
xor U3337 (N_3337,In_6,In_962);
and U3338 (N_3338,In_469,In_423);
and U3339 (N_3339,In_875,In_592);
or U3340 (N_3340,In_815,In_628);
nor U3341 (N_3341,In_406,In_193);
nor U3342 (N_3342,In_79,In_725);
and U3343 (N_3343,In_928,In_868);
nand U3344 (N_3344,In_125,In_680);
and U3345 (N_3345,In_692,In_864);
nor U3346 (N_3346,In_194,In_579);
or U3347 (N_3347,In_608,In_289);
nor U3348 (N_3348,In_844,In_655);
nor U3349 (N_3349,In_36,In_564);
and U3350 (N_3350,In_579,In_36);
and U3351 (N_3351,In_0,In_921);
and U3352 (N_3352,In_390,In_93);
nor U3353 (N_3353,In_765,In_312);
and U3354 (N_3354,In_570,In_282);
nor U3355 (N_3355,In_348,In_254);
nor U3356 (N_3356,In_93,In_996);
nor U3357 (N_3357,In_952,In_855);
and U3358 (N_3358,In_382,In_66);
or U3359 (N_3359,In_858,In_602);
and U3360 (N_3360,In_655,In_865);
nor U3361 (N_3361,In_26,In_898);
or U3362 (N_3362,In_921,In_233);
or U3363 (N_3363,In_460,In_114);
and U3364 (N_3364,In_62,In_623);
nor U3365 (N_3365,In_757,In_690);
nor U3366 (N_3366,In_13,In_123);
nor U3367 (N_3367,In_128,In_792);
and U3368 (N_3368,In_960,In_481);
nor U3369 (N_3369,In_188,In_851);
and U3370 (N_3370,In_174,In_805);
and U3371 (N_3371,In_840,In_349);
nor U3372 (N_3372,In_348,In_52);
nand U3373 (N_3373,In_323,In_252);
nand U3374 (N_3374,In_769,In_32);
or U3375 (N_3375,In_572,In_64);
and U3376 (N_3376,In_838,In_470);
nor U3377 (N_3377,In_994,In_137);
or U3378 (N_3378,In_121,In_411);
xnor U3379 (N_3379,In_560,In_90);
and U3380 (N_3380,In_216,In_203);
nor U3381 (N_3381,In_295,In_813);
or U3382 (N_3382,In_117,In_558);
nor U3383 (N_3383,In_534,In_356);
nor U3384 (N_3384,In_383,In_294);
nor U3385 (N_3385,In_561,In_803);
and U3386 (N_3386,In_322,In_464);
and U3387 (N_3387,In_220,In_439);
and U3388 (N_3388,In_136,In_973);
nor U3389 (N_3389,In_517,In_963);
and U3390 (N_3390,In_328,In_436);
nor U3391 (N_3391,In_433,In_591);
nor U3392 (N_3392,In_395,In_53);
nand U3393 (N_3393,In_379,In_841);
or U3394 (N_3394,In_495,In_757);
and U3395 (N_3395,In_158,In_829);
nand U3396 (N_3396,In_304,In_783);
and U3397 (N_3397,In_962,In_725);
nand U3398 (N_3398,In_338,In_978);
or U3399 (N_3399,In_20,In_793);
and U3400 (N_3400,In_582,In_841);
nand U3401 (N_3401,In_255,In_452);
nand U3402 (N_3402,In_421,In_309);
nor U3403 (N_3403,In_966,In_145);
or U3404 (N_3404,In_576,In_334);
or U3405 (N_3405,In_427,In_380);
or U3406 (N_3406,In_63,In_574);
or U3407 (N_3407,In_376,In_760);
nand U3408 (N_3408,In_719,In_506);
and U3409 (N_3409,In_397,In_716);
and U3410 (N_3410,In_896,In_590);
nand U3411 (N_3411,In_268,In_54);
or U3412 (N_3412,In_52,In_888);
or U3413 (N_3413,In_653,In_43);
or U3414 (N_3414,In_685,In_65);
and U3415 (N_3415,In_154,In_377);
nor U3416 (N_3416,In_618,In_261);
nor U3417 (N_3417,In_695,In_535);
nand U3418 (N_3418,In_291,In_836);
and U3419 (N_3419,In_545,In_986);
nand U3420 (N_3420,In_913,In_848);
nor U3421 (N_3421,In_533,In_782);
or U3422 (N_3422,In_377,In_370);
nand U3423 (N_3423,In_561,In_893);
or U3424 (N_3424,In_530,In_52);
nand U3425 (N_3425,In_807,In_489);
nor U3426 (N_3426,In_406,In_456);
and U3427 (N_3427,In_412,In_943);
or U3428 (N_3428,In_159,In_219);
and U3429 (N_3429,In_453,In_190);
nand U3430 (N_3430,In_738,In_634);
nand U3431 (N_3431,In_406,In_653);
and U3432 (N_3432,In_125,In_585);
or U3433 (N_3433,In_518,In_521);
nand U3434 (N_3434,In_492,In_429);
nand U3435 (N_3435,In_716,In_97);
nor U3436 (N_3436,In_536,In_807);
nor U3437 (N_3437,In_608,In_277);
nor U3438 (N_3438,In_228,In_629);
or U3439 (N_3439,In_523,In_681);
xnor U3440 (N_3440,In_279,In_468);
or U3441 (N_3441,In_124,In_150);
or U3442 (N_3442,In_613,In_549);
and U3443 (N_3443,In_139,In_614);
nor U3444 (N_3444,In_896,In_874);
or U3445 (N_3445,In_361,In_473);
or U3446 (N_3446,In_975,In_137);
nor U3447 (N_3447,In_743,In_330);
or U3448 (N_3448,In_797,In_135);
and U3449 (N_3449,In_787,In_347);
or U3450 (N_3450,In_781,In_906);
or U3451 (N_3451,In_43,In_779);
or U3452 (N_3452,In_13,In_991);
or U3453 (N_3453,In_177,In_579);
and U3454 (N_3454,In_347,In_600);
nor U3455 (N_3455,In_274,In_577);
nor U3456 (N_3456,In_416,In_566);
or U3457 (N_3457,In_307,In_806);
and U3458 (N_3458,In_621,In_469);
nand U3459 (N_3459,In_91,In_613);
nand U3460 (N_3460,In_561,In_954);
xnor U3461 (N_3461,In_511,In_902);
nand U3462 (N_3462,In_974,In_588);
and U3463 (N_3463,In_57,In_393);
nand U3464 (N_3464,In_902,In_667);
nand U3465 (N_3465,In_905,In_120);
or U3466 (N_3466,In_758,In_8);
nand U3467 (N_3467,In_148,In_595);
and U3468 (N_3468,In_404,In_483);
nand U3469 (N_3469,In_229,In_891);
nor U3470 (N_3470,In_330,In_167);
and U3471 (N_3471,In_77,In_243);
nand U3472 (N_3472,In_686,In_829);
or U3473 (N_3473,In_42,In_780);
nand U3474 (N_3474,In_148,In_466);
or U3475 (N_3475,In_173,In_343);
and U3476 (N_3476,In_211,In_72);
or U3477 (N_3477,In_400,In_944);
nor U3478 (N_3478,In_149,In_344);
nand U3479 (N_3479,In_332,In_513);
or U3480 (N_3480,In_907,In_143);
nor U3481 (N_3481,In_891,In_489);
and U3482 (N_3482,In_869,In_619);
or U3483 (N_3483,In_469,In_879);
nand U3484 (N_3484,In_296,In_942);
nor U3485 (N_3485,In_85,In_218);
nand U3486 (N_3486,In_242,In_608);
nor U3487 (N_3487,In_682,In_771);
and U3488 (N_3488,In_53,In_487);
nand U3489 (N_3489,In_692,In_518);
and U3490 (N_3490,In_475,In_770);
nor U3491 (N_3491,In_423,In_432);
or U3492 (N_3492,In_891,In_599);
nand U3493 (N_3493,In_207,In_72);
nand U3494 (N_3494,In_370,In_564);
or U3495 (N_3495,In_520,In_823);
nor U3496 (N_3496,In_132,In_328);
and U3497 (N_3497,In_837,In_327);
nand U3498 (N_3498,In_675,In_433);
nor U3499 (N_3499,In_7,In_181);
nand U3500 (N_3500,In_123,In_298);
and U3501 (N_3501,In_411,In_459);
or U3502 (N_3502,In_30,In_51);
nor U3503 (N_3503,In_9,In_623);
or U3504 (N_3504,In_376,In_781);
and U3505 (N_3505,In_943,In_983);
nand U3506 (N_3506,In_409,In_750);
or U3507 (N_3507,In_184,In_355);
nand U3508 (N_3508,In_508,In_726);
nand U3509 (N_3509,In_620,In_955);
nand U3510 (N_3510,In_457,In_616);
or U3511 (N_3511,In_237,In_984);
or U3512 (N_3512,In_444,In_21);
and U3513 (N_3513,In_189,In_314);
nor U3514 (N_3514,In_13,In_30);
nand U3515 (N_3515,In_733,In_749);
and U3516 (N_3516,In_819,In_366);
nand U3517 (N_3517,In_276,In_861);
or U3518 (N_3518,In_832,In_52);
nand U3519 (N_3519,In_249,In_183);
nand U3520 (N_3520,In_485,In_172);
or U3521 (N_3521,In_46,In_456);
nand U3522 (N_3522,In_676,In_902);
and U3523 (N_3523,In_476,In_255);
xnor U3524 (N_3524,In_638,In_53);
or U3525 (N_3525,In_514,In_277);
and U3526 (N_3526,In_96,In_618);
nor U3527 (N_3527,In_992,In_202);
nand U3528 (N_3528,In_45,In_615);
and U3529 (N_3529,In_557,In_199);
nand U3530 (N_3530,In_847,In_322);
nand U3531 (N_3531,In_932,In_947);
xor U3532 (N_3532,In_901,In_41);
or U3533 (N_3533,In_396,In_453);
nor U3534 (N_3534,In_271,In_730);
and U3535 (N_3535,In_531,In_32);
nor U3536 (N_3536,In_699,In_381);
or U3537 (N_3537,In_172,In_584);
or U3538 (N_3538,In_662,In_57);
nand U3539 (N_3539,In_345,In_217);
and U3540 (N_3540,In_451,In_383);
and U3541 (N_3541,In_910,In_541);
nand U3542 (N_3542,In_529,In_813);
or U3543 (N_3543,In_205,In_386);
nand U3544 (N_3544,In_585,In_21);
and U3545 (N_3545,In_501,In_815);
or U3546 (N_3546,In_623,In_687);
or U3547 (N_3547,In_937,In_152);
or U3548 (N_3548,In_45,In_559);
and U3549 (N_3549,In_611,In_56);
nand U3550 (N_3550,In_330,In_70);
and U3551 (N_3551,In_950,In_940);
nand U3552 (N_3552,In_4,In_974);
and U3553 (N_3553,In_198,In_351);
and U3554 (N_3554,In_174,In_834);
and U3555 (N_3555,In_44,In_16);
and U3556 (N_3556,In_40,In_416);
and U3557 (N_3557,In_988,In_125);
nor U3558 (N_3558,In_281,In_424);
or U3559 (N_3559,In_621,In_492);
nor U3560 (N_3560,In_860,In_330);
nor U3561 (N_3561,In_377,In_206);
nand U3562 (N_3562,In_335,In_859);
and U3563 (N_3563,In_128,In_447);
and U3564 (N_3564,In_909,In_469);
nor U3565 (N_3565,In_670,In_419);
nor U3566 (N_3566,In_345,In_690);
nor U3567 (N_3567,In_446,In_164);
nor U3568 (N_3568,In_483,In_372);
or U3569 (N_3569,In_744,In_969);
nor U3570 (N_3570,In_222,In_919);
or U3571 (N_3571,In_43,In_742);
nor U3572 (N_3572,In_866,In_43);
nand U3573 (N_3573,In_655,In_102);
nor U3574 (N_3574,In_221,In_527);
or U3575 (N_3575,In_437,In_118);
nor U3576 (N_3576,In_174,In_783);
nand U3577 (N_3577,In_186,In_841);
nor U3578 (N_3578,In_199,In_833);
and U3579 (N_3579,In_914,In_606);
nand U3580 (N_3580,In_947,In_731);
nand U3581 (N_3581,In_127,In_945);
or U3582 (N_3582,In_960,In_485);
nor U3583 (N_3583,In_475,In_979);
nor U3584 (N_3584,In_20,In_749);
nand U3585 (N_3585,In_151,In_986);
nor U3586 (N_3586,In_466,In_431);
nor U3587 (N_3587,In_718,In_224);
and U3588 (N_3588,In_659,In_601);
nor U3589 (N_3589,In_381,In_494);
or U3590 (N_3590,In_67,In_348);
nor U3591 (N_3591,In_852,In_904);
nand U3592 (N_3592,In_659,In_475);
or U3593 (N_3593,In_627,In_667);
nand U3594 (N_3594,In_567,In_359);
and U3595 (N_3595,In_73,In_719);
or U3596 (N_3596,In_271,In_375);
or U3597 (N_3597,In_801,In_539);
and U3598 (N_3598,In_856,In_42);
and U3599 (N_3599,In_769,In_737);
and U3600 (N_3600,In_526,In_456);
nor U3601 (N_3601,In_747,In_902);
and U3602 (N_3602,In_99,In_844);
nor U3603 (N_3603,In_470,In_57);
nand U3604 (N_3604,In_250,In_195);
nand U3605 (N_3605,In_793,In_463);
nor U3606 (N_3606,In_920,In_581);
nor U3607 (N_3607,In_377,In_478);
nand U3608 (N_3608,In_45,In_402);
or U3609 (N_3609,In_5,In_967);
and U3610 (N_3610,In_608,In_838);
nor U3611 (N_3611,In_811,In_491);
nand U3612 (N_3612,In_274,In_544);
nand U3613 (N_3613,In_386,In_556);
nand U3614 (N_3614,In_454,In_892);
nand U3615 (N_3615,In_365,In_672);
xnor U3616 (N_3616,In_350,In_221);
or U3617 (N_3617,In_365,In_213);
or U3618 (N_3618,In_109,In_729);
and U3619 (N_3619,In_341,In_601);
nand U3620 (N_3620,In_625,In_873);
nor U3621 (N_3621,In_98,In_210);
nor U3622 (N_3622,In_360,In_322);
nand U3623 (N_3623,In_577,In_455);
or U3624 (N_3624,In_279,In_570);
and U3625 (N_3625,In_137,In_801);
nor U3626 (N_3626,In_95,In_857);
nor U3627 (N_3627,In_109,In_665);
or U3628 (N_3628,In_475,In_210);
nor U3629 (N_3629,In_232,In_712);
and U3630 (N_3630,In_483,In_423);
and U3631 (N_3631,In_24,In_109);
and U3632 (N_3632,In_422,In_774);
and U3633 (N_3633,In_492,In_728);
or U3634 (N_3634,In_894,In_811);
nand U3635 (N_3635,In_888,In_466);
nand U3636 (N_3636,In_537,In_804);
or U3637 (N_3637,In_339,In_677);
nand U3638 (N_3638,In_986,In_195);
or U3639 (N_3639,In_269,In_684);
nand U3640 (N_3640,In_152,In_286);
nor U3641 (N_3641,In_982,In_547);
or U3642 (N_3642,In_473,In_944);
nor U3643 (N_3643,In_419,In_229);
nor U3644 (N_3644,In_243,In_606);
nand U3645 (N_3645,In_744,In_113);
and U3646 (N_3646,In_795,In_658);
nand U3647 (N_3647,In_801,In_848);
or U3648 (N_3648,In_634,In_786);
and U3649 (N_3649,In_947,In_197);
nand U3650 (N_3650,In_205,In_501);
nand U3651 (N_3651,In_320,In_56);
nor U3652 (N_3652,In_550,In_225);
xor U3653 (N_3653,In_625,In_327);
xor U3654 (N_3654,In_592,In_616);
nand U3655 (N_3655,In_486,In_642);
nor U3656 (N_3656,In_442,In_390);
nand U3657 (N_3657,In_271,In_834);
nand U3658 (N_3658,In_499,In_219);
and U3659 (N_3659,In_326,In_186);
and U3660 (N_3660,In_480,In_700);
nand U3661 (N_3661,In_378,In_710);
nor U3662 (N_3662,In_522,In_49);
and U3663 (N_3663,In_401,In_719);
nor U3664 (N_3664,In_517,In_532);
nor U3665 (N_3665,In_746,In_848);
nand U3666 (N_3666,In_51,In_437);
and U3667 (N_3667,In_399,In_137);
nor U3668 (N_3668,In_757,In_770);
nor U3669 (N_3669,In_492,In_776);
nor U3670 (N_3670,In_14,In_143);
or U3671 (N_3671,In_264,In_457);
nor U3672 (N_3672,In_531,In_397);
or U3673 (N_3673,In_178,In_381);
nand U3674 (N_3674,In_214,In_370);
and U3675 (N_3675,In_479,In_558);
nand U3676 (N_3676,In_654,In_158);
and U3677 (N_3677,In_619,In_349);
nand U3678 (N_3678,In_303,In_196);
nand U3679 (N_3679,In_428,In_14);
nand U3680 (N_3680,In_387,In_394);
or U3681 (N_3681,In_746,In_424);
and U3682 (N_3682,In_408,In_853);
nor U3683 (N_3683,In_338,In_906);
or U3684 (N_3684,In_636,In_898);
nor U3685 (N_3685,In_357,In_867);
nor U3686 (N_3686,In_723,In_213);
nor U3687 (N_3687,In_12,In_927);
xor U3688 (N_3688,In_967,In_845);
and U3689 (N_3689,In_293,In_516);
nand U3690 (N_3690,In_562,In_270);
nand U3691 (N_3691,In_266,In_126);
nand U3692 (N_3692,In_256,In_953);
and U3693 (N_3693,In_289,In_692);
nor U3694 (N_3694,In_138,In_510);
and U3695 (N_3695,In_116,In_318);
nor U3696 (N_3696,In_108,In_48);
nor U3697 (N_3697,In_732,In_935);
nand U3698 (N_3698,In_488,In_104);
or U3699 (N_3699,In_601,In_489);
and U3700 (N_3700,In_643,In_908);
or U3701 (N_3701,In_830,In_588);
and U3702 (N_3702,In_614,In_682);
nor U3703 (N_3703,In_531,In_398);
nor U3704 (N_3704,In_821,In_351);
and U3705 (N_3705,In_170,In_481);
and U3706 (N_3706,In_354,In_393);
nor U3707 (N_3707,In_94,In_966);
nor U3708 (N_3708,In_717,In_315);
nand U3709 (N_3709,In_972,In_999);
and U3710 (N_3710,In_500,In_454);
or U3711 (N_3711,In_287,In_868);
and U3712 (N_3712,In_33,In_447);
or U3713 (N_3713,In_438,In_601);
or U3714 (N_3714,In_491,In_328);
nand U3715 (N_3715,In_773,In_361);
xnor U3716 (N_3716,In_561,In_457);
nand U3717 (N_3717,In_326,In_605);
nand U3718 (N_3718,In_481,In_566);
nor U3719 (N_3719,In_881,In_488);
nor U3720 (N_3720,In_610,In_455);
nor U3721 (N_3721,In_789,In_836);
and U3722 (N_3722,In_622,In_185);
or U3723 (N_3723,In_47,In_452);
and U3724 (N_3724,In_827,In_125);
or U3725 (N_3725,In_797,In_833);
or U3726 (N_3726,In_387,In_337);
and U3727 (N_3727,In_327,In_707);
nand U3728 (N_3728,In_780,In_36);
nor U3729 (N_3729,In_509,In_443);
and U3730 (N_3730,In_43,In_821);
or U3731 (N_3731,In_128,In_280);
or U3732 (N_3732,In_845,In_595);
nor U3733 (N_3733,In_744,In_830);
or U3734 (N_3734,In_973,In_443);
nand U3735 (N_3735,In_418,In_656);
or U3736 (N_3736,In_979,In_454);
and U3737 (N_3737,In_27,In_723);
nand U3738 (N_3738,In_294,In_532);
nand U3739 (N_3739,In_175,In_957);
and U3740 (N_3740,In_168,In_443);
nor U3741 (N_3741,In_461,In_475);
and U3742 (N_3742,In_442,In_662);
or U3743 (N_3743,In_882,In_672);
nor U3744 (N_3744,In_583,In_856);
or U3745 (N_3745,In_459,In_119);
and U3746 (N_3746,In_20,In_356);
and U3747 (N_3747,In_256,In_480);
or U3748 (N_3748,In_21,In_212);
and U3749 (N_3749,In_678,In_734);
nor U3750 (N_3750,In_66,In_207);
nand U3751 (N_3751,In_251,In_60);
nor U3752 (N_3752,In_751,In_579);
or U3753 (N_3753,In_166,In_960);
xor U3754 (N_3754,In_959,In_256);
and U3755 (N_3755,In_239,In_615);
and U3756 (N_3756,In_705,In_410);
nor U3757 (N_3757,In_793,In_762);
and U3758 (N_3758,In_921,In_420);
or U3759 (N_3759,In_278,In_234);
nand U3760 (N_3760,In_473,In_935);
nor U3761 (N_3761,In_116,In_829);
nand U3762 (N_3762,In_18,In_715);
nand U3763 (N_3763,In_931,In_175);
nand U3764 (N_3764,In_401,In_464);
and U3765 (N_3765,In_147,In_282);
and U3766 (N_3766,In_271,In_294);
and U3767 (N_3767,In_276,In_630);
nor U3768 (N_3768,In_138,In_765);
or U3769 (N_3769,In_136,In_132);
nor U3770 (N_3770,In_337,In_898);
nor U3771 (N_3771,In_249,In_13);
nor U3772 (N_3772,In_302,In_953);
or U3773 (N_3773,In_277,In_212);
or U3774 (N_3774,In_972,In_660);
or U3775 (N_3775,In_976,In_132);
nand U3776 (N_3776,In_40,In_594);
or U3777 (N_3777,In_674,In_220);
nor U3778 (N_3778,In_192,In_137);
nand U3779 (N_3779,In_928,In_855);
nor U3780 (N_3780,In_175,In_883);
nor U3781 (N_3781,In_918,In_358);
nand U3782 (N_3782,In_859,In_383);
and U3783 (N_3783,In_922,In_88);
and U3784 (N_3784,In_404,In_529);
and U3785 (N_3785,In_49,In_205);
nor U3786 (N_3786,In_424,In_994);
xnor U3787 (N_3787,In_27,In_331);
and U3788 (N_3788,In_579,In_798);
xor U3789 (N_3789,In_894,In_983);
nand U3790 (N_3790,In_471,In_420);
and U3791 (N_3791,In_921,In_663);
and U3792 (N_3792,In_779,In_673);
or U3793 (N_3793,In_768,In_790);
nor U3794 (N_3794,In_734,In_846);
xor U3795 (N_3795,In_965,In_929);
nand U3796 (N_3796,In_723,In_183);
nor U3797 (N_3797,In_322,In_264);
nor U3798 (N_3798,In_314,In_433);
nand U3799 (N_3799,In_606,In_601);
and U3800 (N_3800,In_455,In_474);
and U3801 (N_3801,In_934,In_131);
nand U3802 (N_3802,In_160,In_655);
nand U3803 (N_3803,In_729,In_702);
and U3804 (N_3804,In_554,In_673);
or U3805 (N_3805,In_906,In_7);
or U3806 (N_3806,In_60,In_263);
nor U3807 (N_3807,In_164,In_493);
nand U3808 (N_3808,In_499,In_414);
nand U3809 (N_3809,In_623,In_862);
and U3810 (N_3810,In_116,In_17);
nor U3811 (N_3811,In_524,In_346);
and U3812 (N_3812,In_957,In_856);
nor U3813 (N_3813,In_656,In_239);
xnor U3814 (N_3814,In_204,In_221);
or U3815 (N_3815,In_454,In_394);
nand U3816 (N_3816,In_403,In_770);
or U3817 (N_3817,In_615,In_658);
and U3818 (N_3818,In_447,In_844);
or U3819 (N_3819,In_506,In_858);
or U3820 (N_3820,In_59,In_539);
nand U3821 (N_3821,In_242,In_238);
nor U3822 (N_3822,In_462,In_292);
nor U3823 (N_3823,In_14,In_953);
nand U3824 (N_3824,In_731,In_812);
nand U3825 (N_3825,In_767,In_340);
nand U3826 (N_3826,In_39,In_990);
nor U3827 (N_3827,In_295,In_982);
nor U3828 (N_3828,In_69,In_711);
nor U3829 (N_3829,In_929,In_480);
nand U3830 (N_3830,In_51,In_886);
or U3831 (N_3831,In_640,In_628);
nor U3832 (N_3832,In_890,In_287);
nand U3833 (N_3833,In_740,In_772);
nand U3834 (N_3834,In_145,In_603);
xnor U3835 (N_3835,In_757,In_318);
nand U3836 (N_3836,In_989,In_389);
nand U3837 (N_3837,In_471,In_479);
nor U3838 (N_3838,In_346,In_156);
nand U3839 (N_3839,In_146,In_835);
or U3840 (N_3840,In_566,In_552);
nand U3841 (N_3841,In_940,In_602);
and U3842 (N_3842,In_237,In_915);
nand U3843 (N_3843,In_486,In_118);
and U3844 (N_3844,In_291,In_46);
and U3845 (N_3845,In_153,In_66);
nand U3846 (N_3846,In_872,In_121);
nor U3847 (N_3847,In_204,In_906);
and U3848 (N_3848,In_241,In_34);
nor U3849 (N_3849,In_130,In_118);
nor U3850 (N_3850,In_999,In_123);
or U3851 (N_3851,In_598,In_593);
nor U3852 (N_3852,In_46,In_731);
nand U3853 (N_3853,In_195,In_590);
or U3854 (N_3854,In_158,In_184);
nor U3855 (N_3855,In_339,In_92);
and U3856 (N_3856,In_236,In_622);
or U3857 (N_3857,In_728,In_990);
nor U3858 (N_3858,In_266,In_392);
nand U3859 (N_3859,In_362,In_527);
nand U3860 (N_3860,In_344,In_266);
or U3861 (N_3861,In_775,In_888);
or U3862 (N_3862,In_996,In_605);
nor U3863 (N_3863,In_91,In_942);
and U3864 (N_3864,In_640,In_509);
or U3865 (N_3865,In_119,In_58);
or U3866 (N_3866,In_542,In_75);
nand U3867 (N_3867,In_883,In_984);
and U3868 (N_3868,In_930,In_276);
nand U3869 (N_3869,In_429,In_760);
and U3870 (N_3870,In_331,In_100);
nor U3871 (N_3871,In_892,In_25);
nor U3872 (N_3872,In_156,In_95);
and U3873 (N_3873,In_507,In_937);
nand U3874 (N_3874,In_327,In_793);
nand U3875 (N_3875,In_69,In_935);
nand U3876 (N_3876,In_423,In_349);
nor U3877 (N_3877,In_944,In_517);
and U3878 (N_3878,In_662,In_212);
and U3879 (N_3879,In_182,In_752);
and U3880 (N_3880,In_610,In_906);
nand U3881 (N_3881,In_210,In_753);
and U3882 (N_3882,In_904,In_282);
nand U3883 (N_3883,In_780,In_237);
nor U3884 (N_3884,In_268,In_963);
nand U3885 (N_3885,In_398,In_649);
nand U3886 (N_3886,In_164,In_988);
xor U3887 (N_3887,In_878,In_976);
nor U3888 (N_3888,In_889,In_397);
and U3889 (N_3889,In_942,In_882);
nand U3890 (N_3890,In_397,In_570);
and U3891 (N_3891,In_686,In_350);
or U3892 (N_3892,In_412,In_985);
nand U3893 (N_3893,In_480,In_406);
or U3894 (N_3894,In_344,In_12);
xor U3895 (N_3895,In_484,In_790);
nand U3896 (N_3896,In_358,In_491);
and U3897 (N_3897,In_376,In_805);
and U3898 (N_3898,In_279,In_228);
and U3899 (N_3899,In_376,In_968);
and U3900 (N_3900,In_835,In_100);
and U3901 (N_3901,In_146,In_614);
or U3902 (N_3902,In_395,In_598);
nor U3903 (N_3903,In_525,In_354);
nor U3904 (N_3904,In_502,In_856);
or U3905 (N_3905,In_886,In_905);
or U3906 (N_3906,In_902,In_736);
and U3907 (N_3907,In_316,In_699);
nor U3908 (N_3908,In_823,In_944);
and U3909 (N_3909,In_289,In_567);
or U3910 (N_3910,In_144,In_432);
and U3911 (N_3911,In_740,In_155);
nand U3912 (N_3912,In_284,In_119);
nand U3913 (N_3913,In_601,In_635);
or U3914 (N_3914,In_864,In_253);
or U3915 (N_3915,In_404,In_23);
and U3916 (N_3916,In_576,In_154);
nand U3917 (N_3917,In_959,In_617);
nand U3918 (N_3918,In_691,In_942);
xor U3919 (N_3919,In_931,In_300);
nor U3920 (N_3920,In_578,In_161);
and U3921 (N_3921,In_95,In_299);
nor U3922 (N_3922,In_486,In_954);
or U3923 (N_3923,In_811,In_391);
or U3924 (N_3924,In_716,In_139);
or U3925 (N_3925,In_379,In_627);
or U3926 (N_3926,In_30,In_780);
and U3927 (N_3927,In_740,In_343);
and U3928 (N_3928,In_173,In_5);
xor U3929 (N_3929,In_62,In_956);
or U3930 (N_3930,In_111,In_449);
or U3931 (N_3931,In_827,In_134);
or U3932 (N_3932,In_106,In_927);
nor U3933 (N_3933,In_757,In_65);
nor U3934 (N_3934,In_927,In_226);
nand U3935 (N_3935,In_252,In_169);
or U3936 (N_3936,In_365,In_125);
nor U3937 (N_3937,In_748,In_263);
or U3938 (N_3938,In_617,In_264);
nand U3939 (N_3939,In_943,In_931);
and U3940 (N_3940,In_91,In_768);
nor U3941 (N_3941,In_654,In_262);
or U3942 (N_3942,In_734,In_589);
or U3943 (N_3943,In_962,In_618);
nand U3944 (N_3944,In_170,In_832);
nand U3945 (N_3945,In_227,In_873);
or U3946 (N_3946,In_790,In_562);
nor U3947 (N_3947,In_232,In_102);
and U3948 (N_3948,In_588,In_481);
nand U3949 (N_3949,In_895,In_320);
or U3950 (N_3950,In_925,In_201);
nand U3951 (N_3951,In_569,In_86);
nand U3952 (N_3952,In_716,In_435);
or U3953 (N_3953,In_20,In_571);
or U3954 (N_3954,In_987,In_373);
and U3955 (N_3955,In_410,In_814);
xor U3956 (N_3956,In_300,In_3);
xor U3957 (N_3957,In_663,In_47);
nor U3958 (N_3958,In_720,In_276);
nor U3959 (N_3959,In_271,In_424);
nand U3960 (N_3960,In_112,In_617);
nand U3961 (N_3961,In_742,In_514);
xnor U3962 (N_3962,In_318,In_633);
and U3963 (N_3963,In_367,In_514);
nand U3964 (N_3964,In_702,In_484);
nand U3965 (N_3965,In_803,In_89);
nor U3966 (N_3966,In_793,In_230);
or U3967 (N_3967,In_4,In_261);
nor U3968 (N_3968,In_101,In_774);
and U3969 (N_3969,In_333,In_107);
nand U3970 (N_3970,In_413,In_727);
nand U3971 (N_3971,In_76,In_805);
or U3972 (N_3972,In_231,In_142);
nand U3973 (N_3973,In_156,In_86);
or U3974 (N_3974,In_594,In_215);
and U3975 (N_3975,In_878,In_681);
nor U3976 (N_3976,In_128,In_190);
xnor U3977 (N_3977,In_572,In_416);
and U3978 (N_3978,In_770,In_18);
nor U3979 (N_3979,In_482,In_571);
nand U3980 (N_3980,In_293,In_943);
and U3981 (N_3981,In_625,In_582);
nor U3982 (N_3982,In_238,In_450);
nand U3983 (N_3983,In_675,In_930);
nor U3984 (N_3984,In_363,In_495);
and U3985 (N_3985,In_613,In_979);
and U3986 (N_3986,In_601,In_454);
or U3987 (N_3987,In_661,In_980);
and U3988 (N_3988,In_50,In_582);
nand U3989 (N_3989,In_701,In_628);
nand U3990 (N_3990,In_675,In_649);
and U3991 (N_3991,In_888,In_974);
nor U3992 (N_3992,In_949,In_507);
nor U3993 (N_3993,In_879,In_608);
nor U3994 (N_3994,In_41,In_997);
or U3995 (N_3995,In_599,In_865);
or U3996 (N_3996,In_799,In_281);
nor U3997 (N_3997,In_914,In_38);
nand U3998 (N_3998,In_781,In_236);
nor U3999 (N_3999,In_117,In_582);
xnor U4000 (N_4000,In_818,In_339);
nor U4001 (N_4001,In_946,In_964);
and U4002 (N_4002,In_895,In_195);
and U4003 (N_4003,In_851,In_493);
and U4004 (N_4004,In_643,In_160);
nand U4005 (N_4005,In_574,In_418);
or U4006 (N_4006,In_109,In_105);
or U4007 (N_4007,In_272,In_642);
nand U4008 (N_4008,In_357,In_226);
nand U4009 (N_4009,In_705,In_169);
nand U4010 (N_4010,In_187,In_335);
or U4011 (N_4011,In_402,In_557);
nand U4012 (N_4012,In_261,In_574);
and U4013 (N_4013,In_707,In_454);
nor U4014 (N_4014,In_30,In_31);
or U4015 (N_4015,In_783,In_386);
nand U4016 (N_4016,In_649,In_898);
or U4017 (N_4017,In_747,In_570);
xor U4018 (N_4018,In_36,In_379);
nand U4019 (N_4019,In_547,In_603);
and U4020 (N_4020,In_654,In_37);
and U4021 (N_4021,In_269,In_333);
and U4022 (N_4022,In_935,In_454);
and U4023 (N_4023,In_910,In_873);
or U4024 (N_4024,In_605,In_484);
nand U4025 (N_4025,In_835,In_989);
and U4026 (N_4026,In_429,In_245);
or U4027 (N_4027,In_198,In_709);
and U4028 (N_4028,In_790,In_12);
or U4029 (N_4029,In_401,In_462);
or U4030 (N_4030,In_279,In_755);
nand U4031 (N_4031,In_546,In_748);
nor U4032 (N_4032,In_882,In_243);
and U4033 (N_4033,In_437,In_507);
and U4034 (N_4034,In_807,In_777);
nand U4035 (N_4035,In_222,In_586);
nor U4036 (N_4036,In_506,In_301);
nand U4037 (N_4037,In_480,In_782);
and U4038 (N_4038,In_111,In_777);
nor U4039 (N_4039,In_271,In_950);
nor U4040 (N_4040,In_585,In_906);
and U4041 (N_4041,In_145,In_508);
nand U4042 (N_4042,In_396,In_821);
and U4043 (N_4043,In_854,In_104);
nor U4044 (N_4044,In_847,In_325);
nor U4045 (N_4045,In_685,In_227);
nor U4046 (N_4046,In_580,In_243);
nor U4047 (N_4047,In_835,In_673);
and U4048 (N_4048,In_216,In_365);
nor U4049 (N_4049,In_111,In_723);
and U4050 (N_4050,In_739,In_843);
and U4051 (N_4051,In_296,In_769);
xnor U4052 (N_4052,In_520,In_184);
nand U4053 (N_4053,In_126,In_698);
nand U4054 (N_4054,In_4,In_721);
nor U4055 (N_4055,In_656,In_806);
nand U4056 (N_4056,In_493,In_21);
or U4057 (N_4057,In_622,In_938);
or U4058 (N_4058,In_875,In_191);
and U4059 (N_4059,In_511,In_900);
nand U4060 (N_4060,In_957,In_253);
or U4061 (N_4061,In_25,In_320);
and U4062 (N_4062,In_791,In_450);
and U4063 (N_4063,In_868,In_686);
and U4064 (N_4064,In_335,In_662);
nor U4065 (N_4065,In_246,In_623);
nand U4066 (N_4066,In_636,In_515);
nand U4067 (N_4067,In_576,In_728);
or U4068 (N_4068,In_694,In_254);
nand U4069 (N_4069,In_640,In_544);
and U4070 (N_4070,In_188,In_754);
xor U4071 (N_4071,In_356,In_680);
nand U4072 (N_4072,In_725,In_431);
or U4073 (N_4073,In_533,In_317);
and U4074 (N_4074,In_11,In_367);
and U4075 (N_4075,In_597,In_516);
or U4076 (N_4076,In_467,In_100);
and U4077 (N_4077,In_877,In_158);
nand U4078 (N_4078,In_330,In_336);
or U4079 (N_4079,In_469,In_143);
nor U4080 (N_4080,In_783,In_638);
or U4081 (N_4081,In_250,In_965);
or U4082 (N_4082,In_357,In_377);
nand U4083 (N_4083,In_170,In_831);
nand U4084 (N_4084,In_176,In_303);
and U4085 (N_4085,In_558,In_326);
or U4086 (N_4086,In_319,In_134);
nand U4087 (N_4087,In_851,In_839);
nand U4088 (N_4088,In_868,In_69);
nand U4089 (N_4089,In_730,In_448);
or U4090 (N_4090,In_890,In_552);
or U4091 (N_4091,In_31,In_541);
and U4092 (N_4092,In_505,In_699);
nand U4093 (N_4093,In_937,In_686);
nor U4094 (N_4094,In_560,In_529);
nor U4095 (N_4095,In_605,In_135);
nor U4096 (N_4096,In_687,In_285);
and U4097 (N_4097,In_169,In_517);
nor U4098 (N_4098,In_229,In_629);
nor U4099 (N_4099,In_595,In_245);
or U4100 (N_4100,In_584,In_743);
xor U4101 (N_4101,In_661,In_984);
or U4102 (N_4102,In_295,In_425);
or U4103 (N_4103,In_694,In_620);
nand U4104 (N_4104,In_915,In_163);
xnor U4105 (N_4105,In_955,In_865);
nor U4106 (N_4106,In_651,In_21);
and U4107 (N_4107,In_196,In_202);
and U4108 (N_4108,In_194,In_42);
and U4109 (N_4109,In_426,In_851);
and U4110 (N_4110,In_223,In_749);
and U4111 (N_4111,In_610,In_282);
and U4112 (N_4112,In_929,In_194);
nand U4113 (N_4113,In_635,In_456);
nor U4114 (N_4114,In_12,In_768);
or U4115 (N_4115,In_291,In_87);
nor U4116 (N_4116,In_869,In_205);
and U4117 (N_4117,In_879,In_954);
and U4118 (N_4118,In_71,In_982);
nand U4119 (N_4119,In_539,In_647);
nor U4120 (N_4120,In_413,In_427);
and U4121 (N_4121,In_156,In_347);
or U4122 (N_4122,In_402,In_550);
or U4123 (N_4123,In_942,In_728);
nand U4124 (N_4124,In_560,In_726);
or U4125 (N_4125,In_519,In_874);
and U4126 (N_4126,In_833,In_12);
nor U4127 (N_4127,In_174,In_261);
nand U4128 (N_4128,In_23,In_493);
nand U4129 (N_4129,In_768,In_362);
and U4130 (N_4130,In_324,In_100);
or U4131 (N_4131,In_656,In_328);
nand U4132 (N_4132,In_174,In_845);
nand U4133 (N_4133,In_60,In_138);
or U4134 (N_4134,In_443,In_595);
xor U4135 (N_4135,In_513,In_161);
or U4136 (N_4136,In_390,In_995);
and U4137 (N_4137,In_321,In_47);
nor U4138 (N_4138,In_987,In_572);
nor U4139 (N_4139,In_989,In_946);
xor U4140 (N_4140,In_941,In_489);
nor U4141 (N_4141,In_226,In_907);
nand U4142 (N_4142,In_85,In_954);
nor U4143 (N_4143,In_244,In_863);
nor U4144 (N_4144,In_412,In_971);
nand U4145 (N_4145,In_623,In_136);
nand U4146 (N_4146,In_989,In_478);
nand U4147 (N_4147,In_580,In_702);
nor U4148 (N_4148,In_154,In_232);
nand U4149 (N_4149,In_802,In_178);
nand U4150 (N_4150,In_720,In_489);
nand U4151 (N_4151,In_159,In_357);
nor U4152 (N_4152,In_654,In_356);
or U4153 (N_4153,In_174,In_746);
and U4154 (N_4154,In_632,In_227);
nand U4155 (N_4155,In_831,In_889);
and U4156 (N_4156,In_429,In_501);
nor U4157 (N_4157,In_131,In_796);
nand U4158 (N_4158,In_735,In_201);
nor U4159 (N_4159,In_296,In_275);
or U4160 (N_4160,In_709,In_913);
nor U4161 (N_4161,In_299,In_422);
nand U4162 (N_4162,In_437,In_347);
nand U4163 (N_4163,In_394,In_479);
nand U4164 (N_4164,In_606,In_685);
nor U4165 (N_4165,In_382,In_928);
and U4166 (N_4166,In_616,In_856);
nor U4167 (N_4167,In_695,In_45);
and U4168 (N_4168,In_53,In_144);
or U4169 (N_4169,In_382,In_349);
or U4170 (N_4170,In_726,In_604);
and U4171 (N_4171,In_81,In_505);
or U4172 (N_4172,In_746,In_471);
nor U4173 (N_4173,In_790,In_644);
nor U4174 (N_4174,In_721,In_115);
nand U4175 (N_4175,In_807,In_635);
or U4176 (N_4176,In_881,In_166);
nand U4177 (N_4177,In_472,In_814);
nand U4178 (N_4178,In_983,In_573);
and U4179 (N_4179,In_290,In_874);
nor U4180 (N_4180,In_228,In_18);
nor U4181 (N_4181,In_148,In_886);
or U4182 (N_4182,In_668,In_688);
nor U4183 (N_4183,In_943,In_148);
or U4184 (N_4184,In_308,In_196);
and U4185 (N_4185,In_900,In_292);
or U4186 (N_4186,In_589,In_967);
and U4187 (N_4187,In_379,In_550);
or U4188 (N_4188,In_306,In_61);
nor U4189 (N_4189,In_761,In_834);
or U4190 (N_4190,In_672,In_998);
or U4191 (N_4191,In_936,In_882);
and U4192 (N_4192,In_140,In_143);
or U4193 (N_4193,In_158,In_503);
nor U4194 (N_4194,In_622,In_153);
or U4195 (N_4195,In_715,In_141);
and U4196 (N_4196,In_675,In_355);
and U4197 (N_4197,In_466,In_693);
nor U4198 (N_4198,In_107,In_131);
and U4199 (N_4199,In_344,In_494);
nand U4200 (N_4200,In_472,In_931);
nor U4201 (N_4201,In_382,In_683);
nand U4202 (N_4202,In_918,In_0);
xor U4203 (N_4203,In_725,In_786);
nor U4204 (N_4204,In_975,In_384);
nor U4205 (N_4205,In_595,In_312);
and U4206 (N_4206,In_568,In_938);
nor U4207 (N_4207,In_301,In_703);
nor U4208 (N_4208,In_432,In_632);
or U4209 (N_4209,In_388,In_467);
nand U4210 (N_4210,In_683,In_809);
xnor U4211 (N_4211,In_96,In_402);
nor U4212 (N_4212,In_399,In_377);
nand U4213 (N_4213,In_724,In_248);
nand U4214 (N_4214,In_600,In_318);
nor U4215 (N_4215,In_805,In_876);
or U4216 (N_4216,In_537,In_704);
or U4217 (N_4217,In_607,In_316);
nand U4218 (N_4218,In_862,In_481);
nand U4219 (N_4219,In_213,In_496);
or U4220 (N_4220,In_500,In_831);
or U4221 (N_4221,In_287,In_29);
nand U4222 (N_4222,In_623,In_636);
xor U4223 (N_4223,In_293,In_688);
nor U4224 (N_4224,In_530,In_380);
nand U4225 (N_4225,In_143,In_646);
nand U4226 (N_4226,In_402,In_222);
and U4227 (N_4227,In_906,In_41);
nand U4228 (N_4228,In_551,In_894);
nand U4229 (N_4229,In_4,In_353);
nor U4230 (N_4230,In_258,In_67);
and U4231 (N_4231,In_971,In_959);
and U4232 (N_4232,In_32,In_186);
nand U4233 (N_4233,In_453,In_449);
or U4234 (N_4234,In_949,In_5);
nor U4235 (N_4235,In_126,In_168);
nor U4236 (N_4236,In_57,In_451);
or U4237 (N_4237,In_528,In_227);
nand U4238 (N_4238,In_848,In_166);
nand U4239 (N_4239,In_715,In_509);
nand U4240 (N_4240,In_701,In_303);
or U4241 (N_4241,In_111,In_492);
or U4242 (N_4242,In_354,In_447);
or U4243 (N_4243,In_163,In_233);
nor U4244 (N_4244,In_454,In_148);
and U4245 (N_4245,In_335,In_280);
nand U4246 (N_4246,In_786,In_877);
nor U4247 (N_4247,In_107,In_228);
nand U4248 (N_4248,In_185,In_660);
and U4249 (N_4249,In_706,In_104);
and U4250 (N_4250,In_608,In_297);
nor U4251 (N_4251,In_960,In_226);
or U4252 (N_4252,In_451,In_710);
and U4253 (N_4253,In_284,In_855);
nor U4254 (N_4254,In_407,In_343);
nand U4255 (N_4255,In_459,In_945);
and U4256 (N_4256,In_60,In_912);
nor U4257 (N_4257,In_958,In_34);
or U4258 (N_4258,In_155,In_145);
or U4259 (N_4259,In_430,In_779);
or U4260 (N_4260,In_863,In_327);
nand U4261 (N_4261,In_612,In_123);
and U4262 (N_4262,In_406,In_82);
nor U4263 (N_4263,In_632,In_858);
and U4264 (N_4264,In_32,In_95);
nand U4265 (N_4265,In_807,In_936);
or U4266 (N_4266,In_625,In_627);
or U4267 (N_4267,In_344,In_946);
or U4268 (N_4268,In_762,In_270);
or U4269 (N_4269,In_898,In_846);
or U4270 (N_4270,In_149,In_105);
nor U4271 (N_4271,In_128,In_592);
nand U4272 (N_4272,In_272,In_105);
or U4273 (N_4273,In_980,In_398);
or U4274 (N_4274,In_304,In_203);
and U4275 (N_4275,In_844,In_618);
nor U4276 (N_4276,In_493,In_168);
nor U4277 (N_4277,In_133,In_900);
or U4278 (N_4278,In_768,In_880);
nor U4279 (N_4279,In_753,In_764);
nand U4280 (N_4280,In_574,In_374);
nor U4281 (N_4281,In_43,In_296);
or U4282 (N_4282,In_645,In_819);
nor U4283 (N_4283,In_925,In_581);
and U4284 (N_4284,In_849,In_833);
nor U4285 (N_4285,In_283,In_642);
nand U4286 (N_4286,In_575,In_100);
nand U4287 (N_4287,In_265,In_309);
nor U4288 (N_4288,In_497,In_492);
or U4289 (N_4289,In_730,In_790);
nand U4290 (N_4290,In_981,In_779);
nor U4291 (N_4291,In_773,In_777);
nor U4292 (N_4292,In_129,In_236);
and U4293 (N_4293,In_928,In_991);
and U4294 (N_4294,In_196,In_136);
and U4295 (N_4295,In_422,In_761);
nor U4296 (N_4296,In_682,In_163);
nor U4297 (N_4297,In_870,In_936);
and U4298 (N_4298,In_626,In_394);
or U4299 (N_4299,In_595,In_741);
or U4300 (N_4300,In_340,In_539);
nor U4301 (N_4301,In_102,In_556);
and U4302 (N_4302,In_197,In_345);
nor U4303 (N_4303,In_508,In_200);
and U4304 (N_4304,In_379,In_922);
or U4305 (N_4305,In_491,In_865);
nand U4306 (N_4306,In_362,In_699);
and U4307 (N_4307,In_344,In_857);
or U4308 (N_4308,In_528,In_840);
and U4309 (N_4309,In_784,In_737);
xor U4310 (N_4310,In_172,In_144);
or U4311 (N_4311,In_234,In_777);
or U4312 (N_4312,In_672,In_880);
or U4313 (N_4313,In_207,In_399);
nor U4314 (N_4314,In_703,In_9);
nand U4315 (N_4315,In_945,In_658);
nor U4316 (N_4316,In_144,In_503);
nor U4317 (N_4317,In_471,In_67);
and U4318 (N_4318,In_462,In_968);
or U4319 (N_4319,In_583,In_600);
nand U4320 (N_4320,In_119,In_839);
or U4321 (N_4321,In_907,In_342);
nor U4322 (N_4322,In_358,In_490);
or U4323 (N_4323,In_807,In_448);
or U4324 (N_4324,In_921,In_552);
nor U4325 (N_4325,In_473,In_1);
and U4326 (N_4326,In_256,In_335);
nand U4327 (N_4327,In_361,In_74);
or U4328 (N_4328,In_381,In_942);
or U4329 (N_4329,In_945,In_215);
and U4330 (N_4330,In_320,In_946);
or U4331 (N_4331,In_904,In_209);
nor U4332 (N_4332,In_711,In_355);
or U4333 (N_4333,In_357,In_501);
and U4334 (N_4334,In_855,In_895);
nand U4335 (N_4335,In_526,In_627);
and U4336 (N_4336,In_743,In_319);
and U4337 (N_4337,In_241,In_695);
and U4338 (N_4338,In_622,In_457);
or U4339 (N_4339,In_601,In_953);
xor U4340 (N_4340,In_25,In_491);
nand U4341 (N_4341,In_191,In_628);
nor U4342 (N_4342,In_202,In_525);
nor U4343 (N_4343,In_279,In_392);
nor U4344 (N_4344,In_30,In_697);
or U4345 (N_4345,In_860,In_412);
or U4346 (N_4346,In_141,In_437);
or U4347 (N_4347,In_986,In_946);
and U4348 (N_4348,In_680,In_769);
nand U4349 (N_4349,In_410,In_960);
nand U4350 (N_4350,In_658,In_609);
and U4351 (N_4351,In_87,In_459);
and U4352 (N_4352,In_560,In_906);
and U4353 (N_4353,In_11,In_444);
nor U4354 (N_4354,In_417,In_969);
or U4355 (N_4355,In_516,In_926);
nor U4356 (N_4356,In_74,In_876);
nor U4357 (N_4357,In_770,In_971);
nand U4358 (N_4358,In_764,In_710);
nand U4359 (N_4359,In_66,In_974);
or U4360 (N_4360,In_351,In_986);
nor U4361 (N_4361,In_430,In_149);
and U4362 (N_4362,In_911,In_143);
or U4363 (N_4363,In_159,In_300);
or U4364 (N_4364,In_491,In_981);
and U4365 (N_4365,In_882,In_590);
nor U4366 (N_4366,In_611,In_981);
and U4367 (N_4367,In_293,In_510);
nor U4368 (N_4368,In_664,In_791);
or U4369 (N_4369,In_235,In_925);
nand U4370 (N_4370,In_458,In_274);
and U4371 (N_4371,In_61,In_320);
nand U4372 (N_4372,In_907,In_11);
and U4373 (N_4373,In_259,In_278);
or U4374 (N_4374,In_327,In_134);
and U4375 (N_4375,In_373,In_249);
nor U4376 (N_4376,In_719,In_373);
or U4377 (N_4377,In_866,In_859);
and U4378 (N_4378,In_892,In_445);
nand U4379 (N_4379,In_740,In_467);
nor U4380 (N_4380,In_522,In_356);
nand U4381 (N_4381,In_991,In_439);
nor U4382 (N_4382,In_898,In_886);
nand U4383 (N_4383,In_899,In_172);
and U4384 (N_4384,In_516,In_923);
and U4385 (N_4385,In_299,In_423);
nor U4386 (N_4386,In_824,In_449);
xor U4387 (N_4387,In_697,In_825);
nand U4388 (N_4388,In_65,In_205);
or U4389 (N_4389,In_6,In_871);
or U4390 (N_4390,In_810,In_477);
or U4391 (N_4391,In_430,In_850);
and U4392 (N_4392,In_221,In_460);
nand U4393 (N_4393,In_329,In_537);
or U4394 (N_4394,In_633,In_55);
or U4395 (N_4395,In_778,In_298);
or U4396 (N_4396,In_42,In_346);
xnor U4397 (N_4397,In_417,In_269);
and U4398 (N_4398,In_288,In_366);
or U4399 (N_4399,In_248,In_569);
and U4400 (N_4400,In_954,In_910);
or U4401 (N_4401,In_926,In_312);
and U4402 (N_4402,In_350,In_581);
and U4403 (N_4403,In_980,In_130);
and U4404 (N_4404,In_819,In_101);
nand U4405 (N_4405,In_617,In_999);
nand U4406 (N_4406,In_224,In_155);
and U4407 (N_4407,In_556,In_332);
or U4408 (N_4408,In_49,In_558);
nor U4409 (N_4409,In_876,In_430);
nand U4410 (N_4410,In_517,In_495);
nor U4411 (N_4411,In_59,In_287);
xor U4412 (N_4412,In_858,In_409);
and U4413 (N_4413,In_65,In_666);
or U4414 (N_4414,In_627,In_204);
or U4415 (N_4415,In_450,In_568);
and U4416 (N_4416,In_356,In_779);
nor U4417 (N_4417,In_875,In_951);
and U4418 (N_4418,In_510,In_576);
and U4419 (N_4419,In_713,In_92);
or U4420 (N_4420,In_913,In_854);
and U4421 (N_4421,In_269,In_777);
nor U4422 (N_4422,In_663,In_39);
or U4423 (N_4423,In_760,In_754);
and U4424 (N_4424,In_910,In_72);
nand U4425 (N_4425,In_938,In_193);
nor U4426 (N_4426,In_109,In_9);
nand U4427 (N_4427,In_744,In_718);
nor U4428 (N_4428,In_915,In_734);
nor U4429 (N_4429,In_981,In_190);
nand U4430 (N_4430,In_300,In_928);
nor U4431 (N_4431,In_581,In_42);
nand U4432 (N_4432,In_676,In_266);
xor U4433 (N_4433,In_978,In_377);
or U4434 (N_4434,In_663,In_783);
nand U4435 (N_4435,In_842,In_744);
nor U4436 (N_4436,In_474,In_313);
or U4437 (N_4437,In_22,In_927);
nor U4438 (N_4438,In_428,In_329);
and U4439 (N_4439,In_472,In_995);
nor U4440 (N_4440,In_510,In_794);
and U4441 (N_4441,In_83,In_605);
nand U4442 (N_4442,In_105,In_872);
nor U4443 (N_4443,In_156,In_774);
nand U4444 (N_4444,In_649,In_57);
or U4445 (N_4445,In_470,In_916);
or U4446 (N_4446,In_376,In_621);
and U4447 (N_4447,In_186,In_926);
nor U4448 (N_4448,In_374,In_32);
or U4449 (N_4449,In_601,In_199);
or U4450 (N_4450,In_83,In_751);
nor U4451 (N_4451,In_791,In_853);
nand U4452 (N_4452,In_184,In_778);
or U4453 (N_4453,In_783,In_324);
or U4454 (N_4454,In_797,In_825);
nor U4455 (N_4455,In_968,In_119);
and U4456 (N_4456,In_941,In_274);
nor U4457 (N_4457,In_324,In_439);
nand U4458 (N_4458,In_512,In_242);
and U4459 (N_4459,In_577,In_403);
nor U4460 (N_4460,In_35,In_504);
and U4461 (N_4461,In_500,In_177);
and U4462 (N_4462,In_774,In_772);
nand U4463 (N_4463,In_125,In_794);
nand U4464 (N_4464,In_17,In_51);
and U4465 (N_4465,In_800,In_741);
nand U4466 (N_4466,In_208,In_854);
and U4467 (N_4467,In_2,In_479);
and U4468 (N_4468,In_560,In_245);
nor U4469 (N_4469,In_858,In_556);
nor U4470 (N_4470,In_779,In_385);
nand U4471 (N_4471,In_242,In_284);
nand U4472 (N_4472,In_74,In_689);
or U4473 (N_4473,In_136,In_791);
nor U4474 (N_4474,In_185,In_232);
nor U4475 (N_4475,In_854,In_1);
nand U4476 (N_4476,In_269,In_410);
or U4477 (N_4477,In_677,In_894);
or U4478 (N_4478,In_528,In_183);
nand U4479 (N_4479,In_723,In_441);
or U4480 (N_4480,In_862,In_432);
nor U4481 (N_4481,In_182,In_401);
or U4482 (N_4482,In_731,In_532);
and U4483 (N_4483,In_538,In_706);
or U4484 (N_4484,In_720,In_348);
and U4485 (N_4485,In_446,In_514);
or U4486 (N_4486,In_44,In_781);
and U4487 (N_4487,In_761,In_747);
or U4488 (N_4488,In_965,In_153);
and U4489 (N_4489,In_196,In_918);
or U4490 (N_4490,In_88,In_320);
or U4491 (N_4491,In_109,In_218);
nor U4492 (N_4492,In_450,In_232);
and U4493 (N_4493,In_57,In_14);
nand U4494 (N_4494,In_613,In_359);
or U4495 (N_4495,In_103,In_632);
nand U4496 (N_4496,In_785,In_123);
and U4497 (N_4497,In_350,In_10);
and U4498 (N_4498,In_422,In_229);
or U4499 (N_4499,In_539,In_427);
and U4500 (N_4500,In_73,In_759);
or U4501 (N_4501,In_190,In_264);
and U4502 (N_4502,In_360,In_499);
nor U4503 (N_4503,In_165,In_250);
or U4504 (N_4504,In_725,In_183);
nand U4505 (N_4505,In_473,In_286);
or U4506 (N_4506,In_412,In_171);
or U4507 (N_4507,In_385,In_848);
nand U4508 (N_4508,In_361,In_165);
nand U4509 (N_4509,In_175,In_988);
nand U4510 (N_4510,In_375,In_888);
and U4511 (N_4511,In_980,In_318);
and U4512 (N_4512,In_381,In_37);
or U4513 (N_4513,In_742,In_518);
or U4514 (N_4514,In_930,In_324);
nor U4515 (N_4515,In_173,In_458);
nand U4516 (N_4516,In_917,In_311);
and U4517 (N_4517,In_577,In_894);
and U4518 (N_4518,In_683,In_209);
nand U4519 (N_4519,In_613,In_833);
xnor U4520 (N_4520,In_191,In_125);
and U4521 (N_4521,In_71,In_550);
nor U4522 (N_4522,In_263,In_488);
or U4523 (N_4523,In_954,In_446);
and U4524 (N_4524,In_981,In_520);
or U4525 (N_4525,In_547,In_275);
and U4526 (N_4526,In_391,In_230);
or U4527 (N_4527,In_252,In_113);
or U4528 (N_4528,In_473,In_595);
or U4529 (N_4529,In_358,In_163);
nor U4530 (N_4530,In_259,In_659);
nand U4531 (N_4531,In_33,In_985);
or U4532 (N_4532,In_429,In_136);
nand U4533 (N_4533,In_41,In_893);
nand U4534 (N_4534,In_997,In_245);
or U4535 (N_4535,In_741,In_121);
nor U4536 (N_4536,In_417,In_335);
or U4537 (N_4537,In_703,In_706);
xnor U4538 (N_4538,In_460,In_615);
nor U4539 (N_4539,In_366,In_808);
or U4540 (N_4540,In_512,In_770);
or U4541 (N_4541,In_124,In_911);
nand U4542 (N_4542,In_497,In_673);
nand U4543 (N_4543,In_716,In_799);
and U4544 (N_4544,In_8,In_67);
or U4545 (N_4545,In_851,In_88);
nor U4546 (N_4546,In_476,In_804);
nor U4547 (N_4547,In_816,In_681);
and U4548 (N_4548,In_920,In_828);
or U4549 (N_4549,In_546,In_2);
nor U4550 (N_4550,In_480,In_270);
or U4551 (N_4551,In_519,In_631);
or U4552 (N_4552,In_880,In_892);
and U4553 (N_4553,In_999,In_635);
or U4554 (N_4554,In_248,In_930);
and U4555 (N_4555,In_590,In_109);
nor U4556 (N_4556,In_552,In_194);
or U4557 (N_4557,In_303,In_551);
nand U4558 (N_4558,In_541,In_256);
nor U4559 (N_4559,In_997,In_125);
nand U4560 (N_4560,In_890,In_755);
nand U4561 (N_4561,In_592,In_347);
and U4562 (N_4562,In_753,In_157);
nand U4563 (N_4563,In_605,In_296);
nand U4564 (N_4564,In_15,In_150);
and U4565 (N_4565,In_108,In_760);
xnor U4566 (N_4566,In_517,In_653);
and U4567 (N_4567,In_220,In_97);
nor U4568 (N_4568,In_980,In_20);
nor U4569 (N_4569,In_422,In_957);
nor U4570 (N_4570,In_742,In_65);
and U4571 (N_4571,In_789,In_395);
nor U4572 (N_4572,In_888,In_809);
nand U4573 (N_4573,In_514,In_401);
or U4574 (N_4574,In_927,In_988);
and U4575 (N_4575,In_847,In_781);
or U4576 (N_4576,In_975,In_782);
nand U4577 (N_4577,In_70,In_224);
nand U4578 (N_4578,In_484,In_739);
or U4579 (N_4579,In_569,In_563);
nor U4580 (N_4580,In_740,In_826);
and U4581 (N_4581,In_232,In_467);
nor U4582 (N_4582,In_352,In_141);
and U4583 (N_4583,In_78,In_998);
or U4584 (N_4584,In_248,In_63);
nor U4585 (N_4585,In_417,In_457);
nand U4586 (N_4586,In_555,In_122);
and U4587 (N_4587,In_572,In_316);
or U4588 (N_4588,In_794,In_15);
and U4589 (N_4589,In_890,In_929);
nand U4590 (N_4590,In_434,In_492);
nand U4591 (N_4591,In_45,In_780);
or U4592 (N_4592,In_763,In_373);
nand U4593 (N_4593,In_667,In_137);
and U4594 (N_4594,In_880,In_753);
or U4595 (N_4595,In_996,In_240);
or U4596 (N_4596,In_552,In_979);
nor U4597 (N_4597,In_446,In_869);
nand U4598 (N_4598,In_811,In_347);
nor U4599 (N_4599,In_584,In_557);
nor U4600 (N_4600,In_943,In_574);
nand U4601 (N_4601,In_766,In_647);
nor U4602 (N_4602,In_760,In_451);
or U4603 (N_4603,In_871,In_105);
and U4604 (N_4604,In_567,In_406);
nand U4605 (N_4605,In_213,In_500);
nand U4606 (N_4606,In_468,In_88);
nand U4607 (N_4607,In_700,In_264);
or U4608 (N_4608,In_19,In_553);
and U4609 (N_4609,In_966,In_337);
and U4610 (N_4610,In_244,In_540);
nor U4611 (N_4611,In_887,In_774);
or U4612 (N_4612,In_710,In_160);
and U4613 (N_4613,In_773,In_176);
and U4614 (N_4614,In_13,In_810);
and U4615 (N_4615,In_871,In_673);
nor U4616 (N_4616,In_352,In_920);
nor U4617 (N_4617,In_846,In_610);
nand U4618 (N_4618,In_648,In_162);
nor U4619 (N_4619,In_35,In_925);
or U4620 (N_4620,In_905,In_641);
nor U4621 (N_4621,In_492,In_214);
or U4622 (N_4622,In_810,In_696);
nand U4623 (N_4623,In_36,In_888);
nor U4624 (N_4624,In_357,In_374);
and U4625 (N_4625,In_385,In_86);
nand U4626 (N_4626,In_609,In_169);
nor U4627 (N_4627,In_341,In_418);
nor U4628 (N_4628,In_159,In_50);
nor U4629 (N_4629,In_893,In_527);
nor U4630 (N_4630,In_855,In_321);
and U4631 (N_4631,In_110,In_58);
or U4632 (N_4632,In_91,In_149);
and U4633 (N_4633,In_520,In_461);
and U4634 (N_4634,In_282,In_670);
and U4635 (N_4635,In_724,In_882);
nor U4636 (N_4636,In_295,In_909);
and U4637 (N_4637,In_972,In_978);
nand U4638 (N_4638,In_40,In_351);
nor U4639 (N_4639,In_474,In_984);
nor U4640 (N_4640,In_406,In_874);
nand U4641 (N_4641,In_257,In_822);
and U4642 (N_4642,In_452,In_505);
nand U4643 (N_4643,In_686,In_675);
or U4644 (N_4644,In_106,In_693);
or U4645 (N_4645,In_490,In_79);
and U4646 (N_4646,In_395,In_654);
or U4647 (N_4647,In_61,In_679);
or U4648 (N_4648,In_830,In_974);
nor U4649 (N_4649,In_441,In_681);
or U4650 (N_4650,In_210,In_978);
and U4651 (N_4651,In_823,In_99);
nand U4652 (N_4652,In_991,In_380);
or U4653 (N_4653,In_466,In_286);
xnor U4654 (N_4654,In_216,In_994);
nand U4655 (N_4655,In_925,In_192);
nand U4656 (N_4656,In_141,In_463);
and U4657 (N_4657,In_573,In_589);
and U4658 (N_4658,In_643,In_89);
nand U4659 (N_4659,In_488,In_97);
nor U4660 (N_4660,In_93,In_506);
or U4661 (N_4661,In_514,In_645);
and U4662 (N_4662,In_881,In_619);
and U4663 (N_4663,In_553,In_95);
nor U4664 (N_4664,In_704,In_334);
nor U4665 (N_4665,In_995,In_888);
nor U4666 (N_4666,In_53,In_249);
nand U4667 (N_4667,In_426,In_537);
nor U4668 (N_4668,In_424,In_440);
nor U4669 (N_4669,In_184,In_708);
nand U4670 (N_4670,In_662,In_783);
and U4671 (N_4671,In_419,In_62);
or U4672 (N_4672,In_186,In_168);
nor U4673 (N_4673,In_840,In_419);
nor U4674 (N_4674,In_297,In_549);
nor U4675 (N_4675,In_95,In_109);
nor U4676 (N_4676,In_588,In_85);
nor U4677 (N_4677,In_556,In_215);
nor U4678 (N_4678,In_588,In_140);
or U4679 (N_4679,In_309,In_453);
or U4680 (N_4680,In_62,In_435);
or U4681 (N_4681,In_278,In_13);
xor U4682 (N_4682,In_44,In_40);
and U4683 (N_4683,In_444,In_438);
and U4684 (N_4684,In_996,In_748);
or U4685 (N_4685,In_196,In_945);
or U4686 (N_4686,In_300,In_333);
or U4687 (N_4687,In_984,In_166);
or U4688 (N_4688,In_740,In_53);
xnor U4689 (N_4689,In_932,In_884);
or U4690 (N_4690,In_282,In_417);
or U4691 (N_4691,In_430,In_542);
or U4692 (N_4692,In_758,In_748);
nor U4693 (N_4693,In_182,In_54);
nand U4694 (N_4694,In_96,In_179);
and U4695 (N_4695,In_165,In_523);
nor U4696 (N_4696,In_667,In_793);
or U4697 (N_4697,In_133,In_531);
nand U4698 (N_4698,In_83,In_433);
nor U4699 (N_4699,In_605,In_888);
and U4700 (N_4700,In_837,In_4);
and U4701 (N_4701,In_303,In_800);
xor U4702 (N_4702,In_496,In_533);
nor U4703 (N_4703,In_175,In_892);
and U4704 (N_4704,In_127,In_625);
or U4705 (N_4705,In_126,In_48);
nor U4706 (N_4706,In_720,In_109);
and U4707 (N_4707,In_802,In_886);
or U4708 (N_4708,In_338,In_556);
or U4709 (N_4709,In_610,In_963);
xor U4710 (N_4710,In_10,In_290);
and U4711 (N_4711,In_855,In_666);
nor U4712 (N_4712,In_2,In_181);
nor U4713 (N_4713,In_523,In_750);
nand U4714 (N_4714,In_238,In_118);
nor U4715 (N_4715,In_789,In_547);
nor U4716 (N_4716,In_344,In_90);
and U4717 (N_4717,In_808,In_228);
and U4718 (N_4718,In_923,In_902);
or U4719 (N_4719,In_62,In_786);
nor U4720 (N_4720,In_221,In_385);
nand U4721 (N_4721,In_936,In_351);
and U4722 (N_4722,In_663,In_490);
nand U4723 (N_4723,In_192,In_164);
nand U4724 (N_4724,In_444,In_949);
or U4725 (N_4725,In_363,In_651);
nor U4726 (N_4726,In_334,In_27);
nand U4727 (N_4727,In_2,In_404);
nand U4728 (N_4728,In_940,In_224);
xnor U4729 (N_4729,In_797,In_754);
and U4730 (N_4730,In_261,In_823);
or U4731 (N_4731,In_310,In_428);
nand U4732 (N_4732,In_880,In_346);
nor U4733 (N_4733,In_442,In_287);
or U4734 (N_4734,In_56,In_470);
nor U4735 (N_4735,In_90,In_75);
xor U4736 (N_4736,In_610,In_946);
nand U4737 (N_4737,In_524,In_995);
nand U4738 (N_4738,In_267,In_71);
nand U4739 (N_4739,In_451,In_264);
and U4740 (N_4740,In_126,In_372);
and U4741 (N_4741,In_30,In_578);
or U4742 (N_4742,In_519,In_397);
or U4743 (N_4743,In_978,In_38);
and U4744 (N_4744,In_937,In_602);
or U4745 (N_4745,In_534,In_969);
and U4746 (N_4746,In_448,In_615);
nand U4747 (N_4747,In_522,In_651);
nand U4748 (N_4748,In_262,In_547);
and U4749 (N_4749,In_824,In_372);
and U4750 (N_4750,In_335,In_657);
or U4751 (N_4751,In_48,In_467);
nand U4752 (N_4752,In_404,In_424);
and U4753 (N_4753,In_651,In_294);
and U4754 (N_4754,In_278,In_182);
nand U4755 (N_4755,In_309,In_693);
nor U4756 (N_4756,In_389,In_200);
and U4757 (N_4757,In_368,In_450);
nand U4758 (N_4758,In_792,In_104);
nor U4759 (N_4759,In_220,In_383);
or U4760 (N_4760,In_613,In_94);
nor U4761 (N_4761,In_43,In_552);
nand U4762 (N_4762,In_416,In_778);
xnor U4763 (N_4763,In_271,In_465);
xor U4764 (N_4764,In_795,In_376);
and U4765 (N_4765,In_8,In_70);
nand U4766 (N_4766,In_576,In_634);
nand U4767 (N_4767,In_629,In_824);
nor U4768 (N_4768,In_946,In_332);
nor U4769 (N_4769,In_967,In_855);
nand U4770 (N_4770,In_654,In_914);
and U4771 (N_4771,In_509,In_449);
nor U4772 (N_4772,In_575,In_864);
or U4773 (N_4773,In_973,In_181);
and U4774 (N_4774,In_665,In_966);
and U4775 (N_4775,In_694,In_883);
nand U4776 (N_4776,In_262,In_385);
and U4777 (N_4777,In_720,In_440);
or U4778 (N_4778,In_169,In_36);
nor U4779 (N_4779,In_523,In_238);
nand U4780 (N_4780,In_592,In_296);
xor U4781 (N_4781,In_113,In_527);
nor U4782 (N_4782,In_534,In_369);
or U4783 (N_4783,In_730,In_778);
nor U4784 (N_4784,In_664,In_185);
nor U4785 (N_4785,In_974,In_852);
and U4786 (N_4786,In_52,In_879);
or U4787 (N_4787,In_48,In_338);
and U4788 (N_4788,In_413,In_948);
or U4789 (N_4789,In_694,In_930);
and U4790 (N_4790,In_682,In_152);
nand U4791 (N_4791,In_959,In_575);
and U4792 (N_4792,In_615,In_124);
nor U4793 (N_4793,In_844,In_496);
and U4794 (N_4794,In_442,In_48);
nor U4795 (N_4795,In_826,In_584);
or U4796 (N_4796,In_524,In_986);
nor U4797 (N_4797,In_639,In_502);
or U4798 (N_4798,In_888,In_392);
nor U4799 (N_4799,In_800,In_404);
and U4800 (N_4800,In_417,In_649);
or U4801 (N_4801,In_885,In_978);
and U4802 (N_4802,In_82,In_346);
or U4803 (N_4803,In_329,In_777);
and U4804 (N_4804,In_326,In_580);
nand U4805 (N_4805,In_122,In_650);
or U4806 (N_4806,In_621,In_198);
xnor U4807 (N_4807,In_985,In_289);
and U4808 (N_4808,In_428,In_547);
or U4809 (N_4809,In_71,In_932);
and U4810 (N_4810,In_76,In_207);
nand U4811 (N_4811,In_272,In_945);
nand U4812 (N_4812,In_35,In_146);
nor U4813 (N_4813,In_517,In_932);
nand U4814 (N_4814,In_130,In_20);
nor U4815 (N_4815,In_546,In_561);
nor U4816 (N_4816,In_675,In_605);
or U4817 (N_4817,In_861,In_68);
nor U4818 (N_4818,In_476,In_907);
or U4819 (N_4819,In_208,In_64);
and U4820 (N_4820,In_721,In_311);
and U4821 (N_4821,In_389,In_341);
nand U4822 (N_4822,In_981,In_962);
nor U4823 (N_4823,In_846,In_111);
or U4824 (N_4824,In_502,In_231);
or U4825 (N_4825,In_407,In_89);
or U4826 (N_4826,In_109,In_873);
nand U4827 (N_4827,In_305,In_808);
nor U4828 (N_4828,In_280,In_959);
xor U4829 (N_4829,In_70,In_126);
nor U4830 (N_4830,In_583,In_739);
or U4831 (N_4831,In_496,In_988);
or U4832 (N_4832,In_146,In_348);
nand U4833 (N_4833,In_968,In_617);
or U4834 (N_4834,In_640,In_12);
or U4835 (N_4835,In_849,In_66);
and U4836 (N_4836,In_725,In_945);
or U4837 (N_4837,In_665,In_115);
and U4838 (N_4838,In_332,In_216);
nor U4839 (N_4839,In_149,In_579);
and U4840 (N_4840,In_190,In_305);
and U4841 (N_4841,In_501,In_324);
and U4842 (N_4842,In_355,In_201);
nor U4843 (N_4843,In_554,In_646);
and U4844 (N_4844,In_481,In_516);
and U4845 (N_4845,In_930,In_154);
and U4846 (N_4846,In_235,In_384);
nand U4847 (N_4847,In_102,In_314);
nand U4848 (N_4848,In_991,In_462);
nor U4849 (N_4849,In_465,In_176);
nand U4850 (N_4850,In_144,In_418);
nand U4851 (N_4851,In_441,In_927);
and U4852 (N_4852,In_413,In_328);
or U4853 (N_4853,In_565,In_329);
nand U4854 (N_4854,In_436,In_825);
and U4855 (N_4855,In_306,In_421);
or U4856 (N_4856,In_593,In_909);
nor U4857 (N_4857,In_129,In_582);
or U4858 (N_4858,In_905,In_980);
and U4859 (N_4859,In_133,In_65);
or U4860 (N_4860,In_136,In_397);
nand U4861 (N_4861,In_137,In_218);
and U4862 (N_4862,In_251,In_216);
and U4863 (N_4863,In_496,In_877);
and U4864 (N_4864,In_357,In_64);
or U4865 (N_4865,In_69,In_172);
or U4866 (N_4866,In_401,In_730);
nor U4867 (N_4867,In_698,In_737);
and U4868 (N_4868,In_278,In_201);
and U4869 (N_4869,In_480,In_425);
and U4870 (N_4870,In_549,In_918);
or U4871 (N_4871,In_763,In_919);
and U4872 (N_4872,In_974,In_253);
nand U4873 (N_4873,In_94,In_268);
and U4874 (N_4874,In_742,In_248);
nand U4875 (N_4875,In_925,In_426);
nor U4876 (N_4876,In_840,In_993);
and U4877 (N_4877,In_92,In_492);
nand U4878 (N_4878,In_647,In_179);
nor U4879 (N_4879,In_691,In_718);
nor U4880 (N_4880,In_433,In_424);
nor U4881 (N_4881,In_355,In_58);
or U4882 (N_4882,In_243,In_539);
nor U4883 (N_4883,In_806,In_995);
nor U4884 (N_4884,In_812,In_813);
or U4885 (N_4885,In_825,In_25);
nor U4886 (N_4886,In_696,In_161);
or U4887 (N_4887,In_398,In_293);
nor U4888 (N_4888,In_252,In_809);
nor U4889 (N_4889,In_79,In_545);
or U4890 (N_4890,In_216,In_768);
nor U4891 (N_4891,In_878,In_915);
xor U4892 (N_4892,In_696,In_215);
or U4893 (N_4893,In_951,In_628);
or U4894 (N_4894,In_504,In_12);
nand U4895 (N_4895,In_600,In_445);
nand U4896 (N_4896,In_319,In_866);
and U4897 (N_4897,In_895,In_552);
or U4898 (N_4898,In_37,In_342);
xnor U4899 (N_4899,In_600,In_895);
nand U4900 (N_4900,In_688,In_189);
nand U4901 (N_4901,In_878,In_806);
nand U4902 (N_4902,In_532,In_611);
or U4903 (N_4903,In_892,In_926);
or U4904 (N_4904,In_429,In_773);
or U4905 (N_4905,In_978,In_495);
and U4906 (N_4906,In_530,In_795);
and U4907 (N_4907,In_962,In_768);
and U4908 (N_4908,In_36,In_977);
and U4909 (N_4909,In_128,In_382);
nor U4910 (N_4910,In_172,In_360);
or U4911 (N_4911,In_745,In_241);
or U4912 (N_4912,In_263,In_302);
and U4913 (N_4913,In_424,In_621);
nor U4914 (N_4914,In_885,In_145);
and U4915 (N_4915,In_269,In_345);
or U4916 (N_4916,In_622,In_578);
and U4917 (N_4917,In_435,In_589);
nor U4918 (N_4918,In_716,In_635);
nor U4919 (N_4919,In_146,In_77);
xnor U4920 (N_4920,In_298,In_859);
or U4921 (N_4921,In_674,In_235);
nor U4922 (N_4922,In_196,In_674);
nor U4923 (N_4923,In_802,In_816);
and U4924 (N_4924,In_429,In_748);
and U4925 (N_4925,In_390,In_332);
and U4926 (N_4926,In_749,In_615);
xnor U4927 (N_4927,In_514,In_804);
nand U4928 (N_4928,In_568,In_218);
and U4929 (N_4929,In_869,In_873);
and U4930 (N_4930,In_653,In_294);
nand U4931 (N_4931,In_716,In_47);
or U4932 (N_4932,In_659,In_310);
or U4933 (N_4933,In_183,In_299);
and U4934 (N_4934,In_965,In_284);
nor U4935 (N_4935,In_399,In_178);
and U4936 (N_4936,In_15,In_344);
nand U4937 (N_4937,In_431,In_722);
or U4938 (N_4938,In_103,In_991);
nor U4939 (N_4939,In_304,In_34);
and U4940 (N_4940,In_705,In_753);
and U4941 (N_4941,In_719,In_91);
and U4942 (N_4942,In_33,In_295);
and U4943 (N_4943,In_483,In_168);
or U4944 (N_4944,In_607,In_121);
or U4945 (N_4945,In_831,In_122);
and U4946 (N_4946,In_906,In_528);
nand U4947 (N_4947,In_213,In_131);
nor U4948 (N_4948,In_579,In_82);
nor U4949 (N_4949,In_739,In_755);
nor U4950 (N_4950,In_452,In_292);
and U4951 (N_4951,In_529,In_31);
nor U4952 (N_4952,In_823,In_521);
nand U4953 (N_4953,In_918,In_618);
nor U4954 (N_4954,In_695,In_263);
and U4955 (N_4955,In_262,In_256);
nand U4956 (N_4956,In_917,In_324);
nand U4957 (N_4957,In_431,In_793);
nor U4958 (N_4958,In_904,In_625);
nand U4959 (N_4959,In_145,In_383);
or U4960 (N_4960,In_784,In_486);
nor U4961 (N_4961,In_552,In_831);
nor U4962 (N_4962,In_956,In_276);
or U4963 (N_4963,In_189,In_856);
nand U4964 (N_4964,In_23,In_855);
nor U4965 (N_4965,In_177,In_468);
or U4966 (N_4966,In_771,In_40);
xor U4967 (N_4967,In_807,In_503);
and U4968 (N_4968,In_140,In_159);
or U4969 (N_4969,In_936,In_287);
or U4970 (N_4970,In_652,In_973);
nor U4971 (N_4971,In_20,In_738);
and U4972 (N_4972,In_314,In_13);
nor U4973 (N_4973,In_669,In_14);
and U4974 (N_4974,In_485,In_427);
nor U4975 (N_4975,In_982,In_507);
or U4976 (N_4976,In_592,In_766);
and U4977 (N_4977,In_191,In_491);
and U4978 (N_4978,In_200,In_789);
and U4979 (N_4979,In_487,In_562);
nor U4980 (N_4980,In_145,In_400);
nor U4981 (N_4981,In_847,In_514);
and U4982 (N_4982,In_122,In_195);
or U4983 (N_4983,In_481,In_56);
nor U4984 (N_4984,In_586,In_506);
or U4985 (N_4985,In_426,In_25);
nand U4986 (N_4986,In_535,In_220);
nand U4987 (N_4987,In_828,In_378);
nor U4988 (N_4988,In_318,In_988);
and U4989 (N_4989,In_647,In_118);
nand U4990 (N_4990,In_983,In_132);
nand U4991 (N_4991,In_480,In_853);
or U4992 (N_4992,In_89,In_426);
or U4993 (N_4993,In_19,In_303);
nand U4994 (N_4994,In_151,In_849);
and U4995 (N_4995,In_181,In_72);
nor U4996 (N_4996,In_959,In_663);
nand U4997 (N_4997,In_545,In_299);
nand U4998 (N_4998,In_8,In_59);
or U4999 (N_4999,In_788,In_840);
or U5000 (N_5000,N_3218,N_921);
nor U5001 (N_5001,N_3301,N_3862);
nand U5002 (N_5002,N_751,N_4632);
nand U5003 (N_5003,N_2726,N_4103);
or U5004 (N_5004,N_2557,N_461);
nor U5005 (N_5005,N_4593,N_4022);
nor U5006 (N_5006,N_1359,N_2598);
and U5007 (N_5007,N_4469,N_1188);
nand U5008 (N_5008,N_3485,N_3474);
and U5009 (N_5009,N_2425,N_3466);
nor U5010 (N_5010,N_1297,N_4783);
or U5011 (N_5011,N_1876,N_3510);
and U5012 (N_5012,N_974,N_4064);
and U5013 (N_5013,N_2717,N_3507);
nand U5014 (N_5014,N_4974,N_22);
nor U5015 (N_5015,N_4088,N_1226);
nand U5016 (N_5016,N_2753,N_372);
or U5017 (N_5017,N_3942,N_1323);
nand U5018 (N_5018,N_651,N_3045);
or U5019 (N_5019,N_4289,N_4570);
or U5020 (N_5020,N_452,N_2264);
xor U5021 (N_5021,N_1854,N_322);
xor U5022 (N_5022,N_4118,N_3578);
nor U5023 (N_5023,N_715,N_4466);
nor U5024 (N_5024,N_3201,N_4923);
nand U5025 (N_5025,N_3969,N_3882);
and U5026 (N_5026,N_62,N_1241);
nor U5027 (N_5027,N_3864,N_2581);
or U5028 (N_5028,N_1106,N_2786);
nand U5029 (N_5029,N_1170,N_1908);
nor U5030 (N_5030,N_2061,N_2049);
nor U5031 (N_5031,N_1368,N_3567);
nand U5032 (N_5032,N_2545,N_2779);
and U5033 (N_5033,N_3340,N_3194);
and U5034 (N_5034,N_4502,N_4488);
or U5035 (N_5035,N_2743,N_273);
nor U5036 (N_5036,N_2923,N_160);
or U5037 (N_5037,N_4935,N_2102);
or U5038 (N_5038,N_4395,N_4737);
nor U5039 (N_5039,N_519,N_4730);
or U5040 (N_5040,N_1577,N_822);
or U5041 (N_5041,N_1335,N_4879);
and U5042 (N_5042,N_2064,N_3150);
nand U5043 (N_5043,N_4333,N_4508);
nand U5044 (N_5044,N_2813,N_758);
or U5045 (N_5045,N_128,N_4965);
or U5046 (N_5046,N_4963,N_1589);
nand U5047 (N_5047,N_3160,N_2600);
nand U5048 (N_5048,N_809,N_136);
nand U5049 (N_5049,N_1729,N_3285);
nand U5050 (N_5050,N_3399,N_3792);
or U5051 (N_5051,N_48,N_4304);
nand U5052 (N_5052,N_574,N_1538);
nor U5053 (N_5053,N_1806,N_3946);
nand U5054 (N_5054,N_4751,N_2835);
nor U5055 (N_5055,N_1635,N_537);
nor U5056 (N_5056,N_707,N_3910);
nor U5057 (N_5057,N_3761,N_3759);
nor U5058 (N_5058,N_4769,N_158);
nand U5059 (N_5059,N_3609,N_4249);
and U5060 (N_5060,N_3962,N_3282);
and U5061 (N_5061,N_4072,N_2501);
and U5062 (N_5062,N_238,N_1351);
and U5063 (N_5063,N_2550,N_4049);
nand U5064 (N_5064,N_1303,N_2088);
nand U5065 (N_5065,N_3770,N_4738);
nor U5066 (N_5066,N_956,N_4749);
or U5067 (N_5067,N_1531,N_2213);
nor U5068 (N_5068,N_4375,N_2334);
and U5069 (N_5069,N_451,N_2420);
or U5070 (N_5070,N_996,N_4552);
nor U5071 (N_5071,N_4,N_2597);
nor U5072 (N_5072,N_3491,N_2380);
nand U5073 (N_5073,N_343,N_3621);
or U5074 (N_5074,N_3806,N_2273);
or U5075 (N_5075,N_4201,N_1301);
or U5076 (N_5076,N_4227,N_1572);
or U5077 (N_5077,N_79,N_3065);
and U5078 (N_5078,N_251,N_3290);
and U5079 (N_5079,N_1344,N_472);
and U5080 (N_5080,N_468,N_3648);
nand U5081 (N_5081,N_2169,N_4712);
nor U5082 (N_5082,N_412,N_1040);
nand U5083 (N_5083,N_3941,N_4438);
and U5084 (N_5084,N_620,N_1867);
nand U5085 (N_5085,N_1025,N_2027);
or U5086 (N_5086,N_1332,N_4131);
and U5087 (N_5087,N_3549,N_660);
nor U5088 (N_5088,N_2943,N_635);
nand U5089 (N_5089,N_4157,N_4804);
and U5090 (N_5090,N_4484,N_89);
nand U5091 (N_5091,N_1083,N_1071);
nor U5092 (N_5092,N_3357,N_465);
and U5093 (N_5093,N_4145,N_3619);
and U5094 (N_5094,N_4826,N_2792);
or U5095 (N_5095,N_3914,N_2447);
or U5096 (N_5096,N_843,N_323);
and U5097 (N_5097,N_4808,N_3623);
or U5098 (N_5098,N_723,N_1666);
and U5099 (N_5099,N_3719,N_4128);
nand U5100 (N_5100,N_554,N_4903);
nor U5101 (N_5101,N_733,N_2082);
nor U5102 (N_5102,N_3622,N_3812);
nand U5103 (N_5103,N_1425,N_3456);
and U5104 (N_5104,N_1243,N_1742);
or U5105 (N_5105,N_1848,N_3269);
or U5106 (N_5106,N_1043,N_3950);
xnor U5107 (N_5107,N_4220,N_963);
nor U5108 (N_5108,N_4899,N_233);
and U5109 (N_5109,N_1735,N_2113);
nand U5110 (N_5110,N_1197,N_1761);
nand U5111 (N_5111,N_2708,N_3557);
or U5112 (N_5112,N_152,N_4631);
nor U5113 (N_5113,N_1095,N_1843);
and U5114 (N_5114,N_1861,N_3084);
and U5115 (N_5115,N_3935,N_4196);
and U5116 (N_5116,N_835,N_2278);
nor U5117 (N_5117,N_109,N_3645);
or U5118 (N_5118,N_420,N_3722);
nand U5119 (N_5119,N_3035,N_703);
or U5120 (N_5120,N_2349,N_553);
or U5121 (N_5121,N_2220,N_609);
xor U5122 (N_5122,N_1556,N_2153);
nand U5123 (N_5123,N_3392,N_4212);
nor U5124 (N_5124,N_1107,N_4541);
nand U5125 (N_5125,N_202,N_1820);
and U5126 (N_5126,N_2868,N_3344);
or U5127 (N_5127,N_1795,N_4746);
and U5128 (N_5128,N_3815,N_788);
or U5129 (N_5129,N_339,N_2491);
nor U5130 (N_5130,N_4867,N_4688);
nor U5131 (N_5131,N_4087,N_2133);
nand U5132 (N_5132,N_4098,N_1331);
and U5133 (N_5133,N_1783,N_3189);
and U5134 (N_5134,N_534,N_767);
or U5135 (N_5135,N_1553,N_3682);
xor U5136 (N_5136,N_4277,N_63);
nand U5137 (N_5137,N_414,N_1775);
nor U5138 (N_5138,N_1349,N_1967);
nand U5139 (N_5139,N_1129,N_4959);
nand U5140 (N_5140,N_2343,N_4398);
nand U5141 (N_5141,N_2266,N_380);
nor U5142 (N_5142,N_2787,N_1453);
nand U5143 (N_5143,N_4079,N_3059);
or U5144 (N_5144,N_2670,N_244);
nor U5145 (N_5145,N_4012,N_4601);
or U5146 (N_5146,N_561,N_416);
nor U5147 (N_5147,N_287,N_4710);
and U5148 (N_5148,N_4448,N_123);
or U5149 (N_5149,N_2444,N_909);
nand U5150 (N_5150,N_845,N_493);
or U5151 (N_5151,N_4810,N_2734);
nand U5152 (N_5152,N_3056,N_2657);
and U5153 (N_5153,N_4319,N_440);
nor U5154 (N_5154,N_2852,N_1264);
or U5155 (N_5155,N_2148,N_2970);
xnor U5156 (N_5156,N_3709,N_4458);
or U5157 (N_5157,N_4345,N_4793);
nor U5158 (N_5158,N_1618,N_1058);
and U5159 (N_5159,N_4456,N_3402);
nor U5160 (N_5160,N_2988,N_2874);
nand U5161 (N_5161,N_2079,N_607);
nand U5162 (N_5162,N_1838,N_2050);
and U5163 (N_5163,N_826,N_2941);
nor U5164 (N_5164,N_3366,N_3968);
or U5165 (N_5165,N_3369,N_3013);
and U5166 (N_5166,N_4885,N_1702);
and U5167 (N_5167,N_3877,N_1602);
or U5168 (N_5168,N_2015,N_975);
nor U5169 (N_5169,N_4347,N_4270);
and U5170 (N_5170,N_3880,N_4567);
nor U5171 (N_5171,N_4150,N_56);
nand U5172 (N_5172,N_3727,N_1657);
xnor U5173 (N_5173,N_959,N_4482);
xnor U5174 (N_5174,N_1113,N_833);
nand U5175 (N_5175,N_3793,N_3554);
nor U5176 (N_5176,N_4256,N_2283);
nand U5177 (N_5177,N_4801,N_922);
and U5178 (N_5178,N_2924,N_759);
or U5179 (N_5179,N_4332,N_4207);
and U5180 (N_5180,N_2442,N_4405);
nor U5181 (N_5181,N_1953,N_364);
nor U5182 (N_5182,N_3795,N_2480);
nand U5183 (N_5183,N_4120,N_1490);
nand U5184 (N_5184,N_2257,N_1026);
or U5185 (N_5185,N_391,N_3071);
nor U5186 (N_5186,N_4619,N_491);
or U5187 (N_5187,N_1777,N_1669);
nand U5188 (N_5188,N_898,N_2910);
nand U5189 (N_5189,N_3909,N_2508);
nor U5190 (N_5190,N_3390,N_1146);
or U5191 (N_5191,N_2593,N_13);
or U5192 (N_5192,N_2231,N_1562);
nor U5193 (N_5193,N_1916,N_917);
nor U5194 (N_5194,N_3429,N_1765);
and U5195 (N_5195,N_3317,N_2976);
nor U5196 (N_5196,N_215,N_3790);
or U5197 (N_5197,N_3106,N_1703);
nand U5198 (N_5198,N_1151,N_641);
or U5199 (N_5199,N_4327,N_1055);
nor U5200 (N_5200,N_3169,N_4317);
nor U5201 (N_5201,N_786,N_1380);
nand U5202 (N_5202,N_3611,N_3257);
or U5203 (N_5203,N_823,N_442);
nor U5204 (N_5204,N_270,N_4984);
nor U5205 (N_5205,N_2732,N_4537);
and U5206 (N_5206,N_4994,N_814);
nor U5207 (N_5207,N_1542,N_3827);
or U5208 (N_5208,N_3565,N_4866);
nand U5209 (N_5209,N_3731,N_4446);
or U5210 (N_5210,N_2221,N_2100);
nor U5211 (N_5211,N_4063,N_1520);
or U5212 (N_5212,N_508,N_1634);
nor U5213 (N_5213,N_1017,N_2030);
and U5214 (N_5214,N_2496,N_2002);
and U5215 (N_5215,N_1858,N_2471);
and U5216 (N_5216,N_512,N_634);
nand U5217 (N_5217,N_4968,N_1688);
or U5218 (N_5218,N_565,N_3261);
nand U5219 (N_5219,N_1596,N_3679);
and U5220 (N_5220,N_588,N_3772);
nor U5221 (N_5221,N_4158,N_3075);
nor U5222 (N_5222,N_1003,N_3175);
nand U5223 (N_5223,N_3416,N_4384);
and U5224 (N_5224,N_131,N_4136);
nor U5225 (N_5225,N_1700,N_3388);
nand U5226 (N_5226,N_2437,N_2504);
nor U5227 (N_5227,N_1200,N_67);
nand U5228 (N_5228,N_4286,N_4013);
nor U5229 (N_5229,N_2093,N_1924);
nand U5230 (N_5230,N_648,N_1884);
nor U5231 (N_5231,N_1825,N_4873);
nand U5232 (N_5232,N_3547,N_3669);
nor U5233 (N_5233,N_2429,N_1552);
and U5234 (N_5234,N_3769,N_4206);
and U5235 (N_5235,N_1169,N_3353);
or U5236 (N_5236,N_2675,N_216);
and U5237 (N_5237,N_2531,N_901);
nor U5238 (N_5238,N_2003,N_1519);
or U5239 (N_5239,N_2710,N_1006);
nand U5240 (N_5240,N_4926,N_298);
nor U5241 (N_5241,N_4178,N_122);
and U5242 (N_5242,N_3744,N_326);
and U5243 (N_5243,N_3384,N_2189);
nand U5244 (N_5244,N_3265,N_606);
nand U5245 (N_5245,N_2206,N_1438);
or U5246 (N_5246,N_3568,N_201);
and U5247 (N_5247,N_503,N_3575);
and U5248 (N_5248,N_4652,N_1082);
or U5249 (N_5249,N_1550,N_66);
nor U5250 (N_5250,N_107,N_2387);
and U5251 (N_5251,N_4915,N_2532);
xnor U5252 (N_5252,N_1222,N_2633);
nor U5253 (N_5253,N_894,N_1649);
or U5254 (N_5254,N_77,N_713);
nand U5255 (N_5255,N_4720,N_4023);
or U5256 (N_5256,N_837,N_1679);
nand U5257 (N_5257,N_3019,N_1746);
nor U5258 (N_5258,N_3143,N_3440);
and U5259 (N_5259,N_2951,N_3514);
nor U5260 (N_5260,N_1752,N_489);
or U5261 (N_5261,N_576,N_2669);
or U5262 (N_5262,N_3330,N_133);
and U5263 (N_5263,N_163,N_4371);
or U5264 (N_5264,N_138,N_612);
nor U5265 (N_5265,N_4388,N_3320);
nand U5266 (N_5266,N_1855,N_882);
nand U5267 (N_5267,N_2952,N_4330);
or U5268 (N_5268,N_692,N_2929);
or U5269 (N_5269,N_3347,N_1460);
nand U5270 (N_5270,N_3208,N_3741);
nand U5271 (N_5271,N_4889,N_1032);
and U5272 (N_5272,N_4556,N_1633);
or U5273 (N_5273,N_3158,N_2366);
xor U5274 (N_5274,N_2954,N_3241);
nor U5275 (N_5275,N_1617,N_4230);
and U5276 (N_5276,N_591,N_1153);
nand U5277 (N_5277,N_2573,N_4465);
nand U5278 (N_5278,N_399,N_3156);
and U5279 (N_5279,N_4831,N_3982);
or U5280 (N_5280,N_1590,N_3328);
nand U5281 (N_5281,N_4768,N_4346);
nor U5282 (N_5282,N_1944,N_4147);
nor U5283 (N_5283,N_437,N_754);
nand U5284 (N_5284,N_3073,N_1039);
nor U5285 (N_5285,N_2311,N_1404);
and U5286 (N_5286,N_4082,N_3725);
nand U5287 (N_5287,N_2772,N_830);
or U5288 (N_5288,N_3524,N_1511);
nor U5289 (N_5289,N_302,N_4638);
nand U5290 (N_5290,N_1636,N_3028);
nand U5291 (N_5291,N_1336,N_4154);
nand U5292 (N_5292,N_3453,N_4499);
and U5293 (N_5293,N_2288,N_987);
nand U5294 (N_5294,N_2018,N_1893);
nand U5295 (N_5295,N_1698,N_2078);
nor U5296 (N_5296,N_2276,N_4297);
or U5297 (N_5297,N_2932,N_2737);
or U5298 (N_5298,N_1972,N_1427);
nand U5299 (N_5299,N_4264,N_2121);
nand U5300 (N_5300,N_303,N_1644);
xnor U5301 (N_5301,N_1112,N_4790);
or U5302 (N_5302,N_4534,N_895);
and U5303 (N_5303,N_4721,N_1677);
and U5304 (N_5304,N_2660,N_772);
and U5305 (N_5305,N_4503,N_2497);
and U5306 (N_5306,N_3949,N_4957);
nor U5307 (N_5307,N_2468,N_2596);
and U5308 (N_5308,N_3837,N_3386);
and U5309 (N_5309,N_577,N_3368);
or U5310 (N_5310,N_4139,N_299);
xnor U5311 (N_5311,N_4126,N_3182);
or U5312 (N_5312,N_2484,N_3253);
and U5313 (N_5313,N_4054,N_2367);
nand U5314 (N_5314,N_633,N_2004);
and U5315 (N_5315,N_3526,N_3487);
nor U5316 (N_5316,N_2423,N_3764);
nand U5317 (N_5317,N_778,N_3615);
or U5318 (N_5318,N_4180,N_1218);
nand U5319 (N_5319,N_3960,N_2449);
xor U5320 (N_5320,N_1047,N_3591);
and U5321 (N_5321,N_2255,N_639);
or U5322 (N_5322,N_1873,N_225);
or U5323 (N_5323,N_3986,N_3464);
nor U5324 (N_5324,N_661,N_3696);
nor U5325 (N_5325,N_4301,N_3225);
and U5326 (N_5326,N_327,N_3472);
and U5327 (N_5327,N_3650,N_1706);
or U5328 (N_5328,N_3054,N_1551);
nand U5329 (N_5329,N_4603,N_1262);
nor U5330 (N_5330,N_535,N_3801);
nand U5331 (N_5331,N_3102,N_2940);
and U5332 (N_5332,N_4548,N_258);
xor U5333 (N_5333,N_1137,N_1952);
nand U5334 (N_5334,N_2135,N_3447);
nor U5335 (N_5335,N_4102,N_3604);
nand U5336 (N_5336,N_2540,N_2385);
nor U5337 (N_5337,N_4165,N_1849);
and U5338 (N_5338,N_3420,N_4151);
nand U5339 (N_5339,N_272,N_3496);
and U5340 (N_5340,N_3367,N_3715);
nor U5341 (N_5341,N_2486,N_965);
and U5342 (N_5342,N_3270,N_4622);
and U5343 (N_5343,N_4573,N_2871);
nor U5344 (N_5344,N_4191,N_1583);
nor U5345 (N_5345,N_390,N_4676);
nand U5346 (N_5346,N_4618,N_3873);
nand U5347 (N_5347,N_2167,N_3096);
or U5348 (N_5348,N_3064,N_1318);
or U5349 (N_5349,N_3625,N_739);
nor U5350 (N_5350,N_4862,N_1997);
nor U5351 (N_5351,N_4365,N_3083);
or U5352 (N_5352,N_4861,N_1670);
nor U5353 (N_5353,N_3435,N_2321);
and U5354 (N_5354,N_117,N_3842);
nor U5355 (N_5355,N_2766,N_2464);
and U5356 (N_5356,N_4017,N_517);
nor U5357 (N_5357,N_546,N_1048);
and U5358 (N_5358,N_173,N_1182);
and U5359 (N_5359,N_1105,N_4539);
nand U5360 (N_5360,N_4640,N_2780);
and U5361 (N_5361,N_4169,N_149);
and U5362 (N_5362,N_3778,N_3661);
nand U5363 (N_5363,N_2158,N_3569);
nor U5364 (N_5364,N_1672,N_262);
or U5365 (N_5365,N_1483,N_1371);
or U5366 (N_5366,N_1465,N_590);
and U5367 (N_5367,N_3900,N_3652);
xnor U5368 (N_5368,N_698,N_4172);
and U5369 (N_5369,N_3897,N_2705);
nor U5370 (N_5370,N_3766,N_4991);
nand U5371 (N_5371,N_3867,N_3785);
nand U5372 (N_5372,N_3959,N_1183);
xor U5373 (N_5373,N_2277,N_2930);
nand U5374 (N_5374,N_899,N_2275);
nor U5375 (N_5375,N_4988,N_2977);
nor U5376 (N_5376,N_548,N_3562);
nand U5377 (N_5377,N_2006,N_1998);
and U5378 (N_5378,N_1288,N_969);
xnor U5379 (N_5379,N_1831,N_1066);
nor U5380 (N_5380,N_3999,N_4918);
or U5381 (N_5381,N_1664,N_3180);
and U5382 (N_5382,N_1886,N_1127);
or U5383 (N_5383,N_2627,N_3932);
nor U5384 (N_5384,N_530,N_397);
and U5385 (N_5385,N_387,N_335);
nand U5386 (N_5386,N_860,N_3058);
or U5387 (N_5387,N_3295,N_1304);
and U5388 (N_5388,N_2274,N_3044);
xnor U5389 (N_5389,N_4479,N_1466);
nor U5390 (N_5390,N_4759,N_2237);
nor U5391 (N_5391,N_4413,N_453);
nand U5392 (N_5392,N_3039,N_1193);
and U5393 (N_5393,N_19,N_3040);
or U5394 (N_5394,N_3275,N_2562);
nand U5395 (N_5395,N_3841,N_4524);
nor U5396 (N_5396,N_3574,N_1533);
nand U5397 (N_5397,N_1035,N_2363);
nand U5398 (N_5398,N_4050,N_1444);
and U5399 (N_5399,N_1949,N_4450);
nand U5400 (N_5400,N_4391,N_1513);
and U5401 (N_5401,N_4745,N_433);
or U5402 (N_5402,N_2267,N_168);
nor U5403 (N_5403,N_818,N_1);
nand U5404 (N_5404,N_1126,N_4124);
or U5405 (N_5405,N_1823,N_3442);
and U5406 (N_5406,N_4084,N_3890);
nand U5407 (N_5407,N_219,N_2042);
and U5408 (N_5408,N_1203,N_804);
nor U5409 (N_5409,N_3432,N_3237);
nor U5410 (N_5410,N_873,N_2760);
nand U5411 (N_5411,N_647,N_968);
nand U5412 (N_5412,N_3259,N_3281);
or U5413 (N_5413,N_2984,N_1272);
nand U5414 (N_5414,N_4040,N_3674);
or U5415 (N_5415,N_2348,N_2033);
nor U5416 (N_5416,N_3082,N_2552);
or U5417 (N_5417,N_4161,N_3885);
nor U5418 (N_5418,N_3541,N_2375);
nor U5419 (N_5419,N_2535,N_4441);
nand U5420 (N_5420,N_1646,N_4774);
nor U5421 (N_5421,N_1291,N_3400);
nand U5422 (N_5422,N_745,N_2691);
nor U5423 (N_5423,N_3355,N_3427);
and U5424 (N_5424,N_3371,N_3919);
or U5425 (N_5425,N_2488,N_2605);
and U5426 (N_5426,N_1611,N_2163);
or U5427 (N_5427,N_3707,N_1324);
and U5428 (N_5428,N_1956,N_1383);
nand U5429 (N_5429,N_2067,N_3660);
or U5430 (N_5430,N_4892,N_3140);
nand U5431 (N_5431,N_304,N_4000);
or U5432 (N_5432,N_3691,N_324);
and U5433 (N_5433,N_3459,N_3752);
xor U5434 (N_5434,N_815,N_3947);
nand U5435 (N_5435,N_3703,N_34);
and U5436 (N_5436,N_4007,N_2564);
or U5437 (N_5437,N_1704,N_875);
or U5438 (N_5438,N_24,N_2178);
or U5439 (N_5439,N_2115,N_3336);
or U5440 (N_5440,N_2697,N_3678);
nand U5441 (N_5441,N_4372,N_4644);
and U5442 (N_5442,N_3186,N_3803);
and U5443 (N_5443,N_3874,N_1196);
nand U5444 (N_5444,N_631,N_470);
nor U5445 (N_5445,N_2320,N_1198);
nor U5446 (N_5446,N_1960,N_2060);
or U5447 (N_5447,N_1311,N_4516);
or U5448 (N_5448,N_1049,N_1534);
or U5449 (N_5449,N_2522,N_4529);
nand U5450 (N_5450,N_520,N_1434);
nor U5451 (N_5451,N_1092,N_350);
or U5452 (N_5452,N_2809,N_4341);
nor U5453 (N_5453,N_1504,N_3298);
nor U5454 (N_5454,N_4527,N_1367);
and U5455 (N_5455,N_2920,N_2238);
and U5456 (N_5456,N_3513,N_2136);
nor U5457 (N_5457,N_3405,N_3504);
nor U5458 (N_5458,N_3230,N_1179);
nand U5459 (N_5459,N_3878,N_3256);
nor U5460 (N_5460,N_753,N_2979);
xor U5461 (N_5461,N_3178,N_277);
and U5462 (N_5462,N_106,N_690);
or U5463 (N_5463,N_2401,N_3583);
nand U5464 (N_5464,N_781,N_4369);
and U5465 (N_5465,N_4995,N_3219);
nor U5466 (N_5466,N_4075,N_4351);
and U5467 (N_5467,N_1452,N_1292);
nand U5468 (N_5468,N_348,N_3346);
nand U5469 (N_5469,N_992,N_4753);
xor U5470 (N_5470,N_3776,N_3791);
or U5471 (N_5471,N_4668,N_4684);
or U5472 (N_5472,N_3060,N_2197);
or U5473 (N_5473,N_4123,N_2877);
nor U5474 (N_5474,N_1966,N_2895);
nor U5475 (N_5475,N_1308,N_4357);
nor U5476 (N_5476,N_11,N_3970);
nand U5477 (N_5477,N_742,N_4173);
nand U5478 (N_5478,N_83,N_1115);
nand U5479 (N_5479,N_115,N_1213);
nor U5480 (N_5480,N_1437,N_730);
xor U5481 (N_5481,N_913,N_1525);
and U5482 (N_5482,N_3086,N_3217);
nor U5483 (N_5483,N_3104,N_916);
nand U5484 (N_5484,N_1441,N_926);
nor U5485 (N_5485,N_4325,N_1374);
nand U5486 (N_5486,N_4675,N_1537);
nor U5487 (N_5487,N_583,N_4069);
nand U5488 (N_5488,N_4133,N_4170);
and U5489 (N_5489,N_1424,N_4600);
or U5490 (N_5490,N_1718,N_572);
nand U5491 (N_5491,N_3198,N_876);
nor U5492 (N_5492,N_2559,N_4893);
or U5493 (N_5493,N_3740,N_3103);
and U5494 (N_5494,N_4002,N_4758);
or U5495 (N_5495,N_1109,N_3005);
and U5496 (N_5496,N_3988,N_935);
nand U5497 (N_5497,N_2201,N_2107);
nand U5498 (N_5498,N_2771,N_886);
or U5499 (N_5499,N_2541,N_4510);
or U5500 (N_5500,N_2602,N_2399);
or U5501 (N_5501,N_2196,N_4789);
nor U5502 (N_5502,N_756,N_1809);
nand U5503 (N_5503,N_105,N_2473);
or U5504 (N_5504,N_1856,N_2495);
nand U5505 (N_5505,N_4842,N_2180);
nor U5506 (N_5506,N_4665,N_4038);
xor U5507 (N_5507,N_1217,N_1265);
nand U5508 (N_5508,N_1751,N_3659);
nand U5509 (N_5509,N_4740,N_1089);
xnor U5510 (N_5510,N_4559,N_4097);
nand U5511 (N_5511,N_810,N_1457);
or U5512 (N_5512,N_2137,N_3961);
nand U5513 (N_5513,N_4318,N_3642);
and U5514 (N_5514,N_2204,N_4925);
and U5515 (N_5515,N_1135,N_1599);
or U5516 (N_5516,N_1945,N_1484);
or U5517 (N_5517,N_1632,N_2489);
xor U5518 (N_5518,N_1393,N_2007);
nor U5519 (N_5519,N_4344,N_990);
and U5520 (N_5520,N_2776,N_1912);
and U5521 (N_5521,N_2020,N_4896);
nand U5522 (N_5522,N_1894,N_3220);
nand U5523 (N_5523,N_1240,N_1724);
and U5524 (N_5524,N_2626,N_2892);
nor U5525 (N_5525,N_538,N_1470);
or U5526 (N_5526,N_1046,N_3193);
or U5527 (N_5527,N_3244,N_906);
nand U5528 (N_5528,N_1509,N_602);
and U5529 (N_5529,N_3859,N_1619);
and U5530 (N_5530,N_4697,N_344);
and U5531 (N_5531,N_880,N_4838);
nor U5532 (N_5532,N_986,N_1645);
or U5533 (N_5533,N_626,N_2156);
and U5534 (N_5534,N_1660,N_4074);
and U5535 (N_5535,N_2099,N_960);
nor U5536 (N_5536,N_4846,N_3992);
nor U5537 (N_5537,N_3843,N_3907);
and U5538 (N_5538,N_54,N_4581);
nand U5539 (N_5539,N_338,N_3538);
nor U5540 (N_5540,N_4673,N_3047);
nand U5541 (N_5541,N_449,N_3467);
nor U5542 (N_5542,N_4694,N_991);
nor U5543 (N_5543,N_4816,N_3543);
or U5544 (N_5544,N_75,N_4755);
and U5545 (N_5545,N_236,N_2112);
nor U5546 (N_5546,N_3138,N_3135);
xnor U5547 (N_5547,N_3533,N_890);
nand U5548 (N_5548,N_1536,N_3098);
nor U5549 (N_5549,N_2476,N_2808);
nand U5550 (N_5550,N_4518,N_30);
nand U5551 (N_5551,N_4427,N_151);
nor U5552 (N_5552,N_857,N_3302);
nor U5553 (N_5553,N_1505,N_2788);
and U5554 (N_5554,N_1248,N_1920);
and U5555 (N_5555,N_1630,N_891);
and U5556 (N_5556,N_3584,N_2680);
and U5557 (N_5557,N_2448,N_2721);
or U5558 (N_5558,N_2542,N_1896);
and U5559 (N_5559,N_2900,N_3836);
xor U5560 (N_5560,N_4791,N_1699);
or U5561 (N_5561,N_752,N_487);
and U5562 (N_5562,N_1012,N_4685);
nor U5563 (N_5563,N_2667,N_719);
and U5564 (N_5564,N_3974,N_2641);
xor U5565 (N_5565,N_1869,N_3729);
nand U5566 (N_5566,N_223,N_4282);
nor U5567 (N_5567,N_4628,N_1587);
nor U5568 (N_5568,N_1910,N_1363);
or U5569 (N_5569,N_1766,N_1093);
or U5570 (N_5570,N_2948,N_180);
or U5571 (N_5571,N_3278,N_2461);
and U5572 (N_5572,N_2499,N_4033);
or U5573 (N_5573,N_3249,N_127);
or U5574 (N_5574,N_4606,N_2939);
nand U5575 (N_5575,N_1352,N_1022);
or U5576 (N_5576,N_1889,N_741);
or U5577 (N_5577,N_2707,N_2256);
and U5578 (N_5578,N_4423,N_2029);
or U5579 (N_5579,N_1481,N_3594);
nor U5580 (N_5580,N_2720,N_4526);
and U5581 (N_5581,N_4961,N_142);
nor U5582 (N_5582,N_4034,N_3306);
or U5583 (N_5583,N_3687,N_4627);
and U5584 (N_5584,N_435,N_1643);
nand U5585 (N_5585,N_4511,N_4979);
nand U5586 (N_5586,N_2730,N_879);
and U5587 (N_5587,N_1340,N_4176);
or U5588 (N_5588,N_2314,N_531);
nand U5589 (N_5589,N_1013,N_912);
and U5590 (N_5590,N_1733,N_3503);
nand U5591 (N_5591,N_3706,N_4175);
nor U5592 (N_5592,N_1171,N_907);
nand U5593 (N_5593,N_3711,N_4835);
nor U5594 (N_5594,N_3667,N_2785);
or U5595 (N_5595,N_2377,N_3068);
or U5596 (N_5596,N_289,N_2512);
nand U5597 (N_5597,N_4980,N_3279);
nor U5598 (N_5598,N_3164,N_3255);
and U5599 (N_5599,N_625,N_764);
or U5600 (N_5600,N_1494,N_4268);
nand U5601 (N_5601,N_1637,N_834);
or U5602 (N_5602,N_4617,N_4026);
and U5603 (N_5603,N_4661,N_4240);
and U5604 (N_5604,N_2190,N_4315);
nor U5605 (N_5605,N_363,N_16);
nor U5606 (N_5606,N_950,N_1697);
nor U5607 (N_5607,N_4397,N_4140);
nand U5608 (N_5608,N_4592,N_4431);
and U5609 (N_5609,N_4945,N_4967);
and U5610 (N_5610,N_4822,N_51);
or U5611 (N_5611,N_1651,N_2427);
nand U5612 (N_5612,N_2834,N_675);
nor U5613 (N_5613,N_1345,N_3321);
and U5614 (N_5614,N_1691,N_1813);
or U5615 (N_5615,N_584,N_819);
or U5616 (N_5616,N_953,N_2432);
and U5617 (N_5617,N_3902,N_1933);
nor U5618 (N_5618,N_3777,N_2807);
xor U5619 (N_5619,N_4800,N_1571);
or U5620 (N_5620,N_2368,N_3922);
nor U5621 (N_5621,N_1300,N_4238);
nor U5622 (N_5622,N_3665,N_4155);
and U5623 (N_5623,N_3937,N_700);
or U5624 (N_5624,N_2373,N_1118);
and U5625 (N_5625,N_4202,N_2635);
and U5626 (N_5626,N_2569,N_3522);
nand U5627 (N_5627,N_2594,N_4797);
or U5628 (N_5628,N_1832,N_4860);
nor U5629 (N_5629,N_4922,N_858);
nand U5630 (N_5630,N_2563,N_382);
nand U5631 (N_5631,N_3597,N_1435);
and U5632 (N_5632,N_3954,N_1125);
and U5633 (N_5633,N_1946,N_1067);
or U5634 (N_5634,N_2783,N_3751);
nor U5635 (N_5635,N_2854,N_2964);
or U5636 (N_5636,N_4387,N_4251);
and U5637 (N_5637,N_706,N_727);
nor U5638 (N_5638,N_4636,N_1150);
nand U5639 (N_5639,N_1687,N_2173);
nor U5640 (N_5640,N_3500,N_3101);
or U5641 (N_5641,N_4306,N_434);
or U5642 (N_5642,N_4761,N_3893);
and U5643 (N_5643,N_920,N_1707);
or U5644 (N_5644,N_3117,N_2567);
or U5645 (N_5645,N_4574,N_1541);
nand U5646 (N_5646,N_2339,N_1499);
nand U5647 (N_5647,N_1756,N_2700);
nor U5648 (N_5648,N_3489,N_2915);
nand U5649 (N_5649,N_4189,N_2400);
nor U5650 (N_5650,N_17,N_2200);
nand U5651 (N_5651,N_1251,N_3134);
and U5652 (N_5652,N_1007,N_650);
nand U5653 (N_5653,N_1951,N_154);
nand U5654 (N_5654,N_259,N_654);
or U5655 (N_5655,N_4642,N_4285);
or U5656 (N_5656,N_3417,N_1267);
nand U5657 (N_5657,N_2165,N_523);
and U5658 (N_5658,N_39,N_697);
nand U5659 (N_5659,N_1527,N_3157);
nand U5660 (N_5660,N_2182,N_3161);
nor U5661 (N_5661,N_2784,N_3262);
or U5662 (N_5662,N_1502,N_2819);
or U5663 (N_5663,N_3990,N_3199);
or U5664 (N_5664,N_4578,N_2590);
and U5665 (N_5665,N_2301,N_952);
and U5666 (N_5666,N_2799,N_4210);
nand U5667 (N_5667,N_785,N_1430);
nand U5668 (N_5668,N_184,N_3518);
or U5669 (N_5669,N_3601,N_4451);
xor U5670 (N_5670,N_3415,N_4702);
and U5671 (N_5671,N_2850,N_3976);
and U5672 (N_5672,N_4930,N_3539);
nand U5673 (N_5673,N_1398,N_4895);
nand U5674 (N_5674,N_2413,N_2472);
nor U5675 (N_5675,N_1963,N_1907);
nor U5676 (N_5676,N_3258,N_2162);
nor U5677 (N_5677,N_4402,N_2847);
nand U5678 (N_5678,N_1904,N_4382);
nor U5679 (N_5679,N_3532,N_3042);
xnor U5680 (N_5680,N_2736,N_4942);
or U5681 (N_5681,N_2232,N_4208);
xor U5682 (N_5682,N_1192,N_2996);
or U5683 (N_5683,N_844,N_1554);
and U5684 (N_5684,N_869,N_1338);
nor U5685 (N_5685,N_4489,N_1623);
nand U5686 (N_5686,N_3046,N_3644);
and U5687 (N_5687,N_3197,N_4009);
or U5688 (N_5688,N_3001,N_361);
nand U5689 (N_5689,N_4514,N_2722);
and U5690 (N_5690,N_2233,N_3536);
nand U5691 (N_5691,N_4300,N_1320);
xor U5692 (N_5692,N_1266,N_1540);
nand U5693 (N_5693,N_710,N_643);
nor U5694 (N_5694,N_2487,N_2800);
and U5695 (N_5695,N_3166,N_808);
nor U5696 (N_5696,N_3573,N_2687);
and U5697 (N_5697,N_1467,N_1787);
nand U5698 (N_5698,N_1252,N_3738);
nand U5699 (N_5699,N_27,N_2709);
or U5700 (N_5700,N_954,N_2409);
or U5701 (N_5701,N_3196,N_411);
and U5702 (N_5702,N_477,N_2582);
nand U5703 (N_5703,N_2207,N_4312);
nand U5704 (N_5704,N_2553,N_1516);
nand U5705 (N_5705,N_2530,N_3593);
nor U5706 (N_5706,N_3312,N_1165);
nor U5707 (N_5707,N_998,N_265);
nor U5708 (N_5708,N_4679,N_3204);
nand U5709 (N_5709,N_4643,N_4505);
nand U5710 (N_5710,N_2069,N_1286);
or U5711 (N_5711,N_3233,N_4030);
and U5712 (N_5712,N_1803,N_1898);
and U5713 (N_5713,N_2815,N_2778);
nand U5714 (N_5714,N_3308,N_1913);
or U5715 (N_5715,N_4159,N_1350);
and U5716 (N_5716,N_3957,N_3779);
and U5717 (N_5717,N_3737,N_4198);
nor U5718 (N_5718,N_3657,N_832);
nor U5719 (N_5719,N_2947,N_2728);
or U5720 (N_5720,N_4543,N_3069);
or U5721 (N_5721,N_1027,N_2175);
and U5722 (N_5722,N_3352,N_4805);
and U5723 (N_5723,N_904,N_2685);
or U5724 (N_5724,N_278,N_3465);
or U5725 (N_5725,N_4259,N_2191);
xnor U5726 (N_5726,N_3067,N_3050);
nand U5727 (N_5727,N_540,N_2992);
nand U5728 (N_5728,N_4241,N_2995);
and U5729 (N_5729,N_2518,N_2599);
and U5730 (N_5730,N_1957,N_3359);
or U5731 (N_5731,N_4607,N_1711);
or U5732 (N_5732,N_4782,N_852);
and U5733 (N_5733,N_2284,N_4817);
and U5734 (N_5734,N_1033,N_2052);
nor U5735 (N_5735,N_787,N_3699);
or U5736 (N_5736,N_1705,N_3868);
nand U5737 (N_5737,N_228,N_4635);
nand U5738 (N_5738,N_1405,N_3426);
nor U5739 (N_5739,N_1010,N_2051);
nand U5740 (N_5740,N_2205,N_4031);
nor U5741 (N_5741,N_1784,N_1221);
nor U5742 (N_5742,N_2089,N_1408);
and U5743 (N_5743,N_2319,N_3494);
nor U5744 (N_5744,N_3232,N_2406);
and U5745 (N_5745,N_3863,N_2682);
nand U5746 (N_5746,N_276,N_4616);
or U5747 (N_5747,N_1369,N_4024);
or U5748 (N_5748,N_1674,N_80);
and U5749 (N_5749,N_2584,N_357);
or U5750 (N_5750,N_2229,N_2899);
nor U5751 (N_5751,N_829,N_2978);
nand U5752 (N_5752,N_2362,N_3356);
nor U5753 (N_5753,N_3553,N_3207);
or U5754 (N_5754,N_3525,N_888);
nand U5755 (N_5755,N_120,N_356);
or U5756 (N_5756,N_1215,N_896);
and U5757 (N_5757,N_2379,N_1391);
or U5758 (N_5758,N_4338,N_2802);
or U5759 (N_5759,N_7,N_4436);
nand U5760 (N_5760,N_902,N_3438);
or U5761 (N_5761,N_2333,N_4778);
or U5762 (N_5762,N_4827,N_2898);
nand U5763 (N_5763,N_1487,N_861);
or U5764 (N_5764,N_208,N_1223);
or U5765 (N_5765,N_3482,N_4214);
nor U5766 (N_5766,N_365,N_4468);
nand U5767 (N_5767,N_455,N_578);
nor U5768 (N_5768,N_3153,N_58);
xnor U5769 (N_5769,N_4531,N_1415);
nor U5770 (N_5770,N_599,N_3109);
and U5771 (N_5771,N_3462,N_1296);
or U5772 (N_5772,N_3423,N_526);
nor U5773 (N_5773,N_4305,N_4594);
nor U5774 (N_5774,N_307,N_1544);
xnor U5775 (N_5775,N_3690,N_2625);
and U5776 (N_5776,N_3120,N_766);
nor U5777 (N_5777,N_4244,N_708);
and U5778 (N_5778,N_498,N_337);
or U5779 (N_5779,N_21,N_1138);
and U5780 (N_5780,N_1725,N_2063);
and U5781 (N_5781,N_1339,N_2094);
and U5782 (N_5782,N_981,N_1469);
and U5783 (N_5783,N_2937,N_1713);
nand U5784 (N_5784,N_3333,N_509);
nand U5785 (N_5785,N_462,N_3452);
nand U5786 (N_5786,N_3283,N_2934);
xnor U5787 (N_5787,N_3631,N_4711);
or U5788 (N_5788,N_4236,N_1759);
nand U5789 (N_5789,N_3587,N_4560);
nand U5790 (N_5790,N_1567,N_1407);
and U5791 (N_5791,N_1496,N_3763);
or U5792 (N_5792,N_181,N_938);
or U5793 (N_5793,N_2103,N_1372);
nor U5794 (N_5794,N_29,N_738);
nand U5795 (N_5795,N_3409,N_4071);
and U5796 (N_5796,N_4366,N_32);
or U5797 (N_5797,N_1719,N_667);
nand U5798 (N_5798,N_4334,N_593);
nor U5799 (N_5799,N_2887,N_4856);
or U5800 (N_5800,N_4847,N_1841);
and U5801 (N_5801,N_1727,N_2748);
and U5802 (N_5802,N_267,N_1720);
nor U5803 (N_5803,N_1019,N_4955);
nor U5804 (N_5804,N_4844,N_724);
xor U5805 (N_5805,N_4597,N_3546);
or U5806 (N_5806,N_958,N_2492);
nor U5807 (N_5807,N_2011,N_1638);
and U5808 (N_5808,N_3603,N_1431);
nand U5809 (N_5809,N_239,N_2671);
nand U5810 (N_5810,N_192,N_4478);
nand U5811 (N_5811,N_2282,N_2095);
nand U5812 (N_5812,N_1827,N_760);
nand U5813 (N_5813,N_2546,N_1476);
nand U5814 (N_5814,N_3748,N_4356);
nor U5815 (N_5815,N_2259,N_4584);
and U5816 (N_5816,N_97,N_147);
and U5817 (N_5817,N_1594,N_3984);
and U5818 (N_5818,N_3991,N_709);
nor U5819 (N_5819,N_4442,N_2134);
or U5820 (N_5820,N_4686,N_1557);
nand U5821 (N_5821,N_2938,N_4973);
or U5822 (N_5822,N_3350,N_384);
nor U5823 (N_5823,N_1175,N_4485);
nand U5824 (N_5824,N_329,N_4512);
nand U5825 (N_5825,N_1835,N_4887);
nand U5826 (N_5826,N_4951,N_4396);
nand U5827 (N_5827,N_28,N_4096);
nand U5828 (N_5828,N_134,N_1401);
or U5829 (N_5829,N_1822,N_3339);
and U5830 (N_5830,N_4149,N_2746);
nor U5831 (N_5831,N_1736,N_881);
and U5832 (N_5832,N_183,N_2053);
nor U5833 (N_5833,N_4435,N_4373);
or U5834 (N_5834,N_1354,N_1927);
and U5835 (N_5835,N_3647,N_2818);
nor U5836 (N_5836,N_4536,N_4390);
and U5837 (N_5837,N_268,N_2210);
or U5838 (N_5838,N_2001,N_2604);
and U5839 (N_5839,N_1863,N_1478);
and U5840 (N_5840,N_966,N_4274);
or U5841 (N_5841,N_1280,N_4443);
nor U5842 (N_5842,N_2610,N_2132);
nand U5843 (N_5843,N_4806,N_2653);
nor U5844 (N_5844,N_4342,N_3662);
nor U5845 (N_5845,N_1947,N_989);
and U5846 (N_5846,N_628,N_1942);
and U5847 (N_5847,N_2389,N_14);
nand U5848 (N_5848,N_4716,N_2620);
or U5849 (N_5849,N_3181,N_883);
and U5850 (N_5850,N_3151,N_408);
nand U5851 (N_5851,N_2853,N_401);
or U5852 (N_5852,N_3338,N_821);
nor U5853 (N_5853,N_197,N_1610);
and U5854 (N_5854,N_2214,N_3720);
and U5855 (N_5855,N_2265,N_4062);
or U5856 (N_5856,N_2836,N_2616);
or U5857 (N_5857,N_3956,N_1906);
or U5858 (N_5858,N_4998,N_1445);
nor U5859 (N_5859,N_3917,N_474);
or U5860 (N_5860,N_3030,N_2485);
or U5861 (N_5861,N_2096,N_2617);
nor U5862 (N_5862,N_3263,N_3499);
nor U5863 (N_5863,N_20,N_78);
and U5864 (N_5864,N_831,N_4771);
or U5865 (N_5865,N_1984,N_1382);
and U5866 (N_5866,N_1501,N_2860);
nand U5867 (N_5867,N_2549,N_1754);
nor U5868 (N_5868,N_1604,N_4598);
xor U5869 (N_5869,N_2208,N_3299);
or U5870 (N_5870,N_1974,N_4743);
nand U5871 (N_5871,N_2285,N_3857);
nor U5872 (N_5872,N_1885,N_3108);
and U5873 (N_5873,N_1686,N_893);
or U5874 (N_5874,N_176,N_3805);
and U5875 (N_5875,N_4765,N_378);
nor U5876 (N_5876,N_4378,N_1325);
nand U5877 (N_5877,N_4615,N_3814);
or U5878 (N_5878,N_4420,N_1529);
nand U5879 (N_5879,N_373,N_3571);
nor U5880 (N_5880,N_4564,N_351);
or U5881 (N_5881,N_3971,N_1322);
nor U5882 (N_5882,N_1448,N_4354);
and U5883 (N_5883,N_3183,N_4876);
nand U5884 (N_5884,N_1269,N_3797);
nand U5885 (N_5885,N_3879,N_2644);
or U5886 (N_5886,N_3403,N_3443);
and U5887 (N_5887,N_250,N_4141);
or U5888 (N_5888,N_2500,N_3130);
or U5889 (N_5889,N_1714,N_4381);
or U5890 (N_5890,N_2092,N_424);
nand U5891 (N_5891,N_560,N_4353);
or U5892 (N_5892,N_985,N_4515);
nand U5893 (N_5893,N_3951,N_889);
and U5894 (N_5894,N_2452,N_1355);
or U5895 (N_5895,N_2477,N_206);
nand U5896 (N_5896,N_783,N_3478);
or U5897 (N_5897,N_3558,N_980);
and U5898 (N_5898,N_2073,N_2827);
nand U5899 (N_5899,N_1734,N_4493);
xor U5900 (N_5900,N_218,N_3332);
nand U5901 (N_5901,N_2843,N_2026);
and U5902 (N_5902,N_3114,N_668);
nand U5903 (N_5903,N_3505,N_1036);
or U5904 (N_5904,N_3294,N_1462);
nand U5905 (N_5905,N_1103,N_488);
nand U5906 (N_5906,N_3870,N_3017);
nor U5907 (N_5907,N_1991,N_1053);
nor U5908 (N_5908,N_1409,N_332);
nand U5909 (N_5909,N_1123,N_4042);
and U5910 (N_5910,N_1302,N_3052);
or U5911 (N_5911,N_3079,N_3926);
nand U5912 (N_5912,N_4744,N_1185);
and U5913 (N_5913,N_2645,N_288);
or U5914 (N_5914,N_1001,N_42);
and U5915 (N_5915,N_3903,N_359);
and U5916 (N_5916,N_693,N_1819);
or U5917 (N_5917,N_2603,N_1479);
nand U5918 (N_5918,N_1456,N_235);
nand U5919 (N_5919,N_1034,N_3586);
xnor U5920 (N_5920,N_1764,N_4784);
nor U5921 (N_5921,N_436,N_458);
nand U5922 (N_5922,N_1936,N_2122);
or U5923 (N_5923,N_1807,N_1675);
nor U5924 (N_5924,N_3639,N_4474);
nor U5925 (N_5925,N_3928,N_2634);
or U5926 (N_5926,N_521,N_98);
and U5927 (N_5927,N_2960,N_379);
nor U5928 (N_5928,N_1167,N_3948);
nor U5929 (N_5929,N_4188,N_4848);
nor U5930 (N_5930,N_2460,N_4407);
nor U5931 (N_5931,N_3329,N_2036);
and U5932 (N_5932,N_1285,N_71);
nand U5933 (N_5933,N_1037,N_3326);
and U5934 (N_5934,N_1615,N_1261);
or U5935 (N_5935,N_2969,N_3242);
or U5936 (N_5936,N_292,N_3431);
nor U5937 (N_5937,N_4779,N_3498);
and U5938 (N_5938,N_3418,N_3936);
xor U5939 (N_5939,N_1124,N_282);
or U5940 (N_5940,N_3886,N_3906);
nor U5941 (N_5941,N_3072,N_2739);
nand U5942 (N_5942,N_2662,N_824);
nand U5943 (N_5943,N_2828,N_2085);
nor U5944 (N_5944,N_2989,N_3643);
nor U5945 (N_5945,N_4001,N_3126);
nand U5946 (N_5946,N_4106,N_43);
or U5947 (N_5947,N_3572,N_1609);
nand U5948 (N_5948,N_776,N_3385);
or U5949 (N_5949,N_4936,N_1426);
and U5950 (N_5950,N_88,N_2885);
and U5951 (N_5951,N_1753,N_2798);
nor U5952 (N_5952,N_2575,N_2548);
and U5953 (N_5953,N_3798,N_544);
nand U5954 (N_5954,N_4752,N_4379);
nor U5955 (N_5955,N_2515,N_4611);
nor U5956 (N_5956,N_3407,N_1459);
or U5957 (N_5957,N_280,N_504);
nand U5958 (N_5958,N_704,N_1000);
and U5959 (N_5959,N_4693,N_1422);
or U5960 (N_5960,N_4775,N_430);
or U5961 (N_5961,N_2514,N_3668);
and U5962 (N_5962,N_286,N_3074);
or U5963 (N_5963,N_1247,N_2765);
and U5964 (N_5964,N_1988,N_393);
nand U5965 (N_5965,N_4225,N_3983);
and U5966 (N_5966,N_539,N_846);
nand U5967 (N_5967,N_1143,N_4956);
and U5968 (N_5968,N_4582,N_1605);
or U5969 (N_5969,N_2629,N_301);
nand U5970 (N_5970,N_3461,N_3335);
or U5971 (N_5971,N_1229,N_2554);
or U5972 (N_5972,N_3425,N_266);
and U5973 (N_5973,N_604,N_2370);
nand U5974 (N_5974,N_50,N_877);
or U5975 (N_5975,N_2529,N_4649);
or U5976 (N_5976,N_2975,N_3486);
nand U5977 (N_5977,N_269,N_2639);
or U5978 (N_5978,N_2507,N_4185);
or U5979 (N_5979,N_971,N_1358);
nor U5980 (N_5980,N_1121,N_1722);
nand U5981 (N_5981,N_2801,N_4105);
nor U5982 (N_5982,N_932,N_685);
nand U5983 (N_5983,N_84,N_406);
nand U5984 (N_5984,N_1500,N_3112);
and U5985 (N_5985,N_3325,N_1458);
nor U5986 (N_5986,N_1573,N_1246);
nor U5987 (N_5987,N_4507,N_1845);
or U5988 (N_5988,N_2914,N_3471);
and U5989 (N_5989,N_2750,N_1160);
nor U5990 (N_5990,N_849,N_2431);
nor U5991 (N_5991,N_4003,N_716);
or U5992 (N_5992,N_4987,N_203);
or U5993 (N_5993,N_1085,N_3148);
nand U5994 (N_5994,N_3009,N_2656);
or U5995 (N_5995,N_3819,N_3972);
nand U5996 (N_5996,N_1159,N_1316);
or U5997 (N_5997,N_2712,N_260);
and U5998 (N_5998,N_1728,N_2747);
or U5999 (N_5999,N_3853,N_3179);
nor U6000 (N_6000,N_4999,N_2234);
nor U6001 (N_6001,N_4832,N_1954);
nand U6002 (N_6002,N_4855,N_1879);
and U6003 (N_6003,N_4361,N_3348);
nor U6004 (N_6004,N_2615,N_3437);
and U6005 (N_6005,N_4027,N_290);
and U6006 (N_6006,N_191,N_3414);
or U6007 (N_6007,N_3226,N_1943);
nand U6008 (N_6008,N_1802,N_2544);
nor U6009 (N_6009,N_2754,N_4840);
nand U6010 (N_6010,N_2408,N_4331);
and U6011 (N_6011,N_1909,N_146);
nand U6012 (N_6012,N_1507,N_3274);
or U6013 (N_6013,N_744,N_3955);
or U6014 (N_6014,N_3272,N_2896);
or U6015 (N_6015,N_2878,N_4051);
nand U6016 (N_6016,N_4795,N_2337);
or U6017 (N_6017,N_200,N_2858);
or U6018 (N_6018,N_4047,N_2568);
nand U6019 (N_6019,N_4586,N_1673);
nand U6020 (N_6020,N_4544,N_4950);
and U6021 (N_6021,N_3094,N_3799);
or U6022 (N_6022,N_4046,N_4815);
or U6023 (N_6023,N_1740,N_4715);
nand U6024 (N_6024,N_4368,N_4246);
nand U6025 (N_6025,N_4181,N_903);
nor U6026 (N_6026,N_1413,N_3782);
or U6027 (N_6027,N_3780,N_1833);
and U6028 (N_6028,N_4913,N_3834);
nor U6029 (N_6029,N_2411,N_2821);
xor U6030 (N_6030,N_4972,N_652);
or U6031 (N_6031,N_4750,N_4293);
nor U6032 (N_6032,N_4811,N_2955);
or U6033 (N_6033,N_2715,N_1814);
nand U6034 (N_6034,N_1360,N_4641);
or U6035 (N_6035,N_1493,N_983);
nand U6036 (N_6036,N_4219,N_2211);
nand U6037 (N_6037,N_4709,N_3817);
and U6038 (N_6038,N_3528,N_3755);
or U6039 (N_6039,N_2829,N_4059);
nand U6040 (N_6040,N_4056,N_4585);
or U6041 (N_6041,N_1341,N_4019);
nor U6042 (N_6042,N_2462,N_476);
nor U6043 (N_6043,N_3627,N_939);
or U6044 (N_6044,N_195,N_4932);
and U6045 (N_6045,N_828,N_855);
and U6046 (N_6046,N_1767,N_3908);
nand U6047 (N_6047,N_4943,N_864);
nand U6048 (N_6048,N_1811,N_3023);
and U6049 (N_6049,N_2945,N_3376);
nor U6050 (N_6050,N_4271,N_2193);
nand U6051 (N_6051,N_838,N_1808);
or U6052 (N_6052,N_640,N_4812);
nand U6053 (N_6053,N_1975,N_910);
and U6054 (N_6054,N_2623,N_4590);
or U6055 (N_6055,N_2478,N_1865);
and U6056 (N_6056,N_2402,N_1878);
nor U6057 (N_6057,N_3202,N_2727);
or U6058 (N_6058,N_2647,N_3610);
xor U6059 (N_6059,N_2463,N_4298);
xor U6060 (N_6060,N_2066,N_961);
or U6061 (N_6061,N_3869,N_4850);
or U6062 (N_6062,N_1081,N_970);
nand U6063 (N_6063,N_475,N_4993);
and U6064 (N_6064,N_111,N_1120);
xor U6065 (N_6065,N_3187,N_140);
nor U6066 (N_6066,N_4360,N_1931);
and U6067 (N_6067,N_210,N_3239);
and U6068 (N_6068,N_137,N_4890);
nand U6069 (N_6069,N_571,N_2738);
nand U6070 (N_6070,N_3977,N_3015);
and U6071 (N_6071,N_2181,N_3760);
or U6072 (N_6072,N_3891,N_4722);
nor U6073 (N_6073,N_4269,N_1601);
or U6074 (N_6074,N_3310,N_2711);
and U6075 (N_6075,N_2300,N_4119);
nand U6076 (N_6076,N_1805,N_749);
xor U6077 (N_6077,N_2246,N_496);
or U6078 (N_6078,N_3304,N_2879);
or U6079 (N_6079,N_4522,N_1317);
or U6080 (N_6080,N_279,N_4869);
and U6081 (N_6081,N_559,N_2047);
nand U6082 (N_6082,N_4883,N_1710);
nand U6083 (N_6083,N_4646,N_1781);
xnor U6084 (N_6084,N_4143,N_2290);
and U6085 (N_6085,N_614,N_516);
and U6086 (N_6086,N_2681,N_4818);
nor U6087 (N_6087,N_3724,N_4283);
and U6088 (N_6088,N_3925,N_2927);
nor U6089 (N_6089,N_2312,N_2723);
or U6090 (N_6090,N_4445,N_2294);
or U6091 (N_6091,N_3404,N_2005);
or U6092 (N_6092,N_1928,N_3783);
nand U6093 (N_6093,N_396,N_3031);
nor U6094 (N_6094,N_3319,N_885);
nand U6095 (N_6095,N_3041,N_2849);
or U6096 (N_6096,N_1696,N_3292);
nand U6097 (N_6097,N_1874,N_1512);
or U6098 (N_6098,N_1480,N_4610);
or U6099 (N_6099,N_3736,N_3492);
nand U6100 (N_6100,N_2901,N_3624);
nor U6101 (N_6101,N_4323,N_240);
nand U6102 (N_6102,N_4645,N_494);
nor U6103 (N_6103,N_4362,N_3675);
nor U6104 (N_6104,N_1812,N_214);
and U6105 (N_6105,N_2672,N_4086);
and U6106 (N_6106,N_4914,N_2904);
xnor U6107 (N_6107,N_3314,N_3635);
and U6108 (N_6108,N_3688,N_2882);
xnor U6109 (N_6109,N_547,N_3953);
or U6110 (N_6110,N_415,N_2994);
or U6111 (N_6111,N_4569,N_3246);
or U6112 (N_6112,N_4599,N_4523);
or U6113 (N_6113,N_2140,N_3614);
and U6114 (N_6114,N_0,N_3714);
or U6115 (N_6115,N_1362,N_1187);
nand U6116 (N_6116,N_2142,N_2601);
xor U6117 (N_6117,N_1968,N_3224);
and U6118 (N_6118,N_2987,N_1062);
nor U6119 (N_6119,N_1695,N_3383);
nor U6120 (N_6120,N_2381,N_736);
nand U6121 (N_6121,N_96,N_377);
nor U6122 (N_6122,N_3307,N_1373);
and U6123 (N_6123,N_144,N_1989);
xnor U6124 (N_6124,N_4053,N_4877);
or U6125 (N_6125,N_4113,N_2322);
and U6126 (N_6126,N_4898,N_3716);
nor U6127 (N_6127,N_699,N_2903);
or U6128 (N_6128,N_3360,N_3579);
nor U6129 (N_6129,N_2174,N_688);
and U6130 (N_6130,N_2944,N_1498);
and U6131 (N_6131,N_659,N_1970);
nand U6132 (N_6132,N_3396,N_1790);
nand U6133 (N_6133,N_3343,N_3318);
or U6134 (N_6134,N_2146,N_4905);
or U6135 (N_6135,N_1029,N_3739);
or U6136 (N_6136,N_4248,N_95);
xor U6137 (N_6137,N_4112,N_4328);
or U6138 (N_6138,N_4623,N_2905);
nand U6139 (N_6139,N_3284,N_245);
or U6140 (N_6140,N_291,N_1847);
and U6141 (N_6141,N_1941,N_1021);
nand U6142 (N_6142,N_1041,N_3481);
and U6143 (N_6143,N_1955,N_1653);
nor U6144 (N_6144,N_315,N_1581);
and U6145 (N_6145,N_4052,N_644);
nand U6146 (N_6146,N_2304,N_2008);
or U6147 (N_6147,N_1996,N_4389);
nand U6148 (N_6148,N_948,N_1818);
nor U6149 (N_6149,N_3630,N_851);
and U6150 (N_6150,N_4377,N_3750);
nor U6151 (N_6151,N_3147,N_1853);
nor U6152 (N_6152,N_2812,N_4909);
and U6153 (N_6153,N_124,N_4205);
nand U6154 (N_6154,N_1575,N_3705);
nor U6155 (N_6155,N_3723,N_2253);
nand U6156 (N_6156,N_4813,N_2228);
or U6157 (N_6157,N_1190,N_1826);
and U6158 (N_6158,N_1597,N_4470);
or U6159 (N_6159,N_2713,N_1486);
nand U6160 (N_6160,N_3252,N_1312);
xor U6161 (N_6161,N_1794,N_3989);
or U6162 (N_6162,N_2317,N_2417);
or U6163 (N_6163,N_1621,N_422);
xnor U6164 (N_6164,N_59,N_423);
nand U6165 (N_6165,N_4187,N_3933);
nor U6166 (N_6166,N_3555,N_1983);
and U6167 (N_6167,N_4107,N_4359);
and U6168 (N_6168,N_4177,N_1348);
and U6169 (N_6169,N_1627,N_816);
and U6170 (N_6170,N_4910,N_3243);
and U6171 (N_6171,N_595,N_1390);
or U6172 (N_6172,N_2833,N_4741);
xor U6173 (N_6173,N_2663,N_768);
nand U6174 (N_6174,N_859,N_3033);
nand U6175 (N_6175,N_4222,N_575);
nor U6176 (N_6176,N_12,N_2145);
and U6177 (N_6177,N_1094,N_1521);
nor U6178 (N_6178,N_1976,N_2551);
nand U6179 (N_6179,N_663,N_404);
or U6180 (N_6180,N_1168,N_1676);
or U6181 (N_6181,N_867,N_3155);
nor U6182 (N_6182,N_579,N_4284);
nand U6183 (N_6183,N_1563,N_765);
nand U6184 (N_6184,N_944,N_656);
or U6185 (N_6185,N_771,N_2125);
or U6186 (N_6186,N_4834,N_2740);
and U6187 (N_6187,N_1681,N_4513);
nand U6188 (N_6188,N_3502,N_511);
and U6189 (N_6189,N_2386,N_2543);
xor U6190 (N_6190,N_114,N_314);
nand U6191 (N_6191,N_740,N_4520);
and U6192 (N_6192,N_623,N_2607);
or U6193 (N_6193,N_3616,N_3544);
or U6194 (N_6194,N_4558,N_3113);
nand U6195 (N_6195,N_469,N_825);
nand U6196 (N_6196,N_3866,N_9);
and U6197 (N_6197,N_2365,N_1449);
nand U6198 (N_6198,N_3892,N_2757);
or U6199 (N_6199,N_2292,N_2781);
nand U6200 (N_6200,N_2865,N_802);
or U6201 (N_6201,N_3479,N_220);
and U6202 (N_6202,N_1224,N_949);
and U6203 (N_6203,N_102,N_732);
or U6204 (N_6204,N_2676,N_1314);
nand U6205 (N_6205,N_976,N_1990);
or U6206 (N_6206,N_402,N_1546);
and U6207 (N_6207,N_3004,N_4650);
or U6208 (N_6208,N_4707,N_321);
and U6209 (N_6209,N_2440,N_3381);
nor U6210 (N_6210,N_4604,N_1543);
or U6211 (N_6211,N_3280,N_1329);
or U6212 (N_6212,N_2382,N_2579);
or U6213 (N_6213,N_4014,N_2245);
and U6214 (N_6214,N_924,N_3773);
and U6215 (N_6215,N_3912,N_1157);
nor U6216 (N_6216,N_3527,N_2106);
or U6217 (N_6217,N_513,N_3666);
nor U6218 (N_6218,N_132,N_1347);
nor U6219 (N_6219,N_2185,N_4029);
and U6220 (N_6220,N_2764,N_4852);
nand U6221 (N_6221,N_4713,N_3771);
and U6222 (N_6222,N_4085,N_2186);
or U6223 (N_6223,N_712,N_2816);
nor U6224 (N_6224,N_3831,N_4902);
and U6225 (N_6225,N_3168,N_2538);
or U6226 (N_6226,N_1661,N_2446);
or U6227 (N_6227,N_2469,N_2524);
nor U6228 (N_6228,N_4242,N_3095);
nand U6229 (N_6229,N_2152,N_69);
or U6230 (N_6230,N_2908,N_4996);
or U6231 (N_6231,N_945,N_1829);
nand U6232 (N_6232,N_358,N_4823);
nand U6233 (N_6233,N_1779,N_4433);
nor U6234 (N_6234,N_3828,N_479);
or U6235 (N_6235,N_3742,N_1439);
and U6236 (N_6236,N_4865,N_347);
and U6237 (N_6237,N_1386,N_2128);
nor U6238 (N_6238,N_3322,N_4303);
xor U6239 (N_6239,N_3018,N_3629);
and U6240 (N_6240,N_454,N_3931);
or U6241 (N_6241,N_2661,N_1100);
nor U6242 (N_6242,N_3264,N_4504);
xor U6243 (N_6243,N_2794,N_4928);
and U6244 (N_6244,N_4408,N_3581);
and U6245 (N_6245,N_611,N_1258);
and U6246 (N_6246,N_3458,N_330);
nand U6247 (N_6247,N_2880,N_3331);
nand U6248 (N_6248,N_283,N_598);
and U6249 (N_6249,N_3080,N_4166);
or U6250 (N_6250,N_3592,N_689);
nor U6251 (N_6251,N_2589,N_1079);
or U6252 (N_6252,N_1073,N_457);
nor U6253 (N_6253,N_1319,N_2547);
and U6254 (N_6254,N_3855,N_172);
or U6255 (N_6255,N_755,N_2482);
or U6256 (N_6256,N_3365,N_4255);
nor U6257 (N_6257,N_1231,N_4561);
nand U6258 (N_6258,N_3470,N_2091);
and U6259 (N_6259,N_2139,N_1009);
and U6260 (N_6260,N_1432,N_4992);
nor U6261 (N_6261,N_3231,N_4762);
nand U6262 (N_6262,N_1139,N_2310);
or U6263 (N_6263,N_4894,N_4519);
or U6264 (N_6264,N_2353,N_471);
nand U6265 (N_6265,N_3449,N_4572);
nor U6266 (N_6266,N_761,N_4048);
nand U6267 (N_6267,N_2733,N_4335);
nor U6268 (N_6268,N_4726,N_726);
nor U6269 (N_6269,N_3641,N_3683);
or U6270 (N_6270,N_4580,N_499);
and U6271 (N_6271,N_4252,N_4015);
nand U6272 (N_6272,N_178,N_2466);
or U6273 (N_6273,N_2313,N_4058);
and U6274 (N_6274,N_1060,N_2510);
nand U6275 (N_6275,N_3626,N_480);
or U6276 (N_6276,N_1260,N_2830);
or U6277 (N_6277,N_1709,N_1102);
nand U6278 (N_6278,N_3938,N_254);
and U6279 (N_6279,N_1815,N_3915);
or U6280 (N_6280,N_4370,N_3297);
nor U6281 (N_6281,N_3125,N_618);
nor U6282 (N_6282,N_2698,N_2347);
nor U6283 (N_6283,N_3898,N_2272);
nor U6284 (N_6284,N_4683,N_284);
and U6285 (N_6285,N_3309,N_3684);
nor U6286 (N_6286,N_1921,N_946);
and U6287 (N_6287,N_421,N_1796);
and U6288 (N_6288,N_2693,N_2613);
nand U6289 (N_6289,N_3846,N_2045);
nand U6290 (N_6290,N_2101,N_2203);
nor U6291 (N_6291,N_4411,N_198);
nand U6292 (N_6292,N_1514,N_2318);
and U6293 (N_6293,N_1134,N_3523);
or U6294 (N_6294,N_3115,N_3920);
and U6295 (N_6295,N_2450,N_850);
and U6296 (N_6296,N_1201,N_3428);
nand U6297 (N_6297,N_4290,N_3123);
and U6298 (N_6298,N_3354,N_4043);
nand U6299 (N_6299,N_3901,N_4595);
nor U6300 (N_6300,N_4653,N_1207);
or U6301 (N_6301,N_1433,N_3216);
xor U6302 (N_6302,N_3685,N_795);
and U6303 (N_6303,N_2863,N_4203);
and U6304 (N_6304,N_551,N_3053);
and U6305 (N_6305,N_1585,N_2742);
nand U6306 (N_6306,N_3756,N_4494);
nor U6307 (N_6307,N_4424,N_2990);
and U6308 (N_6308,N_4473,N_85);
nand U6309 (N_6309,N_4182,N_3475);
xnor U6310 (N_6310,N_2479,N_4579);
nand U6311 (N_6311,N_261,N_466);
or U6312 (N_6312,N_352,N_3865);
or U6313 (N_6313,N_580,N_562);
or U6314 (N_6314,N_130,N_2840);
or U6315 (N_6315,N_2533,N_3535);
or U6316 (N_6316,N_3576,N_2188);
or U6317 (N_6317,N_4630,N_613);
nand U6318 (N_6318,N_4948,N_3612);
and U6319 (N_6319,N_563,N_680);
nand U6320 (N_6320,N_300,N_1087);
nand U6321 (N_6321,N_312,N_1084);
or U6322 (N_6322,N_427,N_4837);
nand U6323 (N_6323,N_1903,N_1940);
nand U6324 (N_6324,N_4137,N_3305);
nand U6325 (N_6325,N_2741,N_1693);
nand U6326 (N_6326,N_2291,N_2537);
nor U6327 (N_6327,N_2022,N_4476);
nand U6328 (N_6328,N_3501,N_4291);
or U6329 (N_6329,N_3191,N_2239);
nor U6330 (N_6330,N_866,N_2144);
and U6331 (N_6331,N_4016,N_182);
nor U6332 (N_6332,N_1206,N_3210);
nor U6333 (N_6333,N_4174,N_702);
or U6334 (N_6334,N_3184,N_4204);
nor U6335 (N_6335,N_3077,N_4944);
xor U6336 (N_6336,N_1315,N_285);
or U6337 (N_6337,N_2724,N_2421);
or U6338 (N_6338,N_1859,N_1624);
and U6339 (N_6339,N_2345,N_459);
and U6340 (N_6340,N_777,N_4055);
and U6341 (N_6341,N_4138,N_2884);
nand U6342 (N_6342,N_3747,N_1517);
nand U6343 (N_6343,N_3512,N_2012);
nor U6344 (N_6344,N_1785,N_3016);
or U6345 (N_6345,N_645,N_4217);
and U6346 (N_6346,N_1925,N_3702);
or U6347 (N_6347,N_570,N_1214);
and U6348 (N_6348,N_2396,N_597);
and U6349 (N_6349,N_2021,N_3493);
nor U6350 (N_6350,N_2806,N_2749);
nor U6351 (N_6351,N_126,N_3658);
xor U6352 (N_6352,N_865,N_2338);
or U6353 (N_6353,N_4718,N_2374);
nand U6354 (N_6354,N_4500,N_1986);
and U6355 (N_6355,N_99,N_3136);
and U6356 (N_6356,N_2775,N_3287);
or U6357 (N_6357,N_3767,N_3651);
or U6358 (N_6358,N_4589,N_2159);
or U6359 (N_6359,N_4637,N_4927);
nand U6360 (N_6360,N_3825,N_811);
nand U6361 (N_6361,N_1178,N_2555);
or U6362 (N_6362,N_1277,N_1477);
or U6363 (N_6363,N_3081,N_1090);
nand U6364 (N_6364,N_3844,N_2703);
and U6365 (N_6365,N_1366,N_121);
and U6366 (N_6366,N_854,N_199);
nand U6367 (N_6367,N_627,N_1902);
nand U6368 (N_6368,N_4958,N_2525);
nand U6369 (N_6369,N_4200,N_194);
nor U6370 (N_6370,N_4881,N_3607);
nand U6371 (N_6371,N_3380,N_3389);
nand U6372 (N_6372,N_4434,N_4886);
and U6373 (N_6373,N_4990,N_1648);
and U6374 (N_6374,N_3026,N_2171);
or U6375 (N_6375,N_1568,N_2059);
nor U6376 (N_6376,N_863,N_2804);
xor U6377 (N_6377,N_2856,N_3940);
nor U6378 (N_6378,N_2302,N_4235);
nand U6379 (N_6379,N_186,N_2692);
nor U6380 (N_6380,N_4280,N_2398);
and U6381 (N_6381,N_1882,N_4545);
nand U6382 (N_6382,N_4455,N_1116);
and U6383 (N_6383,N_2013,N_4337);
nand U6384 (N_6384,N_4608,N_2841);
xor U6385 (N_6385,N_4028,N_3291);
and U6386 (N_6386,N_3710,N_2695);
and U6387 (N_6387,N_1077,N_2074);
nor U6388 (N_6388,N_1712,N_1872);
nor U6389 (N_6389,N_305,N_2331);
nand U6390 (N_6390,N_2678,N_4432);
nand U6391 (N_6391,N_3649,N_2351);
nor U6392 (N_6392,N_1194,N_153);
and U6393 (N_6393,N_1110,N_4908);
or U6394 (N_6394,N_892,N_4247);
or U6395 (N_6395,N_3433,N_3966);
and U6396 (N_6396,N_1189,N_3823);
and U6397 (N_6397,N_2963,N_2395);
nor U6398 (N_6398,N_4754,N_1532);
nand U6399 (N_6399,N_2494,N_2909);
and U6400 (N_6400,N_3395,N_1045);
nand U6401 (N_6401,N_1219,N_3599);
or U6402 (N_6402,N_1772,N_405);
nand U6403 (N_6403,N_779,N_3745);
and U6404 (N_6404,N_908,N_4742);
and U6405 (N_6405,N_1181,N_1450);
or U6406 (N_6406,N_4706,N_1429);
nor U6407 (N_6407,N_1606,N_1631);
nand U6408 (N_6408,N_4179,N_1926);
or U6409 (N_6409,N_497,N_1321);
or U6410 (N_6410,N_2483,N_1891);
nor U6411 (N_6411,N_3595,N_646);
nor U6412 (N_6412,N_1154,N_1642);
or U6413 (N_6413,N_665,N_4296);
nor U6414 (N_6414,N_1236,N_1914);
and U6415 (N_6415,N_3963,N_1443);
nor U6416 (N_6416,N_1570,N_1173);
nand U6417 (N_6417,N_3676,N_10);
nand U6418 (N_6418,N_2357,N_366);
and U6419 (N_6419,N_1184,N_2985);
nand U6420 (N_6420,N_4010,N_2864);
nand U6421 (N_6421,N_3698,N_2793);
or U6422 (N_6422,N_3012,N_257);
or U6423 (N_6423,N_1144,N_4857);
nand U6424 (N_6424,N_3195,N_673);
nand U6425 (N_6425,N_3762,N_4209);
and U6426 (N_6426,N_2773,N_293);
nand U6427 (N_6427,N_3358,N_4036);
or U6428 (N_6428,N_4025,N_3913);
nor U6429 (N_6429,N_2262,N_2759);
nor U6430 (N_6430,N_4350,N_556);
or U6431 (N_6431,N_2024,N_3362);
nand U6432 (N_6432,N_4125,N_3826);
nor U6433 (N_6433,N_4399,N_2855);
and U6434 (N_6434,N_662,N_1708);
nor U6435 (N_6435,N_157,N_1446);
nand U6436 (N_6436,N_2086,N_1682);
nor U6437 (N_6437,N_4757,N_518);
nand U6438 (N_6438,N_3824,N_2034);
nor U6439 (N_6439,N_264,N_3848);
nor U6440 (N_6440,N_3816,N_1897);
nor U6441 (N_6441,N_110,N_2528);
nand U6442 (N_6442,N_596,N_2055);
or U6443 (N_6443,N_1578,N_2108);
or U6444 (N_6444,N_1208,N_4417);
nand U6445 (N_6445,N_426,N_1131);
or U6446 (N_6446,N_125,N_2391);
and U6447 (N_6447,N_2688,N_1334);
nand U6448 (N_6448,N_3796,N_2958);
nand U6449 (N_6449,N_2572,N_928);
and U6450 (N_6450,N_636,N_3967);
or U6451 (N_6451,N_594,N_3145);
nand U6452 (N_6452,N_1929,N_564);
nand U6453 (N_6453,N_4939,N_4836);
and U6454 (N_6454,N_4218,N_1743);
nand U6455 (N_6455,N_1560,N_3010);
nand U6456 (N_6456,N_1973,N_3434);
and U6457 (N_6457,N_2873,N_1030);
or U6458 (N_6458,N_15,N_4634);
nand U6459 (N_6459,N_4975,N_3634);
and U6460 (N_6460,N_4674,N_2745);
xor U6461 (N_6461,N_1922,N_951);
nor U6462 (N_6462,N_2279,N_2424);
and U6463 (N_6463,N_2636,N_2658);
or U6464 (N_6464,N_1436,N_3765);
nor U6465 (N_6465,N_911,N_1442);
nor U6466 (N_6466,N_621,N_1810);
nand U6467 (N_6467,N_1239,N_1211);
or U6468 (N_6468,N_2040,N_64);
nand U6469 (N_6469,N_3097,N_94);
nor U6470 (N_6470,N_1816,N_296);
or U6471 (N_6471,N_177,N_4153);
or U6472 (N_6472,N_4272,N_346);
and U6473 (N_6473,N_2418,N_1620);
nand U6474 (N_6474,N_1629,N_6);
or U6475 (N_6475,N_678,N_3718);
and U6476 (N_6476,N_467,N_4190);
nand U6477 (N_6477,N_3832,N_1343);
nand U6478 (N_6478,N_1004,N_53);
nand U6479 (N_6479,N_248,N_4678);
or U6480 (N_6480,N_1758,N_1559);
nor U6481 (N_6481,N_3245,N_3519);
nor U6482 (N_6482,N_1640,N_3965);
nand U6483 (N_6483,N_3923,N_4461);
and U6484 (N_6484,N_2412,N_757);
nand U6485 (N_6485,N_2767,N_145);
or U6486 (N_6486,N_1330,N_2459);
or U6487 (N_6487,N_2076,N_1044);
and U6488 (N_6488,N_1271,N_1830);
nor U6489 (N_6489,N_311,N_2109);
nand U6490 (N_6490,N_1423,N_4497);
nand U6491 (N_6491,N_4223,N_4521);
nand U6492 (N_6492,N_3695,N_999);
xnor U6493 (N_6493,N_789,N_3810);
nand U6494 (N_6494,N_1639,N_3784);
and U6495 (N_6495,N_1995,N_4954);
and U6496 (N_6496,N_4501,N_4766);
xnor U6497 (N_6497,N_3559,N_4273);
or U6498 (N_6498,N_4110,N_2439);
nor U6499 (N_6499,N_796,N_2457);
and U6500 (N_6500,N_1608,N_2614);
and U6501 (N_6501,N_558,N_484);
nand U6502 (N_6502,N_2519,N_4553);
or U6503 (N_6503,N_4629,N_2054);
and U6504 (N_6504,N_2889,N_1402);
or U6505 (N_6505,N_1524,N_4472);
nand U6506 (N_6506,N_316,N_1999);
nor U6507 (N_6507,N_4414,N_1394);
and U6508 (N_6508,N_947,N_982);
or U6509 (N_6509,N_3273,N_2744);
and U6510 (N_6510,N_1406,N_2848);
nand U6511 (N_6511,N_657,N_92);
nand U6512 (N_6512,N_4163,N_4410);
nor U6513 (N_6513,N_2098,N_3439);
nand U6514 (N_6514,N_2652,N_4736);
and U6515 (N_6515,N_3704,N_3022);
nand U6516 (N_6516,N_1287,N_2138);
xnor U6517 (N_6517,N_3192,N_1774);
nand U6518 (N_6518,N_1014,N_3315);
and U6519 (N_6519,N_143,N_1274);
nor U6520 (N_6520,N_413,N_4566);
and U6521 (N_6521,N_542,N_167);
nor U6522 (N_6522,N_1054,N_4853);
nand U6523 (N_6523,N_4193,N_4279);
nor U6524 (N_6524,N_2696,N_2791);
nand U6525 (N_6525,N_4321,N_3000);
and U6526 (N_6526,N_1395,N_3342);
nand U6527 (N_6527,N_169,N_443);
or U6528 (N_6528,N_4067,N_4563);
and U6529 (N_6529,N_3717,N_4551);
nand U6530 (N_6530,N_385,N_2982);
nand U6531 (N_6531,N_1057,N_4981);
nor U6532 (N_6532,N_4863,N_3632);
nor U6533 (N_6533,N_1647,N_737);
or U6534 (N_6534,N_2242,N_4919);
or U6535 (N_6535,N_748,N_3378);
and U6536 (N_6536,N_1381,N_666);
and U6537 (N_6537,N_211,N_4226);
and U6538 (N_6538,N_919,N_1346);
and U6539 (N_6539,N_4449,N_1156);
and U6540 (N_6540,N_341,N_297);
or U6541 (N_6541,N_3146,N_4117);
nor U6542 (N_6542,N_1163,N_4299);
xnor U6543 (N_6543,N_403,N_1918);
nor U6544 (N_6544,N_207,N_1566);
nor U6545 (N_6545,N_2336,N_1052);
and U6546 (N_6546,N_388,N_2360);
or U6547 (N_6547,N_1204,N_506);
xor U6548 (N_6548,N_2116,N_3176);
nand U6549 (N_6549,N_1971,N_522);
nand U6550 (N_6550,N_994,N_2651);
or U6551 (N_6551,N_3768,N_2445);
and U6552 (N_6552,N_1839,N_1461);
or U6553 (N_6553,N_1576,N_4463);
and U6554 (N_6554,N_229,N_4788);
nand U6555 (N_6555,N_1934,N_3995);
nor U6556 (N_6556,N_4100,N_2706);
or U6557 (N_6557,N_1685,N_3170);
nor U6558 (N_6558,N_2701,N_4677);
nor U6559 (N_6559,N_4506,N_2668);
nor U6560 (N_6560,N_2650,N_232);
and U6561 (N_6561,N_2950,N_4940);
nand U6562 (N_6562,N_3128,N_2677);
or U6563 (N_6563,N_791,N_2991);
and U6564 (N_6564,N_185,N_2886);
nor U6565 (N_6565,N_3671,N_4916);
and U6566 (N_6566,N_345,N_439);
nand U6567 (N_6567,N_4376,N_1038);
and U6568 (N_6568,N_4708,N_1656);
nor U6569 (N_6569,N_2624,N_2039);
and U6570 (N_6570,N_1683,N_139);
nand U6571 (N_6571,N_543,N_1018);
or U6572 (N_6572,N_3495,N_81);
and U6573 (N_6573,N_1762,N_1721);
nor U6574 (N_6574,N_4385,N_4447);
or U6575 (N_6575,N_3633,N_2862);
nor U6576 (N_6576,N_2986,N_1545);
nand U6577 (N_6577,N_1377,N_4322);
nand U6578 (N_6578,N_4492,N_1965);
nand U6579 (N_6579,N_2926,N_3377);
nand U6580 (N_6580,N_3139,N_3838);
nand U6581 (N_6581,N_3861,N_1210);
nand U6582 (N_6582,N_2888,N_4006);
nand U6583 (N_6583,N_3653,N_4920);
and U6584 (N_6584,N_2025,N_3311);
and U6585 (N_6585,N_773,N_4971);
and U6586 (N_6586,N_4243,N_1962);
and U6587 (N_6587,N_1780,N_4825);
or U6588 (N_6588,N_170,N_1020);
nor U6589 (N_6589,N_624,N_3100);
and U6590 (N_6590,N_1295,N_4267);
and U6591 (N_6591,N_4229,N_632);
and U6592 (N_6592,N_4546,N_820);
or U6593 (N_6593,N_2243,N_3905);
and U6594 (N_6594,N_2595,N_3975);
nand U6595 (N_6595,N_4964,N_2316);
or U6596 (N_6596,N_4409,N_1234);
and U6597 (N_6597,N_4670,N_605);
xnor U6598 (N_6598,N_4421,N_2404);
and U6599 (N_6599,N_2323,N_1883);
and U6600 (N_6600,N_3943,N_3758);
nor U6601 (N_6601,N_1117,N_237);
or U6602 (N_6602,N_448,N_4134);
or U6603 (N_6603,N_2729,N_1726);
nand U6604 (N_6604,N_231,N_3884);
nand U6605 (N_6605,N_2419,N_1455);
and U6606 (N_6606,N_4739,N_4363);
and U6607 (N_6607,N_3985,N_1792);
nor U6608 (N_6608,N_840,N_2694);
or U6609 (N_6609,N_221,N_2325);
nor U6610 (N_6610,N_1801,N_4666);
nand U6611 (N_6611,N_398,N_3398);
nor U6612 (N_6612,N_4626,N_2513);
or U6613 (N_6613,N_2126,N_4035);
nor U6614 (N_6614,N_4116,N_1421);
nand U6615 (N_6615,N_2498,N_249);
nand U6616 (N_6616,N_3899,N_774);
nor U6617 (N_6617,N_119,N_722);
nand U6618 (N_6618,N_2305,N_2110);
and U6619 (N_6619,N_319,N_2227);
nand U6620 (N_6620,N_2921,N_3821);
nand U6621 (N_6621,N_3835,N_792);
xor U6622 (N_6622,N_1141,N_1471);
or U6623 (N_6623,N_3221,N_3840);
or U6624 (N_6624,N_3455,N_2394);
nor U6625 (N_6625,N_490,N_2202);
or U6626 (N_6626,N_549,N_3620);
nand U6627 (N_6627,N_1978,N_4734);
nor U6628 (N_6628,N_1773,N_395);
nor U6629 (N_6629,N_2774,N_369);
or U6630 (N_6630,N_37,N_1028);
nand U6631 (N_6631,N_4310,N_2962);
or U6632 (N_6632,N_3205,N_1690);
or U6633 (N_6633,N_3511,N_3924);
and U6634 (N_6634,N_4374,N_4091);
nand U6635 (N_6635,N_2111,N_4819);
or U6636 (N_6636,N_2358,N_747);
nor U6637 (N_6637,N_3605,N_4234);
or U6638 (N_6638,N_4849,N_4682);
nor U6639 (N_6639,N_1738,N_2490);
and U6640 (N_6640,N_967,N_4156);
or U6641 (N_6641,N_2797,N_3590);
or U6642 (N_6642,N_2983,N_2571);
or U6643 (N_6643,N_3002,N_4900);
and U6644 (N_6644,N_3952,N_4672);
nand U6645 (N_6645,N_3144,N_2974);
nand U6646 (N_6646,N_1158,N_3930);
nand U6647 (N_6647,N_1474,N_3889);
or U6648 (N_6648,N_1342,N_4875);
and U6649 (N_6649,N_3066,N_4639);
and U6650 (N_6650,N_2770,N_2925);
and U6651 (N_6651,N_1528,N_4127);
and U6652 (N_6652,N_1561,N_3248);
or U6653 (N_6653,N_4253,N_3177);
nor U6654 (N_6654,N_1412,N_3206);
and U6655 (N_6655,N_936,N_1652);
nand U6656 (N_6656,N_1689,N_1799);
or U6657 (N_6657,N_1111,N_1482);
nand U6658 (N_6658,N_340,N_1595);
and U6659 (N_6659,N_1361,N_4192);
or U6660 (N_6660,N_528,N_2837);
nor U6661 (N_6661,N_1485,N_3227);
or U6662 (N_6662,N_1088,N_4349);
xnor U6663 (N_6663,N_4092,N_3379);
nand U6664 (N_6664,N_4596,N_2315);
nor U6665 (N_6665,N_3849,N_4937);
nand U6666 (N_6666,N_187,N_4888);
or U6667 (N_6667,N_1418,N_701);
nand U6668 (N_6668,N_4633,N_4949);
and U6669 (N_6669,N_4868,N_841);
nor U6670 (N_6670,N_4785,N_3037);
nor U6671 (N_6671,N_1655,N_1428);
and U6672 (N_6672,N_4260,N_1981);
nor U6673 (N_6673,N_4912,N_1798);
or U6674 (N_6674,N_2673,N_3468);
nor U6675 (N_6675,N_642,N_429);
and U6676 (N_6676,N_2361,N_1491);
or U6677 (N_6677,N_4870,N_2252);
nor U6678 (N_6678,N_4820,N_2751);
and U6679 (N_6679,N_3087,N_1895);
or U6680 (N_6680,N_2124,N_456);
and U6681 (N_6681,N_2967,N_3375);
or U6682 (N_6682,N_381,N_3334);
or U6683 (N_6683,N_2359,N_589);
or U6684 (N_6684,N_793,N_4904);
or U6685 (N_6685,N_817,N_18);
nand U6686 (N_6686,N_1199,N_3229);
and U6687 (N_6687,N_527,N_2505);
nor U6688 (N_6688,N_4352,N_4452);
or U6689 (N_6689,N_3266,N_2080);
nor U6690 (N_6690,N_4076,N_419);
and U6691 (N_6691,N_2824,N_1901);
nand U6692 (N_6692,N_4724,N_3490);
nand U6693 (N_6693,N_217,N_1096);
nor U6694 (N_6694,N_1667,N_308);
nor U6695 (N_6695,N_3271,N_4471);
nand U6696 (N_6696,N_2578,N_2465);
nand U6697 (N_6697,N_4004,N_2071);
or U6698 (N_6698,N_3712,N_2838);
and U6699 (N_6699,N_993,N_4135);
or U6700 (N_6700,N_728,N_2608);
and U6701 (N_6701,N_1011,N_637);
nor U6702 (N_6702,N_4845,N_2890);
and U6703 (N_6703,N_2166,N_2068);
or U6704 (N_6704,N_1122,N_2330);
nor U6705 (N_6705,N_2588,N_2817);
nor U6706 (N_6706,N_4555,N_4415);
nor U6707 (N_6707,N_2511,N_1195);
or U6708 (N_6708,N_2931,N_2831);
or U6709 (N_6709,N_252,N_2058);
or U6710 (N_6710,N_1770,N_4211);
or U6711 (N_6711,N_3162,N_1140);
and U6712 (N_6712,N_4329,N_3876);
nand U6713 (N_6713,N_4403,N_3124);
nand U6714 (N_6714,N_2117,N_4609);
nand U6715 (N_6715,N_4756,N_1750);
or U6716 (N_6716,N_2481,N_2390);
nor U6717 (N_6717,N_1273,N_3024);
nand U6718 (N_6718,N_1306,N_4401);
or U6719 (N_6719,N_271,N_4542);
and U6720 (N_6720,N_4648,N_3450);
and U6721 (N_6721,N_4809,N_4763);
nand U6722 (N_6722,N_4733,N_2451);
nand U6723 (N_6723,N_4429,N_2935);
or U6724 (N_6724,N_2949,N_3520);
nand U6725 (N_6725,N_1776,N_4997);
and U6726 (N_6726,N_4020,N_3267);
nor U6727 (N_6727,N_3708,N_4966);
and U6728 (N_6728,N_2619,N_1177);
and U6729 (N_6729,N_2704,N_2378);
xnor U6730 (N_6730,N_2179,N_1939);
nand U6731 (N_6731,N_2536,N_1881);
and U6732 (N_6732,N_4144,N_1626);
nor U6733 (N_6733,N_2699,N_2119);
or U6734 (N_6734,N_3577,N_2014);
and U6735 (N_6735,N_4486,N_868);
and U6736 (N_6736,N_1769,N_862);
nor U6737 (N_6737,N_536,N_4224);
and U6738 (N_6738,N_148,N_2922);
nand U6739 (N_6739,N_2346,N_4917);
or U6740 (N_6740,N_2971,N_4528);
nand U6741 (N_6741,N_2965,N_1923);
nor U6742 (N_6742,N_1911,N_1930);
nor U6743 (N_6743,N_4487,N_4911);
and U6744 (N_6744,N_3361,N_4821);
nor U6745 (N_6745,N_3119,N_3602);
nand U6746 (N_6746,N_2521,N_2308);
nor U6747 (N_6747,N_3732,N_1370);
or U6748 (N_6748,N_3754,N_3235);
and U6749 (N_6749,N_1840,N_2803);
nor U6750 (N_6750,N_3713,N_1416);
nor U6751 (N_6751,N_763,N_3822);
nand U6752 (N_6752,N_1463,N_653);
or U6753 (N_6753,N_984,N_2226);
nand U6754 (N_6754,N_438,N_4309);
nand U6755 (N_6755,N_3421,N_3677);
and U6756 (N_6756,N_4258,N_4530);
nand U6757 (N_6757,N_1917,N_1489);
nor U6758 (N_6758,N_3149,N_3172);
nand U6759 (N_6759,N_3057,N_937);
and U6760 (N_6760,N_4281,N_3804);
nor U6761 (N_6761,N_3373,N_2344);
or U6762 (N_6762,N_3585,N_3542);
xor U6763 (N_6763,N_2942,N_4705);
and U6764 (N_6764,N_318,N_313);
xnor U6765 (N_6765,N_1950,N_3457);
nand U6766 (N_6766,N_4588,N_2805);
nand U6767 (N_6767,N_2155,N_4184);
or U6768 (N_6768,N_2410,N_2434);
nor U6769 (N_6769,N_2157,N_842);
or U6770 (N_6770,N_2307,N_4621);
nor U6771 (N_6771,N_112,N_353);
and U6772 (N_6772,N_696,N_3673);
nor U6773 (N_6773,N_1717,N_1786);
and U6774 (N_6774,N_275,N_1616);
and U6775 (N_6775,N_807,N_2023);
nand U6776 (N_6776,N_243,N_70);
and U6777 (N_6777,N_4428,N_1663);
nor U6778 (N_6778,N_1327,N_4786);
nand U6779 (N_6779,N_979,N_1064);
or U6780 (N_6780,N_446,N_4459);
or U6781 (N_6781,N_495,N_362);
nand U6782 (N_6782,N_1147,N_510);
nor U6783 (N_6783,N_38,N_2956);
and U6784 (N_6784,N_827,N_3313);
nand U6785 (N_6785,N_2150,N_3159);
nor U6786 (N_6786,N_1747,N_884);
or U6787 (N_6787,N_2170,N_2570);
nand U6788 (N_6788,N_1397,N_1069);
or U6789 (N_6789,N_2453,N_1410);
nand U6790 (N_6790,N_3129,N_3300);
or U6791 (N_6791,N_4878,N_3152);
nor U6792 (N_6792,N_162,N_1739);
or U6793 (N_6793,N_3561,N_1600);
xnor U6794 (N_6794,N_4068,N_1376);
nor U6795 (N_6795,N_1614,N_3006);
and U6796 (N_6796,N_1824,N_4663);
nand U6797 (N_6797,N_887,N_1622);
or U6798 (N_6798,N_386,N_1056);
and U6799 (N_6799,N_2795,N_2044);
nor U6800 (N_6800,N_995,N_1959);
nand U6801 (N_6801,N_3883,N_4186);
or U6802 (N_6802,N_2,N_1662);
or U6803 (N_6803,N_2648,N_4404);
or U6804 (N_6804,N_60,N_2164);
or U6805 (N_6805,N_4393,N_806);
nand U6806 (N_6806,N_1658,N_3200);
nand U6807 (N_6807,N_3185,N_2609);
or U6808 (N_6808,N_4953,N_242);
nor U6809 (N_6809,N_4947,N_4656);
xor U6810 (N_6810,N_532,N_3656);
or U6811 (N_6811,N_3394,N_1378);
or U6812 (N_6812,N_2072,N_3540);
nand U6813 (N_6813,N_1024,N_2114);
or U6814 (N_6814,N_2894,N_4907);
nand U6815 (N_6815,N_794,N_103);
or U6816 (N_6816,N_770,N_4457);
nor U6817 (N_6817,N_2782,N_4041);
nand U6818 (N_6818,N_3856,N_1420);
or U6819 (N_6819,N_2017,N_1162);
nand U6820 (N_6820,N_4278,N_3881);
and U6821 (N_6821,N_2075,N_1548);
nor U6822 (N_6822,N_4308,N_872);
nand U6823 (N_6823,N_3895,N_4897);
nor U6824 (N_6824,N_4093,N_3250);
and U6825 (N_6825,N_188,N_4772);
nor U6826 (N_6826,N_1396,N_3473);
and U6827 (N_6827,N_1935,N_4614);
nor U6828 (N_6828,N_4044,N_4314);
nor U6829 (N_6829,N_431,N_2674);
or U6830 (N_6830,N_1042,N_1031);
and U6831 (N_6831,N_1791,N_4307);
and U6832 (N_6832,N_3463,N_1797);
or U6833 (N_6833,N_3174,N_4439);
nor U6834 (N_6834,N_2383,N_2643);
or U6835 (N_6835,N_3142,N_3854);
nand U6836 (N_6836,N_3131,N_1298);
or U6837 (N_6837,N_87,N_4691);
nand U6838 (N_6838,N_33,N_3436);
or U6839 (N_6839,N_4065,N_4073);
nand U6840 (N_6840,N_2534,N_735);
and U6841 (N_6841,N_2820,N_1782);
nor U6842 (N_6842,N_4517,N_3008);
nand U6843 (N_6843,N_3788,N_603);
and U6844 (N_6844,N_3871,N_502);
nor U6845 (N_6845,N_918,N_4660);
nor U6846 (N_6846,N_4394,N_35);
and U6847 (N_6847,N_1692,N_1080);
nand U6848 (N_6848,N_4938,N_4090);
nand U6849 (N_6849,N_658,N_4250);
or U6850 (N_6850,N_1250,N_3664);
nor U6851 (N_6851,N_2293,N_801);
nand U6852 (N_6852,N_3588,N_3007);
nand U6853 (N_6853,N_4985,N_4245);
nor U6854 (N_6854,N_1249,N_649);
nand U6855 (N_6855,N_569,N_444);
nor U6856 (N_6856,N_1259,N_525);
and U6857 (N_6857,N_3618,N_129);
nor U6858 (N_6858,N_1464,N_4554);
and U6859 (N_6859,N_1851,N_4658);
nor U6860 (N_6860,N_2606,N_2846);
nand U6861 (N_6861,N_432,N_878);
or U6862 (N_6862,N_1526,N_2376);
and U6863 (N_6863,N_4509,N_1864);
nor U6864 (N_6864,N_1613,N_1628);
or U6865 (N_6865,N_717,N_3105);
or U6866 (N_6866,N_1290,N_2659);
nand U6867 (N_6867,N_2755,N_2209);
and U6868 (N_6868,N_2867,N_2070);
nor U6869 (N_6869,N_2881,N_3958);
nor U6870 (N_6870,N_2271,N_3945);
nor U6871 (N_6871,N_3032,N_389);
and U6872 (N_6872,N_4257,N_3993);
nor U6873 (N_6873,N_4444,N_1230);
and U6874 (N_6874,N_2435,N_2254);
or U6875 (N_6875,N_2031,N_2260);
nand U6876 (N_6876,N_4231,N_4263);
and U6877 (N_6877,N_2961,N_3163);
or U6878 (N_6878,N_2041,N_3372);
nor U6879 (N_6879,N_3445,N_1174);
nor U6880 (N_6880,N_541,N_3617);
nor U6881 (N_6881,N_2289,N_769);
and U6882 (N_6882,N_4729,N_2768);
nor U6883 (N_6883,N_4577,N_711);
nor U6884 (N_6884,N_686,N_4162);
or U6885 (N_6885,N_3014,N_3469);
and U6886 (N_6886,N_847,N_4094);
nor U6887 (N_6887,N_3268,N_306);
nand U6888 (N_6888,N_328,N_1788);
or U6889 (N_6889,N_65,N_1364);
nor U6890 (N_6890,N_4460,N_2928);
nor U6891 (N_6891,N_3735,N_1964);
nor U6892 (N_6892,N_2364,N_734);
nand U6893 (N_6893,N_2241,N_3918);
or U6894 (N_6894,N_3247,N_4221);
nand U6895 (N_6895,N_721,N_2369);
and U6896 (N_6896,N_2517,N_2143);
nand U6897 (N_6897,N_342,N_3686);
and U6898 (N_6898,N_4418,N_86);
or U6899 (N_6899,N_4343,N_529);
nand U6900 (N_6900,N_2638,N_2105);
and U6901 (N_6901,N_3997,N_2637);
nor U6902 (N_6902,N_3589,N_4477);
nor U6903 (N_6903,N_1846,N_179);
or U6904 (N_6904,N_3516,N_4095);
nor U6905 (N_6905,N_1598,N_2936);
nor U6906 (N_6906,N_2332,N_4576);
nand U6907 (N_6907,N_1757,N_1385);
nor U6908 (N_6908,N_156,N_1403);
and U6909 (N_6909,N_1937,N_3670);
nand U6910 (N_6910,N_3476,N_3580);
and U6911 (N_6911,N_4828,N_674);
and U6912 (N_6912,N_1289,N_1938);
and U6913 (N_6913,N_2851,N_1763);
nand U6914 (N_6914,N_274,N_1212);
and U6915 (N_6915,N_731,N_533);
nor U6916 (N_6916,N_3987,N_3663);
nand U6917 (N_6917,N_3293,N_1357);
and U6918 (N_6918,N_374,N_2244);
nor U6919 (N_6919,N_3055,N_4406);
nor U6920 (N_6920,N_212,N_1804);
or U6921 (N_6921,N_3011,N_367);
and U6922 (N_6922,N_281,N_4792);
nand U6923 (N_6923,N_2268,N_47);
or U6924 (N_6924,N_190,N_90);
and U6925 (N_6925,N_55,N_682);
and U6926 (N_6926,N_460,N_1015);
nor U6927 (N_6927,N_3110,N_2664);
and U6928 (N_6928,N_630,N_671);
and U6929 (N_6929,N_3730,N_3099);
or U6930 (N_6930,N_1253,N_725);
nor U6931 (N_6931,N_2355,N_856);
nor U6932 (N_6932,N_4727,N_4557);
nor U6933 (N_6933,N_4874,N_3749);
or U6934 (N_6934,N_1591,N_371);
and U6935 (N_6935,N_934,N_3051);
and U6936 (N_6936,N_1745,N_4807);
or U6937 (N_6937,N_2580,N_4081);
nor U6938 (N_6938,N_4562,N_2035);
and U6939 (N_6939,N_4723,N_3809);
or U6940 (N_6940,N_4146,N_4699);
nand U6941 (N_6941,N_3118,N_1282);
and U6942 (N_6942,N_4454,N_2384);
and U6943 (N_6943,N_684,N_4764);
and U6944 (N_6944,N_2062,N_1389);
xnor U6945 (N_6945,N_4295,N_677);
nor U6946 (N_6946,N_933,N_629);
or U6947 (N_6947,N_2141,N_4089);
nor U6948 (N_6948,N_1166,N_2861);
or U6949 (N_6949,N_972,N_1870);
or U6950 (N_6950,N_3288,N_1313);
nand U6951 (N_6951,N_4851,N_1958);
and U6952 (N_6952,N_2090,N_2814);
nor U6953 (N_6953,N_1233,N_310);
nor U6954 (N_6954,N_2043,N_4142);
and U6955 (N_6955,N_1592,N_82);
and U6956 (N_6956,N_2341,N_4254);
nand U6957 (N_6957,N_1993,N_1293);
nand U6958 (N_6958,N_253,N_4767);
and U6959 (N_6959,N_2065,N_3916);
xnor U6960 (N_6960,N_3043,N_1625);
nand U6961 (N_6961,N_1715,N_2016);
nor U6962 (N_6962,N_3787,N_874);
or U6963 (N_6963,N_41,N_1299);
nand U6964 (N_6964,N_997,N_1866);
and U6965 (N_6965,N_2415,N_1076);
and U6966 (N_6966,N_619,N_1098);
or U6967 (N_6967,N_1172,N_1050);
nand U6968 (N_6968,N_175,N_4719);
or U6969 (N_6969,N_3111,N_4168);
or U6970 (N_6970,N_1744,N_3980);
or U6971 (N_6971,N_336,N_2883);
and U6972 (N_6972,N_2866,N_392);
nor U6973 (N_6973,N_376,N_1440);
and U6974 (N_6974,N_2556,N_2154);
nor U6975 (N_6975,N_4164,N_4549);
and U6976 (N_6976,N_4152,N_4872);
nand U6977 (N_6977,N_4101,N_2422);
nand U6978 (N_6978,N_418,N_4550);
and U6979 (N_6979,N_973,N_799);
and U6980 (N_6980,N_4781,N_2902);
or U6981 (N_6981,N_3406,N_1399);
nor U6982 (N_6982,N_492,N_3324);
nand U6983 (N_6983,N_601,N_2187);
nor U6984 (N_6984,N_4777,N_486);
nand U6985 (N_6985,N_171,N_3786);
or U6986 (N_6986,N_581,N_3370);
or U6987 (N_6987,N_4864,N_2561);
or U6988 (N_6988,N_655,N_3345);
or U6989 (N_6989,N_3483,N_1209);
nor U6990 (N_6990,N_3374,N_1555);
nand U6991 (N_6991,N_670,N_2223);
nor U6992 (N_6992,N_1091,N_718);
xnor U6993 (N_6993,N_4525,N_3171);
nor U6994 (N_6994,N_1837,N_2666);
or U6995 (N_6995,N_2702,N_4324);
and U6996 (N_6996,N_2019,N_4419);
nand U6997 (N_6997,N_2998,N_3550);
nor U6998 (N_6998,N_2263,N_2576);
nor U6999 (N_6999,N_375,N_2622);
nand U7000 (N_7000,N_4924,N_839);
nor U7001 (N_7001,N_2097,N_3537);
nor U7002 (N_7002,N_3888,N_2371);
nand U7003 (N_7003,N_295,N_2297);
nor U7004 (N_7004,N_2789,N_309);
or U7005 (N_7005,N_4701,N_4647);
or U7006 (N_7006,N_1086,N_2032);
nand U7007 (N_7007,N_3213,N_1579);
and U7008 (N_7008,N_1969,N_2719);
nand U7009 (N_7009,N_942,N_2917);
nor U7010 (N_7010,N_545,N_1255);
nand U7011 (N_7011,N_3807,N_2876);
xnor U7012 (N_7012,N_743,N_1821);
or U7013 (N_7013,N_4183,N_1145);
nor U7014 (N_7014,N_3531,N_3430);
nand U7015 (N_7015,N_317,N_2946);
xor U7016 (N_7016,N_1326,N_1379);
xnor U7017 (N_7017,N_3228,N_1284);
nand U7018 (N_7018,N_4583,N_166);
or U7019 (N_7019,N_4704,N_2118);
xnor U7020 (N_7020,N_2212,N_4773);
nor U7021 (N_7021,N_2842,N_4498);
or U7022 (N_7022,N_3121,N_4662);
nor U7023 (N_7023,N_2335,N_4664);
nor U7024 (N_7024,N_1142,N_3934);
and U7025 (N_7025,N_409,N_3636);
nand U7026 (N_7026,N_2628,N_3872);
nor U7027 (N_7027,N_3038,N_4430);
and U7028 (N_7028,N_1768,N_2428);
xnor U7029 (N_7029,N_3829,N_1417);
or U7030 (N_7030,N_3638,N_683);
and U7031 (N_7031,N_4061,N_2918);
nand U7032 (N_7032,N_1612,N_2642);
and U7033 (N_7033,N_1659,N_2104);
nor U7034 (N_7034,N_2131,N_2458);
or U7035 (N_7035,N_4266,N_4412);
and U7036 (N_7036,N_4311,N_1755);
nand U7037 (N_7037,N_4367,N_2372);
and U7038 (N_7038,N_4669,N_3551);
nand U7039 (N_7039,N_2758,N_2586);
or U7040 (N_7040,N_927,N_3820);
and U7041 (N_7041,N_1539,N_256);
nand U7042 (N_7042,N_4213,N_798);
nand U7043 (N_7043,N_2993,N_1680);
nor U7044 (N_7044,N_174,N_4931);
and U7045 (N_7045,N_2328,N_3833);
nand U7046 (N_7046,N_205,N_1186);
xnor U7047 (N_7047,N_1447,N_3484);
nor U7048 (N_7048,N_1202,N_108);
or U7049 (N_7049,N_4538,N_2340);
nor U7050 (N_7050,N_2217,N_3341);
nand U7051 (N_7051,N_1016,N_1023);
or U7052 (N_7052,N_4933,N_4859);
or U7053 (N_7053,N_294,N_4731);
or U7054 (N_7054,N_3515,N_4659);
nor U7055 (N_7055,N_4483,N_4571);
nor U7056 (N_7056,N_1723,N_1254);
nor U7057 (N_7057,N_1237,N_2630);
nor U7058 (N_7058,N_4262,N_204);
or U7059 (N_7059,N_2654,N_4540);
nor U7060 (N_7060,N_73,N_3929);
or U7061 (N_7061,N_4833,N_1694);
or U7062 (N_7062,N_57,N_4080);
nor U7063 (N_7063,N_2281,N_524);
or U7064 (N_7064,N_3794,N_568);
nor U7065 (N_7065,N_2037,N_4216);
or U7066 (N_7066,N_4970,N_3401);
nand U7067 (N_7067,N_775,N_325);
or U7068 (N_7068,N_2919,N_3036);
or U7069 (N_7069,N_2826,N_3488);
and U7070 (N_7070,N_3133,N_2611);
nand U7071 (N_7071,N_3697,N_2177);
or U7072 (N_7072,N_4070,N_4320);
or U7073 (N_7073,N_4340,N_159);
or U7074 (N_7074,N_3,N_68);
nand U7075 (N_7075,N_3277,N_2822);
and U7076 (N_7076,N_2000,N_1888);
or U7077 (N_7077,N_3240,N_1850);
nand U7078 (N_7078,N_4841,N_2725);
and U7079 (N_7079,N_3894,N_4288);
nand U7080 (N_7080,N_4703,N_3847);
and U7081 (N_7081,N_4480,N_4228);
nand U7082 (N_7082,N_664,N_4839);
nand U7083 (N_7083,N_1510,N_3654);
nor U7084 (N_7084,N_3132,N_93);
and U7085 (N_7085,N_3582,N_4612);
nor U7086 (N_7086,N_1668,N_3165);
and U7087 (N_7087,N_2298,N_2763);
nor U7088 (N_7088,N_1128,N_1065);
and U7089 (N_7089,N_797,N_331);
and U7090 (N_7090,N_4986,N_978);
and U7091 (N_7091,N_2270,N_1257);
nor U7092 (N_7092,N_1948,N_2084);
nand U7093 (N_7093,N_4625,N_2665);
nor U7094 (N_7094,N_3480,N_74);
or U7095 (N_7095,N_1842,N_3063);
or U7096 (N_7096,N_4039,N_2689);
xnor U7097 (N_7097,N_2872,N_1716);
nor U7098 (N_7098,N_3234,N_370);
or U7099 (N_7099,N_3939,N_464);
and U7100 (N_7100,N_1749,N_4496);
nand U7101 (N_7101,N_681,N_2350);
or U7102 (N_7102,N_1650,N_4239);
nor U7103 (N_7103,N_2845,N_4568);
and U7104 (N_7104,N_784,N_3726);
and U7105 (N_7105,N_4037,N_222);
nor U7106 (N_7106,N_1737,N_2046);
and U7107 (N_7107,N_1075,N_3904);
and U7108 (N_7108,N_4108,N_1263);
nand U7109 (N_7109,N_3560,N_263);
xor U7110 (N_7110,N_2056,N_2999);
and U7111 (N_7111,N_955,N_1078);
and U7112 (N_7112,N_694,N_3397);
and U7113 (N_7113,N_1875,N_1244);
nor U7114 (N_7114,N_2566,N_4237);
nor U7115 (N_7115,N_1678,N_4934);
nor U7116 (N_7116,N_2426,N_4495);
and U7117 (N_7117,N_2585,N_4386);
nand U7118 (N_7118,N_2520,N_3850);
or U7119 (N_7119,N_3141,N_2329);
nor U7120 (N_7120,N_3137,N_1588);
nor U7121 (N_7121,N_1497,N_1793);
and U7122 (N_7122,N_1574,N_4882);
nand U7123 (N_7123,N_2251,N_3327);
and U7124 (N_7124,N_1919,N_2618);
or U7125 (N_7125,N_355,N_3700);
nand U7126 (N_7126,N_672,N_2147);
nand U7127 (N_7127,N_790,N_4681);
nand U7128 (N_7128,N_3387,N_2235);
nand U7129 (N_7129,N_1905,N_1242);
and U7130 (N_7130,N_2972,N_1535);
and U7131 (N_7131,N_4983,N_2192);
nor U7132 (N_7132,N_2199,N_4575);
nor U7133 (N_7133,N_638,N_100);
or U7134 (N_7134,N_2250,N_1276);
and U7135 (N_7135,N_1059,N_1074);
nor U7136 (N_7136,N_2299,N_3049);
nand U7137 (N_7137,N_1852,N_4462);
nand U7138 (N_7138,N_585,N_3521);
and U7139 (N_7139,N_501,N_4018);
or U7140 (N_7140,N_2777,N_848);
and U7141 (N_7141,N_1294,N_3497);
or U7142 (N_7142,N_2342,N_2640);
and U7143 (N_7143,N_566,N_964);
or U7144 (N_7144,N_1337,N_481);
nor U7145 (N_7145,N_2455,N_8);
nor U7146 (N_7146,N_4276,N_482);
nand U7147 (N_7147,N_2077,N_800);
nor U7148 (N_7148,N_622,N_61);
nand U7149 (N_7149,N_3800,N_1387);
nor U7150 (N_7150,N_4871,N_447);
nand U7151 (N_7151,N_2752,N_1582);
nand U7152 (N_7152,N_3508,N_2403);
or U7153 (N_7153,N_4261,N_4941);
nand U7154 (N_7154,N_3477,N_1828);
nor U7155 (N_7155,N_3613,N_1771);
nor U7156 (N_7156,N_1468,N_1508);
or U7157 (N_7157,N_1063,N_234);
or U7158 (N_7158,N_4605,N_1730);
or U7159 (N_7159,N_4787,N_3413);
nand U7160 (N_7160,N_1607,N_1005);
nand U7161 (N_7161,N_929,N_1454);
nor U7162 (N_7162,N_4725,N_101);
or U7163 (N_7163,N_4657,N_1278);
nor U7164 (N_7164,N_1256,N_36);
nor U7165 (N_7165,N_2326,N_3289);
nor U7166 (N_7166,N_3746,N_3596);
and U7167 (N_7167,N_4232,N_4122);
nand U7168 (N_7168,N_2194,N_2456);
and U7169 (N_7169,N_2679,N_2731);
nand U7170 (N_7170,N_2857,N_2649);
xnor U7171 (N_7171,N_334,N_52);
nand U7172 (N_7172,N_669,N_4358);
nor U7173 (N_7173,N_45,N_2009);
or U7174 (N_7174,N_2761,N_4695);
nor U7175 (N_7175,N_1356,N_4799);
nand U7176 (N_7176,N_1101,N_213);
nand U7177 (N_7177,N_230,N_3424);
nor U7178 (N_7178,N_2222,N_2953);
nor U7179 (N_7179,N_1994,N_2981);
and U7180 (N_7180,N_1164,N_2083);
and U7181 (N_7181,N_3029,N_4946);
nand U7182 (N_7182,N_226,N_3564);
nor U7183 (N_7183,N_2762,N_3509);
and U7184 (N_7184,N_4547,N_2997);
and U7185 (N_7185,N_3818,N_4392);
and U7186 (N_7186,N_871,N_3276);
and U7187 (N_7187,N_803,N_691);
nand U7188 (N_7188,N_4132,N_4803);
nor U7189 (N_7189,N_4929,N_3107);
nor U7190 (N_7190,N_4008,N_4978);
or U7191 (N_7191,N_4130,N_2502);
or U7192 (N_7192,N_3681,N_1176);
nor U7193 (N_7193,N_1982,N_2441);
or U7194 (N_7194,N_4111,N_410);
xnor U7195 (N_7195,N_4794,N_1309);
and U7196 (N_7196,N_1979,N_4698);
nand U7197 (N_7197,N_478,N_4077);
and U7198 (N_7198,N_1741,N_2306);
and U7199 (N_7199,N_320,N_3090);
nand U7200 (N_7200,N_3852,N_441);
or U7201 (N_7201,N_1220,N_1475);
nor U7202 (N_7202,N_2388,N_1915);
and U7203 (N_7203,N_1641,N_394);
nor U7204 (N_7204,N_4854,N_552);
nor U7205 (N_7205,N_3323,N_3998);
nor U7206 (N_7206,N_615,N_2087);
and U7207 (N_7207,N_3529,N_4829);
or U7208 (N_7208,N_2646,N_4066);
nor U7209 (N_7209,N_164,N_1860);
or U7210 (N_7210,N_2443,N_555);
or U7211 (N_7211,N_2577,N_2057);
nand U7212 (N_7212,N_1133,N_224);
or U7213 (N_7213,N_4215,N_3858);
nor U7214 (N_7214,N_1270,N_2973);
or U7215 (N_7215,N_3441,N_3203);
or U7216 (N_7216,N_1392,N_3209);
nand U7217 (N_7217,N_161,N_2933);
or U7218 (N_7218,N_1684,N_962);
nand U7219 (N_7219,N_1275,N_4287);
and U7220 (N_7220,N_4770,N_4490);
and U7221 (N_7221,N_3875,N_3689);
and U7222 (N_7222,N_1155,N_3363);
nor U7223 (N_7223,N_3789,N_3296);
nand U7224 (N_7224,N_3721,N_4426);
nand U7225 (N_7225,N_1748,N_3337);
nand U7226 (N_7226,N_1701,N_3927);
and U7227 (N_7227,N_2258,N_676);
nand U7228 (N_7228,N_1503,N_897);
and U7229 (N_7229,N_2393,N_31);
xnor U7230 (N_7230,N_2151,N_1108);
nand U7231 (N_7231,N_76,N_914);
nand U7232 (N_7232,N_3860,N_1857);
or U7233 (N_7233,N_3190,N_3628);
and U7234 (N_7234,N_1191,N_4078);
or U7235 (N_7235,N_428,N_1665);
or U7236 (N_7236,N_4275,N_2897);
or U7237 (N_7237,N_3448,N_3545);
nor U7238 (N_7238,N_1789,N_941);
or U7239 (N_7239,N_550,N_3410);
nand U7240 (N_7240,N_2249,N_2123);
nand U7241 (N_7241,N_2240,N_3419);
or U7242 (N_7242,N_4780,N_923);
nand U7243 (N_7243,N_2261,N_1961);
or U7244 (N_7244,N_3887,N_3364);
and U7245 (N_7245,N_4083,N_1365);
or U7246 (N_7246,N_587,N_2236);
and U7247 (N_7247,N_1900,N_3563);
nor U7248 (N_7248,N_2869,N_3608);
nand U7249 (N_7249,N_2526,N_4292);
or U7250 (N_7250,N_1817,N_26);
and U7251 (N_7251,N_2523,N_1473);
and U7252 (N_7252,N_705,N_2130);
xnor U7253 (N_7253,N_940,N_4171);
nand U7254 (N_7254,N_2823,N_4565);
xnor U7255 (N_7255,N_1130,N_2354);
nor U7256 (N_7256,N_3089,N_2295);
nand U7257 (N_7257,N_40,N_4416);
xor U7258 (N_7258,N_2183,N_943);
nand U7259 (N_7259,N_247,N_1148);
or U7260 (N_7260,N_1569,N_4960);
nand U7261 (N_7261,N_2810,N_4129);
nand U7262 (N_7262,N_445,N_3743);
nand U7263 (N_7263,N_4690,N_2129);
nand U7264 (N_7264,N_1530,N_3672);
nand U7265 (N_7265,N_4194,N_3173);
nor U7266 (N_7266,N_2269,N_2309);
and U7267 (N_7267,N_4491,N_750);
or U7268 (N_7268,N_3808,N_4748);
nand U7269 (N_7269,N_104,N_1518);
nor U7270 (N_7270,N_3994,N_3637);
nor U7271 (N_7271,N_515,N_3655);
and U7272 (N_7272,N_1451,N_2230);
and U7273 (N_7273,N_2416,N_4989);
or U7274 (N_7274,N_2839,N_2906);
or U7275 (N_7275,N_1586,N_1887);
and U7276 (N_7276,N_1932,N_417);
nand U7277 (N_7277,N_3020,N_3640);
nand U7278 (N_7278,N_2509,N_2397);
nand U7279 (N_7279,N_116,N_507);
and U7280 (N_7280,N_3349,N_2120);
xor U7281 (N_7281,N_246,N_1778);
nand U7282 (N_7282,N_3303,N_4348);
nor U7283 (N_7283,N_3839,N_3085);
nand U7284 (N_7284,N_2028,N_4160);
nor U7285 (N_7285,N_4680,N_91);
nand U7286 (N_7286,N_4671,N_3911);
nand U7287 (N_7287,N_4233,N_3548);
or U7288 (N_7288,N_4977,N_1564);
or U7289 (N_7289,N_988,N_49);
nand U7290 (N_7290,N_2198,N_1228);
and U7291 (N_7291,N_3251,N_25);
nor U7292 (N_7292,N_1834,N_1227);
or U7293 (N_7293,N_4294,N_714);
and U7294 (N_7294,N_2832,N_113);
nor U7295 (N_7295,N_2127,N_1268);
nand U7296 (N_7296,N_2558,N_4316);
and U7297 (N_7297,N_925,N_3446);
nand U7298 (N_7298,N_608,N_1836);
nor U7299 (N_7299,N_610,N_2215);
nor U7300 (N_7300,N_3351,N_3167);
and U7301 (N_7301,N_2565,N_1205);
and U7302 (N_7302,N_2467,N_1899);
xnor U7303 (N_7303,N_3733,N_3034);
or U7304 (N_7304,N_4667,N_227);
and U7305 (N_7305,N_1523,N_2735);
nor U7306 (N_7306,N_4982,N_1980);
and U7307 (N_7307,N_1152,N_1279);
or U7308 (N_7308,N_2430,N_2286);
nand U7309 (N_7309,N_4313,N_2859);
or U7310 (N_7310,N_3552,N_1731);
or U7311 (N_7311,N_1400,N_1235);
and U7312 (N_7312,N_4057,N_4355);
or U7313 (N_7313,N_3813,N_3830);
nand U7314 (N_7314,N_695,N_4796);
nor U7315 (N_7315,N_4735,N_1104);
nand U7316 (N_7316,N_150,N_3451);
or U7317 (N_7317,N_189,N_2959);
and U7318 (N_7318,N_4425,N_1411);
nand U7319 (N_7319,N_3212,N_687);
nand U7320 (N_7320,N_4901,N_3517);
nand U7321 (N_7321,N_1119,N_3411);
nor U7322 (N_7322,N_3116,N_1603);
or U7323 (N_7323,N_3127,N_957);
or U7324 (N_7324,N_3964,N_3091);
and U7325 (N_7325,N_567,N_4714);
and U7326 (N_7326,N_4400,N_3646);
or U7327 (N_7327,N_3154,N_425);
or U7328 (N_7328,N_3088,N_2224);
nor U7329 (N_7329,N_333,N_931);
nor U7330 (N_7330,N_977,N_2280);
and U7331 (N_7331,N_2907,N_463);
or U7332 (N_7332,N_72,N_1375);
nor U7333 (N_7333,N_836,N_3062);
nand U7334 (N_7334,N_2980,N_4969);
and U7335 (N_7335,N_2168,N_349);
or U7336 (N_7336,N_1488,N_1549);
or U7337 (N_7337,N_4613,N_1515);
and U7338 (N_7338,N_762,N_2527);
nand U7339 (N_7339,N_255,N_2911);
nor U7340 (N_7340,N_3734,N_2714);
nor U7341 (N_7341,N_1051,N_1868);
or U7342 (N_7342,N_2407,N_3753);
nor U7343 (N_7343,N_2506,N_3382);
nand U7344 (N_7344,N_3692,N_1114);
or U7345 (N_7345,N_3566,N_485);
nand U7346 (N_7346,N_4104,N_1097);
and U7347 (N_7347,N_1419,N_915);
or U7348 (N_7348,N_368,N_1238);
nand U7349 (N_7349,N_2287,N_1992);
nand U7350 (N_7350,N_2160,N_2655);
nand U7351 (N_7351,N_3444,N_4921);
or U7352 (N_7352,N_4624,N_1068);
nand U7353 (N_7353,N_4655,N_4453);
nor U7354 (N_7354,N_2631,N_3598);
or U7355 (N_7355,N_2184,N_2433);
nor U7356 (N_7356,N_505,N_2686);
and U7357 (N_7357,N_1002,N_4717);
nor U7358 (N_7358,N_1760,N_4021);
nand U7359 (N_7359,N_1136,N_2716);
nand U7360 (N_7360,N_4952,N_3802);
nor U7361 (N_7361,N_1977,N_1099);
nor U7362 (N_7362,N_2718,N_1008);
and U7363 (N_7363,N_2811,N_3027);
nand U7364 (N_7364,N_1985,N_4696);
nand U7365 (N_7365,N_1880,N_3422);
nand U7366 (N_7366,N_2324,N_3211);
nand U7367 (N_7367,N_782,N_4732);
and U7368 (N_7368,N_1565,N_780);
nor U7369 (N_7369,N_2796,N_3570);
nor U7370 (N_7370,N_3093,N_3408);
xor U7371 (N_7371,N_4326,N_1132);
or U7372 (N_7372,N_4197,N_5);
or U7373 (N_7373,N_1072,N_4437);
or U7374 (N_7374,N_2621,N_3981);
nand U7375 (N_7375,N_3412,N_3996);
nand U7376 (N_7376,N_3534,N_1506);
nor U7377 (N_7377,N_2690,N_3728);
nor U7378 (N_7378,N_354,N_1892);
and U7379 (N_7379,N_4060,N_3921);
and U7380 (N_7380,N_557,N_3238);
or U7381 (N_7381,N_3215,N_4700);
or U7382 (N_7382,N_1495,N_2844);
nand U7383 (N_7383,N_2825,N_1061);
nand U7384 (N_7384,N_2195,N_1245);
and U7385 (N_7385,N_2769,N_3851);
and U7386 (N_7386,N_241,N_1216);
nand U7387 (N_7387,N_2414,N_2172);
xor U7388 (N_7388,N_473,N_812);
or U7389 (N_7389,N_4467,N_4798);
or U7390 (N_7390,N_1654,N_1558);
and U7391 (N_7391,N_3214,N_3078);
nor U7392 (N_7392,N_4654,N_4011);
nor U7393 (N_7393,N_4976,N_3391);
and U7394 (N_7394,N_4760,N_46);
nor U7395 (N_7395,N_3556,N_2912);
or U7396 (N_7396,N_1180,N_805);
nor U7397 (N_7397,N_1472,N_2296);
nor U7398 (N_7398,N_900,N_4167);
nand U7399 (N_7399,N_3454,N_4602);
and U7400 (N_7400,N_1283,N_4422);
nand U7401 (N_7401,N_3693,N_3775);
xnor U7402 (N_7402,N_4728,N_4843);
xnor U7403 (N_7403,N_746,N_193);
nor U7404 (N_7404,N_853,N_2756);
or U7405 (N_7405,N_2010,N_813);
or U7406 (N_7406,N_2957,N_1307);
nand U7407 (N_7407,N_582,N_3222);
and U7408 (N_7408,N_3122,N_1161);
nand U7409 (N_7409,N_592,N_1800);
nor U7410 (N_7410,N_2875,N_4906);
and U7411 (N_7411,N_4109,N_4199);
nand U7412 (N_7412,N_2503,N_3896);
nor U7413 (N_7413,N_3025,N_4148);
or U7414 (N_7414,N_3757,N_1580);
nand U7415 (N_7415,N_2684,N_1671);
and U7416 (N_7416,N_360,N_3254);
and U7417 (N_7417,N_4776,N_4620);
nand U7418 (N_7418,N_4591,N_483);
and U7419 (N_7419,N_514,N_2893);
and U7420 (N_7420,N_1987,N_3600);
nand U7421 (N_7421,N_2038,N_586);
nand U7422 (N_7422,N_400,N_1492);
nand U7423 (N_7423,N_2612,N_1877);
nor U7424 (N_7424,N_1414,N_2591);
or U7425 (N_7425,N_4380,N_2176);
nand U7426 (N_7426,N_135,N_3506);
nor U7427 (N_7427,N_1310,N_2870);
or U7428 (N_7428,N_3530,N_4440);
nand U7429 (N_7429,N_3048,N_141);
nor U7430 (N_7430,N_4692,N_3811);
nor U7431 (N_7431,N_1232,N_4533);
or U7432 (N_7432,N_1149,N_2048);
or U7433 (N_7433,N_4824,N_2454);
and U7434 (N_7434,N_2916,N_3845);
and U7435 (N_7435,N_4339,N_450);
nand U7436 (N_7436,N_617,N_3973);
nor U7437 (N_7437,N_3223,N_3680);
or U7438 (N_7438,N_1593,N_3774);
nor U7439 (N_7439,N_3944,N_2352);
and U7440 (N_7440,N_2968,N_196);
or U7441 (N_7441,N_2392,N_616);
nor U7442 (N_7442,N_3978,N_2913);
nor U7443 (N_7443,N_2219,N_1732);
or U7444 (N_7444,N_4302,N_2438);
and U7445 (N_7445,N_2303,N_2356);
nand U7446 (N_7446,N_3781,N_3061);
nor U7447 (N_7447,N_1333,N_4814);
and U7448 (N_7448,N_4121,N_2683);
nor U7449 (N_7449,N_1328,N_1522);
or U7450 (N_7450,N_3460,N_2592);
nor U7451 (N_7451,N_679,N_4687);
nor U7452 (N_7452,N_4383,N_1584);
or U7453 (N_7453,N_4884,N_4962);
nor U7454 (N_7454,N_2516,N_3070);
nor U7455 (N_7455,N_1388,N_4336);
or U7456 (N_7456,N_2248,N_118);
nor U7457 (N_7457,N_3003,N_3260);
nor U7458 (N_7458,N_2161,N_383);
and U7459 (N_7459,N_2475,N_1225);
nor U7460 (N_7460,N_2493,N_3979);
or U7461 (N_7461,N_4587,N_2081);
and U7462 (N_7462,N_4045,N_1890);
nor U7463 (N_7463,N_209,N_930);
nor U7464 (N_7464,N_2436,N_1305);
nand U7465 (N_7465,N_2966,N_500);
nand U7466 (N_7466,N_3393,N_4475);
or U7467 (N_7467,N_4532,N_2587);
and U7468 (N_7468,N_600,N_4651);
nand U7469 (N_7469,N_3606,N_4032);
or U7470 (N_7470,N_23,N_155);
and U7471 (N_7471,N_2327,N_4481);
xor U7472 (N_7472,N_573,N_2583);
or U7473 (N_7473,N_4265,N_2891);
and U7474 (N_7474,N_905,N_1281);
nand U7475 (N_7475,N_3092,N_4830);
or U7476 (N_7476,N_2218,N_4364);
nor U7477 (N_7477,N_3701,N_2149);
or U7478 (N_7478,N_4005,N_1844);
xor U7479 (N_7479,N_2574,N_4115);
nor U7480 (N_7480,N_2216,N_4747);
and U7481 (N_7481,N_1353,N_44);
or U7482 (N_7482,N_4099,N_4880);
or U7483 (N_7483,N_2539,N_1871);
and U7484 (N_7484,N_407,N_1547);
nand U7485 (N_7485,N_2247,N_1862);
and U7486 (N_7486,N_3694,N_4802);
nor U7487 (N_7487,N_720,N_729);
nand U7488 (N_7488,N_2405,N_1070);
nor U7489 (N_7489,N_3316,N_2225);
nand U7490 (N_7490,N_4891,N_4114);
and U7491 (N_7491,N_2790,N_2560);
nor U7492 (N_7492,N_165,N_4535);
nor U7493 (N_7493,N_870,N_3286);
or U7494 (N_7494,N_3076,N_3188);
or U7495 (N_7495,N_2632,N_4858);
or U7496 (N_7496,N_4464,N_2470);
and U7497 (N_7497,N_3236,N_1384);
and U7498 (N_7498,N_4689,N_2474);
nand U7499 (N_7499,N_3021,N_4195);
nor U7500 (N_7500,N_400,N_1610);
nand U7501 (N_7501,N_4639,N_3089);
or U7502 (N_7502,N_2862,N_3620);
nand U7503 (N_7503,N_1710,N_3022);
or U7504 (N_7504,N_3635,N_2485);
or U7505 (N_7505,N_2139,N_3209);
nand U7506 (N_7506,N_1111,N_3946);
or U7507 (N_7507,N_4348,N_2951);
nand U7508 (N_7508,N_4633,N_1863);
nor U7509 (N_7509,N_3873,N_1117);
or U7510 (N_7510,N_3942,N_4952);
nor U7511 (N_7511,N_4182,N_4176);
nor U7512 (N_7512,N_2549,N_2931);
nand U7513 (N_7513,N_3093,N_2465);
nor U7514 (N_7514,N_4113,N_546);
and U7515 (N_7515,N_376,N_3235);
or U7516 (N_7516,N_4447,N_1949);
and U7517 (N_7517,N_52,N_2896);
or U7518 (N_7518,N_1677,N_3965);
and U7519 (N_7519,N_1493,N_1008);
or U7520 (N_7520,N_4071,N_264);
nor U7521 (N_7521,N_4661,N_1789);
nand U7522 (N_7522,N_941,N_3625);
nor U7523 (N_7523,N_3399,N_1119);
nor U7524 (N_7524,N_749,N_2792);
nand U7525 (N_7525,N_2772,N_3435);
and U7526 (N_7526,N_2274,N_375);
nand U7527 (N_7527,N_2553,N_1570);
and U7528 (N_7528,N_746,N_261);
nand U7529 (N_7529,N_3422,N_1379);
nor U7530 (N_7530,N_3053,N_3347);
and U7531 (N_7531,N_1938,N_4002);
or U7532 (N_7532,N_1938,N_2225);
xnor U7533 (N_7533,N_2997,N_2140);
nor U7534 (N_7534,N_2277,N_2169);
nor U7535 (N_7535,N_4318,N_3616);
nand U7536 (N_7536,N_622,N_390);
nand U7537 (N_7537,N_809,N_3694);
nor U7538 (N_7538,N_799,N_2460);
or U7539 (N_7539,N_3994,N_3100);
nor U7540 (N_7540,N_606,N_2663);
and U7541 (N_7541,N_1196,N_2989);
or U7542 (N_7542,N_3118,N_2654);
nand U7543 (N_7543,N_4504,N_565);
nor U7544 (N_7544,N_3511,N_1878);
or U7545 (N_7545,N_668,N_4763);
or U7546 (N_7546,N_137,N_3588);
and U7547 (N_7547,N_1679,N_964);
nor U7548 (N_7548,N_3477,N_3883);
or U7549 (N_7549,N_4044,N_3678);
nor U7550 (N_7550,N_139,N_3399);
nor U7551 (N_7551,N_4850,N_686);
nand U7552 (N_7552,N_3889,N_3816);
and U7553 (N_7553,N_1080,N_2828);
xnor U7554 (N_7554,N_3680,N_125);
nor U7555 (N_7555,N_253,N_517);
or U7556 (N_7556,N_450,N_4343);
and U7557 (N_7557,N_1246,N_3666);
or U7558 (N_7558,N_1854,N_4314);
nor U7559 (N_7559,N_2759,N_2976);
nand U7560 (N_7560,N_3691,N_1886);
and U7561 (N_7561,N_3285,N_2923);
nor U7562 (N_7562,N_607,N_3201);
or U7563 (N_7563,N_174,N_1059);
nand U7564 (N_7564,N_1168,N_982);
or U7565 (N_7565,N_4003,N_4038);
or U7566 (N_7566,N_868,N_3737);
xnor U7567 (N_7567,N_4514,N_5);
nor U7568 (N_7568,N_726,N_3564);
nor U7569 (N_7569,N_3735,N_3458);
nor U7570 (N_7570,N_950,N_2399);
nand U7571 (N_7571,N_3034,N_2301);
nor U7572 (N_7572,N_3094,N_4317);
nand U7573 (N_7573,N_2852,N_641);
nand U7574 (N_7574,N_4362,N_3501);
nand U7575 (N_7575,N_948,N_287);
or U7576 (N_7576,N_4239,N_3918);
xnor U7577 (N_7577,N_3551,N_3388);
nand U7578 (N_7578,N_433,N_1317);
and U7579 (N_7579,N_905,N_3396);
nand U7580 (N_7580,N_1990,N_2134);
or U7581 (N_7581,N_1151,N_2477);
nor U7582 (N_7582,N_3009,N_4751);
or U7583 (N_7583,N_883,N_511);
or U7584 (N_7584,N_4812,N_4349);
nand U7585 (N_7585,N_4382,N_3572);
nor U7586 (N_7586,N_1413,N_2893);
nand U7587 (N_7587,N_2547,N_2380);
and U7588 (N_7588,N_22,N_364);
or U7589 (N_7589,N_2932,N_1980);
nand U7590 (N_7590,N_3556,N_4117);
and U7591 (N_7591,N_1553,N_4379);
nor U7592 (N_7592,N_3386,N_390);
nand U7593 (N_7593,N_1777,N_4168);
nand U7594 (N_7594,N_2064,N_3707);
nor U7595 (N_7595,N_3011,N_869);
nand U7596 (N_7596,N_1431,N_2877);
nor U7597 (N_7597,N_421,N_825);
and U7598 (N_7598,N_2334,N_3140);
nor U7599 (N_7599,N_146,N_189);
and U7600 (N_7600,N_2434,N_259);
and U7601 (N_7601,N_1207,N_3804);
or U7602 (N_7602,N_3570,N_2663);
nand U7603 (N_7603,N_1126,N_1984);
and U7604 (N_7604,N_4890,N_4261);
nor U7605 (N_7605,N_3163,N_1179);
and U7606 (N_7606,N_1702,N_1100);
nand U7607 (N_7607,N_3825,N_1712);
or U7608 (N_7608,N_321,N_2734);
nor U7609 (N_7609,N_1516,N_2869);
or U7610 (N_7610,N_1822,N_1497);
nor U7611 (N_7611,N_2828,N_2390);
and U7612 (N_7612,N_2863,N_4417);
or U7613 (N_7613,N_1123,N_4516);
nor U7614 (N_7614,N_4,N_1552);
and U7615 (N_7615,N_2692,N_1568);
nor U7616 (N_7616,N_4123,N_4007);
or U7617 (N_7617,N_1876,N_2903);
nand U7618 (N_7618,N_2614,N_1014);
or U7619 (N_7619,N_942,N_3382);
nor U7620 (N_7620,N_1481,N_979);
nor U7621 (N_7621,N_3528,N_4604);
nand U7622 (N_7622,N_1309,N_4219);
or U7623 (N_7623,N_2027,N_652);
nor U7624 (N_7624,N_4116,N_1767);
nor U7625 (N_7625,N_4391,N_482);
or U7626 (N_7626,N_1528,N_1953);
xor U7627 (N_7627,N_1911,N_2594);
nand U7628 (N_7628,N_3693,N_1960);
nand U7629 (N_7629,N_1487,N_2512);
or U7630 (N_7630,N_1758,N_2154);
nor U7631 (N_7631,N_2676,N_4642);
nor U7632 (N_7632,N_2252,N_1299);
and U7633 (N_7633,N_2525,N_1004);
and U7634 (N_7634,N_2611,N_315);
nor U7635 (N_7635,N_203,N_558);
and U7636 (N_7636,N_2022,N_20);
nand U7637 (N_7637,N_4925,N_2240);
nor U7638 (N_7638,N_2455,N_4435);
or U7639 (N_7639,N_1391,N_2693);
and U7640 (N_7640,N_2303,N_2081);
nor U7641 (N_7641,N_4813,N_677);
xnor U7642 (N_7642,N_3352,N_3754);
nor U7643 (N_7643,N_1106,N_793);
and U7644 (N_7644,N_4696,N_3924);
or U7645 (N_7645,N_3398,N_2263);
nand U7646 (N_7646,N_2507,N_157);
nor U7647 (N_7647,N_253,N_3418);
and U7648 (N_7648,N_4219,N_4546);
nor U7649 (N_7649,N_2105,N_272);
or U7650 (N_7650,N_1162,N_3917);
nand U7651 (N_7651,N_3061,N_1735);
or U7652 (N_7652,N_1480,N_4201);
nand U7653 (N_7653,N_4257,N_2034);
or U7654 (N_7654,N_2163,N_3095);
nand U7655 (N_7655,N_2304,N_737);
nand U7656 (N_7656,N_568,N_2637);
nor U7657 (N_7657,N_4010,N_2396);
xnor U7658 (N_7658,N_4028,N_4115);
or U7659 (N_7659,N_47,N_2801);
and U7660 (N_7660,N_4673,N_3328);
nand U7661 (N_7661,N_1507,N_4804);
or U7662 (N_7662,N_3188,N_2177);
or U7663 (N_7663,N_3857,N_4360);
or U7664 (N_7664,N_3861,N_4261);
nor U7665 (N_7665,N_781,N_2951);
nor U7666 (N_7666,N_1830,N_2377);
nand U7667 (N_7667,N_3216,N_737);
or U7668 (N_7668,N_4205,N_2386);
nor U7669 (N_7669,N_4903,N_2986);
and U7670 (N_7670,N_4567,N_1481);
or U7671 (N_7671,N_2024,N_971);
nor U7672 (N_7672,N_4847,N_814);
nand U7673 (N_7673,N_2964,N_302);
nand U7674 (N_7674,N_4612,N_3507);
nand U7675 (N_7675,N_3814,N_2458);
nor U7676 (N_7676,N_4916,N_566);
nor U7677 (N_7677,N_4620,N_4334);
nor U7678 (N_7678,N_228,N_555);
nand U7679 (N_7679,N_4949,N_515);
nor U7680 (N_7680,N_572,N_4627);
or U7681 (N_7681,N_3376,N_1121);
and U7682 (N_7682,N_1041,N_1243);
nor U7683 (N_7683,N_3270,N_119);
or U7684 (N_7684,N_3781,N_2386);
nor U7685 (N_7685,N_807,N_4224);
nor U7686 (N_7686,N_915,N_1383);
xor U7687 (N_7687,N_3574,N_520);
or U7688 (N_7688,N_2183,N_2240);
nand U7689 (N_7689,N_98,N_1716);
nor U7690 (N_7690,N_3908,N_234);
or U7691 (N_7691,N_2184,N_1571);
and U7692 (N_7692,N_1171,N_4142);
nor U7693 (N_7693,N_1451,N_2928);
nor U7694 (N_7694,N_1027,N_3160);
or U7695 (N_7695,N_854,N_876);
or U7696 (N_7696,N_575,N_4127);
nand U7697 (N_7697,N_3578,N_4124);
xor U7698 (N_7698,N_2257,N_2151);
nand U7699 (N_7699,N_1770,N_176);
nand U7700 (N_7700,N_186,N_2488);
nand U7701 (N_7701,N_4794,N_1440);
or U7702 (N_7702,N_4837,N_4949);
or U7703 (N_7703,N_1658,N_264);
nor U7704 (N_7704,N_764,N_4897);
nand U7705 (N_7705,N_4441,N_2817);
nand U7706 (N_7706,N_4312,N_3074);
and U7707 (N_7707,N_4368,N_623);
or U7708 (N_7708,N_416,N_547);
nor U7709 (N_7709,N_50,N_528);
nor U7710 (N_7710,N_2081,N_1192);
or U7711 (N_7711,N_4853,N_3019);
and U7712 (N_7712,N_3725,N_4701);
nand U7713 (N_7713,N_1541,N_2503);
nand U7714 (N_7714,N_2725,N_4406);
nor U7715 (N_7715,N_3069,N_4398);
nor U7716 (N_7716,N_4418,N_1678);
nor U7717 (N_7717,N_4807,N_3546);
nor U7718 (N_7718,N_1772,N_2268);
and U7719 (N_7719,N_2286,N_4054);
and U7720 (N_7720,N_4597,N_159);
and U7721 (N_7721,N_2453,N_1311);
nor U7722 (N_7722,N_4452,N_980);
nand U7723 (N_7723,N_3174,N_4828);
nor U7724 (N_7724,N_1486,N_1947);
or U7725 (N_7725,N_2644,N_899);
nand U7726 (N_7726,N_2731,N_1363);
nand U7727 (N_7727,N_1498,N_1802);
or U7728 (N_7728,N_1551,N_1853);
and U7729 (N_7729,N_3051,N_988);
or U7730 (N_7730,N_2378,N_145);
nor U7731 (N_7731,N_1104,N_2521);
and U7732 (N_7732,N_3140,N_4972);
nand U7733 (N_7733,N_4953,N_4151);
and U7734 (N_7734,N_914,N_4736);
nand U7735 (N_7735,N_275,N_2940);
and U7736 (N_7736,N_4354,N_1313);
nor U7737 (N_7737,N_2292,N_4438);
nor U7738 (N_7738,N_1248,N_4278);
nand U7739 (N_7739,N_1507,N_2669);
and U7740 (N_7740,N_2531,N_2942);
and U7741 (N_7741,N_3876,N_4091);
or U7742 (N_7742,N_612,N_1672);
and U7743 (N_7743,N_2607,N_936);
nor U7744 (N_7744,N_1186,N_4815);
nor U7745 (N_7745,N_1904,N_1448);
and U7746 (N_7746,N_1680,N_3081);
nand U7747 (N_7747,N_4605,N_4619);
nor U7748 (N_7748,N_4439,N_518);
nor U7749 (N_7749,N_1984,N_4143);
nand U7750 (N_7750,N_2648,N_3512);
nand U7751 (N_7751,N_2677,N_4081);
nor U7752 (N_7752,N_4215,N_921);
nor U7753 (N_7753,N_1447,N_3211);
nand U7754 (N_7754,N_3446,N_805);
xor U7755 (N_7755,N_4091,N_621);
or U7756 (N_7756,N_4428,N_4716);
and U7757 (N_7757,N_4322,N_3603);
nor U7758 (N_7758,N_3289,N_578);
or U7759 (N_7759,N_1323,N_3076);
nand U7760 (N_7760,N_1770,N_4878);
or U7761 (N_7761,N_3880,N_1442);
or U7762 (N_7762,N_2971,N_2408);
nor U7763 (N_7763,N_522,N_3256);
nor U7764 (N_7764,N_3816,N_4091);
nor U7765 (N_7765,N_4597,N_2497);
nor U7766 (N_7766,N_326,N_2375);
nor U7767 (N_7767,N_3889,N_1786);
nand U7768 (N_7768,N_4028,N_3948);
nor U7769 (N_7769,N_1736,N_1617);
nand U7770 (N_7770,N_4507,N_4896);
and U7771 (N_7771,N_3482,N_3898);
nand U7772 (N_7772,N_4456,N_4066);
or U7773 (N_7773,N_345,N_4344);
xor U7774 (N_7774,N_364,N_4092);
nand U7775 (N_7775,N_1716,N_3661);
or U7776 (N_7776,N_3276,N_4378);
nand U7777 (N_7777,N_2854,N_4747);
nand U7778 (N_7778,N_54,N_117);
nor U7779 (N_7779,N_4483,N_4694);
nand U7780 (N_7780,N_1128,N_460);
and U7781 (N_7781,N_4035,N_2971);
or U7782 (N_7782,N_3051,N_4808);
nand U7783 (N_7783,N_3313,N_2787);
nand U7784 (N_7784,N_1771,N_2522);
and U7785 (N_7785,N_3359,N_1511);
nand U7786 (N_7786,N_1405,N_3491);
or U7787 (N_7787,N_3012,N_2809);
or U7788 (N_7788,N_484,N_4421);
and U7789 (N_7789,N_3460,N_4759);
nand U7790 (N_7790,N_3856,N_2053);
nand U7791 (N_7791,N_1476,N_63);
or U7792 (N_7792,N_1189,N_1124);
nand U7793 (N_7793,N_1238,N_870);
nand U7794 (N_7794,N_860,N_581);
or U7795 (N_7795,N_4972,N_1255);
and U7796 (N_7796,N_4387,N_2201);
nand U7797 (N_7797,N_329,N_3838);
nand U7798 (N_7798,N_397,N_794);
nor U7799 (N_7799,N_1528,N_1546);
and U7800 (N_7800,N_871,N_3087);
nand U7801 (N_7801,N_3309,N_1633);
or U7802 (N_7802,N_613,N_2265);
nand U7803 (N_7803,N_2523,N_2901);
or U7804 (N_7804,N_1286,N_3907);
and U7805 (N_7805,N_3254,N_4048);
or U7806 (N_7806,N_4021,N_1510);
nor U7807 (N_7807,N_4083,N_2753);
or U7808 (N_7808,N_1548,N_931);
nor U7809 (N_7809,N_1620,N_1055);
nor U7810 (N_7810,N_359,N_1405);
nand U7811 (N_7811,N_2539,N_4680);
nor U7812 (N_7812,N_2166,N_257);
or U7813 (N_7813,N_271,N_1613);
or U7814 (N_7814,N_3703,N_2808);
nor U7815 (N_7815,N_365,N_4151);
nor U7816 (N_7816,N_2017,N_4449);
nand U7817 (N_7817,N_2283,N_4110);
or U7818 (N_7818,N_2041,N_4223);
nor U7819 (N_7819,N_352,N_3526);
nand U7820 (N_7820,N_4454,N_387);
nand U7821 (N_7821,N_2845,N_1316);
nand U7822 (N_7822,N_1850,N_1467);
nor U7823 (N_7823,N_4147,N_3547);
nand U7824 (N_7824,N_3461,N_2591);
or U7825 (N_7825,N_1882,N_149);
or U7826 (N_7826,N_4609,N_4624);
and U7827 (N_7827,N_2276,N_4751);
nor U7828 (N_7828,N_1572,N_2008);
or U7829 (N_7829,N_1899,N_2794);
and U7830 (N_7830,N_927,N_4119);
nand U7831 (N_7831,N_531,N_4661);
nand U7832 (N_7832,N_487,N_2441);
nand U7833 (N_7833,N_1618,N_3063);
and U7834 (N_7834,N_898,N_1332);
nand U7835 (N_7835,N_4988,N_4141);
nand U7836 (N_7836,N_582,N_2610);
xor U7837 (N_7837,N_2686,N_1871);
and U7838 (N_7838,N_3679,N_1476);
nor U7839 (N_7839,N_4428,N_4077);
nand U7840 (N_7840,N_3740,N_4864);
nand U7841 (N_7841,N_1278,N_4541);
or U7842 (N_7842,N_1212,N_710);
or U7843 (N_7843,N_2412,N_512);
and U7844 (N_7844,N_2021,N_2131);
and U7845 (N_7845,N_3607,N_4953);
or U7846 (N_7846,N_1378,N_480);
and U7847 (N_7847,N_1339,N_4020);
nand U7848 (N_7848,N_4347,N_336);
nor U7849 (N_7849,N_1398,N_1721);
and U7850 (N_7850,N_1128,N_1430);
nor U7851 (N_7851,N_482,N_2123);
nor U7852 (N_7852,N_2943,N_1657);
or U7853 (N_7853,N_3958,N_3464);
nand U7854 (N_7854,N_3501,N_3053);
xor U7855 (N_7855,N_1595,N_3122);
nand U7856 (N_7856,N_4022,N_4033);
nor U7857 (N_7857,N_3126,N_4287);
and U7858 (N_7858,N_713,N_3424);
and U7859 (N_7859,N_410,N_1438);
nand U7860 (N_7860,N_1065,N_1575);
nand U7861 (N_7861,N_3421,N_2660);
nand U7862 (N_7862,N_3799,N_2903);
nand U7863 (N_7863,N_3716,N_1079);
nand U7864 (N_7864,N_3674,N_274);
nor U7865 (N_7865,N_4416,N_3383);
or U7866 (N_7866,N_2296,N_903);
nor U7867 (N_7867,N_1859,N_3805);
nor U7868 (N_7868,N_1074,N_3575);
or U7869 (N_7869,N_679,N_4961);
nand U7870 (N_7870,N_1573,N_4704);
and U7871 (N_7871,N_606,N_2176);
or U7872 (N_7872,N_1197,N_186);
and U7873 (N_7873,N_889,N_303);
nand U7874 (N_7874,N_4192,N_1687);
or U7875 (N_7875,N_4775,N_3863);
or U7876 (N_7876,N_123,N_816);
nor U7877 (N_7877,N_1479,N_1099);
or U7878 (N_7878,N_827,N_2116);
and U7879 (N_7879,N_2709,N_3486);
nand U7880 (N_7880,N_2160,N_1322);
nand U7881 (N_7881,N_2858,N_3892);
and U7882 (N_7882,N_2513,N_1344);
or U7883 (N_7883,N_31,N_3895);
nor U7884 (N_7884,N_1573,N_3820);
or U7885 (N_7885,N_3870,N_4252);
or U7886 (N_7886,N_2216,N_2601);
nand U7887 (N_7887,N_2534,N_3862);
nand U7888 (N_7888,N_3647,N_1213);
nor U7889 (N_7889,N_672,N_1535);
or U7890 (N_7890,N_3212,N_3337);
nand U7891 (N_7891,N_1495,N_4416);
and U7892 (N_7892,N_1758,N_2720);
or U7893 (N_7893,N_563,N_4545);
nand U7894 (N_7894,N_4662,N_1246);
and U7895 (N_7895,N_3401,N_3842);
nand U7896 (N_7896,N_3829,N_1776);
and U7897 (N_7897,N_3748,N_197);
nor U7898 (N_7898,N_555,N_2223);
nand U7899 (N_7899,N_1739,N_3301);
and U7900 (N_7900,N_571,N_1442);
and U7901 (N_7901,N_2996,N_2489);
and U7902 (N_7902,N_4980,N_226);
nor U7903 (N_7903,N_1195,N_1319);
nand U7904 (N_7904,N_1655,N_1018);
nand U7905 (N_7905,N_150,N_960);
and U7906 (N_7906,N_4971,N_4026);
nor U7907 (N_7907,N_2033,N_175);
or U7908 (N_7908,N_3579,N_1275);
nor U7909 (N_7909,N_3381,N_3609);
xor U7910 (N_7910,N_4434,N_3030);
nand U7911 (N_7911,N_56,N_2677);
nand U7912 (N_7912,N_4462,N_3796);
nand U7913 (N_7913,N_2520,N_3073);
nor U7914 (N_7914,N_3395,N_1400);
nand U7915 (N_7915,N_4289,N_1195);
or U7916 (N_7916,N_643,N_2321);
and U7917 (N_7917,N_4858,N_734);
nand U7918 (N_7918,N_1183,N_2941);
nor U7919 (N_7919,N_3827,N_1254);
nor U7920 (N_7920,N_792,N_946);
and U7921 (N_7921,N_802,N_773);
and U7922 (N_7922,N_2308,N_4537);
and U7923 (N_7923,N_4641,N_2603);
or U7924 (N_7924,N_4223,N_1703);
and U7925 (N_7925,N_243,N_4956);
and U7926 (N_7926,N_994,N_3522);
nor U7927 (N_7927,N_2223,N_1240);
nor U7928 (N_7928,N_2493,N_2519);
and U7929 (N_7929,N_3868,N_1966);
or U7930 (N_7930,N_1232,N_3231);
and U7931 (N_7931,N_162,N_3903);
nand U7932 (N_7932,N_4241,N_1203);
and U7933 (N_7933,N_4482,N_4088);
and U7934 (N_7934,N_2705,N_543);
and U7935 (N_7935,N_3282,N_1766);
nor U7936 (N_7936,N_148,N_231);
nand U7937 (N_7937,N_2922,N_1456);
and U7938 (N_7938,N_4646,N_22);
nand U7939 (N_7939,N_4470,N_2484);
nor U7940 (N_7940,N_462,N_1759);
and U7941 (N_7941,N_4931,N_4713);
and U7942 (N_7942,N_2995,N_236);
nand U7943 (N_7943,N_875,N_3759);
or U7944 (N_7944,N_1267,N_1670);
nand U7945 (N_7945,N_3172,N_1255);
and U7946 (N_7946,N_4197,N_1294);
and U7947 (N_7947,N_3920,N_3356);
nor U7948 (N_7948,N_4617,N_3011);
xor U7949 (N_7949,N_3499,N_4476);
nor U7950 (N_7950,N_2543,N_3652);
nor U7951 (N_7951,N_830,N_3107);
and U7952 (N_7952,N_1787,N_2120);
or U7953 (N_7953,N_975,N_1415);
nand U7954 (N_7954,N_4239,N_4182);
or U7955 (N_7955,N_420,N_4508);
nor U7956 (N_7956,N_1295,N_538);
and U7957 (N_7957,N_1177,N_120);
nand U7958 (N_7958,N_101,N_1507);
and U7959 (N_7959,N_4220,N_3045);
nand U7960 (N_7960,N_3287,N_4829);
nor U7961 (N_7961,N_4094,N_815);
or U7962 (N_7962,N_3635,N_1000);
or U7963 (N_7963,N_4028,N_1816);
nor U7964 (N_7964,N_4867,N_2062);
nand U7965 (N_7965,N_2857,N_1204);
or U7966 (N_7966,N_4901,N_1405);
and U7967 (N_7967,N_1656,N_1677);
nand U7968 (N_7968,N_1359,N_3603);
nand U7969 (N_7969,N_4446,N_3495);
and U7970 (N_7970,N_4902,N_1792);
nor U7971 (N_7971,N_2335,N_3650);
nand U7972 (N_7972,N_2030,N_1904);
or U7973 (N_7973,N_2438,N_2576);
and U7974 (N_7974,N_1722,N_2563);
or U7975 (N_7975,N_4957,N_543);
and U7976 (N_7976,N_1639,N_633);
and U7977 (N_7977,N_781,N_530);
nor U7978 (N_7978,N_4464,N_3654);
or U7979 (N_7979,N_2648,N_79);
and U7980 (N_7980,N_4912,N_1964);
nand U7981 (N_7981,N_2028,N_2733);
and U7982 (N_7982,N_4415,N_1571);
nor U7983 (N_7983,N_1973,N_86);
nor U7984 (N_7984,N_3818,N_1849);
or U7985 (N_7985,N_3436,N_987);
nor U7986 (N_7986,N_3533,N_2352);
and U7987 (N_7987,N_1059,N_2802);
or U7988 (N_7988,N_526,N_4397);
nor U7989 (N_7989,N_1464,N_1429);
or U7990 (N_7990,N_2937,N_62);
or U7991 (N_7991,N_73,N_2273);
nand U7992 (N_7992,N_4551,N_648);
nor U7993 (N_7993,N_2974,N_2155);
and U7994 (N_7994,N_648,N_4030);
or U7995 (N_7995,N_4730,N_2568);
nor U7996 (N_7996,N_2322,N_864);
and U7997 (N_7997,N_137,N_2521);
nor U7998 (N_7998,N_1412,N_4713);
and U7999 (N_7999,N_2556,N_125);
or U8000 (N_8000,N_2244,N_4946);
or U8001 (N_8001,N_1170,N_1161);
and U8002 (N_8002,N_4122,N_4845);
nor U8003 (N_8003,N_4791,N_3521);
and U8004 (N_8004,N_4312,N_1292);
and U8005 (N_8005,N_1920,N_1585);
nor U8006 (N_8006,N_4438,N_1395);
or U8007 (N_8007,N_1740,N_3708);
nand U8008 (N_8008,N_1853,N_1132);
nand U8009 (N_8009,N_1717,N_123);
nor U8010 (N_8010,N_1949,N_1588);
or U8011 (N_8011,N_512,N_2189);
or U8012 (N_8012,N_3737,N_3113);
nor U8013 (N_8013,N_4518,N_569);
xnor U8014 (N_8014,N_3709,N_4789);
nor U8015 (N_8015,N_262,N_1910);
nand U8016 (N_8016,N_2197,N_2420);
and U8017 (N_8017,N_4406,N_3286);
and U8018 (N_8018,N_4322,N_992);
nand U8019 (N_8019,N_3452,N_1533);
nand U8020 (N_8020,N_3069,N_4890);
or U8021 (N_8021,N_2371,N_155);
and U8022 (N_8022,N_4503,N_2690);
and U8023 (N_8023,N_3785,N_4334);
nand U8024 (N_8024,N_2612,N_3348);
xnor U8025 (N_8025,N_4708,N_3493);
nor U8026 (N_8026,N_1288,N_3853);
and U8027 (N_8027,N_2925,N_4777);
nand U8028 (N_8028,N_3216,N_2803);
and U8029 (N_8029,N_247,N_3406);
nor U8030 (N_8030,N_3467,N_3945);
and U8031 (N_8031,N_1271,N_3902);
or U8032 (N_8032,N_2884,N_4163);
and U8033 (N_8033,N_4218,N_2400);
nor U8034 (N_8034,N_61,N_966);
or U8035 (N_8035,N_4304,N_4894);
and U8036 (N_8036,N_1761,N_2973);
nand U8037 (N_8037,N_1405,N_1205);
nand U8038 (N_8038,N_3712,N_3179);
and U8039 (N_8039,N_1298,N_1275);
nor U8040 (N_8040,N_3731,N_646);
or U8041 (N_8041,N_266,N_1939);
and U8042 (N_8042,N_64,N_811);
and U8043 (N_8043,N_2045,N_657);
nor U8044 (N_8044,N_4666,N_3693);
or U8045 (N_8045,N_1053,N_2559);
and U8046 (N_8046,N_4107,N_2640);
nor U8047 (N_8047,N_246,N_3836);
or U8048 (N_8048,N_238,N_3075);
and U8049 (N_8049,N_1987,N_22);
nand U8050 (N_8050,N_1702,N_4459);
nand U8051 (N_8051,N_1911,N_3269);
or U8052 (N_8052,N_3295,N_1835);
nand U8053 (N_8053,N_616,N_325);
xnor U8054 (N_8054,N_2588,N_1866);
or U8055 (N_8055,N_3133,N_4028);
xor U8056 (N_8056,N_3747,N_2454);
nand U8057 (N_8057,N_1630,N_1407);
or U8058 (N_8058,N_2050,N_1937);
nand U8059 (N_8059,N_361,N_18);
and U8060 (N_8060,N_568,N_1620);
nand U8061 (N_8061,N_3304,N_3668);
nor U8062 (N_8062,N_1792,N_1833);
or U8063 (N_8063,N_605,N_2919);
nand U8064 (N_8064,N_4203,N_711);
xor U8065 (N_8065,N_1424,N_3457);
or U8066 (N_8066,N_4135,N_737);
nand U8067 (N_8067,N_1427,N_4721);
nand U8068 (N_8068,N_4585,N_37);
nor U8069 (N_8069,N_1855,N_4271);
nor U8070 (N_8070,N_3962,N_267);
xnor U8071 (N_8071,N_664,N_4605);
and U8072 (N_8072,N_176,N_2910);
nand U8073 (N_8073,N_4409,N_2308);
and U8074 (N_8074,N_1073,N_4378);
nor U8075 (N_8075,N_2845,N_2594);
or U8076 (N_8076,N_2121,N_3911);
or U8077 (N_8077,N_3572,N_679);
nor U8078 (N_8078,N_4602,N_3911);
nor U8079 (N_8079,N_3924,N_2647);
nand U8080 (N_8080,N_2212,N_3794);
nor U8081 (N_8081,N_4730,N_707);
nor U8082 (N_8082,N_4436,N_2246);
nor U8083 (N_8083,N_4365,N_1940);
nor U8084 (N_8084,N_2166,N_1581);
or U8085 (N_8085,N_3771,N_4964);
and U8086 (N_8086,N_2874,N_4773);
or U8087 (N_8087,N_1012,N_976);
and U8088 (N_8088,N_4310,N_4519);
nor U8089 (N_8089,N_1731,N_4947);
or U8090 (N_8090,N_698,N_1277);
nand U8091 (N_8091,N_1728,N_4093);
or U8092 (N_8092,N_3654,N_2194);
nand U8093 (N_8093,N_13,N_944);
nand U8094 (N_8094,N_1767,N_4434);
or U8095 (N_8095,N_3309,N_2055);
and U8096 (N_8096,N_4368,N_1838);
and U8097 (N_8097,N_3530,N_2238);
nand U8098 (N_8098,N_2293,N_2200);
or U8099 (N_8099,N_919,N_4262);
nor U8100 (N_8100,N_3232,N_4285);
or U8101 (N_8101,N_2797,N_1747);
nor U8102 (N_8102,N_2841,N_2087);
nand U8103 (N_8103,N_1761,N_2984);
nor U8104 (N_8104,N_4973,N_812);
and U8105 (N_8105,N_1155,N_2479);
nor U8106 (N_8106,N_2887,N_1825);
or U8107 (N_8107,N_3338,N_3433);
and U8108 (N_8108,N_2073,N_3835);
or U8109 (N_8109,N_1505,N_4148);
nor U8110 (N_8110,N_2603,N_4344);
nand U8111 (N_8111,N_99,N_4013);
nor U8112 (N_8112,N_874,N_1038);
and U8113 (N_8113,N_1557,N_4100);
nor U8114 (N_8114,N_4594,N_4449);
and U8115 (N_8115,N_1894,N_3276);
nor U8116 (N_8116,N_1880,N_2970);
or U8117 (N_8117,N_3882,N_4602);
and U8118 (N_8118,N_3717,N_3684);
nor U8119 (N_8119,N_3383,N_2839);
nand U8120 (N_8120,N_1840,N_3843);
and U8121 (N_8121,N_455,N_3508);
and U8122 (N_8122,N_936,N_1778);
or U8123 (N_8123,N_4204,N_4847);
or U8124 (N_8124,N_755,N_3494);
or U8125 (N_8125,N_349,N_2130);
nor U8126 (N_8126,N_525,N_2767);
nor U8127 (N_8127,N_2986,N_2164);
or U8128 (N_8128,N_598,N_3573);
nand U8129 (N_8129,N_3674,N_2017);
nand U8130 (N_8130,N_2225,N_4966);
and U8131 (N_8131,N_3918,N_1194);
nand U8132 (N_8132,N_4612,N_989);
and U8133 (N_8133,N_579,N_467);
and U8134 (N_8134,N_1104,N_3080);
and U8135 (N_8135,N_3501,N_885);
or U8136 (N_8136,N_1062,N_642);
nor U8137 (N_8137,N_242,N_4280);
and U8138 (N_8138,N_1905,N_4474);
or U8139 (N_8139,N_2744,N_864);
nor U8140 (N_8140,N_63,N_2264);
and U8141 (N_8141,N_2993,N_2229);
nor U8142 (N_8142,N_3231,N_102);
nor U8143 (N_8143,N_1415,N_1387);
nand U8144 (N_8144,N_3461,N_293);
or U8145 (N_8145,N_4813,N_1617);
or U8146 (N_8146,N_2527,N_891);
nand U8147 (N_8147,N_3265,N_3307);
xnor U8148 (N_8148,N_3266,N_1508);
and U8149 (N_8149,N_792,N_341);
nand U8150 (N_8150,N_4823,N_2398);
or U8151 (N_8151,N_395,N_4953);
nor U8152 (N_8152,N_2691,N_3977);
and U8153 (N_8153,N_581,N_3257);
and U8154 (N_8154,N_4412,N_2421);
nor U8155 (N_8155,N_167,N_3599);
nor U8156 (N_8156,N_514,N_3406);
and U8157 (N_8157,N_1709,N_3119);
nor U8158 (N_8158,N_4149,N_1538);
and U8159 (N_8159,N_3314,N_3002);
nor U8160 (N_8160,N_4520,N_3909);
nand U8161 (N_8161,N_547,N_1490);
or U8162 (N_8162,N_4591,N_727);
and U8163 (N_8163,N_2993,N_2954);
nor U8164 (N_8164,N_37,N_4145);
nor U8165 (N_8165,N_2517,N_382);
nand U8166 (N_8166,N_1173,N_2188);
and U8167 (N_8167,N_4783,N_1473);
nand U8168 (N_8168,N_2164,N_1369);
nand U8169 (N_8169,N_971,N_283);
nor U8170 (N_8170,N_736,N_1701);
nand U8171 (N_8171,N_883,N_2961);
nor U8172 (N_8172,N_4262,N_4899);
and U8173 (N_8173,N_4864,N_1909);
and U8174 (N_8174,N_1905,N_4127);
nand U8175 (N_8175,N_4542,N_4285);
nand U8176 (N_8176,N_1005,N_4909);
nor U8177 (N_8177,N_3368,N_1077);
nor U8178 (N_8178,N_1396,N_3551);
nor U8179 (N_8179,N_1249,N_3260);
and U8180 (N_8180,N_152,N_1489);
and U8181 (N_8181,N_2882,N_1891);
and U8182 (N_8182,N_2572,N_2699);
nand U8183 (N_8183,N_2335,N_1827);
and U8184 (N_8184,N_3578,N_2051);
nor U8185 (N_8185,N_3379,N_4345);
nand U8186 (N_8186,N_3085,N_1845);
nand U8187 (N_8187,N_2326,N_3335);
nand U8188 (N_8188,N_1679,N_3995);
and U8189 (N_8189,N_282,N_504);
or U8190 (N_8190,N_3586,N_2116);
and U8191 (N_8191,N_4288,N_46);
nand U8192 (N_8192,N_4234,N_4390);
and U8193 (N_8193,N_4707,N_2032);
nand U8194 (N_8194,N_2886,N_1616);
and U8195 (N_8195,N_1431,N_2150);
nand U8196 (N_8196,N_2833,N_3219);
nor U8197 (N_8197,N_863,N_1153);
or U8198 (N_8198,N_4998,N_3284);
nor U8199 (N_8199,N_2458,N_4873);
or U8200 (N_8200,N_388,N_4294);
and U8201 (N_8201,N_3093,N_2094);
nor U8202 (N_8202,N_4494,N_3609);
nand U8203 (N_8203,N_31,N_3000);
nor U8204 (N_8204,N_4985,N_4108);
nand U8205 (N_8205,N_337,N_4875);
nor U8206 (N_8206,N_3479,N_2992);
nor U8207 (N_8207,N_4883,N_3809);
and U8208 (N_8208,N_371,N_4074);
or U8209 (N_8209,N_330,N_3802);
and U8210 (N_8210,N_223,N_1888);
nor U8211 (N_8211,N_3843,N_206);
or U8212 (N_8212,N_841,N_1263);
and U8213 (N_8213,N_4246,N_1150);
or U8214 (N_8214,N_748,N_1649);
or U8215 (N_8215,N_3333,N_3497);
nor U8216 (N_8216,N_2586,N_3299);
nor U8217 (N_8217,N_4366,N_3048);
and U8218 (N_8218,N_3813,N_1458);
or U8219 (N_8219,N_2443,N_1594);
and U8220 (N_8220,N_745,N_4799);
or U8221 (N_8221,N_4986,N_2733);
xor U8222 (N_8222,N_689,N_1771);
xor U8223 (N_8223,N_3465,N_2713);
and U8224 (N_8224,N_4240,N_3513);
and U8225 (N_8225,N_2326,N_2748);
or U8226 (N_8226,N_1130,N_1013);
or U8227 (N_8227,N_3511,N_2356);
nand U8228 (N_8228,N_1809,N_2471);
or U8229 (N_8229,N_4579,N_2929);
nand U8230 (N_8230,N_1291,N_1900);
nand U8231 (N_8231,N_4983,N_3377);
nor U8232 (N_8232,N_2886,N_3982);
nand U8233 (N_8233,N_1204,N_3115);
nand U8234 (N_8234,N_333,N_2193);
nor U8235 (N_8235,N_3487,N_2484);
and U8236 (N_8236,N_1426,N_229);
nor U8237 (N_8237,N_4995,N_381);
and U8238 (N_8238,N_4045,N_593);
nor U8239 (N_8239,N_2256,N_4545);
and U8240 (N_8240,N_1814,N_256);
or U8241 (N_8241,N_2233,N_4243);
nor U8242 (N_8242,N_1008,N_3500);
or U8243 (N_8243,N_2900,N_3510);
nor U8244 (N_8244,N_1997,N_660);
and U8245 (N_8245,N_2865,N_2584);
nand U8246 (N_8246,N_917,N_3179);
or U8247 (N_8247,N_2182,N_3879);
nand U8248 (N_8248,N_3558,N_3309);
and U8249 (N_8249,N_2126,N_1548);
nor U8250 (N_8250,N_3407,N_1580);
or U8251 (N_8251,N_4398,N_2993);
and U8252 (N_8252,N_1448,N_823);
nor U8253 (N_8253,N_3189,N_3483);
and U8254 (N_8254,N_3139,N_1507);
nand U8255 (N_8255,N_1839,N_4273);
nor U8256 (N_8256,N_1393,N_3599);
nand U8257 (N_8257,N_1427,N_1254);
or U8258 (N_8258,N_3436,N_3876);
or U8259 (N_8259,N_1714,N_435);
or U8260 (N_8260,N_3603,N_2052);
and U8261 (N_8261,N_4527,N_2543);
nor U8262 (N_8262,N_4219,N_2068);
or U8263 (N_8263,N_1563,N_2531);
nor U8264 (N_8264,N_1576,N_2556);
xor U8265 (N_8265,N_960,N_375);
nand U8266 (N_8266,N_898,N_1775);
nand U8267 (N_8267,N_1152,N_1602);
or U8268 (N_8268,N_1212,N_1989);
and U8269 (N_8269,N_889,N_1188);
or U8270 (N_8270,N_264,N_332);
xor U8271 (N_8271,N_212,N_4361);
nand U8272 (N_8272,N_3151,N_4320);
and U8273 (N_8273,N_1533,N_2667);
nand U8274 (N_8274,N_938,N_3515);
or U8275 (N_8275,N_2284,N_2655);
and U8276 (N_8276,N_4504,N_3623);
nor U8277 (N_8277,N_2882,N_2572);
nand U8278 (N_8278,N_1646,N_3170);
and U8279 (N_8279,N_2914,N_3304);
nand U8280 (N_8280,N_1848,N_867);
and U8281 (N_8281,N_1799,N_1251);
and U8282 (N_8282,N_2144,N_135);
and U8283 (N_8283,N_4554,N_2053);
and U8284 (N_8284,N_4145,N_2564);
nand U8285 (N_8285,N_3926,N_259);
and U8286 (N_8286,N_1757,N_1144);
xnor U8287 (N_8287,N_3242,N_1770);
nand U8288 (N_8288,N_2264,N_3212);
nand U8289 (N_8289,N_1639,N_4202);
nor U8290 (N_8290,N_3227,N_403);
nor U8291 (N_8291,N_1921,N_913);
and U8292 (N_8292,N_3647,N_2495);
nor U8293 (N_8293,N_445,N_563);
nor U8294 (N_8294,N_13,N_2603);
nor U8295 (N_8295,N_1010,N_973);
or U8296 (N_8296,N_2324,N_4915);
or U8297 (N_8297,N_1466,N_3033);
nor U8298 (N_8298,N_3412,N_3137);
nand U8299 (N_8299,N_3079,N_19);
and U8300 (N_8300,N_2904,N_1106);
nand U8301 (N_8301,N_1642,N_2046);
or U8302 (N_8302,N_1483,N_1361);
or U8303 (N_8303,N_2816,N_2097);
nand U8304 (N_8304,N_2538,N_4730);
nor U8305 (N_8305,N_3226,N_2241);
nand U8306 (N_8306,N_4104,N_2299);
and U8307 (N_8307,N_1210,N_1216);
and U8308 (N_8308,N_4351,N_2778);
nand U8309 (N_8309,N_258,N_913);
and U8310 (N_8310,N_1854,N_2480);
nand U8311 (N_8311,N_996,N_4982);
nor U8312 (N_8312,N_1139,N_3702);
nor U8313 (N_8313,N_129,N_911);
nand U8314 (N_8314,N_2841,N_2487);
nor U8315 (N_8315,N_2492,N_2117);
nor U8316 (N_8316,N_3879,N_4681);
xor U8317 (N_8317,N_2843,N_4624);
nand U8318 (N_8318,N_4867,N_1134);
and U8319 (N_8319,N_2988,N_4589);
nand U8320 (N_8320,N_1312,N_966);
and U8321 (N_8321,N_1377,N_3258);
and U8322 (N_8322,N_3354,N_4084);
nand U8323 (N_8323,N_1772,N_1047);
or U8324 (N_8324,N_2547,N_1049);
nor U8325 (N_8325,N_2369,N_500);
nor U8326 (N_8326,N_4503,N_481);
nor U8327 (N_8327,N_1122,N_3656);
or U8328 (N_8328,N_44,N_1913);
or U8329 (N_8329,N_197,N_4966);
nor U8330 (N_8330,N_4712,N_2778);
nor U8331 (N_8331,N_2935,N_4003);
nand U8332 (N_8332,N_310,N_4578);
and U8333 (N_8333,N_1037,N_2005);
nor U8334 (N_8334,N_4301,N_250);
nor U8335 (N_8335,N_573,N_263);
nand U8336 (N_8336,N_1088,N_485);
nand U8337 (N_8337,N_2239,N_3727);
or U8338 (N_8338,N_3989,N_3504);
nor U8339 (N_8339,N_3241,N_4175);
and U8340 (N_8340,N_4852,N_1355);
nor U8341 (N_8341,N_1384,N_2079);
nand U8342 (N_8342,N_1882,N_4974);
or U8343 (N_8343,N_1628,N_2106);
nand U8344 (N_8344,N_3135,N_2995);
nand U8345 (N_8345,N_1899,N_3863);
xnor U8346 (N_8346,N_2583,N_3389);
and U8347 (N_8347,N_1607,N_4678);
and U8348 (N_8348,N_3230,N_2929);
nand U8349 (N_8349,N_670,N_2595);
nand U8350 (N_8350,N_3099,N_3638);
or U8351 (N_8351,N_955,N_1771);
and U8352 (N_8352,N_764,N_1382);
and U8353 (N_8353,N_1618,N_3823);
and U8354 (N_8354,N_4671,N_696);
or U8355 (N_8355,N_207,N_1443);
nor U8356 (N_8356,N_2534,N_3451);
or U8357 (N_8357,N_3822,N_1965);
nor U8358 (N_8358,N_4434,N_3820);
or U8359 (N_8359,N_2624,N_403);
or U8360 (N_8360,N_3062,N_3748);
and U8361 (N_8361,N_2569,N_3601);
nor U8362 (N_8362,N_207,N_3061);
nand U8363 (N_8363,N_3542,N_1817);
nor U8364 (N_8364,N_4232,N_2416);
xnor U8365 (N_8365,N_4986,N_2547);
nor U8366 (N_8366,N_1642,N_3507);
or U8367 (N_8367,N_4959,N_4087);
nand U8368 (N_8368,N_4561,N_2067);
nand U8369 (N_8369,N_3253,N_3617);
nand U8370 (N_8370,N_177,N_4899);
nand U8371 (N_8371,N_642,N_1440);
and U8372 (N_8372,N_732,N_2538);
and U8373 (N_8373,N_1227,N_2111);
nand U8374 (N_8374,N_1732,N_983);
or U8375 (N_8375,N_279,N_1961);
nor U8376 (N_8376,N_4579,N_143);
nor U8377 (N_8377,N_4495,N_3377);
nand U8378 (N_8378,N_4204,N_4249);
or U8379 (N_8379,N_4126,N_568);
nand U8380 (N_8380,N_1126,N_899);
nand U8381 (N_8381,N_2665,N_4242);
or U8382 (N_8382,N_3199,N_3440);
or U8383 (N_8383,N_1708,N_928);
nor U8384 (N_8384,N_2995,N_4607);
and U8385 (N_8385,N_2739,N_3016);
or U8386 (N_8386,N_4451,N_3888);
and U8387 (N_8387,N_4800,N_2676);
or U8388 (N_8388,N_2432,N_4315);
nor U8389 (N_8389,N_4484,N_264);
or U8390 (N_8390,N_1877,N_1123);
or U8391 (N_8391,N_1943,N_429);
and U8392 (N_8392,N_2549,N_4996);
nand U8393 (N_8393,N_4864,N_1798);
nor U8394 (N_8394,N_203,N_3994);
nor U8395 (N_8395,N_3277,N_4007);
nor U8396 (N_8396,N_3399,N_3105);
and U8397 (N_8397,N_134,N_1235);
nand U8398 (N_8398,N_4402,N_3824);
nor U8399 (N_8399,N_3787,N_2828);
nor U8400 (N_8400,N_825,N_2924);
nand U8401 (N_8401,N_947,N_3992);
nand U8402 (N_8402,N_2168,N_2469);
nand U8403 (N_8403,N_2740,N_4926);
and U8404 (N_8404,N_2388,N_1188);
and U8405 (N_8405,N_292,N_3450);
nand U8406 (N_8406,N_3266,N_4181);
or U8407 (N_8407,N_3643,N_3657);
and U8408 (N_8408,N_3648,N_3383);
nor U8409 (N_8409,N_2210,N_188);
nand U8410 (N_8410,N_559,N_3444);
nor U8411 (N_8411,N_2681,N_1487);
nand U8412 (N_8412,N_1415,N_2088);
nand U8413 (N_8413,N_160,N_1359);
nor U8414 (N_8414,N_4467,N_1898);
xnor U8415 (N_8415,N_324,N_1064);
nor U8416 (N_8416,N_1926,N_3368);
nor U8417 (N_8417,N_3486,N_432);
or U8418 (N_8418,N_2291,N_3073);
or U8419 (N_8419,N_4117,N_4016);
and U8420 (N_8420,N_3888,N_2983);
nor U8421 (N_8421,N_840,N_4271);
nand U8422 (N_8422,N_3173,N_3755);
or U8423 (N_8423,N_1021,N_622);
nand U8424 (N_8424,N_838,N_1208);
nor U8425 (N_8425,N_4516,N_1666);
nor U8426 (N_8426,N_4161,N_4122);
or U8427 (N_8427,N_235,N_4470);
or U8428 (N_8428,N_2201,N_1300);
and U8429 (N_8429,N_3307,N_3629);
and U8430 (N_8430,N_3955,N_1763);
xnor U8431 (N_8431,N_2082,N_1464);
and U8432 (N_8432,N_372,N_1341);
and U8433 (N_8433,N_4045,N_766);
nor U8434 (N_8434,N_92,N_3341);
nor U8435 (N_8435,N_546,N_39);
or U8436 (N_8436,N_1296,N_4470);
and U8437 (N_8437,N_2753,N_2825);
nor U8438 (N_8438,N_171,N_1360);
nand U8439 (N_8439,N_4543,N_3652);
or U8440 (N_8440,N_3707,N_1780);
nand U8441 (N_8441,N_3153,N_1453);
and U8442 (N_8442,N_4242,N_3077);
nor U8443 (N_8443,N_1523,N_3005);
nor U8444 (N_8444,N_984,N_2453);
nand U8445 (N_8445,N_4763,N_1452);
nor U8446 (N_8446,N_3740,N_3699);
nor U8447 (N_8447,N_718,N_3404);
or U8448 (N_8448,N_1278,N_4658);
and U8449 (N_8449,N_2674,N_546);
or U8450 (N_8450,N_1525,N_899);
nor U8451 (N_8451,N_4663,N_1414);
nor U8452 (N_8452,N_2870,N_269);
or U8453 (N_8453,N_114,N_2924);
and U8454 (N_8454,N_1353,N_1318);
nor U8455 (N_8455,N_1394,N_3434);
and U8456 (N_8456,N_130,N_2453);
or U8457 (N_8457,N_1554,N_3026);
nor U8458 (N_8458,N_1478,N_207);
nor U8459 (N_8459,N_4988,N_4251);
or U8460 (N_8460,N_11,N_476);
or U8461 (N_8461,N_2136,N_1483);
or U8462 (N_8462,N_1264,N_2368);
nand U8463 (N_8463,N_2442,N_1268);
xnor U8464 (N_8464,N_1829,N_2341);
xnor U8465 (N_8465,N_549,N_3466);
xnor U8466 (N_8466,N_1039,N_4474);
nor U8467 (N_8467,N_3253,N_2751);
nor U8468 (N_8468,N_1484,N_327);
or U8469 (N_8469,N_3126,N_2973);
nand U8470 (N_8470,N_3886,N_1653);
nor U8471 (N_8471,N_4296,N_2331);
nor U8472 (N_8472,N_4769,N_85);
or U8473 (N_8473,N_268,N_525);
or U8474 (N_8474,N_4738,N_1573);
nand U8475 (N_8475,N_2800,N_4336);
or U8476 (N_8476,N_1221,N_4148);
nor U8477 (N_8477,N_2587,N_2680);
or U8478 (N_8478,N_1770,N_4158);
nor U8479 (N_8479,N_2068,N_3235);
or U8480 (N_8480,N_4411,N_2312);
and U8481 (N_8481,N_1936,N_3150);
or U8482 (N_8482,N_4837,N_3877);
and U8483 (N_8483,N_4273,N_1299);
and U8484 (N_8484,N_881,N_4641);
and U8485 (N_8485,N_461,N_475);
nor U8486 (N_8486,N_1298,N_2189);
or U8487 (N_8487,N_447,N_72);
and U8488 (N_8488,N_4382,N_855);
nor U8489 (N_8489,N_265,N_403);
xor U8490 (N_8490,N_2385,N_3037);
or U8491 (N_8491,N_2796,N_3954);
nand U8492 (N_8492,N_938,N_3872);
and U8493 (N_8493,N_3071,N_2486);
nand U8494 (N_8494,N_4186,N_3875);
nor U8495 (N_8495,N_2172,N_2219);
or U8496 (N_8496,N_2320,N_1572);
nor U8497 (N_8497,N_2579,N_943);
and U8498 (N_8498,N_479,N_3397);
and U8499 (N_8499,N_3579,N_1974);
or U8500 (N_8500,N_2622,N_1505);
or U8501 (N_8501,N_4727,N_4337);
nand U8502 (N_8502,N_159,N_3040);
xor U8503 (N_8503,N_4864,N_4022);
or U8504 (N_8504,N_3688,N_645);
nand U8505 (N_8505,N_2265,N_1389);
and U8506 (N_8506,N_4328,N_3433);
or U8507 (N_8507,N_543,N_4795);
or U8508 (N_8508,N_1567,N_2331);
nor U8509 (N_8509,N_1012,N_3030);
nand U8510 (N_8510,N_4050,N_2346);
and U8511 (N_8511,N_3805,N_750);
nor U8512 (N_8512,N_785,N_346);
and U8513 (N_8513,N_2570,N_2930);
or U8514 (N_8514,N_2051,N_4708);
and U8515 (N_8515,N_982,N_4437);
nand U8516 (N_8516,N_4643,N_214);
nor U8517 (N_8517,N_2540,N_3131);
nor U8518 (N_8518,N_1173,N_596);
and U8519 (N_8519,N_1902,N_2327);
nand U8520 (N_8520,N_644,N_1964);
or U8521 (N_8521,N_2255,N_440);
nor U8522 (N_8522,N_2279,N_4872);
nand U8523 (N_8523,N_109,N_3981);
nand U8524 (N_8524,N_1566,N_4369);
nor U8525 (N_8525,N_4085,N_3559);
nand U8526 (N_8526,N_2313,N_3955);
and U8527 (N_8527,N_490,N_62);
nand U8528 (N_8528,N_304,N_2776);
or U8529 (N_8529,N_2264,N_341);
nor U8530 (N_8530,N_2876,N_2615);
nand U8531 (N_8531,N_345,N_625);
or U8532 (N_8532,N_2843,N_3780);
nand U8533 (N_8533,N_786,N_2743);
nand U8534 (N_8534,N_3998,N_1651);
and U8535 (N_8535,N_2153,N_4297);
nor U8536 (N_8536,N_3057,N_4756);
or U8537 (N_8537,N_4962,N_4117);
nand U8538 (N_8538,N_2086,N_1363);
nand U8539 (N_8539,N_570,N_4728);
and U8540 (N_8540,N_3513,N_431);
or U8541 (N_8541,N_4194,N_1952);
or U8542 (N_8542,N_250,N_1384);
nand U8543 (N_8543,N_1543,N_3487);
and U8544 (N_8544,N_3403,N_4493);
nor U8545 (N_8545,N_1401,N_3615);
and U8546 (N_8546,N_4602,N_3147);
or U8547 (N_8547,N_3731,N_3123);
and U8548 (N_8548,N_2273,N_1433);
or U8549 (N_8549,N_1491,N_3275);
xor U8550 (N_8550,N_582,N_2255);
or U8551 (N_8551,N_2492,N_4398);
nand U8552 (N_8552,N_3778,N_4691);
nor U8553 (N_8553,N_113,N_1708);
or U8554 (N_8554,N_2497,N_891);
nand U8555 (N_8555,N_3147,N_1576);
nor U8556 (N_8556,N_4098,N_632);
or U8557 (N_8557,N_2032,N_4568);
and U8558 (N_8558,N_2460,N_953);
nand U8559 (N_8559,N_4621,N_92);
nand U8560 (N_8560,N_231,N_4445);
nand U8561 (N_8561,N_2046,N_3830);
or U8562 (N_8562,N_4982,N_966);
nor U8563 (N_8563,N_140,N_1095);
xor U8564 (N_8564,N_3928,N_212);
nand U8565 (N_8565,N_3996,N_4732);
and U8566 (N_8566,N_4122,N_4462);
and U8567 (N_8567,N_4793,N_891);
or U8568 (N_8568,N_2606,N_1358);
and U8569 (N_8569,N_3181,N_3120);
and U8570 (N_8570,N_2214,N_4836);
nor U8571 (N_8571,N_4924,N_4949);
and U8572 (N_8572,N_3746,N_4820);
nor U8573 (N_8573,N_1683,N_2451);
and U8574 (N_8574,N_3182,N_732);
nand U8575 (N_8575,N_1136,N_4732);
nor U8576 (N_8576,N_3427,N_539);
or U8577 (N_8577,N_2858,N_3669);
or U8578 (N_8578,N_3917,N_3487);
nand U8579 (N_8579,N_1463,N_4920);
nor U8580 (N_8580,N_1386,N_3126);
nor U8581 (N_8581,N_4004,N_4362);
nor U8582 (N_8582,N_4724,N_688);
nand U8583 (N_8583,N_4497,N_2795);
nand U8584 (N_8584,N_3775,N_3402);
or U8585 (N_8585,N_1181,N_2009);
or U8586 (N_8586,N_178,N_2540);
nand U8587 (N_8587,N_4741,N_383);
nand U8588 (N_8588,N_37,N_3765);
nor U8589 (N_8589,N_1174,N_869);
nand U8590 (N_8590,N_278,N_222);
nor U8591 (N_8591,N_2819,N_3306);
or U8592 (N_8592,N_1731,N_881);
and U8593 (N_8593,N_1912,N_1020);
nor U8594 (N_8594,N_1037,N_2875);
nand U8595 (N_8595,N_3376,N_1874);
xor U8596 (N_8596,N_4407,N_3498);
or U8597 (N_8597,N_543,N_3299);
nand U8598 (N_8598,N_2847,N_3509);
and U8599 (N_8599,N_52,N_4802);
and U8600 (N_8600,N_485,N_1977);
or U8601 (N_8601,N_1266,N_4927);
nand U8602 (N_8602,N_2423,N_1066);
and U8603 (N_8603,N_2729,N_508);
and U8604 (N_8604,N_1854,N_2120);
nand U8605 (N_8605,N_223,N_885);
nor U8606 (N_8606,N_3763,N_4698);
and U8607 (N_8607,N_4154,N_1264);
nand U8608 (N_8608,N_4713,N_435);
nand U8609 (N_8609,N_1987,N_1525);
nor U8610 (N_8610,N_2698,N_3908);
nand U8611 (N_8611,N_184,N_4811);
or U8612 (N_8612,N_3003,N_4490);
and U8613 (N_8613,N_2394,N_2984);
nand U8614 (N_8614,N_3016,N_1736);
and U8615 (N_8615,N_2956,N_3323);
nor U8616 (N_8616,N_615,N_4262);
xnor U8617 (N_8617,N_292,N_3661);
nand U8618 (N_8618,N_4895,N_3118);
nand U8619 (N_8619,N_362,N_3397);
or U8620 (N_8620,N_2491,N_2196);
nand U8621 (N_8621,N_3430,N_3915);
nor U8622 (N_8622,N_4604,N_1004);
nand U8623 (N_8623,N_3731,N_1387);
and U8624 (N_8624,N_4647,N_637);
and U8625 (N_8625,N_3992,N_1424);
or U8626 (N_8626,N_4892,N_4364);
xor U8627 (N_8627,N_973,N_4907);
nand U8628 (N_8628,N_4251,N_2931);
and U8629 (N_8629,N_3737,N_4344);
and U8630 (N_8630,N_4564,N_956);
and U8631 (N_8631,N_55,N_1275);
and U8632 (N_8632,N_2370,N_4215);
nor U8633 (N_8633,N_1499,N_945);
or U8634 (N_8634,N_2221,N_3089);
nor U8635 (N_8635,N_1440,N_1116);
and U8636 (N_8636,N_1310,N_78);
nand U8637 (N_8637,N_4436,N_146);
nor U8638 (N_8638,N_2020,N_4701);
or U8639 (N_8639,N_3550,N_310);
or U8640 (N_8640,N_2959,N_3491);
nor U8641 (N_8641,N_1111,N_2196);
nor U8642 (N_8642,N_2688,N_3173);
or U8643 (N_8643,N_1184,N_744);
nor U8644 (N_8644,N_97,N_479);
nor U8645 (N_8645,N_4741,N_2570);
and U8646 (N_8646,N_3249,N_3028);
nand U8647 (N_8647,N_0,N_3849);
and U8648 (N_8648,N_688,N_1597);
nor U8649 (N_8649,N_238,N_3913);
nand U8650 (N_8650,N_3081,N_4599);
nand U8651 (N_8651,N_2964,N_1808);
and U8652 (N_8652,N_2545,N_1313);
nor U8653 (N_8653,N_2704,N_2591);
nand U8654 (N_8654,N_169,N_3584);
nand U8655 (N_8655,N_4984,N_4566);
nor U8656 (N_8656,N_4772,N_1077);
and U8657 (N_8657,N_1584,N_935);
nor U8658 (N_8658,N_567,N_3868);
nor U8659 (N_8659,N_3846,N_63);
and U8660 (N_8660,N_425,N_4722);
nand U8661 (N_8661,N_1827,N_3265);
or U8662 (N_8662,N_3901,N_813);
nor U8663 (N_8663,N_2892,N_3425);
nor U8664 (N_8664,N_4058,N_3859);
and U8665 (N_8665,N_164,N_2705);
nor U8666 (N_8666,N_3535,N_722);
nor U8667 (N_8667,N_1545,N_3555);
and U8668 (N_8668,N_3683,N_2310);
nand U8669 (N_8669,N_3080,N_2559);
nand U8670 (N_8670,N_919,N_2707);
or U8671 (N_8671,N_4971,N_3916);
and U8672 (N_8672,N_2598,N_4661);
or U8673 (N_8673,N_1698,N_3969);
xnor U8674 (N_8674,N_3940,N_3720);
nor U8675 (N_8675,N_814,N_1320);
or U8676 (N_8676,N_4492,N_894);
nor U8677 (N_8677,N_3983,N_82);
and U8678 (N_8678,N_3234,N_3861);
nor U8679 (N_8679,N_3673,N_1274);
nor U8680 (N_8680,N_1756,N_4429);
xor U8681 (N_8681,N_2478,N_4074);
nor U8682 (N_8682,N_4966,N_1721);
and U8683 (N_8683,N_3626,N_3561);
and U8684 (N_8684,N_2089,N_3268);
nand U8685 (N_8685,N_1624,N_337);
nand U8686 (N_8686,N_493,N_3839);
nand U8687 (N_8687,N_2590,N_3623);
nand U8688 (N_8688,N_2236,N_4800);
nand U8689 (N_8689,N_850,N_486);
or U8690 (N_8690,N_3363,N_845);
or U8691 (N_8691,N_521,N_4656);
or U8692 (N_8692,N_318,N_633);
or U8693 (N_8693,N_3407,N_253);
and U8694 (N_8694,N_1766,N_3271);
and U8695 (N_8695,N_470,N_1791);
and U8696 (N_8696,N_1626,N_154);
nor U8697 (N_8697,N_3230,N_4481);
nand U8698 (N_8698,N_1081,N_1186);
or U8699 (N_8699,N_960,N_3425);
xnor U8700 (N_8700,N_1746,N_4561);
and U8701 (N_8701,N_4943,N_4838);
nor U8702 (N_8702,N_4863,N_487);
or U8703 (N_8703,N_1419,N_4664);
and U8704 (N_8704,N_4659,N_205);
and U8705 (N_8705,N_3292,N_3818);
nor U8706 (N_8706,N_3490,N_1477);
or U8707 (N_8707,N_4717,N_3098);
or U8708 (N_8708,N_2114,N_2749);
nor U8709 (N_8709,N_1253,N_878);
nand U8710 (N_8710,N_3679,N_3429);
and U8711 (N_8711,N_2021,N_4583);
and U8712 (N_8712,N_4925,N_3406);
or U8713 (N_8713,N_4131,N_513);
or U8714 (N_8714,N_2155,N_1770);
or U8715 (N_8715,N_4802,N_426);
nand U8716 (N_8716,N_1427,N_4240);
or U8717 (N_8717,N_1485,N_2621);
and U8718 (N_8718,N_3760,N_1550);
xnor U8719 (N_8719,N_1266,N_369);
nor U8720 (N_8720,N_3408,N_4904);
nand U8721 (N_8721,N_1529,N_294);
nor U8722 (N_8722,N_2858,N_3752);
nand U8723 (N_8723,N_420,N_117);
and U8724 (N_8724,N_3065,N_4877);
and U8725 (N_8725,N_3456,N_332);
nor U8726 (N_8726,N_2936,N_2390);
nor U8727 (N_8727,N_4225,N_3253);
or U8728 (N_8728,N_4459,N_3358);
or U8729 (N_8729,N_2321,N_1067);
and U8730 (N_8730,N_4073,N_4614);
nor U8731 (N_8731,N_1316,N_3357);
nor U8732 (N_8732,N_4580,N_4468);
and U8733 (N_8733,N_4503,N_302);
nand U8734 (N_8734,N_3487,N_2912);
or U8735 (N_8735,N_2244,N_3265);
and U8736 (N_8736,N_148,N_4190);
and U8737 (N_8737,N_3462,N_1402);
xor U8738 (N_8738,N_2178,N_3742);
nand U8739 (N_8739,N_4450,N_430);
or U8740 (N_8740,N_3496,N_2742);
and U8741 (N_8741,N_841,N_4278);
nor U8742 (N_8742,N_43,N_3269);
nor U8743 (N_8743,N_4389,N_978);
nand U8744 (N_8744,N_4430,N_1696);
nor U8745 (N_8745,N_2228,N_1675);
nor U8746 (N_8746,N_2661,N_600);
nand U8747 (N_8747,N_3637,N_1150);
nand U8748 (N_8748,N_1237,N_314);
and U8749 (N_8749,N_4818,N_1102);
nand U8750 (N_8750,N_209,N_3660);
and U8751 (N_8751,N_1828,N_2175);
nor U8752 (N_8752,N_4021,N_2158);
or U8753 (N_8753,N_4176,N_52);
and U8754 (N_8754,N_2081,N_2228);
and U8755 (N_8755,N_3808,N_738);
nor U8756 (N_8756,N_4449,N_2153);
nand U8757 (N_8757,N_4918,N_1732);
or U8758 (N_8758,N_685,N_3299);
or U8759 (N_8759,N_2915,N_2610);
nor U8760 (N_8760,N_27,N_1995);
and U8761 (N_8761,N_314,N_4591);
nand U8762 (N_8762,N_1591,N_56);
nor U8763 (N_8763,N_2243,N_2555);
or U8764 (N_8764,N_3964,N_4891);
nand U8765 (N_8765,N_263,N_2638);
and U8766 (N_8766,N_2204,N_1490);
and U8767 (N_8767,N_4051,N_4987);
nand U8768 (N_8768,N_74,N_4431);
or U8769 (N_8769,N_4409,N_1772);
and U8770 (N_8770,N_1500,N_1584);
nor U8771 (N_8771,N_2422,N_4678);
nand U8772 (N_8772,N_1813,N_4635);
nand U8773 (N_8773,N_2863,N_1053);
nand U8774 (N_8774,N_2589,N_442);
nand U8775 (N_8775,N_4067,N_119);
and U8776 (N_8776,N_4776,N_91);
nor U8777 (N_8777,N_2964,N_404);
or U8778 (N_8778,N_277,N_2111);
nand U8779 (N_8779,N_4978,N_3941);
nand U8780 (N_8780,N_418,N_1529);
or U8781 (N_8781,N_110,N_1154);
nor U8782 (N_8782,N_2595,N_4114);
nand U8783 (N_8783,N_918,N_2830);
and U8784 (N_8784,N_1247,N_4740);
and U8785 (N_8785,N_1999,N_1797);
or U8786 (N_8786,N_4170,N_2533);
and U8787 (N_8787,N_3395,N_4719);
or U8788 (N_8788,N_4262,N_1380);
or U8789 (N_8789,N_4374,N_3142);
and U8790 (N_8790,N_2791,N_756);
or U8791 (N_8791,N_2569,N_4633);
or U8792 (N_8792,N_1735,N_2679);
nand U8793 (N_8793,N_4401,N_1900);
or U8794 (N_8794,N_1981,N_4184);
and U8795 (N_8795,N_2245,N_4707);
and U8796 (N_8796,N_1415,N_3475);
and U8797 (N_8797,N_283,N_1196);
nor U8798 (N_8798,N_568,N_4267);
nor U8799 (N_8799,N_378,N_4921);
nand U8800 (N_8800,N_388,N_4039);
nor U8801 (N_8801,N_2464,N_3010);
and U8802 (N_8802,N_3289,N_2800);
or U8803 (N_8803,N_1288,N_2081);
xor U8804 (N_8804,N_4379,N_1876);
or U8805 (N_8805,N_627,N_3250);
nor U8806 (N_8806,N_2862,N_109);
or U8807 (N_8807,N_4197,N_710);
and U8808 (N_8808,N_4034,N_2375);
nor U8809 (N_8809,N_3561,N_1579);
nand U8810 (N_8810,N_1347,N_2645);
or U8811 (N_8811,N_31,N_3272);
xnor U8812 (N_8812,N_3209,N_4900);
nand U8813 (N_8813,N_1967,N_2176);
and U8814 (N_8814,N_1575,N_932);
nor U8815 (N_8815,N_67,N_4638);
and U8816 (N_8816,N_1400,N_4744);
and U8817 (N_8817,N_3232,N_1109);
nand U8818 (N_8818,N_4409,N_4445);
nor U8819 (N_8819,N_4613,N_1160);
and U8820 (N_8820,N_955,N_1509);
and U8821 (N_8821,N_3675,N_2493);
or U8822 (N_8822,N_2264,N_3859);
nand U8823 (N_8823,N_2554,N_4504);
nor U8824 (N_8824,N_3804,N_3284);
nand U8825 (N_8825,N_2534,N_3537);
nor U8826 (N_8826,N_1660,N_3786);
or U8827 (N_8827,N_160,N_4140);
and U8828 (N_8828,N_3118,N_1495);
nor U8829 (N_8829,N_1134,N_2648);
and U8830 (N_8830,N_714,N_2606);
and U8831 (N_8831,N_1820,N_2563);
and U8832 (N_8832,N_3314,N_308);
or U8833 (N_8833,N_4588,N_533);
and U8834 (N_8834,N_3962,N_2022);
or U8835 (N_8835,N_4780,N_4442);
nor U8836 (N_8836,N_3755,N_2709);
nand U8837 (N_8837,N_3908,N_2279);
xor U8838 (N_8838,N_1537,N_2347);
nor U8839 (N_8839,N_2760,N_714);
and U8840 (N_8840,N_3562,N_4076);
and U8841 (N_8841,N_1620,N_3804);
or U8842 (N_8842,N_1374,N_3588);
or U8843 (N_8843,N_4943,N_2377);
and U8844 (N_8844,N_4225,N_1051);
xnor U8845 (N_8845,N_715,N_3023);
or U8846 (N_8846,N_2728,N_1899);
nor U8847 (N_8847,N_2920,N_3367);
or U8848 (N_8848,N_4474,N_469);
nand U8849 (N_8849,N_428,N_165);
and U8850 (N_8850,N_4319,N_17);
nor U8851 (N_8851,N_1099,N_4509);
nand U8852 (N_8852,N_1411,N_3546);
nor U8853 (N_8853,N_2163,N_502);
and U8854 (N_8854,N_860,N_2282);
and U8855 (N_8855,N_2956,N_4533);
xor U8856 (N_8856,N_564,N_2601);
and U8857 (N_8857,N_3750,N_3757);
nand U8858 (N_8858,N_3043,N_4853);
nor U8859 (N_8859,N_2084,N_4892);
or U8860 (N_8860,N_1994,N_1750);
nor U8861 (N_8861,N_1575,N_4133);
nor U8862 (N_8862,N_2893,N_3065);
nand U8863 (N_8863,N_3330,N_3580);
or U8864 (N_8864,N_726,N_1536);
or U8865 (N_8865,N_894,N_3739);
nor U8866 (N_8866,N_1166,N_4433);
or U8867 (N_8867,N_2982,N_4810);
and U8868 (N_8868,N_1033,N_1813);
nand U8869 (N_8869,N_801,N_971);
nor U8870 (N_8870,N_1596,N_3729);
and U8871 (N_8871,N_3704,N_1899);
or U8872 (N_8872,N_4957,N_2784);
nor U8873 (N_8873,N_934,N_2533);
and U8874 (N_8874,N_4998,N_4435);
and U8875 (N_8875,N_294,N_4416);
and U8876 (N_8876,N_530,N_1605);
xor U8877 (N_8877,N_1230,N_1210);
nand U8878 (N_8878,N_1528,N_4631);
or U8879 (N_8879,N_3259,N_3813);
nor U8880 (N_8880,N_4989,N_1012);
nand U8881 (N_8881,N_2315,N_2470);
and U8882 (N_8882,N_4118,N_1166);
nand U8883 (N_8883,N_257,N_4164);
or U8884 (N_8884,N_3946,N_1288);
nand U8885 (N_8885,N_4859,N_414);
nor U8886 (N_8886,N_3435,N_3461);
nand U8887 (N_8887,N_1223,N_3307);
nor U8888 (N_8888,N_1825,N_664);
or U8889 (N_8889,N_1887,N_1200);
and U8890 (N_8890,N_1129,N_3276);
nor U8891 (N_8891,N_961,N_2600);
xnor U8892 (N_8892,N_2742,N_3461);
and U8893 (N_8893,N_4547,N_4507);
and U8894 (N_8894,N_3883,N_2797);
nand U8895 (N_8895,N_2106,N_1995);
or U8896 (N_8896,N_2855,N_518);
nor U8897 (N_8897,N_3794,N_2720);
or U8898 (N_8898,N_4910,N_2047);
or U8899 (N_8899,N_1543,N_170);
nor U8900 (N_8900,N_658,N_222);
or U8901 (N_8901,N_1423,N_292);
and U8902 (N_8902,N_1914,N_2450);
and U8903 (N_8903,N_845,N_2764);
nand U8904 (N_8904,N_3528,N_2351);
nor U8905 (N_8905,N_476,N_3534);
nand U8906 (N_8906,N_3955,N_1795);
nand U8907 (N_8907,N_441,N_2147);
nand U8908 (N_8908,N_3166,N_552);
nor U8909 (N_8909,N_1230,N_1415);
and U8910 (N_8910,N_3363,N_4042);
nor U8911 (N_8911,N_3146,N_1729);
or U8912 (N_8912,N_965,N_3415);
and U8913 (N_8913,N_4840,N_3444);
nand U8914 (N_8914,N_4058,N_1280);
and U8915 (N_8915,N_4303,N_4937);
or U8916 (N_8916,N_3990,N_4072);
nand U8917 (N_8917,N_3734,N_2471);
nor U8918 (N_8918,N_1686,N_4313);
nand U8919 (N_8919,N_4467,N_4454);
nor U8920 (N_8920,N_1560,N_387);
or U8921 (N_8921,N_4843,N_3404);
nand U8922 (N_8922,N_1587,N_857);
and U8923 (N_8923,N_1738,N_65);
nor U8924 (N_8924,N_3504,N_3711);
xnor U8925 (N_8925,N_4013,N_3431);
nor U8926 (N_8926,N_4421,N_478);
nor U8927 (N_8927,N_1081,N_3169);
or U8928 (N_8928,N_4866,N_1071);
nand U8929 (N_8929,N_997,N_3312);
nand U8930 (N_8930,N_323,N_761);
nor U8931 (N_8931,N_4016,N_3537);
or U8932 (N_8932,N_4325,N_3089);
xor U8933 (N_8933,N_670,N_206);
nor U8934 (N_8934,N_4260,N_2062);
or U8935 (N_8935,N_4398,N_329);
and U8936 (N_8936,N_970,N_2309);
or U8937 (N_8937,N_1380,N_3260);
nand U8938 (N_8938,N_2486,N_1739);
and U8939 (N_8939,N_2468,N_650);
nor U8940 (N_8940,N_732,N_623);
nand U8941 (N_8941,N_2315,N_2532);
xor U8942 (N_8942,N_3941,N_514);
nand U8943 (N_8943,N_1356,N_4082);
nand U8944 (N_8944,N_1022,N_2844);
and U8945 (N_8945,N_3907,N_1176);
nand U8946 (N_8946,N_3245,N_3957);
nand U8947 (N_8947,N_4098,N_1778);
nand U8948 (N_8948,N_473,N_4580);
nand U8949 (N_8949,N_2006,N_1228);
and U8950 (N_8950,N_3895,N_1832);
or U8951 (N_8951,N_2977,N_625);
or U8952 (N_8952,N_910,N_3832);
nor U8953 (N_8953,N_1697,N_4908);
nor U8954 (N_8954,N_3499,N_2324);
or U8955 (N_8955,N_2508,N_280);
nor U8956 (N_8956,N_2798,N_4763);
nand U8957 (N_8957,N_2700,N_1797);
and U8958 (N_8958,N_1273,N_2269);
and U8959 (N_8959,N_1317,N_4910);
and U8960 (N_8960,N_1630,N_4414);
nor U8961 (N_8961,N_1955,N_2173);
nand U8962 (N_8962,N_929,N_879);
or U8963 (N_8963,N_3090,N_1986);
nand U8964 (N_8964,N_1811,N_1955);
nor U8965 (N_8965,N_2699,N_615);
nand U8966 (N_8966,N_3395,N_3341);
and U8967 (N_8967,N_2645,N_2779);
nand U8968 (N_8968,N_4174,N_3312);
nor U8969 (N_8969,N_2053,N_3665);
xor U8970 (N_8970,N_206,N_4345);
nor U8971 (N_8971,N_1752,N_1359);
or U8972 (N_8972,N_1400,N_1579);
or U8973 (N_8973,N_269,N_1959);
or U8974 (N_8974,N_2131,N_4464);
nor U8975 (N_8975,N_4440,N_4214);
nor U8976 (N_8976,N_4082,N_4286);
nand U8977 (N_8977,N_2217,N_1505);
xnor U8978 (N_8978,N_2407,N_4479);
nand U8979 (N_8979,N_4939,N_1349);
and U8980 (N_8980,N_1517,N_1874);
nand U8981 (N_8981,N_1368,N_4157);
nor U8982 (N_8982,N_4594,N_1348);
nand U8983 (N_8983,N_392,N_4470);
or U8984 (N_8984,N_2381,N_2181);
nand U8985 (N_8985,N_2213,N_1263);
nand U8986 (N_8986,N_4178,N_232);
and U8987 (N_8987,N_2180,N_4858);
or U8988 (N_8988,N_2364,N_1632);
nor U8989 (N_8989,N_1376,N_115);
xnor U8990 (N_8990,N_241,N_956);
or U8991 (N_8991,N_897,N_3881);
and U8992 (N_8992,N_4739,N_1025);
or U8993 (N_8993,N_1235,N_710);
or U8994 (N_8994,N_508,N_2879);
and U8995 (N_8995,N_916,N_88);
and U8996 (N_8996,N_2858,N_4606);
nor U8997 (N_8997,N_198,N_3992);
nor U8998 (N_8998,N_3876,N_3777);
nand U8999 (N_8999,N_3178,N_3336);
nand U9000 (N_9000,N_4357,N_2785);
and U9001 (N_9001,N_865,N_1182);
or U9002 (N_9002,N_4732,N_4171);
or U9003 (N_9003,N_1988,N_2291);
nand U9004 (N_9004,N_467,N_1055);
and U9005 (N_9005,N_1601,N_4274);
or U9006 (N_9006,N_1333,N_2932);
nor U9007 (N_9007,N_3375,N_648);
and U9008 (N_9008,N_4576,N_4316);
and U9009 (N_9009,N_121,N_4990);
nor U9010 (N_9010,N_333,N_2969);
or U9011 (N_9011,N_4466,N_2626);
or U9012 (N_9012,N_4910,N_4781);
nor U9013 (N_9013,N_1080,N_4645);
nand U9014 (N_9014,N_4394,N_2754);
nand U9015 (N_9015,N_4029,N_451);
nand U9016 (N_9016,N_3603,N_4903);
nand U9017 (N_9017,N_3153,N_1226);
xnor U9018 (N_9018,N_3931,N_248);
nand U9019 (N_9019,N_336,N_4594);
nor U9020 (N_9020,N_614,N_4578);
nand U9021 (N_9021,N_1498,N_2528);
and U9022 (N_9022,N_3582,N_875);
nand U9023 (N_9023,N_520,N_3093);
and U9024 (N_9024,N_4008,N_634);
or U9025 (N_9025,N_1065,N_2662);
or U9026 (N_9026,N_4660,N_3373);
and U9027 (N_9027,N_3136,N_4553);
nand U9028 (N_9028,N_4831,N_1781);
nor U9029 (N_9029,N_2472,N_3887);
nor U9030 (N_9030,N_2274,N_4485);
nand U9031 (N_9031,N_4823,N_7);
or U9032 (N_9032,N_1608,N_2222);
nor U9033 (N_9033,N_2438,N_642);
or U9034 (N_9034,N_666,N_4604);
or U9035 (N_9035,N_1632,N_477);
and U9036 (N_9036,N_2726,N_733);
nand U9037 (N_9037,N_3563,N_2639);
and U9038 (N_9038,N_1389,N_1921);
and U9039 (N_9039,N_2221,N_1857);
or U9040 (N_9040,N_2261,N_334);
and U9041 (N_9041,N_2734,N_1703);
and U9042 (N_9042,N_1239,N_4769);
nand U9043 (N_9043,N_520,N_1092);
nor U9044 (N_9044,N_4707,N_4822);
or U9045 (N_9045,N_2831,N_4696);
xnor U9046 (N_9046,N_3714,N_4657);
or U9047 (N_9047,N_3843,N_4884);
nand U9048 (N_9048,N_4003,N_2879);
nand U9049 (N_9049,N_4993,N_2459);
nand U9050 (N_9050,N_4658,N_1270);
xor U9051 (N_9051,N_3765,N_231);
nand U9052 (N_9052,N_2177,N_4827);
nand U9053 (N_9053,N_2334,N_4086);
and U9054 (N_9054,N_4872,N_4154);
nand U9055 (N_9055,N_550,N_1089);
nand U9056 (N_9056,N_3978,N_2537);
nand U9057 (N_9057,N_3382,N_1246);
or U9058 (N_9058,N_3434,N_3895);
xor U9059 (N_9059,N_415,N_4486);
nor U9060 (N_9060,N_4177,N_4335);
nor U9061 (N_9061,N_2348,N_759);
nor U9062 (N_9062,N_815,N_2562);
nor U9063 (N_9063,N_3562,N_258);
nor U9064 (N_9064,N_3765,N_4925);
or U9065 (N_9065,N_17,N_512);
nor U9066 (N_9066,N_1222,N_1919);
nor U9067 (N_9067,N_1979,N_1330);
nand U9068 (N_9068,N_914,N_1475);
nor U9069 (N_9069,N_3073,N_1687);
nand U9070 (N_9070,N_1700,N_168);
or U9071 (N_9071,N_884,N_2351);
and U9072 (N_9072,N_647,N_941);
and U9073 (N_9073,N_561,N_1656);
or U9074 (N_9074,N_3334,N_457);
or U9075 (N_9075,N_1153,N_4044);
or U9076 (N_9076,N_1764,N_2300);
nor U9077 (N_9077,N_906,N_1930);
nand U9078 (N_9078,N_1901,N_2251);
nor U9079 (N_9079,N_359,N_2522);
or U9080 (N_9080,N_4168,N_3105);
and U9081 (N_9081,N_2227,N_850);
nand U9082 (N_9082,N_4606,N_4724);
or U9083 (N_9083,N_1746,N_2683);
nor U9084 (N_9084,N_245,N_4167);
nor U9085 (N_9085,N_3702,N_949);
nor U9086 (N_9086,N_3950,N_4105);
nand U9087 (N_9087,N_4244,N_3516);
or U9088 (N_9088,N_728,N_1187);
or U9089 (N_9089,N_3427,N_449);
and U9090 (N_9090,N_1094,N_871);
and U9091 (N_9091,N_1327,N_3033);
nand U9092 (N_9092,N_2085,N_4946);
or U9093 (N_9093,N_2485,N_1850);
nor U9094 (N_9094,N_2231,N_4796);
and U9095 (N_9095,N_943,N_3970);
nor U9096 (N_9096,N_2073,N_4955);
nor U9097 (N_9097,N_4663,N_3671);
nand U9098 (N_9098,N_3400,N_2050);
nand U9099 (N_9099,N_228,N_4812);
nor U9100 (N_9100,N_1012,N_2308);
nor U9101 (N_9101,N_1307,N_2583);
or U9102 (N_9102,N_4080,N_23);
and U9103 (N_9103,N_1098,N_1213);
xnor U9104 (N_9104,N_47,N_560);
and U9105 (N_9105,N_4524,N_1448);
nor U9106 (N_9106,N_1059,N_3977);
or U9107 (N_9107,N_1523,N_4571);
and U9108 (N_9108,N_2496,N_3185);
nor U9109 (N_9109,N_3921,N_1834);
xnor U9110 (N_9110,N_1760,N_491);
or U9111 (N_9111,N_3038,N_741);
nor U9112 (N_9112,N_3368,N_2921);
or U9113 (N_9113,N_3023,N_623);
nor U9114 (N_9114,N_3125,N_3186);
nor U9115 (N_9115,N_4579,N_2209);
nand U9116 (N_9116,N_2268,N_2331);
and U9117 (N_9117,N_3015,N_1266);
nand U9118 (N_9118,N_904,N_2514);
nor U9119 (N_9119,N_1498,N_650);
or U9120 (N_9120,N_1211,N_3896);
nand U9121 (N_9121,N_1681,N_2476);
and U9122 (N_9122,N_341,N_2220);
and U9123 (N_9123,N_1438,N_2035);
or U9124 (N_9124,N_371,N_4001);
nand U9125 (N_9125,N_442,N_1096);
nor U9126 (N_9126,N_1506,N_2204);
or U9127 (N_9127,N_4949,N_500);
nand U9128 (N_9128,N_2510,N_2012);
and U9129 (N_9129,N_4934,N_2673);
and U9130 (N_9130,N_2709,N_4717);
or U9131 (N_9131,N_4075,N_398);
or U9132 (N_9132,N_391,N_2450);
nand U9133 (N_9133,N_3401,N_2325);
and U9134 (N_9134,N_983,N_4925);
and U9135 (N_9135,N_1474,N_2159);
nand U9136 (N_9136,N_1426,N_879);
and U9137 (N_9137,N_2539,N_294);
nor U9138 (N_9138,N_3864,N_3792);
and U9139 (N_9139,N_4630,N_2386);
or U9140 (N_9140,N_563,N_402);
nor U9141 (N_9141,N_443,N_1924);
nor U9142 (N_9142,N_2266,N_3842);
or U9143 (N_9143,N_2154,N_229);
and U9144 (N_9144,N_4677,N_3000);
or U9145 (N_9145,N_3496,N_3299);
xor U9146 (N_9146,N_2219,N_3117);
and U9147 (N_9147,N_2842,N_4895);
and U9148 (N_9148,N_3560,N_867);
nand U9149 (N_9149,N_4164,N_723);
or U9150 (N_9150,N_4181,N_4256);
nor U9151 (N_9151,N_3023,N_3905);
or U9152 (N_9152,N_717,N_618);
nor U9153 (N_9153,N_1846,N_676);
nor U9154 (N_9154,N_2959,N_20);
nand U9155 (N_9155,N_4257,N_4977);
and U9156 (N_9156,N_3383,N_940);
nand U9157 (N_9157,N_3555,N_3855);
nand U9158 (N_9158,N_3785,N_4866);
xnor U9159 (N_9159,N_1508,N_2220);
nor U9160 (N_9160,N_1171,N_285);
or U9161 (N_9161,N_3274,N_128);
or U9162 (N_9162,N_4012,N_2610);
or U9163 (N_9163,N_3077,N_4527);
and U9164 (N_9164,N_1285,N_2190);
or U9165 (N_9165,N_4184,N_357);
or U9166 (N_9166,N_530,N_4318);
or U9167 (N_9167,N_1784,N_4564);
or U9168 (N_9168,N_781,N_50);
nor U9169 (N_9169,N_313,N_4935);
nand U9170 (N_9170,N_3308,N_3800);
nor U9171 (N_9171,N_1754,N_547);
nor U9172 (N_9172,N_2387,N_3085);
or U9173 (N_9173,N_2993,N_3176);
nor U9174 (N_9174,N_3912,N_4441);
nor U9175 (N_9175,N_3398,N_4261);
nand U9176 (N_9176,N_3770,N_2398);
nand U9177 (N_9177,N_2438,N_234);
nor U9178 (N_9178,N_4003,N_2099);
nor U9179 (N_9179,N_1852,N_1630);
nand U9180 (N_9180,N_4882,N_253);
and U9181 (N_9181,N_1763,N_1628);
and U9182 (N_9182,N_1921,N_38);
nand U9183 (N_9183,N_4317,N_2017);
nand U9184 (N_9184,N_2249,N_4610);
nand U9185 (N_9185,N_4643,N_4809);
nor U9186 (N_9186,N_4311,N_819);
or U9187 (N_9187,N_875,N_3383);
and U9188 (N_9188,N_1055,N_2479);
or U9189 (N_9189,N_3388,N_2282);
nand U9190 (N_9190,N_3774,N_4674);
nor U9191 (N_9191,N_3448,N_4209);
or U9192 (N_9192,N_4290,N_4026);
nor U9193 (N_9193,N_1325,N_2749);
nand U9194 (N_9194,N_4457,N_1817);
nand U9195 (N_9195,N_4728,N_2482);
or U9196 (N_9196,N_740,N_2759);
or U9197 (N_9197,N_3347,N_1100);
and U9198 (N_9198,N_2151,N_3189);
nor U9199 (N_9199,N_3147,N_4880);
and U9200 (N_9200,N_4155,N_2416);
nand U9201 (N_9201,N_2552,N_3822);
and U9202 (N_9202,N_3796,N_547);
or U9203 (N_9203,N_2764,N_40);
nor U9204 (N_9204,N_1789,N_2496);
and U9205 (N_9205,N_1221,N_2250);
nor U9206 (N_9206,N_734,N_865);
nand U9207 (N_9207,N_4059,N_3867);
nand U9208 (N_9208,N_4531,N_3791);
nand U9209 (N_9209,N_3470,N_1413);
nor U9210 (N_9210,N_2267,N_992);
or U9211 (N_9211,N_3437,N_3134);
nand U9212 (N_9212,N_512,N_1508);
nand U9213 (N_9213,N_319,N_3002);
and U9214 (N_9214,N_2472,N_209);
nand U9215 (N_9215,N_1948,N_1236);
nand U9216 (N_9216,N_883,N_2346);
nand U9217 (N_9217,N_1609,N_1391);
or U9218 (N_9218,N_251,N_4509);
nand U9219 (N_9219,N_647,N_3872);
nand U9220 (N_9220,N_276,N_4646);
nor U9221 (N_9221,N_4990,N_3625);
or U9222 (N_9222,N_72,N_2678);
or U9223 (N_9223,N_3788,N_4078);
nand U9224 (N_9224,N_3567,N_2626);
nand U9225 (N_9225,N_2048,N_1909);
nor U9226 (N_9226,N_3793,N_3165);
or U9227 (N_9227,N_3923,N_4118);
and U9228 (N_9228,N_4822,N_353);
nor U9229 (N_9229,N_168,N_1147);
and U9230 (N_9230,N_4914,N_125);
nand U9231 (N_9231,N_1850,N_4817);
or U9232 (N_9232,N_575,N_3228);
or U9233 (N_9233,N_4515,N_1243);
nand U9234 (N_9234,N_1660,N_3313);
or U9235 (N_9235,N_3861,N_93);
nor U9236 (N_9236,N_3595,N_2119);
or U9237 (N_9237,N_1838,N_983);
or U9238 (N_9238,N_3251,N_1703);
and U9239 (N_9239,N_2179,N_1360);
or U9240 (N_9240,N_2269,N_1077);
nand U9241 (N_9241,N_967,N_2263);
nor U9242 (N_9242,N_4382,N_1365);
or U9243 (N_9243,N_4124,N_1088);
and U9244 (N_9244,N_2886,N_2497);
nand U9245 (N_9245,N_1136,N_1225);
and U9246 (N_9246,N_1627,N_1013);
and U9247 (N_9247,N_3704,N_2288);
nor U9248 (N_9248,N_3658,N_543);
nor U9249 (N_9249,N_4354,N_2169);
nor U9250 (N_9250,N_2023,N_3963);
xnor U9251 (N_9251,N_3316,N_64);
or U9252 (N_9252,N_1610,N_436);
and U9253 (N_9253,N_2672,N_4535);
and U9254 (N_9254,N_757,N_1955);
nand U9255 (N_9255,N_1914,N_4137);
nand U9256 (N_9256,N_340,N_1931);
xnor U9257 (N_9257,N_4069,N_1150);
and U9258 (N_9258,N_1200,N_1137);
and U9259 (N_9259,N_3551,N_1318);
nand U9260 (N_9260,N_3664,N_4481);
or U9261 (N_9261,N_147,N_1273);
xnor U9262 (N_9262,N_4437,N_3475);
and U9263 (N_9263,N_1411,N_3622);
nor U9264 (N_9264,N_1579,N_4858);
and U9265 (N_9265,N_1791,N_3010);
nor U9266 (N_9266,N_3183,N_3513);
or U9267 (N_9267,N_2571,N_927);
nor U9268 (N_9268,N_4688,N_762);
and U9269 (N_9269,N_1006,N_466);
nand U9270 (N_9270,N_3709,N_4493);
and U9271 (N_9271,N_1698,N_2636);
or U9272 (N_9272,N_282,N_4641);
and U9273 (N_9273,N_3711,N_3406);
nor U9274 (N_9274,N_2806,N_4279);
or U9275 (N_9275,N_2986,N_1578);
nor U9276 (N_9276,N_520,N_1127);
and U9277 (N_9277,N_550,N_3995);
nand U9278 (N_9278,N_3042,N_996);
or U9279 (N_9279,N_1142,N_4280);
or U9280 (N_9280,N_4752,N_279);
nor U9281 (N_9281,N_1814,N_3733);
nand U9282 (N_9282,N_3756,N_3935);
or U9283 (N_9283,N_339,N_2616);
nor U9284 (N_9284,N_3911,N_1727);
and U9285 (N_9285,N_4379,N_4195);
nand U9286 (N_9286,N_123,N_1541);
and U9287 (N_9287,N_1991,N_4357);
nor U9288 (N_9288,N_4168,N_2946);
nand U9289 (N_9289,N_1179,N_15);
nor U9290 (N_9290,N_1404,N_4069);
nor U9291 (N_9291,N_3625,N_2590);
nand U9292 (N_9292,N_3612,N_1609);
and U9293 (N_9293,N_809,N_4243);
nand U9294 (N_9294,N_4434,N_2367);
nand U9295 (N_9295,N_145,N_1320);
or U9296 (N_9296,N_1147,N_209);
or U9297 (N_9297,N_4778,N_2804);
nor U9298 (N_9298,N_1248,N_1870);
nand U9299 (N_9299,N_3889,N_870);
nand U9300 (N_9300,N_218,N_3438);
and U9301 (N_9301,N_3949,N_1032);
or U9302 (N_9302,N_1693,N_3410);
nand U9303 (N_9303,N_794,N_2458);
nor U9304 (N_9304,N_4319,N_2620);
and U9305 (N_9305,N_1996,N_2901);
nand U9306 (N_9306,N_2197,N_3210);
nand U9307 (N_9307,N_1849,N_1259);
or U9308 (N_9308,N_4032,N_2316);
nor U9309 (N_9309,N_2835,N_738);
or U9310 (N_9310,N_2819,N_294);
or U9311 (N_9311,N_3926,N_2776);
nor U9312 (N_9312,N_635,N_2518);
nor U9313 (N_9313,N_4186,N_370);
nor U9314 (N_9314,N_1973,N_4781);
nand U9315 (N_9315,N_4107,N_2045);
and U9316 (N_9316,N_570,N_922);
nand U9317 (N_9317,N_4600,N_1060);
nand U9318 (N_9318,N_4065,N_229);
nor U9319 (N_9319,N_4933,N_4397);
and U9320 (N_9320,N_3822,N_4056);
or U9321 (N_9321,N_2041,N_605);
and U9322 (N_9322,N_4445,N_490);
nor U9323 (N_9323,N_4429,N_2733);
or U9324 (N_9324,N_3121,N_655);
and U9325 (N_9325,N_1011,N_4068);
or U9326 (N_9326,N_3135,N_2314);
nor U9327 (N_9327,N_4954,N_983);
and U9328 (N_9328,N_227,N_1755);
nor U9329 (N_9329,N_2743,N_192);
and U9330 (N_9330,N_4561,N_3809);
or U9331 (N_9331,N_253,N_2112);
nand U9332 (N_9332,N_1029,N_888);
nand U9333 (N_9333,N_1549,N_95);
or U9334 (N_9334,N_883,N_2662);
nand U9335 (N_9335,N_4666,N_4453);
nand U9336 (N_9336,N_4595,N_2060);
and U9337 (N_9337,N_654,N_401);
or U9338 (N_9338,N_2588,N_2848);
nor U9339 (N_9339,N_3888,N_1849);
or U9340 (N_9340,N_3559,N_275);
nor U9341 (N_9341,N_2881,N_1411);
nand U9342 (N_9342,N_2709,N_1567);
and U9343 (N_9343,N_95,N_2519);
nor U9344 (N_9344,N_898,N_6);
or U9345 (N_9345,N_2664,N_1004);
nand U9346 (N_9346,N_3621,N_1552);
nor U9347 (N_9347,N_3168,N_1210);
nand U9348 (N_9348,N_2977,N_1623);
nand U9349 (N_9349,N_2834,N_814);
and U9350 (N_9350,N_4742,N_3189);
and U9351 (N_9351,N_1022,N_418);
and U9352 (N_9352,N_1093,N_1336);
nand U9353 (N_9353,N_3850,N_3082);
nand U9354 (N_9354,N_1426,N_1906);
and U9355 (N_9355,N_2816,N_1879);
or U9356 (N_9356,N_1689,N_3444);
xnor U9357 (N_9357,N_955,N_1744);
nand U9358 (N_9358,N_1559,N_647);
nor U9359 (N_9359,N_1039,N_2933);
or U9360 (N_9360,N_1142,N_4798);
or U9361 (N_9361,N_1761,N_2457);
or U9362 (N_9362,N_3935,N_195);
nand U9363 (N_9363,N_3259,N_4238);
and U9364 (N_9364,N_1744,N_3095);
or U9365 (N_9365,N_790,N_1584);
or U9366 (N_9366,N_927,N_4565);
or U9367 (N_9367,N_534,N_2893);
nand U9368 (N_9368,N_3800,N_2953);
nor U9369 (N_9369,N_1249,N_2747);
or U9370 (N_9370,N_1270,N_2405);
nor U9371 (N_9371,N_2229,N_2038);
or U9372 (N_9372,N_802,N_4242);
nand U9373 (N_9373,N_1058,N_908);
or U9374 (N_9374,N_4509,N_2695);
nor U9375 (N_9375,N_1558,N_1693);
nor U9376 (N_9376,N_1919,N_2717);
and U9377 (N_9377,N_1651,N_1419);
or U9378 (N_9378,N_3565,N_2376);
and U9379 (N_9379,N_3423,N_3539);
nand U9380 (N_9380,N_3226,N_2330);
or U9381 (N_9381,N_599,N_949);
nor U9382 (N_9382,N_1818,N_3025);
and U9383 (N_9383,N_1008,N_2680);
nand U9384 (N_9384,N_2288,N_3827);
or U9385 (N_9385,N_3856,N_276);
or U9386 (N_9386,N_2560,N_1127);
nand U9387 (N_9387,N_4295,N_4951);
or U9388 (N_9388,N_1350,N_74);
or U9389 (N_9389,N_3500,N_504);
nand U9390 (N_9390,N_1174,N_36);
and U9391 (N_9391,N_4421,N_2899);
or U9392 (N_9392,N_740,N_3600);
nor U9393 (N_9393,N_2325,N_410);
nor U9394 (N_9394,N_2167,N_1354);
or U9395 (N_9395,N_2078,N_4856);
or U9396 (N_9396,N_2104,N_34);
nor U9397 (N_9397,N_4033,N_138);
xor U9398 (N_9398,N_1549,N_3707);
nand U9399 (N_9399,N_4442,N_2377);
nor U9400 (N_9400,N_331,N_1338);
nor U9401 (N_9401,N_1542,N_486);
nor U9402 (N_9402,N_4568,N_689);
nor U9403 (N_9403,N_553,N_3655);
and U9404 (N_9404,N_3125,N_1087);
or U9405 (N_9405,N_172,N_791);
or U9406 (N_9406,N_4876,N_4003);
nor U9407 (N_9407,N_446,N_2572);
xor U9408 (N_9408,N_2255,N_1558);
nor U9409 (N_9409,N_174,N_2513);
nand U9410 (N_9410,N_3272,N_3231);
nand U9411 (N_9411,N_1208,N_2080);
or U9412 (N_9412,N_2399,N_514);
nand U9413 (N_9413,N_1242,N_2147);
or U9414 (N_9414,N_1422,N_1548);
and U9415 (N_9415,N_675,N_3398);
nand U9416 (N_9416,N_1801,N_1312);
and U9417 (N_9417,N_248,N_1173);
nor U9418 (N_9418,N_2987,N_4435);
nand U9419 (N_9419,N_1244,N_3369);
nor U9420 (N_9420,N_4520,N_2156);
xor U9421 (N_9421,N_2230,N_2517);
xor U9422 (N_9422,N_4961,N_3363);
xnor U9423 (N_9423,N_395,N_649);
or U9424 (N_9424,N_1525,N_741);
or U9425 (N_9425,N_2896,N_4634);
or U9426 (N_9426,N_1542,N_4335);
nand U9427 (N_9427,N_339,N_2661);
and U9428 (N_9428,N_3881,N_3654);
and U9429 (N_9429,N_3233,N_672);
and U9430 (N_9430,N_2186,N_1548);
or U9431 (N_9431,N_228,N_1652);
nand U9432 (N_9432,N_1483,N_374);
and U9433 (N_9433,N_1801,N_1123);
nor U9434 (N_9434,N_3143,N_3694);
xnor U9435 (N_9435,N_507,N_4098);
nand U9436 (N_9436,N_2007,N_325);
and U9437 (N_9437,N_2385,N_1178);
or U9438 (N_9438,N_829,N_2374);
nor U9439 (N_9439,N_2168,N_1227);
nor U9440 (N_9440,N_1728,N_2375);
nor U9441 (N_9441,N_4560,N_2949);
nor U9442 (N_9442,N_635,N_3750);
or U9443 (N_9443,N_2844,N_4081);
or U9444 (N_9444,N_2778,N_1669);
or U9445 (N_9445,N_98,N_3024);
xor U9446 (N_9446,N_164,N_425);
nor U9447 (N_9447,N_3791,N_20);
or U9448 (N_9448,N_3266,N_932);
nand U9449 (N_9449,N_1108,N_4846);
and U9450 (N_9450,N_1924,N_3021);
nor U9451 (N_9451,N_4252,N_4463);
and U9452 (N_9452,N_1625,N_348);
and U9453 (N_9453,N_4538,N_212);
nand U9454 (N_9454,N_2523,N_1652);
or U9455 (N_9455,N_620,N_3062);
nor U9456 (N_9456,N_851,N_3694);
and U9457 (N_9457,N_3790,N_3445);
nand U9458 (N_9458,N_530,N_3141);
nand U9459 (N_9459,N_4940,N_23);
or U9460 (N_9460,N_4677,N_2095);
or U9461 (N_9461,N_2518,N_4994);
nor U9462 (N_9462,N_15,N_3789);
nand U9463 (N_9463,N_4722,N_2887);
nor U9464 (N_9464,N_3559,N_60);
nand U9465 (N_9465,N_476,N_156);
nor U9466 (N_9466,N_3772,N_3375);
or U9467 (N_9467,N_1239,N_399);
nor U9468 (N_9468,N_3056,N_3169);
or U9469 (N_9469,N_1987,N_3643);
nand U9470 (N_9470,N_4484,N_2975);
or U9471 (N_9471,N_553,N_4033);
nor U9472 (N_9472,N_3375,N_2004);
or U9473 (N_9473,N_2978,N_2815);
and U9474 (N_9474,N_4746,N_3423);
nor U9475 (N_9475,N_4624,N_4109);
nor U9476 (N_9476,N_4405,N_4052);
nand U9477 (N_9477,N_253,N_174);
or U9478 (N_9478,N_4783,N_2152);
or U9479 (N_9479,N_3896,N_3946);
or U9480 (N_9480,N_1662,N_2577);
nor U9481 (N_9481,N_1141,N_4225);
nand U9482 (N_9482,N_2248,N_3156);
or U9483 (N_9483,N_392,N_4494);
nand U9484 (N_9484,N_1487,N_6);
nand U9485 (N_9485,N_1000,N_3719);
nor U9486 (N_9486,N_2910,N_1144);
nand U9487 (N_9487,N_3888,N_1228);
or U9488 (N_9488,N_1493,N_3135);
or U9489 (N_9489,N_3463,N_4893);
or U9490 (N_9490,N_208,N_139);
or U9491 (N_9491,N_1977,N_2528);
and U9492 (N_9492,N_527,N_3091);
nand U9493 (N_9493,N_1710,N_1753);
or U9494 (N_9494,N_2005,N_2101);
nor U9495 (N_9495,N_1951,N_4922);
nor U9496 (N_9496,N_4970,N_3402);
nor U9497 (N_9497,N_1886,N_3790);
or U9498 (N_9498,N_432,N_1420);
or U9499 (N_9499,N_4068,N_2873);
nand U9500 (N_9500,N_157,N_1524);
nor U9501 (N_9501,N_669,N_4169);
and U9502 (N_9502,N_1666,N_4898);
nor U9503 (N_9503,N_3698,N_2417);
nor U9504 (N_9504,N_2055,N_1087);
and U9505 (N_9505,N_419,N_3153);
or U9506 (N_9506,N_3983,N_4536);
nand U9507 (N_9507,N_67,N_2538);
nor U9508 (N_9508,N_1330,N_4759);
nor U9509 (N_9509,N_1287,N_441);
and U9510 (N_9510,N_4467,N_3714);
nand U9511 (N_9511,N_2502,N_2241);
nand U9512 (N_9512,N_202,N_2011);
nand U9513 (N_9513,N_1244,N_1195);
or U9514 (N_9514,N_452,N_572);
nand U9515 (N_9515,N_4714,N_163);
or U9516 (N_9516,N_3099,N_4855);
nand U9517 (N_9517,N_40,N_2880);
or U9518 (N_9518,N_715,N_2021);
or U9519 (N_9519,N_38,N_297);
nor U9520 (N_9520,N_3569,N_3164);
nand U9521 (N_9521,N_3931,N_1522);
or U9522 (N_9522,N_3031,N_2242);
and U9523 (N_9523,N_4804,N_3478);
nand U9524 (N_9524,N_3912,N_598);
and U9525 (N_9525,N_438,N_4598);
nand U9526 (N_9526,N_662,N_3988);
nand U9527 (N_9527,N_2684,N_3490);
nor U9528 (N_9528,N_2791,N_930);
and U9529 (N_9529,N_2674,N_393);
and U9530 (N_9530,N_2746,N_1276);
nor U9531 (N_9531,N_977,N_3114);
and U9532 (N_9532,N_4524,N_1895);
or U9533 (N_9533,N_3648,N_3709);
and U9534 (N_9534,N_693,N_2458);
and U9535 (N_9535,N_3591,N_4749);
nand U9536 (N_9536,N_3434,N_4921);
nor U9537 (N_9537,N_4122,N_98);
nor U9538 (N_9538,N_4574,N_1650);
nand U9539 (N_9539,N_4152,N_3662);
nor U9540 (N_9540,N_4443,N_1924);
or U9541 (N_9541,N_4543,N_797);
or U9542 (N_9542,N_954,N_3452);
and U9543 (N_9543,N_3109,N_4230);
or U9544 (N_9544,N_4658,N_4985);
and U9545 (N_9545,N_1805,N_4972);
nand U9546 (N_9546,N_3730,N_1841);
and U9547 (N_9547,N_2226,N_4918);
nor U9548 (N_9548,N_3087,N_3688);
nor U9549 (N_9549,N_3262,N_4482);
nand U9550 (N_9550,N_4648,N_3462);
and U9551 (N_9551,N_2952,N_521);
nor U9552 (N_9552,N_4802,N_4301);
or U9553 (N_9553,N_4728,N_3986);
nand U9554 (N_9554,N_1996,N_4154);
and U9555 (N_9555,N_1573,N_1922);
or U9556 (N_9556,N_638,N_3337);
nor U9557 (N_9557,N_4837,N_4595);
or U9558 (N_9558,N_2677,N_1029);
nand U9559 (N_9559,N_2362,N_3021);
and U9560 (N_9560,N_2257,N_2171);
and U9561 (N_9561,N_2417,N_1447);
nor U9562 (N_9562,N_1103,N_4126);
and U9563 (N_9563,N_1261,N_3097);
nor U9564 (N_9564,N_4180,N_1249);
and U9565 (N_9565,N_4653,N_424);
and U9566 (N_9566,N_4594,N_3366);
or U9567 (N_9567,N_2791,N_2580);
nand U9568 (N_9568,N_4347,N_794);
and U9569 (N_9569,N_2699,N_4568);
and U9570 (N_9570,N_2428,N_2947);
or U9571 (N_9571,N_1179,N_4730);
xor U9572 (N_9572,N_475,N_2739);
or U9573 (N_9573,N_2735,N_409);
or U9574 (N_9574,N_56,N_3168);
nor U9575 (N_9575,N_3754,N_1377);
xor U9576 (N_9576,N_2900,N_127);
nand U9577 (N_9577,N_903,N_3139);
xnor U9578 (N_9578,N_4742,N_3867);
nand U9579 (N_9579,N_2380,N_3590);
nor U9580 (N_9580,N_363,N_3648);
nand U9581 (N_9581,N_2362,N_1871);
nor U9582 (N_9582,N_4481,N_1796);
or U9583 (N_9583,N_3333,N_1601);
or U9584 (N_9584,N_2353,N_4103);
nor U9585 (N_9585,N_4079,N_829);
and U9586 (N_9586,N_1594,N_3674);
and U9587 (N_9587,N_2309,N_2359);
and U9588 (N_9588,N_2000,N_2981);
nor U9589 (N_9589,N_4338,N_2529);
nand U9590 (N_9590,N_1773,N_163);
nand U9591 (N_9591,N_652,N_648);
nand U9592 (N_9592,N_1922,N_3647);
nor U9593 (N_9593,N_1189,N_2947);
and U9594 (N_9594,N_4981,N_4622);
and U9595 (N_9595,N_1964,N_1368);
nor U9596 (N_9596,N_1968,N_2020);
and U9597 (N_9597,N_1761,N_1799);
or U9598 (N_9598,N_110,N_1532);
and U9599 (N_9599,N_3741,N_3141);
or U9600 (N_9600,N_638,N_4097);
and U9601 (N_9601,N_1060,N_3757);
and U9602 (N_9602,N_4928,N_3363);
nand U9603 (N_9603,N_4596,N_419);
and U9604 (N_9604,N_3448,N_3088);
nor U9605 (N_9605,N_2469,N_4645);
or U9606 (N_9606,N_54,N_288);
or U9607 (N_9607,N_1804,N_2688);
nand U9608 (N_9608,N_1771,N_3204);
or U9609 (N_9609,N_4,N_3815);
or U9610 (N_9610,N_602,N_1169);
or U9611 (N_9611,N_2469,N_4747);
nand U9612 (N_9612,N_363,N_3274);
xnor U9613 (N_9613,N_663,N_2366);
nor U9614 (N_9614,N_3000,N_4363);
and U9615 (N_9615,N_285,N_4019);
or U9616 (N_9616,N_4557,N_2633);
or U9617 (N_9617,N_1726,N_4746);
nand U9618 (N_9618,N_2763,N_2296);
or U9619 (N_9619,N_2346,N_1173);
nand U9620 (N_9620,N_2536,N_1280);
nand U9621 (N_9621,N_1832,N_140);
nand U9622 (N_9622,N_3156,N_1646);
and U9623 (N_9623,N_416,N_4568);
nand U9624 (N_9624,N_978,N_858);
nand U9625 (N_9625,N_3121,N_2315);
nor U9626 (N_9626,N_3567,N_4288);
and U9627 (N_9627,N_73,N_4834);
nor U9628 (N_9628,N_2153,N_1205);
nor U9629 (N_9629,N_4371,N_1589);
xnor U9630 (N_9630,N_1509,N_2763);
nor U9631 (N_9631,N_3327,N_3258);
and U9632 (N_9632,N_1661,N_3015);
nor U9633 (N_9633,N_1084,N_1014);
nor U9634 (N_9634,N_56,N_669);
nor U9635 (N_9635,N_536,N_647);
nor U9636 (N_9636,N_2469,N_918);
and U9637 (N_9637,N_4040,N_4386);
or U9638 (N_9638,N_1151,N_3545);
nor U9639 (N_9639,N_525,N_1707);
nand U9640 (N_9640,N_2547,N_3490);
or U9641 (N_9641,N_1792,N_1664);
nor U9642 (N_9642,N_4435,N_3530);
nand U9643 (N_9643,N_2318,N_4154);
and U9644 (N_9644,N_1156,N_420);
nor U9645 (N_9645,N_2273,N_806);
and U9646 (N_9646,N_1180,N_3434);
nand U9647 (N_9647,N_4371,N_2714);
nor U9648 (N_9648,N_2797,N_4290);
nand U9649 (N_9649,N_1474,N_480);
nor U9650 (N_9650,N_3223,N_4791);
and U9651 (N_9651,N_3045,N_310);
and U9652 (N_9652,N_1108,N_963);
nand U9653 (N_9653,N_3407,N_1077);
nor U9654 (N_9654,N_3624,N_2250);
or U9655 (N_9655,N_827,N_4657);
and U9656 (N_9656,N_3175,N_4513);
and U9657 (N_9657,N_4519,N_931);
nand U9658 (N_9658,N_2548,N_4578);
nor U9659 (N_9659,N_4500,N_2747);
or U9660 (N_9660,N_3487,N_448);
and U9661 (N_9661,N_26,N_3912);
nor U9662 (N_9662,N_4740,N_1535);
or U9663 (N_9663,N_4994,N_1325);
nand U9664 (N_9664,N_1545,N_1297);
and U9665 (N_9665,N_4918,N_2346);
nand U9666 (N_9666,N_2790,N_4334);
nor U9667 (N_9667,N_1490,N_2083);
nor U9668 (N_9668,N_3412,N_1960);
and U9669 (N_9669,N_3624,N_1807);
and U9670 (N_9670,N_1215,N_2314);
nand U9671 (N_9671,N_2045,N_35);
and U9672 (N_9672,N_4748,N_3862);
nand U9673 (N_9673,N_1487,N_4335);
and U9674 (N_9674,N_2697,N_3601);
and U9675 (N_9675,N_2828,N_81);
nand U9676 (N_9676,N_4547,N_756);
nand U9677 (N_9677,N_264,N_4532);
and U9678 (N_9678,N_4056,N_4441);
nand U9679 (N_9679,N_3894,N_3322);
nor U9680 (N_9680,N_533,N_1168);
nand U9681 (N_9681,N_3083,N_3138);
and U9682 (N_9682,N_861,N_1180);
xor U9683 (N_9683,N_1134,N_4169);
or U9684 (N_9684,N_1088,N_1065);
nor U9685 (N_9685,N_866,N_4198);
or U9686 (N_9686,N_4425,N_2945);
and U9687 (N_9687,N_4764,N_512);
and U9688 (N_9688,N_2571,N_4025);
nand U9689 (N_9689,N_2655,N_4143);
nand U9690 (N_9690,N_644,N_692);
nor U9691 (N_9691,N_715,N_3058);
or U9692 (N_9692,N_2342,N_2226);
nand U9693 (N_9693,N_173,N_528);
nand U9694 (N_9694,N_4709,N_3486);
nand U9695 (N_9695,N_1108,N_4769);
or U9696 (N_9696,N_3332,N_1856);
xnor U9697 (N_9697,N_2007,N_4289);
nand U9698 (N_9698,N_1962,N_4146);
nand U9699 (N_9699,N_3803,N_2841);
nand U9700 (N_9700,N_3584,N_766);
nor U9701 (N_9701,N_385,N_2065);
nor U9702 (N_9702,N_3023,N_2248);
or U9703 (N_9703,N_4291,N_1695);
nor U9704 (N_9704,N_2361,N_2580);
and U9705 (N_9705,N_3511,N_2658);
or U9706 (N_9706,N_2880,N_652);
and U9707 (N_9707,N_515,N_302);
and U9708 (N_9708,N_57,N_2295);
or U9709 (N_9709,N_4151,N_1255);
nand U9710 (N_9710,N_1018,N_4795);
and U9711 (N_9711,N_4497,N_2141);
and U9712 (N_9712,N_3433,N_1319);
or U9713 (N_9713,N_2110,N_2595);
nand U9714 (N_9714,N_2890,N_781);
and U9715 (N_9715,N_4355,N_827);
xnor U9716 (N_9716,N_1937,N_3289);
nor U9717 (N_9717,N_1485,N_4083);
nand U9718 (N_9718,N_1372,N_4489);
nand U9719 (N_9719,N_142,N_3942);
or U9720 (N_9720,N_2625,N_2092);
nor U9721 (N_9721,N_3855,N_4987);
and U9722 (N_9722,N_1508,N_208);
nor U9723 (N_9723,N_133,N_806);
nor U9724 (N_9724,N_4646,N_4149);
and U9725 (N_9725,N_3130,N_2769);
or U9726 (N_9726,N_3928,N_4673);
nand U9727 (N_9727,N_4658,N_4889);
nand U9728 (N_9728,N_351,N_4684);
and U9729 (N_9729,N_495,N_2535);
and U9730 (N_9730,N_1145,N_4901);
nand U9731 (N_9731,N_1297,N_4737);
nand U9732 (N_9732,N_1270,N_726);
nor U9733 (N_9733,N_825,N_643);
or U9734 (N_9734,N_4264,N_1970);
and U9735 (N_9735,N_4651,N_3718);
and U9736 (N_9736,N_52,N_3675);
nor U9737 (N_9737,N_2354,N_2255);
nand U9738 (N_9738,N_3445,N_3725);
or U9739 (N_9739,N_2390,N_4559);
nand U9740 (N_9740,N_4905,N_302);
xor U9741 (N_9741,N_3075,N_489);
nor U9742 (N_9742,N_1547,N_3231);
nand U9743 (N_9743,N_3985,N_1623);
nor U9744 (N_9744,N_2091,N_4565);
nand U9745 (N_9745,N_48,N_1346);
or U9746 (N_9746,N_2658,N_2330);
or U9747 (N_9747,N_1630,N_3278);
and U9748 (N_9748,N_1763,N_1207);
and U9749 (N_9749,N_3915,N_2804);
and U9750 (N_9750,N_4655,N_4572);
nor U9751 (N_9751,N_2730,N_4347);
or U9752 (N_9752,N_558,N_1246);
or U9753 (N_9753,N_2245,N_3328);
nor U9754 (N_9754,N_2638,N_2163);
nand U9755 (N_9755,N_4391,N_3591);
and U9756 (N_9756,N_910,N_3690);
and U9757 (N_9757,N_556,N_3779);
nor U9758 (N_9758,N_1051,N_208);
nand U9759 (N_9759,N_561,N_3818);
nand U9760 (N_9760,N_4617,N_240);
and U9761 (N_9761,N_19,N_684);
and U9762 (N_9762,N_2778,N_4652);
nor U9763 (N_9763,N_141,N_2863);
and U9764 (N_9764,N_4443,N_600);
or U9765 (N_9765,N_2458,N_326);
and U9766 (N_9766,N_2872,N_3534);
and U9767 (N_9767,N_4663,N_4256);
or U9768 (N_9768,N_1077,N_1486);
or U9769 (N_9769,N_569,N_236);
and U9770 (N_9770,N_4224,N_1595);
nor U9771 (N_9771,N_391,N_1180);
xor U9772 (N_9772,N_3562,N_2779);
or U9773 (N_9773,N_2840,N_3809);
nand U9774 (N_9774,N_780,N_2251);
nand U9775 (N_9775,N_2257,N_3761);
nand U9776 (N_9776,N_2690,N_854);
nor U9777 (N_9777,N_58,N_4631);
or U9778 (N_9778,N_4000,N_1780);
nor U9779 (N_9779,N_2835,N_868);
or U9780 (N_9780,N_2000,N_1511);
nor U9781 (N_9781,N_3215,N_1595);
nand U9782 (N_9782,N_453,N_2015);
nor U9783 (N_9783,N_3979,N_1184);
nor U9784 (N_9784,N_3212,N_3273);
or U9785 (N_9785,N_4428,N_492);
nand U9786 (N_9786,N_1137,N_3631);
xor U9787 (N_9787,N_437,N_2371);
and U9788 (N_9788,N_3703,N_3689);
or U9789 (N_9789,N_1655,N_2261);
nand U9790 (N_9790,N_791,N_431);
or U9791 (N_9791,N_4278,N_2513);
and U9792 (N_9792,N_2580,N_1208);
nand U9793 (N_9793,N_2639,N_2845);
nand U9794 (N_9794,N_2464,N_2017);
and U9795 (N_9795,N_3566,N_1086);
nand U9796 (N_9796,N_3145,N_2045);
or U9797 (N_9797,N_1973,N_4435);
and U9798 (N_9798,N_294,N_4848);
or U9799 (N_9799,N_342,N_3130);
nor U9800 (N_9800,N_563,N_3387);
nor U9801 (N_9801,N_568,N_1495);
nor U9802 (N_9802,N_2024,N_2183);
or U9803 (N_9803,N_4249,N_3528);
nor U9804 (N_9804,N_2766,N_3529);
nand U9805 (N_9805,N_3086,N_3289);
nand U9806 (N_9806,N_2433,N_880);
nand U9807 (N_9807,N_937,N_2807);
or U9808 (N_9808,N_1389,N_647);
or U9809 (N_9809,N_4331,N_1503);
and U9810 (N_9810,N_378,N_1757);
or U9811 (N_9811,N_4914,N_4002);
nand U9812 (N_9812,N_2332,N_3173);
and U9813 (N_9813,N_4446,N_409);
nand U9814 (N_9814,N_1417,N_3550);
nor U9815 (N_9815,N_2288,N_1186);
nor U9816 (N_9816,N_3497,N_2523);
or U9817 (N_9817,N_4374,N_2180);
and U9818 (N_9818,N_2899,N_3285);
nor U9819 (N_9819,N_2077,N_992);
nor U9820 (N_9820,N_2614,N_3927);
and U9821 (N_9821,N_4975,N_2124);
nand U9822 (N_9822,N_4399,N_2000);
nand U9823 (N_9823,N_343,N_3364);
and U9824 (N_9824,N_3291,N_1169);
nor U9825 (N_9825,N_2406,N_2962);
nor U9826 (N_9826,N_3362,N_3571);
nor U9827 (N_9827,N_2021,N_1780);
nor U9828 (N_9828,N_2144,N_449);
and U9829 (N_9829,N_29,N_2374);
and U9830 (N_9830,N_2425,N_4943);
or U9831 (N_9831,N_2891,N_4005);
nor U9832 (N_9832,N_2671,N_2700);
nor U9833 (N_9833,N_4748,N_4786);
or U9834 (N_9834,N_4763,N_2714);
and U9835 (N_9835,N_1387,N_821);
nand U9836 (N_9836,N_3016,N_4436);
and U9837 (N_9837,N_3942,N_2287);
nand U9838 (N_9838,N_3600,N_3184);
nand U9839 (N_9839,N_806,N_2367);
nor U9840 (N_9840,N_2810,N_1228);
and U9841 (N_9841,N_3279,N_252);
or U9842 (N_9842,N_4038,N_356);
nand U9843 (N_9843,N_4818,N_1130);
nor U9844 (N_9844,N_4041,N_445);
nand U9845 (N_9845,N_824,N_4993);
and U9846 (N_9846,N_3905,N_4764);
nor U9847 (N_9847,N_580,N_3358);
or U9848 (N_9848,N_4132,N_1442);
and U9849 (N_9849,N_4135,N_3825);
or U9850 (N_9850,N_1768,N_4258);
or U9851 (N_9851,N_4959,N_2103);
and U9852 (N_9852,N_4306,N_3844);
nand U9853 (N_9853,N_5,N_2984);
and U9854 (N_9854,N_520,N_2130);
nand U9855 (N_9855,N_1338,N_4404);
nand U9856 (N_9856,N_2777,N_4004);
nor U9857 (N_9857,N_3857,N_3476);
nor U9858 (N_9858,N_31,N_4657);
and U9859 (N_9859,N_2386,N_894);
and U9860 (N_9860,N_1869,N_3433);
or U9861 (N_9861,N_771,N_3453);
nand U9862 (N_9862,N_43,N_2931);
or U9863 (N_9863,N_2256,N_1722);
and U9864 (N_9864,N_2665,N_2721);
and U9865 (N_9865,N_115,N_3145);
and U9866 (N_9866,N_204,N_3383);
nand U9867 (N_9867,N_2342,N_697);
nor U9868 (N_9868,N_4068,N_4436);
nor U9869 (N_9869,N_4523,N_319);
and U9870 (N_9870,N_2146,N_1742);
or U9871 (N_9871,N_4636,N_4264);
or U9872 (N_9872,N_4370,N_3170);
nor U9873 (N_9873,N_2073,N_3219);
nand U9874 (N_9874,N_1119,N_1214);
nor U9875 (N_9875,N_14,N_4431);
or U9876 (N_9876,N_1198,N_4873);
xnor U9877 (N_9877,N_2870,N_4634);
and U9878 (N_9878,N_1639,N_3125);
and U9879 (N_9879,N_2797,N_4889);
nor U9880 (N_9880,N_1965,N_2208);
nor U9881 (N_9881,N_3249,N_1644);
nor U9882 (N_9882,N_2846,N_3999);
xor U9883 (N_9883,N_1736,N_4220);
and U9884 (N_9884,N_3184,N_914);
nand U9885 (N_9885,N_1393,N_2223);
xnor U9886 (N_9886,N_4890,N_4628);
nand U9887 (N_9887,N_4802,N_3312);
nor U9888 (N_9888,N_4858,N_3829);
nand U9889 (N_9889,N_572,N_4538);
or U9890 (N_9890,N_4665,N_4752);
and U9891 (N_9891,N_1143,N_1317);
and U9892 (N_9892,N_4269,N_43);
and U9893 (N_9893,N_1160,N_1847);
nor U9894 (N_9894,N_2142,N_2713);
nand U9895 (N_9895,N_4901,N_2620);
nand U9896 (N_9896,N_1658,N_4335);
nor U9897 (N_9897,N_483,N_419);
nand U9898 (N_9898,N_4431,N_315);
nor U9899 (N_9899,N_3007,N_560);
or U9900 (N_9900,N_3653,N_330);
or U9901 (N_9901,N_4608,N_1870);
nand U9902 (N_9902,N_3588,N_2775);
nand U9903 (N_9903,N_3387,N_3339);
xor U9904 (N_9904,N_2020,N_2853);
nor U9905 (N_9905,N_2599,N_4010);
nand U9906 (N_9906,N_3791,N_1519);
nand U9907 (N_9907,N_3918,N_259);
or U9908 (N_9908,N_3057,N_3273);
nand U9909 (N_9909,N_1019,N_2523);
nand U9910 (N_9910,N_4217,N_2048);
nor U9911 (N_9911,N_3434,N_3047);
nor U9912 (N_9912,N_3182,N_1814);
nor U9913 (N_9913,N_2260,N_2074);
xnor U9914 (N_9914,N_4590,N_3704);
or U9915 (N_9915,N_4172,N_4003);
or U9916 (N_9916,N_4982,N_4246);
or U9917 (N_9917,N_3549,N_441);
and U9918 (N_9918,N_4751,N_1047);
or U9919 (N_9919,N_1832,N_4499);
or U9920 (N_9920,N_2579,N_1356);
nor U9921 (N_9921,N_3095,N_3692);
and U9922 (N_9922,N_4222,N_2620);
nor U9923 (N_9923,N_2407,N_1966);
nor U9924 (N_9924,N_2581,N_3133);
nand U9925 (N_9925,N_4203,N_3861);
and U9926 (N_9926,N_1199,N_2940);
xnor U9927 (N_9927,N_92,N_4010);
or U9928 (N_9928,N_4740,N_1121);
nor U9929 (N_9929,N_930,N_3235);
nand U9930 (N_9930,N_796,N_2749);
nand U9931 (N_9931,N_1629,N_3128);
or U9932 (N_9932,N_618,N_389);
or U9933 (N_9933,N_758,N_4104);
nor U9934 (N_9934,N_2225,N_3955);
and U9935 (N_9935,N_1955,N_4970);
and U9936 (N_9936,N_4064,N_2415);
nor U9937 (N_9937,N_3650,N_2591);
and U9938 (N_9938,N_4513,N_2788);
nor U9939 (N_9939,N_3389,N_3065);
nand U9940 (N_9940,N_761,N_2354);
nand U9941 (N_9941,N_1881,N_3573);
nor U9942 (N_9942,N_2590,N_2615);
and U9943 (N_9943,N_1954,N_169);
or U9944 (N_9944,N_882,N_2385);
nand U9945 (N_9945,N_1878,N_4711);
nand U9946 (N_9946,N_4904,N_1315);
nor U9947 (N_9947,N_3745,N_4428);
and U9948 (N_9948,N_1620,N_4025);
or U9949 (N_9949,N_779,N_2598);
and U9950 (N_9950,N_1052,N_4414);
and U9951 (N_9951,N_3206,N_3889);
or U9952 (N_9952,N_341,N_715);
or U9953 (N_9953,N_2695,N_1591);
nand U9954 (N_9954,N_4440,N_2236);
nand U9955 (N_9955,N_3749,N_898);
or U9956 (N_9956,N_1569,N_157);
nor U9957 (N_9957,N_3635,N_1729);
nor U9958 (N_9958,N_2471,N_550);
or U9959 (N_9959,N_3471,N_2750);
or U9960 (N_9960,N_438,N_4640);
nor U9961 (N_9961,N_1808,N_4166);
nor U9962 (N_9962,N_2671,N_2608);
and U9963 (N_9963,N_2372,N_1725);
and U9964 (N_9964,N_4227,N_2564);
or U9965 (N_9965,N_414,N_2427);
nor U9966 (N_9966,N_762,N_2536);
and U9967 (N_9967,N_2990,N_507);
nor U9968 (N_9968,N_4559,N_4512);
nand U9969 (N_9969,N_1533,N_468);
nor U9970 (N_9970,N_4741,N_4548);
and U9971 (N_9971,N_4455,N_279);
nor U9972 (N_9972,N_4599,N_4253);
or U9973 (N_9973,N_4858,N_4321);
nand U9974 (N_9974,N_1571,N_4230);
or U9975 (N_9975,N_3738,N_1262);
nand U9976 (N_9976,N_2094,N_2942);
nor U9977 (N_9977,N_4046,N_2242);
or U9978 (N_9978,N_4542,N_1098);
nor U9979 (N_9979,N_4433,N_2385);
or U9980 (N_9980,N_764,N_3088);
xor U9981 (N_9981,N_3474,N_4895);
or U9982 (N_9982,N_1716,N_1275);
nand U9983 (N_9983,N_2333,N_1121);
nor U9984 (N_9984,N_1551,N_3703);
and U9985 (N_9985,N_4384,N_4973);
or U9986 (N_9986,N_2175,N_4052);
and U9987 (N_9987,N_3097,N_1197);
and U9988 (N_9988,N_600,N_950);
nor U9989 (N_9989,N_1373,N_4052);
or U9990 (N_9990,N_498,N_3866);
nor U9991 (N_9991,N_2612,N_2945);
or U9992 (N_9992,N_3916,N_2131);
nand U9993 (N_9993,N_2951,N_1615);
and U9994 (N_9994,N_784,N_3184);
or U9995 (N_9995,N_1636,N_99);
and U9996 (N_9996,N_286,N_524);
nand U9997 (N_9997,N_3117,N_4448);
and U9998 (N_9998,N_3917,N_11);
nand U9999 (N_9999,N_311,N_4874);
nand UO_0 (O_0,N_5102,N_7930);
nor UO_1 (O_1,N_8913,N_5921);
or UO_2 (O_2,N_7416,N_9108);
nand UO_3 (O_3,N_9412,N_5333);
xnor UO_4 (O_4,N_7685,N_9269);
or UO_5 (O_5,N_6215,N_5338);
nand UO_6 (O_6,N_8130,N_6308);
and UO_7 (O_7,N_5538,N_9358);
or UO_8 (O_8,N_8672,N_6531);
or UO_9 (O_9,N_6165,N_8113);
and UO_10 (O_10,N_8204,N_5770);
or UO_11 (O_11,N_6597,N_8151);
or UO_12 (O_12,N_9981,N_5882);
or UO_13 (O_13,N_7436,N_9496);
nor UO_14 (O_14,N_7691,N_7086);
nand UO_15 (O_15,N_5835,N_8694);
xor UO_16 (O_16,N_9676,N_6708);
nor UO_17 (O_17,N_9497,N_9103);
and UO_18 (O_18,N_6617,N_9001);
nor UO_19 (O_19,N_6945,N_9641);
nor UO_20 (O_20,N_9443,N_8363);
and UO_21 (O_21,N_9402,N_8689);
xnor UO_22 (O_22,N_7374,N_7655);
nand UO_23 (O_23,N_7388,N_9891);
nor UO_24 (O_24,N_9219,N_7980);
xnor UO_25 (O_25,N_5091,N_6787);
or UO_26 (O_26,N_6272,N_7471);
nand UO_27 (O_27,N_6565,N_5824);
or UO_28 (O_28,N_7643,N_7236);
nand UO_29 (O_29,N_7078,N_9717);
nand UO_30 (O_30,N_5808,N_5070);
nor UO_31 (O_31,N_5024,N_6784);
or UO_32 (O_32,N_9809,N_6760);
nor UO_33 (O_33,N_7110,N_8926);
and UO_34 (O_34,N_6742,N_9499);
and UO_35 (O_35,N_9617,N_9996);
or UO_36 (O_36,N_9986,N_5236);
or UO_37 (O_37,N_7451,N_6640);
or UO_38 (O_38,N_5879,N_5115);
and UO_39 (O_39,N_6131,N_8166);
and UO_40 (O_40,N_7612,N_5011);
and UO_41 (O_41,N_5419,N_9018);
or UO_42 (O_42,N_8624,N_5677);
nor UO_43 (O_43,N_9045,N_8815);
nand UO_44 (O_44,N_7763,N_5174);
nor UO_45 (O_45,N_8998,N_5249);
and UO_46 (O_46,N_6081,N_5660);
nand UO_47 (O_47,N_8801,N_5001);
nor UO_48 (O_48,N_7143,N_7144);
or UO_49 (O_49,N_7011,N_6044);
xnor UO_50 (O_50,N_8799,N_7058);
nand UO_51 (O_51,N_6070,N_8845);
nand UO_52 (O_52,N_6395,N_6413);
nand UO_53 (O_53,N_8293,N_5943);
nand UO_54 (O_54,N_8723,N_8902);
nor UO_55 (O_55,N_9854,N_6690);
and UO_56 (O_56,N_8663,N_6257);
or UO_57 (O_57,N_6752,N_6851);
or UO_58 (O_58,N_6483,N_5222);
nor UO_59 (O_59,N_7611,N_9249);
nand UO_60 (O_60,N_9738,N_7540);
and UO_61 (O_61,N_8083,N_9245);
xnor UO_62 (O_62,N_7921,N_7813);
nand UO_63 (O_63,N_7102,N_5244);
nor UO_64 (O_64,N_5522,N_6190);
and UO_65 (O_65,N_5811,N_9461);
nor UO_66 (O_66,N_7559,N_9229);
xor UO_67 (O_67,N_6009,N_6360);
nand UO_68 (O_68,N_5080,N_7072);
and UO_69 (O_69,N_5324,N_9916);
nand UO_70 (O_70,N_6829,N_7607);
nand UO_71 (O_71,N_8231,N_7184);
nor UO_72 (O_72,N_5365,N_9863);
nor UO_73 (O_73,N_6814,N_7196);
or UO_74 (O_74,N_9762,N_6125);
and UO_75 (O_75,N_6668,N_5747);
nor UO_76 (O_76,N_6912,N_9642);
or UO_77 (O_77,N_9083,N_9488);
nor UO_78 (O_78,N_9369,N_9519);
and UO_79 (O_79,N_9119,N_9091);
nor UO_80 (O_80,N_9516,N_9743);
or UO_81 (O_81,N_9753,N_9155);
and UO_82 (O_82,N_5175,N_9089);
nand UO_83 (O_83,N_9065,N_6620);
or UO_84 (O_84,N_6260,N_8922);
nor UO_85 (O_85,N_7270,N_6545);
and UO_86 (O_86,N_8659,N_5107);
and UO_87 (O_87,N_8236,N_9677);
nor UO_88 (O_88,N_9475,N_6812);
nor UO_89 (O_89,N_5858,N_6994);
or UO_90 (O_90,N_5966,N_6654);
nand UO_91 (O_91,N_9974,N_5743);
and UO_92 (O_92,N_6628,N_8167);
or UO_93 (O_93,N_6553,N_8911);
nor UO_94 (O_94,N_5006,N_6189);
nand UO_95 (O_95,N_8608,N_9750);
or UO_96 (O_96,N_5823,N_5642);
nor UO_97 (O_97,N_9152,N_5780);
or UO_98 (O_98,N_7588,N_7850);
nand UO_99 (O_99,N_5904,N_5157);
nand UO_100 (O_100,N_6169,N_9137);
or UO_101 (O_101,N_5326,N_6805);
and UO_102 (O_102,N_5438,N_7573);
or UO_103 (O_103,N_9346,N_8310);
and UO_104 (O_104,N_8170,N_6704);
nand UO_105 (O_105,N_9262,N_6033);
or UO_106 (O_106,N_8417,N_5672);
or UO_107 (O_107,N_9212,N_7867);
and UO_108 (O_108,N_9790,N_9841);
and UO_109 (O_109,N_8732,N_6627);
nor UO_110 (O_110,N_8772,N_7729);
or UO_111 (O_111,N_6621,N_7030);
or UO_112 (O_112,N_8557,N_5550);
nand UO_113 (O_113,N_5322,N_7803);
nor UO_114 (O_114,N_5388,N_6476);
nand UO_115 (O_115,N_6614,N_8391);
nor UO_116 (O_116,N_9679,N_6057);
nor UO_117 (O_117,N_7268,N_9701);
and UO_118 (O_118,N_8094,N_8379);
nand UO_119 (O_119,N_9355,N_6132);
or UO_120 (O_120,N_7247,N_6767);
nor UO_121 (O_121,N_9168,N_6422);
or UO_122 (O_122,N_6105,N_6246);
nor UO_123 (O_123,N_9194,N_6468);
nand UO_124 (O_124,N_9541,N_6339);
nand UO_125 (O_125,N_7570,N_7961);
or UO_126 (O_126,N_6035,N_6355);
or UO_127 (O_127,N_6879,N_5878);
or UO_128 (O_128,N_6734,N_6327);
nand UO_129 (O_129,N_8843,N_8014);
or UO_130 (O_130,N_6954,N_9304);
nor UO_131 (O_131,N_6836,N_5826);
or UO_132 (O_132,N_7115,N_9940);
xnor UO_133 (O_133,N_9768,N_9321);
nor UO_134 (O_134,N_5467,N_7764);
and UO_135 (O_135,N_8896,N_5893);
or UO_136 (O_136,N_5217,N_6867);
nor UO_137 (O_137,N_9274,N_7008);
and UO_138 (O_138,N_8467,N_5142);
or UO_139 (O_139,N_7207,N_6645);
and UO_140 (O_140,N_6328,N_6604);
and UO_141 (O_141,N_9786,N_6456);
nand UO_142 (O_142,N_5705,N_7375);
nand UO_143 (O_143,N_5089,N_6801);
nor UO_144 (O_144,N_5674,N_9374);
or UO_145 (O_145,N_5922,N_5171);
and UO_146 (O_146,N_5450,N_5699);
or UO_147 (O_147,N_6968,N_9002);
nand UO_148 (O_148,N_9605,N_8301);
or UO_149 (O_149,N_5487,N_9494);
and UO_150 (O_150,N_9399,N_7034);
nor UO_151 (O_151,N_6644,N_5295);
nor UO_152 (O_152,N_5177,N_8838);
or UO_153 (O_153,N_7628,N_7895);
or UO_154 (O_154,N_6475,N_9156);
nand UO_155 (O_155,N_6925,N_9631);
or UO_156 (O_156,N_8985,N_6126);
nor UO_157 (O_157,N_6003,N_6015);
and UO_158 (O_158,N_9817,N_6709);
and UO_159 (O_159,N_8077,N_8058);
or UO_160 (O_160,N_5393,N_7329);
and UO_161 (O_161,N_8543,N_6243);
nor UO_162 (O_162,N_6554,N_9433);
and UO_163 (O_163,N_6838,N_5636);
and UO_164 (O_164,N_9362,N_9422);
nor UO_165 (O_165,N_5968,N_7593);
or UO_166 (O_166,N_7864,N_9834);
or UO_167 (O_167,N_7299,N_6130);
or UO_168 (O_168,N_6083,N_7314);
and UO_169 (O_169,N_6870,N_5809);
nand UO_170 (O_170,N_6825,N_8386);
xnor UO_171 (O_171,N_7892,N_7448);
nand UO_172 (O_172,N_5300,N_8741);
and UO_173 (O_173,N_7551,N_8459);
xor UO_174 (O_174,N_7185,N_7529);
or UO_175 (O_175,N_7241,N_6445);
and UO_176 (O_176,N_7337,N_5353);
nand UO_177 (O_177,N_7440,N_9059);
nand UO_178 (O_178,N_6205,N_7082);
and UO_179 (O_179,N_9446,N_6529);
nand UO_180 (O_180,N_7336,N_7470);
and UO_181 (O_181,N_5418,N_7784);
and UO_182 (O_182,N_9545,N_9917);
and UO_183 (O_183,N_5383,N_8583);
nor UO_184 (O_184,N_5109,N_7794);
nor UO_185 (O_185,N_7810,N_7477);
nor UO_186 (O_186,N_9153,N_9344);
and UO_187 (O_187,N_5323,N_5122);
nand UO_188 (O_188,N_8376,N_9512);
nor UO_189 (O_189,N_9439,N_6472);
nand UO_190 (O_190,N_6139,N_5130);
and UO_191 (O_191,N_9730,N_9894);
and UO_192 (O_192,N_9534,N_7123);
and UO_193 (O_193,N_6425,N_8773);
nor UO_194 (O_194,N_9359,N_9231);
nor UO_195 (O_195,N_5124,N_6095);
and UO_196 (O_196,N_5013,N_9182);
nand UO_197 (O_197,N_7438,N_8008);
nor UO_198 (O_198,N_6559,N_6290);
nand UO_199 (O_199,N_5870,N_6128);
xor UO_200 (O_200,N_6089,N_9892);
nor UO_201 (O_201,N_7823,N_8532);
nor UO_202 (O_202,N_6262,N_8341);
or UO_203 (O_203,N_9092,N_7390);
xnor UO_204 (O_204,N_5030,N_5817);
and UO_205 (O_205,N_7775,N_7589);
nor UO_206 (O_206,N_5100,N_9813);
nand UO_207 (O_207,N_9339,N_5570);
nor UO_208 (O_208,N_5661,N_5955);
nor UO_209 (O_209,N_5237,N_6098);
or UO_210 (O_210,N_9919,N_7595);
nand UO_211 (O_211,N_5099,N_7974);
and UO_212 (O_212,N_9553,N_6869);
xor UO_213 (O_213,N_9252,N_7317);
or UO_214 (O_214,N_6901,N_6728);
and UO_215 (O_215,N_5709,N_7124);
nand UO_216 (O_216,N_9132,N_6657);
and UO_217 (O_217,N_8273,N_9118);
or UO_218 (O_218,N_5996,N_5377);
and UO_219 (O_219,N_7069,N_9003);
and UO_220 (O_220,N_6878,N_7945);
nand UO_221 (O_221,N_5457,N_8103);
nand UO_222 (O_222,N_8964,N_9409);
nor UO_223 (O_223,N_5216,N_6774);
nor UO_224 (O_224,N_5867,N_5039);
and UO_225 (O_225,N_9131,N_8333);
nor UO_226 (O_226,N_9945,N_8359);
nand UO_227 (O_227,N_5860,N_6052);
and UO_228 (O_228,N_8099,N_8050);
nand UO_229 (O_229,N_7662,N_7792);
or UO_230 (O_230,N_6646,N_7107);
nand UO_231 (O_231,N_5724,N_8511);
nand UO_232 (O_232,N_9026,N_6135);
nor UO_233 (O_233,N_9053,N_8766);
nor UO_234 (O_234,N_5678,N_9959);
or UO_235 (O_235,N_7862,N_9444);
nand UO_236 (O_236,N_6210,N_8397);
nor UO_237 (O_237,N_5206,N_5204);
nor UO_238 (O_238,N_7742,N_6523);
nor UO_239 (O_239,N_5374,N_8404);
and UO_240 (O_240,N_8821,N_5746);
xor UO_241 (O_241,N_6357,N_5977);
and UO_242 (O_242,N_8044,N_9550);
nand UO_243 (O_243,N_8355,N_5992);
nor UO_244 (O_244,N_7488,N_5799);
nand UO_245 (O_245,N_5077,N_6334);
or UO_246 (O_246,N_8952,N_8597);
nor UO_247 (O_247,N_9086,N_5009);
and UO_248 (O_248,N_5573,N_6622);
nor UO_249 (O_249,N_9827,N_9862);
nand UO_250 (O_250,N_9998,N_6772);
nor UO_251 (O_251,N_8161,N_5275);
nand UO_252 (O_252,N_8452,N_8500);
or UO_253 (O_253,N_9174,N_5763);
nor UO_254 (O_254,N_5474,N_5460);
or UO_255 (O_255,N_7884,N_8461);
nand UO_256 (O_256,N_7901,N_8146);
or UO_257 (O_257,N_7800,N_8668);
or UO_258 (O_258,N_9818,N_9203);
and UO_259 (O_259,N_5373,N_9273);
nand UO_260 (O_260,N_5640,N_5126);
xor UO_261 (O_261,N_8975,N_7262);
nor UO_262 (O_262,N_6388,N_9657);
and UO_263 (O_263,N_8762,N_9902);
nor UO_264 (O_264,N_7659,N_8238);
nor UO_265 (O_265,N_6942,N_7172);
and UO_266 (O_266,N_8371,N_9543);
nor UO_267 (O_267,N_5276,N_9463);
or UO_268 (O_268,N_8043,N_6444);
and UO_269 (O_269,N_7905,N_5361);
or UO_270 (O_270,N_6679,N_8610);
or UO_271 (O_271,N_8574,N_8810);
nor UO_272 (O_272,N_6350,N_8639);
and UO_273 (O_273,N_8319,N_7600);
or UO_274 (O_274,N_8742,N_5469);
or UO_275 (O_275,N_7261,N_9610);
or UO_276 (O_276,N_6889,N_8612);
and UO_277 (O_277,N_9146,N_6791);
nor UO_278 (O_278,N_9546,N_6376);
nand UO_279 (O_279,N_9686,N_6658);
nand UO_280 (O_280,N_5164,N_7049);
nand UO_281 (O_281,N_8925,N_5702);
and UO_282 (O_282,N_9139,N_8234);
nand UO_283 (O_283,N_5925,N_7520);
nand UO_284 (O_284,N_7431,N_5987);
and UO_285 (O_285,N_6223,N_6401);
nor UO_286 (O_286,N_6740,N_8060);
or UO_287 (O_287,N_6955,N_9347);
xor UO_288 (O_288,N_6458,N_8786);
nand UO_289 (O_289,N_9885,N_6129);
nor UO_290 (O_290,N_8314,N_8803);
nor UO_291 (O_291,N_5886,N_8826);
nor UO_292 (O_292,N_9825,N_8835);
nand UO_293 (O_293,N_9284,N_5425);
or UO_294 (O_294,N_9232,N_9205);
nand UO_295 (O_295,N_6859,N_8478);
or UO_296 (O_296,N_7796,N_5197);
nor UO_297 (O_297,N_7765,N_8444);
nor UO_298 (O_298,N_5494,N_8136);
and UO_299 (O_299,N_6331,N_8480);
nor UO_300 (O_300,N_9987,N_9125);
or UO_301 (O_301,N_7754,N_5047);
nor UO_302 (O_302,N_8721,N_9082);
nor UO_303 (O_303,N_8448,N_7865);
nor UO_304 (O_304,N_7672,N_8393);
nor UO_305 (O_305,N_8941,N_9434);
or UO_306 (O_306,N_7349,N_7669);
nand UO_307 (O_307,N_6498,N_9529);
nand UO_308 (O_308,N_5371,N_9844);
or UO_309 (O_309,N_9832,N_5914);
nand UO_310 (O_310,N_7826,N_9297);
or UO_311 (O_311,N_6440,N_8981);
nand UO_312 (O_312,N_5631,N_6716);
nand UO_313 (O_313,N_5283,N_5635);
or UO_314 (O_314,N_8795,N_8358);
nor UO_315 (O_315,N_6754,N_8388);
or UO_316 (O_316,N_7780,N_9907);
nand UO_317 (O_317,N_9847,N_8362);
and UO_318 (O_318,N_6244,N_9525);
nand UO_319 (O_319,N_6637,N_8267);
nand UO_320 (O_320,N_7485,N_9848);
nand UO_321 (O_321,N_7205,N_5167);
or UO_322 (O_322,N_7511,N_6963);
nand UO_323 (O_323,N_5211,N_9366);
and UO_324 (O_324,N_6281,N_6564);
nand UO_325 (O_325,N_8777,N_5659);
and UO_326 (O_326,N_7933,N_6178);
nand UO_327 (O_327,N_5583,N_9878);
nor UO_328 (O_328,N_5604,N_8134);
or UO_329 (O_329,N_9333,N_5078);
nor UO_330 (O_330,N_7458,N_5155);
and UO_331 (O_331,N_5725,N_8768);
nand UO_332 (O_332,N_9142,N_5857);
or UO_333 (O_333,N_5213,N_8318);
nand UO_334 (O_334,N_9975,N_8878);
and UO_335 (O_335,N_6071,N_5394);
or UO_336 (O_336,N_8451,N_8097);
and UO_337 (O_337,N_7094,N_9635);
and UO_338 (O_338,N_7041,N_6739);
nand UO_339 (O_339,N_8701,N_7723);
or UO_340 (O_340,N_9332,N_6027);
or UO_341 (O_341,N_5958,N_9719);
nand UO_342 (O_342,N_8651,N_7189);
nand UO_343 (O_343,N_7047,N_5548);
xnor UO_344 (O_344,N_6577,N_6799);
or UO_345 (O_345,N_9382,N_7582);
nand UO_346 (O_346,N_9342,N_6600);
and UO_347 (O_347,N_9031,N_5569);
and UO_348 (O_348,N_8212,N_6750);
nand UO_349 (O_349,N_7635,N_6006);
nor UO_350 (O_350,N_5228,N_9157);
and UO_351 (O_351,N_6624,N_9643);
nand UO_352 (O_352,N_9306,N_7420);
xnor UO_353 (O_353,N_5859,N_8600);
and UO_354 (O_354,N_8122,N_8887);
or UO_355 (O_355,N_7000,N_7234);
or UO_356 (O_356,N_9170,N_9654);
xor UO_357 (O_357,N_9791,N_6714);
xor UO_358 (O_358,N_9705,N_6601);
and UO_359 (O_359,N_5629,N_8085);
nand UO_360 (O_360,N_6359,N_9084);
xnor UO_361 (O_361,N_7820,N_5180);
and UO_362 (O_362,N_7517,N_6944);
nor UO_363 (O_363,N_8104,N_5536);
and UO_364 (O_364,N_9549,N_9624);
or UO_365 (O_365,N_6034,N_8631);
and UO_366 (O_366,N_9783,N_5815);
nor UO_367 (O_367,N_9842,N_7956);
nor UO_368 (O_368,N_8764,N_5287);
or UO_369 (O_369,N_9567,N_9729);
and UO_370 (O_370,N_8549,N_7287);
or UO_371 (O_371,N_8877,N_5482);
and UO_372 (O_372,N_7907,N_9852);
and UO_373 (O_373,N_5931,N_5641);
nand UO_374 (O_374,N_5481,N_7958);
and UO_375 (O_375,N_8670,N_6194);
and UO_376 (O_376,N_5121,N_6305);
or UO_377 (O_377,N_5723,N_6183);
nand UO_378 (O_378,N_7854,N_8797);
nand UO_379 (O_379,N_9619,N_5138);
nor UO_380 (O_380,N_8072,N_7362);
and UO_381 (O_381,N_9370,N_5549);
nor UO_382 (O_382,N_9391,N_8729);
or UO_383 (O_383,N_6462,N_5452);
nand UO_384 (O_384,N_5971,N_8126);
nor UO_385 (O_385,N_9055,N_8185);
or UO_386 (O_386,N_9950,N_5158);
nor UO_387 (O_387,N_8547,N_8957);
nand UO_388 (O_388,N_9353,N_5762);
and UO_389 (O_389,N_7392,N_7461);
nor UO_390 (O_390,N_5579,N_9038);
nand UO_391 (O_391,N_8502,N_8493);
nor UO_392 (O_392,N_6965,N_7146);
or UO_393 (O_393,N_5576,N_6623);
or UO_394 (O_394,N_5719,N_9503);
and UO_395 (O_395,N_6978,N_7577);
nor UO_396 (O_396,N_8935,N_8013);
and UO_397 (O_397,N_7063,N_8372);
or UO_398 (O_398,N_7311,N_8554);
and UO_399 (O_399,N_6802,N_7541);
or UO_400 (O_400,N_5832,N_6478);
nor UO_401 (O_401,N_9966,N_7727);
and UO_402 (O_402,N_7518,N_5691);
nor UO_403 (O_403,N_9363,N_9493);
or UO_404 (O_404,N_8886,N_6186);
or UO_405 (O_405,N_5431,N_7500);
nor UO_406 (O_406,N_8225,N_9239);
nand UO_407 (O_407,N_6108,N_7565);
or UO_408 (O_408,N_9429,N_9487);
and UO_409 (O_409,N_7696,N_8249);
and UO_410 (O_410,N_7935,N_9853);
or UO_411 (O_411,N_8472,N_6489);
or UO_412 (O_412,N_8034,N_7838);
nand UO_413 (O_413,N_5288,N_6151);
nor UO_414 (O_414,N_8984,N_6687);
nand UO_415 (O_415,N_6049,N_6524);
nor UO_416 (O_416,N_7979,N_5471);
nand UO_417 (O_417,N_7563,N_9656);
nor UO_418 (O_418,N_7004,N_6217);
nor UO_419 (O_419,N_8573,N_5301);
and UO_420 (O_420,N_8110,N_7130);
nor UO_421 (O_421,N_7739,N_6797);
nand UO_422 (O_422,N_5706,N_5871);
xnor UO_423 (O_423,N_5403,N_6496);
nor UO_424 (O_424,N_8759,N_7598);
nor UO_425 (O_425,N_5646,N_7028);
and UO_426 (O_426,N_7219,N_9006);
nand UO_427 (O_427,N_6090,N_7339);
and UO_428 (O_428,N_7206,N_7298);
or UO_429 (O_429,N_9835,N_8324);
nor UO_430 (O_430,N_5639,N_7285);
nand UO_431 (O_431,N_6631,N_7626);
nand UO_432 (O_432,N_6710,N_9540);
nor UO_433 (O_433,N_5697,N_9751);
and UO_434 (O_434,N_5653,N_6174);
nand UO_435 (O_435,N_9165,N_5575);
or UO_436 (O_436,N_6193,N_5994);
or UO_437 (O_437,N_5007,N_6741);
nor UO_438 (O_438,N_9517,N_9017);
nor UO_439 (O_439,N_8514,N_7751);
or UO_440 (O_440,N_6147,N_5856);
nand UO_441 (O_441,N_5502,N_7015);
and UO_442 (O_442,N_6252,N_9413);
and UO_443 (O_443,N_8783,N_8295);
xnor UO_444 (O_444,N_7700,N_6284);
or UO_445 (O_445,N_9060,N_8163);
nor UO_446 (O_446,N_5008,N_8010);
or UO_447 (O_447,N_6660,N_7964);
nand UO_448 (O_448,N_7297,N_6168);
nor UO_449 (O_449,N_9187,N_7999);
nand UO_450 (O_450,N_5280,N_5478);
and UO_451 (O_451,N_8428,N_8398);
and UO_452 (O_452,N_6446,N_9872);
and UO_453 (O_453,N_5359,N_6952);
or UO_454 (O_454,N_9670,N_5065);
or UO_455 (O_455,N_8108,N_6439);
xor UO_456 (O_456,N_6214,N_9547);
nor UO_457 (O_457,N_6857,N_8011);
and UO_458 (O_458,N_9754,N_9218);
nor UO_459 (O_459,N_5510,N_6695);
or UO_460 (O_460,N_8971,N_8041);
and UO_461 (O_461,N_6259,N_8778);
nor UO_462 (O_462,N_5045,N_8958);
nor UO_463 (O_463,N_6932,N_9291);
nand UO_464 (O_464,N_5830,N_6776);
or UO_465 (O_465,N_5598,N_8458);
nor UO_466 (O_466,N_6042,N_8872);
and UO_467 (O_467,N_6803,N_8496);
and UO_468 (O_468,N_7399,N_8842);
nor UO_469 (O_469,N_7989,N_7748);
and UO_470 (O_470,N_8177,N_8223);
or UO_471 (O_471,N_5599,N_8062);
nor UO_472 (O_472,N_7567,N_6579);
nor UO_473 (O_473,N_5057,N_6539);
nand UO_474 (O_474,N_8380,N_8447);
nand UO_475 (O_475,N_6557,N_8654);
nand UO_476 (O_476,N_8337,N_9167);
nand UO_477 (O_477,N_6289,N_9352);
and UO_478 (O_478,N_9933,N_8403);
and UO_479 (O_479,N_5546,N_9718);
nand UO_480 (O_480,N_9081,N_5503);
and UO_481 (O_481,N_6573,N_9840);
nor UO_482 (O_482,N_7161,N_5890);
and UO_483 (O_483,N_6023,N_6166);
and UO_484 (O_484,N_9855,N_9068);
or UO_485 (O_485,N_5738,N_8775);
nor UO_486 (O_486,N_7716,N_8748);
nor UO_487 (O_487,N_8237,N_8174);
and UO_488 (O_488,N_9597,N_6022);
and UO_489 (O_489,N_6104,N_6062);
nor UO_490 (O_490,N_6002,N_8196);
nor UO_491 (O_491,N_5517,N_6267);
nand UO_492 (O_492,N_8885,N_7973);
xnor UO_493 (O_493,N_6465,N_7051);
nor UO_494 (O_494,N_7100,N_7957);
or UO_495 (O_495,N_6897,N_7427);
or UO_496 (O_496,N_8120,N_7753);
and UO_497 (O_497,N_7652,N_9178);
nand UO_498 (O_498,N_6699,N_7624);
nand UO_499 (O_499,N_5578,N_9228);
and UO_500 (O_500,N_6661,N_7649);
nor UO_501 (O_501,N_8944,N_9538);
or UO_502 (O_502,N_5028,N_9481);
nor UO_503 (O_503,N_8717,N_8508);
and UO_504 (O_504,N_5755,N_5923);
nor UO_505 (O_505,N_6546,N_9141);
or UO_506 (O_506,N_5416,N_5310);
and UO_507 (O_507,N_9280,N_7323);
nand UO_508 (O_508,N_6997,N_5215);
or UO_509 (O_509,N_8744,N_7983);
nor UO_510 (O_510,N_7195,N_5146);
or UO_511 (O_511,N_7762,N_5504);
nor UO_512 (O_512,N_6029,N_9047);
nor UO_513 (O_513,N_6103,N_6584);
or UO_514 (O_514,N_5243,N_9314);
nand UO_515 (O_515,N_6939,N_6398);
nand UO_516 (O_516,N_6552,N_9238);
nor UO_517 (O_517,N_8870,N_7245);
or UO_518 (O_518,N_7689,N_8469);
nor UO_519 (O_519,N_7068,N_6138);
or UO_520 (O_520,N_9526,N_9161);
nand UO_521 (O_521,N_5477,N_6732);
and UO_522 (O_522,N_5611,N_8009);
nand UO_523 (O_523,N_6650,N_7103);
or UO_524 (O_524,N_8805,N_8284);
or UO_525 (O_525,N_9063,N_9367);
or UO_526 (O_526,N_7188,N_7851);
and UO_527 (O_527,N_7083,N_9169);
xnor UO_528 (O_528,N_6636,N_5509);
nand UO_529 (O_529,N_5978,N_8195);
and UO_530 (O_530,N_7940,N_8264);
nand UO_531 (O_531,N_5563,N_8344);
xnor UO_532 (O_532,N_5372,N_6429);
nand UO_533 (O_533,N_9849,N_6196);
or UO_534 (O_534,N_8831,N_8018);
nand UO_535 (O_535,N_7680,N_9931);
nand UO_536 (O_536,N_6967,N_5543);
nor UO_537 (O_537,N_8630,N_9838);
nand UO_538 (O_538,N_9420,N_6266);
nand UO_539 (O_539,N_6474,N_5730);
xnor UO_540 (O_540,N_8735,N_9015);
nor UO_541 (O_541,N_5590,N_6338);
nand UO_542 (O_542,N_9021,N_6040);
or UO_543 (O_543,N_6093,N_5259);
nor UO_544 (O_544,N_9570,N_8875);
or UO_545 (O_545,N_9162,N_9900);
and UO_546 (O_546,N_9057,N_7531);
nand UO_547 (O_547,N_5033,N_7056);
nand UO_548 (O_548,N_9708,N_7985);
xor UO_549 (O_549,N_7098,N_6972);
and UO_550 (O_550,N_5527,N_6816);
nor UO_551 (O_551,N_8178,N_7804);
and UO_552 (O_552,N_8818,N_8147);
nand UO_553 (O_553,N_9448,N_5897);
and UO_554 (O_554,N_9527,N_6228);
nand UO_555 (O_555,N_8017,N_7858);
nor UO_556 (O_556,N_5220,N_5785);
nand UO_557 (O_557,N_8501,N_9775);
nand UO_558 (O_558,N_7106,N_8712);
nor UO_559 (O_559,N_6826,N_7325);
or UO_560 (O_560,N_5584,N_8145);
nor UO_561 (O_561,N_8304,N_5540);
nor UO_562 (O_562,N_7977,N_8978);
and UO_563 (O_563,N_5818,N_7183);
nor UO_564 (O_564,N_5567,N_6491);
nor UO_565 (O_565,N_8131,N_5245);
nand UO_566 (O_566,N_7080,N_9793);
or UO_567 (O_567,N_5501,N_5076);
nand UO_568 (O_568,N_6815,N_9360);
nor UO_569 (O_569,N_8367,N_6335);
or UO_570 (O_570,N_6510,N_7352);
or UO_571 (O_571,N_9099,N_6255);
or UO_572 (O_572,N_5408,N_6216);
and UO_573 (O_573,N_7487,N_9257);
nor UO_574 (O_574,N_6056,N_7404);
and UO_575 (O_575,N_7164,N_9421);
nand UO_576 (O_576,N_6635,N_7237);
nor UO_577 (O_577,N_8825,N_9076);
nor UO_578 (O_578,N_8640,N_6821);
and UO_579 (O_579,N_7359,N_6583);
or UO_580 (O_580,N_9430,N_8855);
and UO_581 (O_581,N_9992,N_9106);
xnor UO_582 (O_582,N_5680,N_6854);
nor UO_583 (O_583,N_9577,N_7200);
or UO_584 (O_584,N_6833,N_7145);
nor UO_585 (O_585,N_7660,N_6689);
nor UO_586 (O_586,N_8931,N_9311);
nor UO_587 (O_587,N_7277,N_7807);
or UO_588 (O_588,N_5791,N_9225);
and UO_589 (O_589,N_7318,N_7027);
xnor UO_590 (O_590,N_8587,N_6811);
and UO_591 (O_591,N_5050,N_8288);
nand UO_592 (O_592,N_5754,N_5516);
or UO_593 (O_593,N_5272,N_8986);
and UO_594 (O_594,N_6729,N_5294);
nand UO_595 (O_595,N_5402,N_6686);
and UO_596 (O_596,N_9887,N_8435);
xor UO_597 (O_597,N_5473,N_9824);
or UO_598 (O_598,N_6344,N_7613);
or UO_599 (O_599,N_8025,N_7350);
or UO_600 (O_600,N_8261,N_8290);
or UO_601 (O_601,N_9637,N_6014);
and UO_602 (O_602,N_8620,N_6115);
nor UO_603 (O_603,N_5190,N_8248);
and UO_604 (O_604,N_6771,N_6497);
and UO_605 (O_605,N_9890,N_6894);
nand UO_606 (O_606,N_8325,N_8253);
or UO_607 (O_607,N_5991,N_7581);
or UO_608 (O_608,N_9868,N_5376);
and UO_609 (O_609,N_8987,N_5166);
or UO_610 (O_610,N_5081,N_8862);
and UO_611 (O_611,N_8138,N_5348);
nor UO_612 (O_612,N_9723,N_6188);
and UO_613 (O_613,N_6948,N_9601);
or UO_614 (O_614,N_6322,N_9877);
and UO_615 (O_615,N_5453,N_5628);
or UO_616 (O_616,N_7396,N_8497);
or UO_617 (O_617,N_5307,N_5690);
nor UO_618 (O_618,N_9915,N_6986);
or UO_619 (O_619,N_6719,N_7639);
nor UO_620 (O_620,N_8739,N_8117);
xor UO_621 (O_621,N_8946,N_5898);
nand UO_622 (O_622,N_9242,N_6466);
nor UO_623 (O_623,N_7046,N_5002);
or UO_624 (O_624,N_5937,N_8577);
and UO_625 (O_625,N_7125,N_7258);
nor UO_626 (O_626,N_9952,N_9766);
or UO_627 (O_627,N_9953,N_5456);
nor UO_628 (O_628,N_9958,N_8753);
nor UO_629 (O_629,N_9523,N_5414);
nand UO_630 (O_630,N_7126,N_8649);
nand UO_631 (O_631,N_7335,N_9233);
nor UO_632 (O_632,N_7148,N_8883);
nand UO_633 (O_633,N_6117,N_8006);
and UO_634 (O_634,N_9495,N_5685);
and UO_635 (O_635,N_8603,N_6505);
nand UO_636 (O_636,N_5470,N_9310);
and UO_637 (O_637,N_7453,N_7181);
or UO_638 (O_638,N_9810,N_6346);
or UO_639 (O_639,N_8751,N_8107);
and UO_640 (O_640,N_6176,N_8173);
or UO_641 (O_641,N_6431,N_9951);
nor UO_642 (O_642,N_7310,N_9025);
nand UO_643 (O_643,N_7618,N_9687);
or UO_644 (O_644,N_7422,N_9881);
and UO_645 (O_645,N_6480,N_8977);
or UO_646 (O_646,N_7821,N_6481);
or UO_647 (O_647,N_5406,N_5692);
and UO_648 (O_648,N_9943,N_8594);
nand UO_649 (O_649,N_6542,N_5883);
and UO_650 (O_650,N_9508,N_5075);
xnor UO_651 (O_651,N_8351,N_5391);
nand UO_652 (O_652,N_8165,N_5513);
and UO_653 (O_653,N_9075,N_8182);
and UO_654 (O_654,N_6667,N_6933);
nand UO_655 (O_655,N_9285,N_8703);
nand UO_656 (O_656,N_8832,N_8046);
or UO_657 (O_657,N_6835,N_6673);
and UO_658 (O_658,N_7990,N_8437);
or UO_659 (O_659,N_6324,N_7939);
nor UO_660 (O_660,N_7367,N_8320);
xor UO_661 (O_661,N_8410,N_5643);
or UO_662 (O_662,N_5210,N_6038);
nand UO_663 (O_663,N_7141,N_5200);
or UO_664 (O_664,N_7226,N_8598);
and UO_665 (O_665,N_5360,N_6025);
and UO_666 (O_666,N_7139,N_6983);
or UO_667 (O_667,N_6839,N_5693);
nand UO_668 (O_668,N_9771,N_8760);
or UO_669 (O_669,N_7802,N_5980);
and UO_670 (O_670,N_8585,N_9589);
nor UO_671 (O_671,N_5209,N_5430);
nor UO_672 (O_672,N_6459,N_5106);
nand UO_673 (O_673,N_5930,N_8648);
nor UO_674 (O_674,N_9979,N_7142);
nand UO_675 (O_675,N_9357,N_6936);
nand UO_676 (O_676,N_5151,N_9898);
or UO_677 (O_677,N_8124,N_9101);
or UO_678 (O_678,N_9611,N_7906);
nand UO_679 (O_679,N_5498,N_6434);
and UO_680 (O_680,N_7202,N_5814);
nand UO_681 (O_681,N_9436,N_8889);
or UO_682 (O_682,N_5186,N_8851);
or UO_683 (O_683,N_8794,N_6187);
nand UO_684 (O_684,N_9761,N_5565);
nand UO_685 (O_685,N_5582,N_9383);
or UO_686 (O_686,N_9912,N_9560);
nand UO_687 (O_687,N_8405,N_5490);
or UO_688 (O_688,N_6443,N_9948);
or UO_689 (O_689,N_7308,N_7455);
and UO_690 (O_690,N_6288,N_9368);
or UO_691 (O_691,N_7526,N_5435);
nor UO_692 (O_692,N_8230,N_7093);
and UO_693 (O_693,N_5561,N_8357);
and UO_694 (O_694,N_8157,N_7340);
nand UO_695 (O_695,N_7413,N_9442);
nand UO_696 (O_696,N_6769,N_8492);
nand UO_697 (O_697,N_6956,N_6005);
nor UO_698 (O_698,N_9515,N_6314);
nor UO_699 (O_699,N_7720,N_9312);
nand UO_700 (O_700,N_5831,N_8529);
and UO_701 (O_701,N_6184,N_9464);
and UO_702 (O_702,N_5267,N_7411);
nand UO_703 (O_703,N_5038,N_9189);
nand UO_704 (O_704,N_6375,N_9389);
and UO_705 (O_705,N_5954,N_9336);
nor UO_706 (O_706,N_7843,N_5619);
or UO_707 (O_707,N_6924,N_5759);
nand UO_708 (O_708,N_9684,N_6935);
nor UO_709 (O_709,N_7281,N_9795);
nand UO_710 (O_710,N_7966,N_5269);
or UO_711 (O_711,N_6541,N_6079);
or UO_712 (O_712,N_8658,N_6737);
and UO_713 (O_713,N_6682,N_5255);
and UO_714 (O_714,N_8491,N_9160);
and UO_715 (O_715,N_7361,N_9000);
or UO_716 (O_716,N_6930,N_9556);
or UO_717 (O_717,N_9542,N_7348);
nor UO_718 (O_718,N_9685,N_8856);
or UO_719 (O_719,N_9678,N_6863);
and UO_720 (O_720,N_6352,N_5205);
and UO_721 (O_721,N_8915,N_8697);
nor UO_722 (O_722,N_9027,N_7408);
or UO_723 (O_723,N_9417,N_7136);
nor UO_724 (O_724,N_8507,N_7376);
nor UO_725 (O_725,N_9435,N_8693);
xnor UO_726 (O_726,N_5313,N_8681);
nand UO_727 (O_727,N_5606,N_5334);
nor UO_728 (O_728,N_6148,N_6175);
and UO_729 (O_729,N_6946,N_5668);
or UO_730 (O_730,N_9320,N_5772);
and UO_731 (O_731,N_8892,N_9268);
nor UO_732 (O_732,N_6641,N_7912);
nand UO_733 (O_733,N_5173,N_7952);
nor UO_734 (O_734,N_6414,N_9195);
nor UO_735 (O_735,N_6268,N_7721);
nand UO_736 (O_736,N_7707,N_8031);
and UO_737 (O_737,N_7710,N_9069);
nor UO_738 (O_738,N_8348,N_7857);
nor UO_739 (O_739,N_9440,N_8096);
and UO_740 (O_740,N_6325,N_8814);
or UO_741 (O_741,N_8316,N_5184);
nand UO_742 (O_742,N_5945,N_7460);
and UO_743 (O_743,N_7846,N_7831);
nor UO_744 (O_744,N_9787,N_8488);
and UO_745 (O_745,N_5330,N_7341);
nor UO_746 (O_746,N_5074,N_5906);
or UO_747 (O_747,N_8933,N_9133);
and UO_748 (O_748,N_9801,N_6551);
and UO_749 (O_749,N_8949,N_7863);
nand UO_750 (O_750,N_9036,N_5613);
nand UO_751 (O_751,N_7293,N_6582);
nor UO_752 (O_752,N_9323,N_6349);
nand UO_753 (O_753,N_6775,N_6050);
or UO_754 (O_754,N_5202,N_8312);
nor UO_755 (O_755,N_8269,N_8271);
xnor UO_756 (O_756,N_6410,N_6743);
nor UO_757 (O_757,N_9270,N_5603);
and UO_758 (O_758,N_9845,N_9504);
or UO_759 (O_759,N_9043,N_8427);
nor UO_760 (O_760,N_6590,N_5834);
xnor UO_761 (O_761,N_6208,N_5368);
nor UO_762 (O_762,N_8042,N_7849);
xnor UO_763 (O_763,N_7428,N_7668);
nand UO_764 (O_764,N_5123,N_6361);
nor UO_765 (O_765,N_8788,N_9615);
nor UO_766 (O_766,N_5557,N_8037);
nand UO_767 (O_767,N_8463,N_5404);
or UO_768 (O_768,N_7836,N_9478);
or UO_769 (O_769,N_8205,N_5010);
nand UO_770 (O_770,N_7075,N_8308);
nor UO_771 (O_771,N_7366,N_6326);
nand UO_772 (O_772,N_6156,N_9576);
and UO_773 (O_773,N_5223,N_7633);
nor UO_774 (O_774,N_6837,N_6271);
nand UO_775 (O_775,N_7223,N_7770);
nor UO_776 (O_776,N_8686,N_8580);
or UO_777 (O_777,N_6626,N_7510);
or UO_778 (O_778,N_8531,N_9186);
or UO_779 (O_779,N_7280,N_7993);
nor UO_780 (O_780,N_6959,N_6347);
nand UO_781 (O_781,N_7386,N_7437);
and UO_782 (O_782,N_8627,N_7553);
nand UO_783 (O_783,N_8638,N_9914);
or UO_784 (O_784,N_6018,N_8336);
nand UO_785 (O_785,N_5199,N_7430);
or UO_786 (O_786,N_8518,N_6976);
or UO_787 (O_787,N_8030,N_9145);
nor UO_788 (O_788,N_5740,N_7535);
or UO_789 (O_789,N_8976,N_5976);
nand UO_790 (O_790,N_6571,N_5566);
or UO_791 (O_791,N_6064,N_9588);
nand UO_792 (O_792,N_8158,N_8071);
and UO_793 (O_793,N_5447,N_5358);
nor UO_794 (O_794,N_5340,N_9812);
and UO_795 (O_795,N_9010,N_6211);
nor UO_796 (O_796,N_6063,N_8039);
nor UO_797 (O_797,N_8973,N_6379);
nand UO_798 (O_798,N_7452,N_8216);
or UO_799 (O_799,N_7294,N_6399);
nand UO_800 (O_800,N_8282,N_8360);
nand UO_801 (O_801,N_5093,N_7832);
or UO_802 (O_802,N_9938,N_5936);
nor UO_803 (O_803,N_6655,N_7373);
and UO_804 (O_804,N_5686,N_6329);
nand UO_805 (O_805,N_7779,N_9665);
nor UO_806 (O_806,N_5251,N_7552);
and UO_807 (O_807,N_9532,N_9466);
nand UO_808 (O_808,N_9792,N_5734);
and UO_809 (O_809,N_6107,N_8558);
or UO_810 (O_810,N_9064,N_7380);
and UO_811 (O_811,N_6721,N_7016);
xnor UO_812 (O_812,N_7043,N_9005);
and UO_813 (O_813,N_8745,N_6982);
or UO_814 (O_814,N_8483,N_5682);
and UO_815 (O_815,N_8432,N_5306);
or UO_816 (O_816,N_5959,N_7222);
xnor UO_817 (O_817,N_5983,N_7590);
and UO_818 (O_818,N_7941,N_7229);
and UO_819 (O_819,N_6204,N_7300);
nor UO_820 (O_820,N_5426,N_7539);
nor UO_821 (O_821,N_7465,N_5644);
and UO_822 (O_822,N_6696,N_6922);
nor UO_823 (O_823,N_5493,N_7155);
nand UO_824 (O_824,N_7743,N_8526);
or UO_825 (O_825,N_8849,N_6037);
nor UO_826 (O_826,N_8628,N_5120);
and UO_827 (O_827,N_6921,N_7874);
nand UO_828 (O_828,N_5896,N_5083);
xor UO_829 (O_829,N_6011,N_9074);
nor UO_830 (O_830,N_5339,N_8121);
nand UO_831 (O_831,N_6759,N_5900);
nand UO_832 (O_832,N_6382,N_7345);
nor UO_833 (O_833,N_7055,N_6609);
or UO_834 (O_834,N_6818,N_8460);
and UO_835 (O_835,N_7159,N_8682);
nor UO_836 (O_836,N_8841,N_6989);
and UO_837 (O_837,N_5187,N_7827);
or UO_838 (O_838,N_9941,N_8217);
nand UO_839 (O_839,N_6237,N_6424);
or UO_840 (O_840,N_5364,N_5821);
nand UO_841 (O_841,N_5328,N_8313);
xor UO_842 (O_842,N_8567,N_5194);
nor UO_843 (O_843,N_6819,N_5317);
or UO_844 (O_844,N_6102,N_8361);
nor UO_845 (O_845,N_6778,N_6492);
or UO_846 (O_846,N_6852,N_8462);
or UO_847 (O_847,N_9757,N_6926);
and UO_848 (O_848,N_6442,N_8669);
and UO_849 (O_849,N_7506,N_9067);
nand UO_850 (O_850,N_5448,N_6581);
and UO_851 (O_851,N_6763,N_6171);
nand UO_852 (O_852,N_8495,N_8515);
and UO_853 (O_853,N_6162,N_7902);
nor UO_854 (O_854,N_8455,N_9349);
or UO_855 (O_855,N_6302,N_5833);
or UO_856 (O_856,N_6987,N_8450);
and UO_857 (O_857,N_8836,N_7671);
nor UO_858 (O_858,N_9254,N_5344);
or UO_859 (O_859,N_9638,N_8517);
nor UO_860 (O_860,N_6157,N_6957);
or UO_861 (O_861,N_9058,N_6633);
or UO_862 (O_862,N_9282,N_9973);
nand UO_863 (O_863,N_5880,N_7248);
nand UO_864 (O_864,N_8868,N_8141);
and UO_865 (O_865,N_8589,N_5296);
or UO_866 (O_866,N_9626,N_9469);
and UO_867 (O_867,N_6490,N_9348);
xor UO_868 (O_868,N_6218,N_8029);
nand UO_869 (O_869,N_5449,N_6532);
xnor UO_870 (O_870,N_6047,N_9096);
nor UO_871 (O_871,N_8787,N_8416);
nor UO_872 (O_872,N_7524,N_6448);
nand UO_873 (O_873,N_7646,N_8683);
nand UO_874 (O_874,N_6762,N_6416);
or UO_875 (O_875,N_8521,N_5003);
and UO_876 (O_876,N_8137,N_5627);
or UO_877 (O_877,N_9266,N_7233);
or UO_878 (O_878,N_5363,N_5841);
nor UO_879 (O_879,N_9293,N_7284);
or UO_880 (O_880,N_5088,N_6877);
nor UO_881 (O_881,N_8149,N_7704);
nand UO_882 (O_882,N_5367,N_8906);
nor UO_883 (O_883,N_7208,N_6372);
and UO_884 (O_884,N_9078,N_7304);
nor UO_885 (O_885,N_7276,N_9387);
or UO_886 (O_886,N_6397,N_8299);
nor UO_887 (O_887,N_9926,N_9301);
nor UO_888 (O_888,N_6727,N_9895);
nor UO_889 (O_889,N_7274,N_7204);
or UO_890 (O_890,N_5411,N_8572);
and UO_891 (O_891,N_7564,N_8705);
or UO_892 (O_892,N_7423,N_8481);
or UO_893 (O_893,N_9049,N_8101);
nand UO_894 (O_894,N_7953,N_9755);
or UO_895 (O_895,N_6518,N_5104);
and UO_896 (O_896,N_9967,N_6088);
or UO_897 (O_897,N_9731,N_6464);
or UO_898 (O_898,N_8203,N_9376);
nand UO_899 (O_899,N_7631,N_5589);
and UO_900 (O_900,N_7264,N_5903);
nor UO_901 (O_901,N_8934,N_7343);
nand UO_902 (O_902,N_5369,N_6513);
and UO_903 (O_903,N_8401,N_6306);
xor UO_904 (O_904,N_5620,N_9562);
or UO_905 (O_905,N_5915,N_6152);
nor UO_906 (O_906,N_7736,N_8560);
nand UO_907 (O_907,N_9821,N_8189);
nor UO_908 (O_908,N_8260,N_8415);
and UO_909 (O_909,N_5514,N_7419);
and UO_910 (O_910,N_6514,N_6731);
or UO_911 (O_911,N_5073,N_6566);
and UO_912 (O_912,N_5472,N_9797);
or UO_913 (O_913,N_9419,N_5749);
and UO_914 (O_914,N_6371,N_9380);
nand UO_915 (O_915,N_7147,N_8709);
nand UO_916 (O_916,N_8746,N_6745);
nand UO_917 (O_917,N_5341,N_7682);
nand UO_918 (O_918,N_7508,N_9509);
or UO_919 (O_919,N_9837,N_5684);
nor UO_920 (O_920,N_8206,N_5568);
nor UO_921 (O_921,N_6342,N_7883);
and UO_922 (O_922,N_8678,N_8942);
or UO_923 (O_923,N_8402,N_8364);
and UO_924 (O_924,N_7224,N_5193);
nor UO_925 (O_925,N_8876,N_8242);
or UO_926 (O_926,N_8430,N_7873);
and UO_927 (O_927,N_7839,N_8733);
and UO_928 (O_928,N_8930,N_8244);
or UO_929 (O_929,N_6900,N_5544);
or UO_930 (O_930,N_7307,N_9649);
or UO_931 (O_931,N_7745,N_8707);
and UO_932 (O_932,N_7117,N_6880);
or UO_933 (O_933,N_5060,N_7412);
and UO_934 (O_934,N_5554,N_6907);
and UO_935 (O_935,N_8637,N_9234);
and UO_936 (O_936,N_8382,N_5891);
or UO_937 (O_937,N_7353,N_9460);
or UO_938 (O_938,N_7834,N_7490);
or UO_939 (O_939,N_7722,N_6865);
or UO_940 (O_940,N_5183,N_7724);
and UO_941 (O_941,N_7271,N_6538);
or UO_942 (O_942,N_9115,N_8169);
and UO_943 (O_943,N_8001,N_5311);
and UO_944 (O_944,N_6535,N_7194);
and UO_945 (O_945,N_8713,N_9769);
nand UO_946 (O_946,N_9322,N_8700);
nand UO_947 (O_947,N_6084,N_8197);
nand UO_948 (O_948,N_9300,N_9984);
and UO_949 (O_949,N_9211,N_9403);
nor UO_950 (O_950,N_7586,N_7666);
xor UO_951 (O_951,N_7861,N_7869);
nand UO_952 (O_952,N_8383,N_9603);
nor UO_953 (O_953,N_5189,N_7180);
or UO_954 (O_954,N_8160,N_8486);
nand UO_955 (O_955,N_7228,N_5715);
nor UO_956 (O_956,N_6087,N_8421);
or UO_957 (O_957,N_7587,N_5154);
or UO_958 (O_958,N_8909,N_8399);
or UO_959 (O_959,N_6036,N_7240);
or UO_960 (O_960,N_9112,N_8633);
and UO_961 (O_961,N_6606,N_5172);
or UO_962 (O_962,N_9287,N_7459);
nor UO_963 (O_963,N_7400,N_6294);
or UO_964 (O_964,N_6254,N_6643);
or UO_965 (O_965,N_7176,N_8859);
nand UO_966 (O_966,N_8143,N_8431);
nor UO_967 (O_967,N_6630,N_7216);
xor UO_968 (O_968,N_5788,N_5845);
nand UO_969 (O_969,N_5355,N_8334);
xor UO_970 (O_970,N_5286,N_9955);
nor UO_971 (O_971,N_8028,N_8711);
or UO_972 (O_972,N_6479,N_5198);
nand UO_973 (O_973,N_5037,N_7692);
nor UO_974 (O_974,N_6021,N_8626);
or UO_975 (O_975,N_7548,N_7503);
and UO_976 (O_976,N_9210,N_6530);
and UO_977 (O_977,N_6419,N_5035);
nand UO_978 (O_978,N_7741,N_6423);
and UO_979 (O_979,N_6452,N_7574);
or UO_980 (O_980,N_9317,N_9123);
and UO_981 (O_981,N_8307,N_8617);
and UO_982 (O_982,N_6961,N_5912);
or UO_983 (O_983,N_5562,N_8864);
nor UO_984 (O_984,N_8082,N_6124);
nand UO_985 (O_985,N_6781,N_8412);
nand UO_986 (O_986,N_7523,N_9636);
or UO_987 (O_987,N_5564,N_6247);
nor UO_988 (O_988,N_8660,N_5132);
nand UO_989 (O_989,N_6450,N_7640);
or UO_990 (O_990,N_6274,N_6675);
nor UO_991 (O_991,N_8761,N_6144);
and UO_992 (O_992,N_9144,N_5117);
nor UO_993 (O_993,N_7137,N_8005);
nor UO_994 (O_994,N_5507,N_7899);
nor UO_995 (O_995,N_7090,N_9013);
nor UO_996 (O_996,N_9897,N_9271);
nand UO_997 (O_997,N_7812,N_5515);
nand UO_998 (O_998,N_8609,N_6608);
nor UO_999 (O_999,N_9978,N_7385);
and UO_1000 (O_1000,N_5233,N_9477);
nor UO_1001 (O_1001,N_7717,N_8356);
or UO_1002 (O_1002,N_8961,N_5745);
nand UO_1003 (O_1003,N_5840,N_6301);
nand UO_1004 (O_1004,N_6993,N_7866);
or UO_1005 (O_1005,N_9612,N_5145);
or UO_1006 (O_1006,N_7709,N_9586);
or UO_1007 (O_1007,N_9480,N_7886);
nand UO_1008 (O_1008,N_8895,N_8890);
nor UO_1009 (O_1009,N_5948,N_5025);
or UO_1010 (O_1010,N_9428,N_6201);
nor UO_1011 (O_1011,N_9467,N_9468);
nor UO_1012 (O_1012,N_6562,N_7642);
and UO_1013 (O_1013,N_7406,N_8513);
nand UO_1014 (O_1014,N_8525,N_8664);
nor UO_1015 (O_1015,N_6753,N_7238);
or UO_1016 (O_1016,N_5116,N_9758);
or UO_1017 (O_1017,N_7513,N_6735);
nor UO_1018 (O_1018,N_7481,N_7533);
and UO_1019 (O_1019,N_5947,N_8861);
nor UO_1020 (O_1020,N_8969,N_6938);
nand UO_1021 (O_1021,N_8673,N_9693);
nor UO_1022 (O_1022,N_8903,N_7095);
nand UO_1023 (O_1023,N_8438,N_6996);
nor UO_1024 (O_1024,N_7475,N_9632);
and UO_1025 (O_1025,N_5464,N_8118);
and UO_1026 (O_1026,N_7381,N_6256);
and UO_1027 (O_1027,N_6285,N_5837);
and UO_1028 (O_1028,N_6913,N_7173);
nand UO_1029 (O_1029,N_8300,N_9505);
or UO_1030 (O_1030,N_5445,N_7816);
and UO_1031 (O_1031,N_9331,N_7758);
and UO_1032 (O_1032,N_9700,N_8340);
and UO_1033 (O_1033,N_6406,N_7833);
nand UO_1034 (O_1034,N_8498,N_9646);
or UO_1035 (O_1035,N_9260,N_5234);
nor UO_1036 (O_1036,N_8716,N_7734);
nor UO_1037 (O_1037,N_5807,N_6293);
or UO_1038 (O_1038,N_6618,N_9807);
or UO_1039 (O_1039,N_9584,N_6122);
nand UO_1040 (O_1040,N_5389,N_5935);
or UO_1041 (O_1041,N_5385,N_9223);
or UO_1042 (O_1042,N_6421,N_8132);
or UO_1043 (O_1043,N_6312,N_6457);
nand UO_1044 (O_1044,N_5854,N_5497);
nor UO_1045 (O_1045,N_7604,N_5728);
nor UO_1046 (O_1046,N_6467,N_6280);
nor UO_1047 (O_1047,N_6061,N_9286);
nand UO_1048 (O_1048,N_7225,N_8622);
nand UO_1049 (O_1049,N_6950,N_6845);
and UO_1050 (O_1050,N_9255,N_6943);
and UO_1051 (O_1051,N_8918,N_7759);
and UO_1052 (O_1052,N_5461,N_5032);
nand UO_1053 (O_1053,N_6842,N_9384);
nand UO_1054 (O_1054,N_6822,N_9803);
and UO_1055 (O_1055,N_8687,N_7537);
and UO_1056 (O_1056,N_7156,N_6966);
nor UO_1057 (O_1057,N_6962,N_6449);
xor UO_1058 (O_1058,N_5846,N_8426);
nor UO_1059 (O_1059,N_9995,N_8407);
nand UO_1060 (O_1060,N_9695,N_6898);
nor UO_1061 (O_1061,N_9298,N_6874);
nor UO_1062 (O_1062,N_7609,N_5196);
nand UO_1063 (O_1063,N_6477,N_8991);
nor UO_1064 (O_1064,N_9537,N_8737);
and UO_1065 (O_1065,N_8007,N_7583);
nand UO_1066 (O_1066,N_9901,N_8774);
or UO_1067 (O_1067,N_7519,N_8588);
nand UO_1068 (O_1068,N_9566,N_5645);
and UO_1069 (O_1069,N_7661,N_7887);
nor UO_1070 (O_1070,N_6563,N_7674);
or UO_1071 (O_1071,N_6336,N_6984);
nor UO_1072 (O_1072,N_7536,N_5999);
nor UO_1073 (O_1073,N_8586,N_9592);
nor UO_1074 (O_1074,N_9315,N_5454);
and UO_1075 (O_1075,N_5622,N_6885);
nor UO_1076 (O_1076,N_7505,N_5392);
and UO_1077 (O_1077,N_8305,N_7502);
or UO_1078 (O_1078,N_5427,N_6998);
or UO_1079 (O_1079,N_7872,N_9608);
or UO_1080 (O_1080,N_9354,N_6804);
xor UO_1081 (O_1081,N_5708,N_9054);
nor UO_1082 (O_1082,N_9215,N_7542);
nand UO_1083 (O_1083,N_6291,N_9557);
xor UO_1084 (O_1084,N_6619,N_6173);
nand UO_1085 (O_1085,N_5488,N_8411);
nor UO_1086 (O_1086,N_6275,N_5401);
nor UO_1087 (O_1087,N_6078,N_5783);
nor UO_1088 (O_1088,N_9292,N_7031);
or UO_1089 (O_1089,N_8552,N_6094);
nand UO_1090 (O_1090,N_6820,N_9748);
or UO_1091 (O_1091,N_8243,N_7089);
or UO_1092 (O_1092,N_5535,N_8853);
nor UO_1093 (O_1093,N_7774,N_5335);
or UO_1094 (O_1094,N_5552,N_8816);
nor UO_1095 (O_1095,N_7382,N_9644);
or UO_1096 (O_1096,N_8229,N_5972);
nor UO_1097 (O_1097,N_6019,N_8235);
nand UO_1098 (O_1098,N_9935,N_7077);
nor UO_1099 (O_1099,N_5665,N_7688);
xor UO_1100 (O_1100,N_9489,N_5547);
nor UO_1101 (O_1101,N_7992,N_8436);
and UO_1102 (O_1102,N_6999,N_5005);
or UO_1103 (O_1103,N_9850,N_7922);
or UO_1104 (O_1104,N_5140,N_9325);
and UO_1105 (O_1105,N_8179,N_9341);
or UO_1106 (O_1106,N_5034,N_7168);
or UO_1107 (O_1107,N_6534,N_8176);
or UO_1108 (O_1108,N_9535,N_5410);
nand UO_1109 (O_1109,N_6121,N_8089);
nand UO_1110 (O_1110,N_7330,N_6917);
and UO_1111 (O_1111,N_7606,N_5701);
or UO_1112 (O_1112,N_9621,N_8763);
or UO_1113 (O_1113,N_6817,N_5351);
or UO_1114 (O_1114,N_6733,N_8544);
nand UO_1115 (O_1115,N_5433,N_7888);
nand UO_1116 (O_1116,N_7737,N_7603);
nor UO_1117 (O_1117,N_8477,N_9490);
and UO_1118 (O_1118,N_8604,N_7712);
nand UO_1119 (O_1119,N_9544,N_8616);
and UO_1120 (O_1120,N_8190,N_9217);
nor UO_1121 (O_1121,N_5291,N_8068);
or UO_1122 (O_1122,N_8523,N_9253);
nor UO_1123 (O_1123,N_8470,N_7934);
nand UO_1124 (O_1124,N_6871,N_7243);
and UO_1125 (O_1125,N_9030,N_8530);
nor UO_1126 (O_1126,N_6886,N_5825);
and UO_1127 (O_1127,N_7715,N_6790);
and UO_1128 (O_1128,N_5905,N_6722);
or UO_1129 (O_1129,N_5892,N_8955);
xor UO_1130 (O_1130,N_5605,N_8102);
and UO_1131 (O_1131,N_7670,N_8127);
nand UO_1132 (O_1132,N_8180,N_9640);
and UO_1133 (O_1133,N_6296,N_6153);
nor UO_1134 (O_1134,N_7351,N_7575);
nor UO_1135 (O_1135,N_7509,N_9077);
or UO_1136 (O_1136,N_9364,N_8784);
xnor UO_1137 (O_1137,N_5188,N_9121);
nand UO_1138 (O_1138,N_8475,N_8199);
or UO_1139 (O_1139,N_8796,N_6488);
or UO_1140 (O_1140,N_7210,N_6891);
nor UO_1141 (O_1141,N_5271,N_7114);
or UO_1142 (O_1142,N_8718,N_8070);
nand UO_1143 (O_1143,N_8449,N_5950);
nand UO_1144 (O_1144,N_9909,N_6170);
nand UO_1145 (O_1145,N_9438,N_9129);
nor UO_1146 (O_1146,N_7657,N_5812);
and UO_1147 (O_1147,N_9798,N_8429);
nor UO_1148 (O_1148,N_7331,N_6207);
nor UO_1149 (O_1149,N_6206,N_9288);
nor UO_1150 (O_1150,N_8540,N_6681);
nor UO_1151 (O_1151,N_5952,N_8109);
and UO_1152 (O_1152,N_5413,N_8413);
nor UO_1153 (O_1153,N_7085,N_8209);
nor UO_1154 (O_1154,N_9202,N_6091);
or UO_1155 (O_1155,N_5851,N_7835);
and UO_1156 (O_1156,N_5676,N_6780);
and UO_1157 (O_1157,N_5732,N_9281);
and UO_1158 (O_1158,N_9936,N_6586);
nor UO_1159 (O_1159,N_7917,N_9024);
and UO_1160 (O_1160,N_8509,N_6783);
nor UO_1161 (O_1161,N_9248,N_8075);
nand UO_1162 (O_1162,N_5793,N_8387);
and UO_1163 (O_1163,N_5864,N_5465);
nor UO_1164 (O_1164,N_9426,N_9749);
or UO_1165 (O_1165,N_5349,N_6893);
and UO_1166 (O_1166,N_5695,N_8339);
or UO_1167 (O_1167,N_8750,N_5960);
nand UO_1168 (O_1168,N_8066,N_8652);
nand UO_1169 (O_1169,N_5484,N_7528);
and UO_1170 (O_1170,N_5203,N_7842);
and UO_1171 (O_1171,N_5181,N_5592);
nand UO_1172 (O_1172,N_7384,N_6694);
nor UO_1173 (O_1173,N_8710,N_5874);
nand UO_1174 (O_1174,N_6858,N_6903);
or UO_1175 (O_1175,N_6602,N_7319);
or UO_1176 (O_1176,N_7215,N_5500);
nor UO_1177 (O_1177,N_7131,N_9214);
nor UO_1178 (O_1178,N_8822,N_5325);
nand UO_1179 (O_1179,N_7844,N_7496);
nand UO_1180 (O_1180,N_7035,N_9764);
and UO_1181 (O_1181,N_8884,N_7776);
nor UO_1182 (O_1182,N_6454,N_5593);
and UO_1183 (O_1183,N_7246,N_5920);
nor UO_1184 (O_1184,N_9022,N_5451);
nand UO_1185 (O_1185,N_9949,N_8406);
nand UO_1186 (O_1186,N_7442,N_7479);
nor UO_1187 (O_1187,N_7150,N_8317);
nor UO_1188 (O_1188,N_8219,N_6407);
nor UO_1189 (O_1189,N_7057,N_8016);
or UO_1190 (O_1190,N_9087,N_9111);
nand UO_1191 (O_1191,N_5944,N_5395);
nand UO_1192 (O_1192,N_8390,N_8270);
or UO_1193 (O_1193,N_9548,N_8418);
nor UO_1194 (O_1194,N_8392,N_5023);
nor UO_1195 (O_1195,N_7418,N_9816);
nand UO_1196 (O_1196,N_7425,N_5398);
nand UO_1197 (O_1197,N_9456,N_6143);
or UO_1198 (O_1198,N_6227,N_9805);
xor UO_1199 (O_1199,N_9836,N_8211);
nand UO_1200 (O_1200,N_5979,N_5354);
nor UO_1201 (O_1201,N_9602,N_5843);
or UO_1202 (O_1202,N_7221,N_7177);
and UO_1203 (O_1203,N_9008,N_6547);
nand UO_1204 (O_1204,N_8980,N_5670);
and UO_1205 (O_1205,N_6213,N_9451);
and UO_1206 (O_1206,N_5524,N_8067);
nand UO_1207 (O_1207,N_9579,N_6297);
and UO_1208 (O_1208,N_8688,N_6828);
nand UO_1209 (O_1209,N_5873,N_6315);
nand UO_1210 (O_1210,N_9410,N_8164);
nand UO_1211 (O_1211,N_5278,N_6848);
and UO_1212 (O_1212,N_9140,N_8939);
nand UO_1213 (O_1213,N_9727,N_9770);
or UO_1214 (O_1214,N_7976,N_8232);
xnor UO_1215 (O_1215,N_6764,N_5284);
xor UO_1216 (O_1216,N_5266,N_6919);
nand UO_1217 (O_1217,N_7708,N_7122);
nand UO_1218 (O_1218,N_5984,N_8613);
nor UO_1219 (O_1219,N_5806,N_6585);
nor UO_1220 (O_1220,N_8181,N_5409);
and UO_1221 (O_1221,N_8106,N_6995);
and UO_1222 (O_1222,N_9962,N_5437);
and UO_1223 (O_1223,N_6150,N_7771);
and UO_1224 (O_1224,N_8650,N_7363);
nand UO_1225 (O_1225,N_5790,N_7963);
or UO_1226 (O_1226,N_8860,N_8591);
nor UO_1227 (O_1227,N_5650,N_8065);
nor UO_1228 (O_1228,N_7986,N_7617);
nand UO_1229 (O_1229,N_9639,N_8695);
and UO_1230 (O_1230,N_5331,N_9405);
nand UO_1231 (O_1231,N_5137,N_8542);
nand UO_1232 (O_1232,N_5757,N_7473);
and UO_1233 (O_1233,N_6389,N_7108);
or UO_1234 (O_1234,N_5533,N_9014);
or UO_1235 (O_1235,N_7959,N_8601);
or UO_1236 (O_1236,N_7768,N_8756);
nor UO_1237 (O_1237,N_5910,N_5136);
nor UO_1238 (O_1238,N_9784,N_7326);
and UO_1239 (O_1239,N_5263,N_7052);
nor UO_1240 (O_1240,N_7493,N_5658);
nand UO_1241 (O_1241,N_5262,N_5176);
and UO_1242 (O_1242,N_6415,N_6113);
nor UO_1243 (O_1243,N_9088,N_6908);
or UO_1244 (O_1244,N_6086,N_9316);
and UO_1245 (O_1245,N_6855,N_6283);
or UO_1246 (O_1246,N_7483,N_9860);
or UO_1247 (O_1247,N_5382,N_5671);
nor UO_1248 (O_1248,N_9127,N_7165);
nand UO_1249 (O_1249,N_6768,N_9732);
or UO_1250 (O_1250,N_5327,N_8869);
or UO_1251 (O_1251,N_9924,N_6309);
or UO_1252 (O_1252,N_6703,N_8302);
and UO_1253 (O_1253,N_9171,N_8023);
nor UO_1254 (O_1254,N_6508,N_6220);
nand UO_1255 (O_1255,N_6528,N_8015);
or UO_1256 (O_1256,N_5163,N_8002);
and UO_1257 (O_1257,N_7897,N_5321);
nor UO_1258 (O_1258,N_7257,N_9558);
nor UO_1259 (O_1259,N_9741,N_9113);
nor UO_1260 (O_1260,N_5614,N_8054);
and UO_1261 (O_1261,N_5139,N_9150);
or UO_1262 (O_1262,N_9650,N_5962);
or UO_1263 (O_1263,N_6110,N_9050);
nand UO_1264 (O_1264,N_5733,N_9875);
or UO_1265 (O_1265,N_8090,N_6221);
xnor UO_1266 (O_1266,N_7254,N_5689);
or UO_1267 (O_1267,N_9564,N_5352);
nor UO_1268 (O_1268,N_6882,N_8779);
nand UO_1269 (O_1269,N_8893,N_6931);
nor UO_1270 (O_1270,N_8621,N_9864);
nor UO_1271 (O_1271,N_9134,N_5909);
nand UO_1272 (O_1272,N_6120,N_9859);
or UO_1273 (O_1273,N_9691,N_7071);
or UO_1274 (O_1274,N_7855,N_9272);
and UO_1275 (O_1275,N_9385,N_5304);
or UO_1276 (O_1276,N_7059,N_7878);
or UO_1277 (O_1277,N_5717,N_8280);
nand UO_1278 (O_1278,N_9871,N_5610);
nor UO_1279 (O_1279,N_5346,N_9595);
nand UO_1280 (O_1280,N_5347,N_7410);
or UO_1281 (O_1281,N_7480,N_7291);
and UO_1282 (O_1282,N_7039,N_9867);
nand UO_1283 (O_1283,N_9230,N_5722);
and UO_1284 (O_1284,N_7462,N_7576);
nor UO_1285 (O_1285,N_8960,N_7608);
nor UO_1286 (O_1286,N_8378,N_8852);
nand UO_1287 (O_1287,N_8192,N_8924);
nand UO_1288 (O_1288,N_6368,N_9607);
or UO_1289 (O_1289,N_7009,N_9843);
nand UO_1290 (O_1290,N_6773,N_5902);
nor UO_1291 (O_1291,N_9033,N_5170);
nor UO_1292 (O_1292,N_5105,N_7432);
and UO_1293 (O_1293,N_7468,N_6793);
nand UO_1294 (O_1294,N_9681,N_6106);
nand UO_1295 (O_1295,N_8634,N_7620);
nor UO_1296 (O_1296,N_8440,N_9580);
nor UO_1297 (O_1297,N_5118,N_5828);
and UO_1298 (O_1298,N_7320,N_6048);
nand UO_1299 (O_1299,N_5545,N_6755);
or UO_1300 (O_1300,N_7497,N_9046);
or UO_1301 (O_1301,N_8093,N_9513);
nor UO_1302 (O_1302,N_7357,N_7121);
or UO_1303 (O_1303,N_5739,N_9934);
nor UO_1304 (O_1304,N_5782,N_9596);
nor UO_1305 (O_1305,N_7925,N_6503);
xor UO_1306 (O_1306,N_8982,N_8671);
nor UO_1307 (O_1307,N_8330,N_5907);
nand UO_1308 (O_1308,N_5626,N_7286);
and UO_1309 (O_1309,N_7970,N_9007);
and UO_1310 (O_1310,N_8974,N_5534);
and UO_1311 (O_1311,N_5125,N_6625);
or UO_1312 (O_1312,N_9613,N_7190);
and UO_1313 (O_1313,N_5253,N_5779);
nand UO_1314 (O_1314,N_5495,N_6504);
and UO_1315 (O_1315,N_9999,N_8020);
or UO_1316 (O_1316,N_8263,N_8482);
nand UO_1317 (O_1317,N_6794,N_7022);
and UO_1318 (O_1318,N_7026,N_6066);
and UO_1319 (O_1319,N_9124,N_7914);
nor UO_1320 (O_1320,N_5990,N_6981);
or UO_1321 (O_1321,N_5526,N_9672);
nor UO_1322 (O_1322,N_7198,N_5953);
and UO_1323 (O_1323,N_5869,N_8685);
nand UO_1324 (O_1324,N_5742,N_8112);
nand UO_1325 (O_1325,N_7738,N_9415);
and UO_1326 (O_1326,N_6390,N_8139);
nand UO_1327 (O_1327,N_6807,N_7398);
and UO_1328 (O_1328,N_7971,N_7445);
nor UO_1329 (O_1329,N_5633,N_5337);
or UO_1330 (O_1330,N_9338,N_7288);
or UO_1331 (O_1331,N_7160,N_6928);
nand UO_1332 (O_1332,N_7991,N_7911);
and UO_1333 (O_1333,N_6487,N_6909);
nand UO_1334 (O_1334,N_8278,N_9991);
and UO_1335 (O_1335,N_8999,N_9425);
or UO_1336 (O_1336,N_6786,N_9176);
or UO_1337 (O_1337,N_7275,N_8012);
or UO_1338 (O_1338,N_9942,N_5721);
nand UO_1339 (O_1339,N_6765,N_7650);
nand UO_1340 (O_1340,N_7538,N_8563);
xnor UO_1341 (O_1341,N_5608,N_8487);
and UO_1342 (O_1342,N_7664,N_5624);
or UO_1343 (O_1343,N_9484,N_8061);
xnor UO_1344 (O_1344,N_6736,N_5694);
or UO_1345 (O_1345,N_8040,N_9977);
and UO_1346 (O_1346,N_8837,N_6560);
and UO_1347 (O_1347,N_6451,N_5956);
nor UO_1348 (O_1348,N_8254,N_7066);
nor UO_1349 (O_1349,N_7693,N_8615);
nor UO_1350 (O_1350,N_7881,N_5111);
or UO_1351 (O_1351,N_9628,N_5268);
nand UO_1352 (O_1352,N_7967,N_6540);
nand UO_1353 (O_1353,N_5703,N_5056);
nor UO_1354 (O_1354,N_5924,N_6588);
and UO_1355 (O_1355,N_7615,N_8992);
nand UO_1356 (O_1356,N_8704,N_9117);
nor UO_1357 (O_1357,N_6337,N_6073);
and UO_1358 (O_1358,N_8863,N_6561);
nand UO_1359 (O_1359,N_5888,N_9221);
nor UO_1360 (O_1360,N_6556,N_7321);
nor UO_1361 (O_1361,N_9172,N_6788);
nand UO_1362 (O_1362,N_8433,N_8220);
nand UO_1363 (O_1363,N_6884,N_9423);
or UO_1364 (O_1364,N_7890,N_8321);
xnor UO_1365 (O_1365,N_5201,N_9811);
or UO_1366 (O_1366,N_9598,N_5061);
nor UO_1367 (O_1367,N_5231,N_9128);
and UO_1368 (O_1368,N_8551,N_5390);
and UO_1369 (O_1369,N_7965,N_7227);
and UO_1370 (O_1370,N_9307,N_9154);
and UO_1371 (O_1371,N_7766,N_8076);
nor UO_1372 (O_1372,N_9590,N_7037);
nor UO_1373 (O_1373,N_9623,N_7358);
and UO_1374 (O_1374,N_6366,N_5265);
nand UO_1375 (O_1375,N_7740,N_5441);
nand UO_1376 (O_1376,N_9648,N_5378);
and UO_1377 (O_1377,N_7259,N_7749);
nand UO_1378 (O_1378,N_8919,N_8731);
nand UO_1379 (O_1379,N_6548,N_6234);
or UO_1380 (O_1380,N_8983,N_7087);
and UO_1381 (O_1381,N_8506,N_5961);
and UO_1382 (O_1382,N_8806,N_5969);
and UO_1383 (O_1383,N_8874,N_7853);
and UO_1384 (O_1384,N_7327,N_9259);
nor UO_1385 (O_1385,N_9073,N_8665);
and UO_1386 (O_1386,N_9373,N_8623);
nand UO_1387 (O_1387,N_9452,N_6844);
and UO_1388 (O_1388,N_6951,N_5663);
or UO_1389 (O_1389,N_7006,N_8857);
nand UO_1390 (O_1390,N_7778,N_7580);
nand UO_1391 (O_1391,N_8605,N_9457);
nand UO_1392 (O_1392,N_5872,N_7711);
and UO_1393 (O_1393,N_7054,N_7454);
nor UO_1394 (O_1394,N_5518,N_5232);
nand UO_1395 (O_1395,N_5021,N_7435);
nor UO_1396 (O_1396,N_8996,N_5729);
nor UO_1397 (O_1397,N_6333,N_5483);
or UO_1398 (O_1398,N_9216,N_8747);
nand UO_1399 (O_1399,N_6353,N_6656);
and UO_1400 (O_1400,N_8119,N_9044);
nor UO_1401 (O_1401,N_6116,N_8049);
nand UO_1402 (O_1402,N_5768,N_8781);
nand UO_1403 (O_1403,N_6004,N_5748);
nor UO_1404 (O_1404,N_7875,N_9957);
or UO_1405 (O_1405,N_9309,N_9712);
nor UO_1406 (O_1406,N_9163,N_8546);
nand UO_1407 (O_1407,N_6670,N_7414);
xnor UO_1408 (O_1408,N_6576,N_7415);
nor UO_1409 (O_1409,N_6408,N_5919);
nand UO_1410 (O_1410,N_5917,N_5769);
or UO_1411 (O_1411,N_5687,N_9913);
and UO_1412 (O_1412,N_6789,N_7267);
or UO_1413 (O_1413,N_8520,N_5014);
nor UO_1414 (O_1414,N_7023,N_5462);
nand UO_1415 (O_1415,N_6595,N_6340);
or UO_1416 (O_1416,N_9395,N_7220);
nand UO_1417 (O_1417,N_5096,N_8954);
nor UO_1418 (O_1418,N_5758,N_8259);
and UO_1419 (O_1419,N_9569,N_5270);
and UO_1420 (O_1420,N_9394,N_9616);
nand UO_1421 (O_1421,N_9702,N_6868);
nor UO_1422 (O_1422,N_7547,N_8303);
nor UO_1423 (O_1423,N_7097,N_8024);
and UO_1424 (O_1424,N_6941,N_5844);
nor UO_1425 (O_1425,N_6536,N_5053);
or UO_1426 (O_1426,N_9737,N_5884);
and UO_1427 (O_1427,N_9829,N_7446);
nand UO_1428 (O_1428,N_7569,N_7101);
nand UO_1429 (O_1429,N_7342,N_6386);
or UO_1430 (O_1430,N_5279,N_8898);
nor UO_1431 (O_1431,N_9774,N_6300);
nor UO_1432 (O_1432,N_6392,N_7111);
or UO_1433 (O_1433,N_8827,N_6242);
or UO_1434 (O_1434,N_6484,N_7870);
or UO_1435 (O_1435,N_9396,N_8201);
nor UO_1436 (O_1436,N_7073,N_7937);
nand UO_1437 (O_1437,N_6509,N_5696);
or UO_1438 (O_1438,N_5881,N_8566);
nand UO_1439 (O_1439,N_7599,N_9908);
nand UO_1440 (O_1440,N_7191,N_8879);
nand UO_1441 (O_1441,N_9808,N_9130);
nor UO_1442 (O_1442,N_5805,N_5305);
nor UO_1443 (O_1443,N_6832,N_7084);
nor UO_1444 (O_1444,N_9283,N_7309);
and UO_1445 (O_1445,N_8965,N_5588);
nand UO_1446 (O_1446,N_9710,N_6843);
and UO_1447 (O_1447,N_5662,N_5258);
nand UO_1448 (O_1448,N_9583,N_9237);
nor UO_1449 (O_1449,N_9114,N_8274);
and UO_1450 (O_1450,N_9667,N_7393);
nand UO_1451 (O_1451,N_9191,N_9244);
and UO_1452 (O_1452,N_5652,N_6749);
nand UO_1453 (O_1453,N_5901,N_5292);
nor UO_1454 (O_1454,N_7401,N_8840);
xor UO_1455 (O_1455,N_9066,N_9828);
and UO_1456 (O_1456,N_7433,N_9606);
nor UO_1457 (O_1457,N_7507,N_6526);
and UO_1458 (O_1458,N_8596,N_5342);
nor UO_1459 (O_1459,N_5380,N_7504);
or UO_1460 (O_1460,N_6671,N_7684);
nor UO_1461 (O_1461,N_8215,N_6348);
xnor UO_1462 (O_1462,N_5838,N_8098);
nor UO_1463 (O_1463,N_7347,N_7616);
nand UO_1464 (O_1464,N_6077,N_5370);
nand UO_1465 (O_1465,N_9722,N_6747);
nor UO_1466 (O_1466,N_9275,N_8882);
nand UO_1467 (O_1467,N_7444,N_8644);
or UO_1468 (O_1468,N_6258,N_9498);
nor UO_1469 (O_1469,N_7654,N_7903);
nor UO_1470 (O_1470,N_6558,N_8063);
nor UO_1471 (O_1471,N_9192,N_9655);
nor UO_1472 (O_1472,N_5855,N_7278);
nor UO_1473 (O_1473,N_5816,N_5044);
nor UO_1474 (O_1474,N_9381,N_9029);
and UO_1475 (O_1475,N_5439,N_8632);
nand UO_1476 (O_1476,N_7908,N_5601);
nand UO_1477 (O_1477,N_9851,N_8804);
or UO_1478 (O_1478,N_7313,N_8228);
and UO_1479 (O_1479,N_9876,N_8920);
nor UO_1480 (O_1480,N_5097,N_8148);
xor UO_1481 (O_1481,N_7602,N_9659);
nand UO_1482 (O_1482,N_7417,N_9692);
nand UO_1483 (O_1483,N_6700,N_7091);
nand UO_1484 (O_1484,N_6311,N_6354);
xor UO_1485 (O_1485,N_8258,N_7369);
xnor UO_1486 (O_1486,N_8728,N_6374);
or UO_1487 (O_1487,N_6685,N_5314);
nor UO_1488 (O_1488,N_8692,N_9663);
nand UO_1489 (O_1489,N_5819,N_9683);
nor UO_1490 (O_1490,N_8726,N_9767);
xnor UO_1491 (O_1491,N_5055,N_9910);
and UO_1492 (O_1492,N_8048,N_7492);
or UO_1493 (O_1493,N_9080,N_8140);
xnor UO_1494 (O_1494,N_9980,N_6520);
nor UO_1495 (O_1495,N_6404,N_6054);
nor UO_1496 (O_1496,N_5655,N_8286);
nor UO_1497 (O_1497,N_9889,N_9398);
and UO_1498 (O_1498,N_6430,N_7891);
or UO_1499 (O_1499,N_8943,N_6396);
endmodule