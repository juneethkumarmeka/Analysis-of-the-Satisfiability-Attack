module basic_1500_15000_2000_100_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_797,In_415);
xnor U1 (N_1,In_88,In_808);
nor U2 (N_2,In_931,In_522);
nor U3 (N_3,In_1320,In_849);
nand U4 (N_4,In_1352,In_519);
or U5 (N_5,In_403,In_578);
xnor U6 (N_6,In_1262,In_69);
or U7 (N_7,In_795,In_1488);
and U8 (N_8,In_1165,In_641);
nor U9 (N_9,In_92,In_168);
and U10 (N_10,In_251,In_208);
nand U11 (N_11,In_323,In_1004);
or U12 (N_12,In_1167,In_891);
or U13 (N_13,In_650,In_135);
or U14 (N_14,In_957,In_331);
or U15 (N_15,In_1222,In_1483);
and U16 (N_16,In_21,In_62);
nor U17 (N_17,In_357,In_2);
and U18 (N_18,In_827,In_541);
nor U19 (N_19,In_921,In_911);
or U20 (N_20,In_250,In_1146);
xnor U21 (N_21,In_1285,In_1446);
or U22 (N_22,In_1168,In_1407);
nand U23 (N_23,In_637,In_1208);
nand U24 (N_24,In_657,In_432);
or U25 (N_25,In_536,In_1094);
nand U26 (N_26,In_1154,In_1019);
xnor U27 (N_27,In_858,In_1074);
nor U28 (N_28,In_1455,In_400);
nor U29 (N_29,In_527,In_229);
nand U30 (N_30,In_1032,In_475);
nand U31 (N_31,In_1117,In_1387);
xor U32 (N_32,In_1113,In_65);
or U33 (N_33,In_205,In_939);
and U34 (N_34,In_502,In_1489);
or U35 (N_35,In_221,In_620);
or U36 (N_36,In_633,In_873);
xnor U37 (N_37,In_456,In_1394);
xor U38 (N_38,In_1369,In_480);
xnor U39 (N_39,In_362,In_699);
xnor U40 (N_40,In_1422,In_1327);
and U41 (N_41,In_1125,In_215);
nor U42 (N_42,In_387,In_1238);
or U43 (N_43,In_58,In_466);
nand U44 (N_44,In_252,In_1170);
nor U45 (N_45,In_52,In_28);
nor U46 (N_46,In_934,In_1250);
nor U47 (N_47,In_860,In_1034);
xor U48 (N_48,In_241,In_1178);
nand U49 (N_49,In_971,In_1185);
and U50 (N_50,In_568,In_384);
xor U51 (N_51,In_476,In_825);
or U52 (N_52,In_1015,In_870);
xnor U53 (N_53,In_1209,In_978);
nor U54 (N_54,In_1204,In_489);
nand U55 (N_55,In_1196,In_182);
and U56 (N_56,In_467,In_1449);
nand U57 (N_57,In_1467,In_1367);
xnor U58 (N_58,In_1482,In_974);
or U59 (N_59,In_976,In_1368);
or U60 (N_60,In_728,In_1420);
and U61 (N_61,In_1240,In_946);
nand U62 (N_62,In_1150,In_490);
and U63 (N_63,In_837,In_1048);
nor U64 (N_64,In_181,In_410);
and U65 (N_65,In_580,In_1025);
nor U66 (N_66,In_1353,In_523);
and U67 (N_67,In_433,In_555);
or U68 (N_68,In_553,In_360);
xor U69 (N_69,In_64,In_698);
xor U70 (N_70,In_100,In_1014);
nor U71 (N_71,In_932,In_600);
or U72 (N_72,In_347,In_492);
nor U73 (N_73,In_611,In_628);
and U74 (N_74,In_1399,In_1477);
or U75 (N_75,In_1003,In_1129);
nor U76 (N_76,In_140,In_908);
nor U77 (N_77,In_417,In_645);
xor U78 (N_78,In_109,In_816);
or U79 (N_79,In_1149,In_243);
nand U80 (N_80,In_775,In_917);
and U81 (N_81,In_393,In_1249);
or U82 (N_82,In_593,In_1405);
nor U83 (N_83,In_1356,In_1331);
xor U84 (N_84,In_327,In_428);
or U85 (N_85,In_546,In_590);
nor U86 (N_86,In_223,In_558);
and U87 (N_87,In_292,In_719);
or U88 (N_88,In_1417,In_1263);
nor U89 (N_89,In_705,In_226);
and U90 (N_90,In_499,In_701);
nor U91 (N_91,In_1491,In_312);
xnor U92 (N_92,In_582,In_416);
and U93 (N_93,In_570,In_671);
nand U94 (N_94,In_604,In_50);
and U95 (N_95,In_683,In_975);
and U96 (N_96,In_1148,In_867);
or U97 (N_97,In_634,In_144);
or U98 (N_98,In_378,In_1427);
or U99 (N_99,In_794,In_591);
and U100 (N_100,In_550,In_535);
nand U101 (N_101,In_1479,In_1051);
and U102 (N_102,In_1232,In_1342);
xnor U103 (N_103,In_1314,In_1438);
or U104 (N_104,In_1053,In_1036);
or U105 (N_105,In_413,In_183);
or U106 (N_106,In_1084,In_430);
and U107 (N_107,In_1218,In_201);
or U108 (N_108,In_1062,In_1227);
xnor U109 (N_109,In_508,In_624);
nand U110 (N_110,In_329,In_1210);
nor U111 (N_111,In_20,In_713);
xnor U112 (N_112,In_905,In_426);
and U113 (N_113,In_875,In_210);
and U114 (N_114,In_659,In_813);
nand U115 (N_115,In_748,In_147);
and U116 (N_116,In_772,In_836);
nor U117 (N_117,In_1144,In_264);
nor U118 (N_118,In_317,In_740);
xnor U119 (N_119,In_1445,In_708);
and U120 (N_120,In_494,In_1041);
or U121 (N_121,In_254,In_171);
and U122 (N_122,In_1081,In_320);
nand U123 (N_123,In_947,In_75);
or U124 (N_124,In_674,In_1038);
nor U125 (N_125,In_279,In_493);
nor U126 (N_126,In_1323,In_618);
nand U127 (N_127,In_742,In_663);
nor U128 (N_128,In_1079,In_642);
or U129 (N_129,In_782,In_824);
nand U130 (N_130,In_488,In_122);
xor U131 (N_131,In_40,In_124);
or U132 (N_132,In_608,In_167);
xor U133 (N_133,In_1241,In_1);
and U134 (N_134,In_1463,In_1220);
nor U135 (N_135,In_961,In_694);
or U136 (N_136,In_994,In_389);
nor U137 (N_137,In_636,In_512);
nor U138 (N_138,In_1098,In_391);
xor U139 (N_139,In_969,In_1176);
nor U140 (N_140,In_709,In_1305);
and U141 (N_141,In_1137,In_1141);
or U142 (N_142,In_1182,In_814);
nor U143 (N_143,In_599,In_78);
nand U144 (N_144,In_776,In_638);
or U145 (N_145,In_865,In_77);
and U146 (N_146,In_1122,In_1103);
and U147 (N_147,In_392,In_22);
nand U148 (N_148,In_449,In_283);
and U149 (N_149,In_809,In_734);
or U150 (N_150,N_120,In_190);
and U151 (N_151,In_1008,In_1063);
nand U152 (N_152,In_131,In_1310);
and U153 (N_153,In_589,N_49);
nor U154 (N_154,In_528,In_959);
nor U155 (N_155,In_697,In_1092);
or U156 (N_156,In_601,In_1005);
nand U157 (N_157,In_204,In_901);
nand U158 (N_158,In_848,In_1145);
xor U159 (N_159,In_665,In_534);
and U160 (N_160,In_817,In_1085);
nor U161 (N_161,In_1415,In_675);
xnor U162 (N_162,In_1410,In_815);
xnor U163 (N_163,In_273,N_130);
nor U164 (N_164,In_439,In_847);
nand U165 (N_165,In_784,In_635);
or U166 (N_166,In_557,In_1087);
and U167 (N_167,In_105,N_31);
nand U168 (N_168,In_12,In_481);
xnor U169 (N_169,In_197,In_532);
nand U170 (N_170,In_106,In_965);
xnor U171 (N_171,In_861,In_1059);
or U172 (N_172,In_585,N_123);
nand U173 (N_173,In_1118,In_130);
xnor U174 (N_174,In_1006,In_285);
xor U175 (N_175,In_414,In_455);
nor U176 (N_176,In_496,In_1304);
xnor U177 (N_177,In_1212,In_330);
nor U178 (N_178,In_596,In_1105);
nor U179 (N_179,In_244,In_690);
nor U180 (N_180,In_91,In_74);
nand U181 (N_181,In_515,In_1236);
nand U182 (N_182,In_649,N_34);
nand U183 (N_183,N_24,In_343);
xnor U184 (N_184,In_457,In_798);
and U185 (N_185,In_379,In_1200);
and U186 (N_186,In_1264,N_128);
and U187 (N_187,In_318,In_800);
and U188 (N_188,In_517,In_991);
xnor U189 (N_189,In_565,In_306);
or U190 (N_190,In_595,In_857);
and U191 (N_191,In_1409,In_818);
or U192 (N_192,In_364,In_348);
or U193 (N_193,In_380,In_29);
xnor U194 (N_194,In_1043,In_345);
nand U195 (N_195,N_13,In_1357);
or U196 (N_196,In_1026,In_262);
nor U197 (N_197,In_643,In_1276);
nand U198 (N_198,In_670,In_57);
and U199 (N_199,In_1269,In_136);
or U200 (N_200,In_575,In_446);
nand U201 (N_201,In_55,In_117);
nor U202 (N_202,In_929,In_664);
or U203 (N_203,In_1377,In_332);
or U204 (N_204,In_339,In_1365);
nand U205 (N_205,In_1341,In_763);
xnor U206 (N_206,In_371,In_552);
and U207 (N_207,In_463,In_1362);
or U208 (N_208,N_8,N_54);
nand U209 (N_209,In_113,In_491);
xnor U210 (N_210,N_148,In_1309);
nor U211 (N_211,In_1336,In_93);
nand U212 (N_212,In_462,In_443);
xor U213 (N_213,N_46,In_1108);
or U214 (N_214,In_531,In_655);
xor U215 (N_215,In_910,In_166);
nor U216 (N_216,In_654,In_887);
xor U217 (N_217,In_909,In_1132);
nor U218 (N_218,In_896,In_313);
or U219 (N_219,In_186,In_566);
nand U220 (N_220,In_884,In_841);
nand U221 (N_221,In_777,In_354);
and U222 (N_222,N_23,In_1257);
or U223 (N_223,In_988,In_429);
or U224 (N_224,In_53,In_757);
nand U225 (N_225,In_289,In_316);
or U226 (N_226,In_108,In_892);
nor U227 (N_227,In_559,In_823);
xnor U228 (N_228,In_743,In_998);
nor U229 (N_229,In_1239,In_514);
and U230 (N_230,In_471,In_1373);
xnor U231 (N_231,N_15,In_1473);
or U232 (N_232,In_383,In_1009);
or U233 (N_233,In_606,In_504);
xnor U234 (N_234,In_765,In_647);
xnor U235 (N_235,In_274,In_625);
or U236 (N_236,In_1088,In_1308);
nor U237 (N_237,In_1234,In_1030);
and U238 (N_238,In_673,In_1278);
nand U239 (N_239,In_472,N_48);
xor U240 (N_240,In_145,In_394);
xor U241 (N_241,In_1267,In_793);
nor U242 (N_242,In_469,N_39);
nor U243 (N_243,In_1172,In_1237);
or U244 (N_244,In_381,N_144);
nand U245 (N_245,In_34,In_258);
or U246 (N_246,N_113,In_1187);
and U247 (N_247,In_406,In_352);
xnor U248 (N_248,In_882,In_1119);
or U249 (N_249,In_342,In_543);
or U250 (N_250,In_195,In_501);
or U251 (N_251,In_717,In_792);
or U252 (N_252,In_881,In_275);
and U253 (N_253,In_878,In_866);
xor U254 (N_254,In_1364,In_497);
nand U255 (N_255,In_933,In_335);
and U256 (N_256,In_1198,In_483);
xor U257 (N_257,In_1343,In_603);
xor U258 (N_258,In_454,In_1339);
nand U259 (N_259,In_260,In_930);
nor U260 (N_260,In_1421,In_706);
and U261 (N_261,In_588,In_1175);
and U262 (N_262,In_747,In_282);
nand U263 (N_263,In_193,In_453);
or U264 (N_264,In_723,In_1286);
or U265 (N_265,In_1457,N_43);
nor U266 (N_266,In_27,In_160);
and U267 (N_267,In_1181,In_1426);
xnor U268 (N_268,In_1333,In_1465);
nor U269 (N_269,In_288,In_1072);
nand U270 (N_270,In_1192,In_407);
nor U271 (N_271,In_1383,N_115);
xor U272 (N_272,In_177,N_20);
or U273 (N_273,In_1462,In_1090);
and U274 (N_274,In_926,N_62);
or U275 (N_275,In_983,In_1121);
xnor U276 (N_276,In_1490,In_803);
xnor U277 (N_277,In_950,In_24);
xnor U278 (N_278,In_159,In_1423);
xor U279 (N_279,In_894,In_658);
or U280 (N_280,N_67,In_1441);
and U281 (N_281,In_175,In_781);
nand U282 (N_282,In_72,In_1224);
nor U283 (N_283,In_851,In_1280);
xnor U284 (N_284,In_125,In_89);
or U285 (N_285,In_547,In_962);
nor U286 (N_286,In_265,In_322);
nor U287 (N_287,In_987,N_76);
xnor U288 (N_288,In_1416,In_1156);
xnor U289 (N_289,In_1271,In_1425);
or U290 (N_290,In_750,In_1289);
or U291 (N_291,In_902,N_40);
nor U292 (N_292,In_1470,In_738);
and U293 (N_293,In_544,In_1444);
nand U294 (N_294,In_1207,In_1223);
nor U295 (N_295,In_944,In_1406);
nand U296 (N_296,In_778,In_1151);
nand U297 (N_297,In_291,In_1318);
nand U298 (N_298,In_626,In_812);
xor U299 (N_299,In_1114,In_680);
nand U300 (N_300,In_32,In_666);
nor U301 (N_301,In_760,In_725);
nor U302 (N_302,N_223,In_948);
or U303 (N_303,N_121,In_419);
nor U304 (N_304,In_460,In_1066);
nor U305 (N_305,N_82,In_859);
and U306 (N_306,In_754,N_116);
and U307 (N_307,In_188,In_1096);
nand U308 (N_308,In_485,In_1221);
nor U309 (N_309,In_1219,In_39);
and U310 (N_310,N_216,In_679);
or U311 (N_311,In_821,In_1229);
xor U312 (N_312,In_421,In_774);
nor U313 (N_313,In_985,In_1231);
nand U314 (N_314,In_533,In_468);
and U315 (N_315,In_1291,In_368);
xor U316 (N_316,In_1312,In_1055);
and U317 (N_317,In_810,In_257);
and U318 (N_318,N_68,In_925);
and U319 (N_319,In_669,In_744);
or U320 (N_320,In_1329,N_190);
xor U321 (N_321,In_115,In_630);
nor U322 (N_322,In_33,In_386);
and U323 (N_323,N_207,In_79);
xor U324 (N_324,In_1284,N_14);
and U325 (N_325,N_60,In_15);
nand U326 (N_326,In_1018,In_1259);
or U327 (N_327,In_94,In_672);
nand U328 (N_328,In_629,In_337);
or U329 (N_329,In_1017,N_124);
nor U330 (N_330,In_819,In_646);
nand U331 (N_331,In_296,N_66);
nor U332 (N_332,In_1100,N_184);
or U333 (N_333,In_358,In_459);
nor U334 (N_334,In_1296,In_422);
nand U335 (N_335,In_684,In_940);
nor U336 (N_336,In_266,In_294);
and U337 (N_337,In_1251,In_1303);
or U338 (N_338,In_377,In_158);
and U339 (N_339,N_260,In_1130);
and U340 (N_340,N_254,N_234);
nor U341 (N_341,In_1374,In_1325);
or U342 (N_342,In_839,N_210);
and U343 (N_343,In_1474,In_622);
and U344 (N_344,In_1190,N_265);
or U345 (N_345,In_1344,In_268);
or U346 (N_346,In_854,In_325);
xor U347 (N_347,N_75,In_581);
nand U348 (N_348,In_179,N_38);
or U349 (N_349,N_110,In_762);
or U350 (N_350,In_1412,In_1225);
and U351 (N_351,N_140,In_1136);
nor U352 (N_352,In_1272,N_78);
xnor U353 (N_353,N_224,N_199);
xor U354 (N_354,In_1253,N_74);
xor U355 (N_355,In_955,N_73);
and U356 (N_356,In_960,In_990);
and U357 (N_357,In_928,In_1022);
nand U358 (N_358,N_119,In_804);
xor U359 (N_359,In_1177,In_1171);
and U360 (N_360,In_833,In_486);
or U361 (N_361,In_143,In_46);
nand U362 (N_362,In_464,In_949);
or U363 (N_363,In_1452,In_716);
nor U364 (N_364,In_355,In_912);
nand U365 (N_365,In_838,In_1328);
and U366 (N_366,In_977,In_752);
nand U367 (N_367,In_1045,N_232);
and U368 (N_368,In_18,In_324);
xor U369 (N_369,In_1366,In_1469);
nand U370 (N_370,In_1155,In_731);
nand U371 (N_371,In_1195,In_1299);
xor U372 (N_372,In_35,In_1486);
xor U373 (N_373,In_919,In_227);
nand U374 (N_374,In_1307,In_602);
nor U375 (N_375,In_1306,In_548);
or U376 (N_376,In_554,In_290);
nor U377 (N_377,In_104,N_213);
nor U378 (N_378,In_209,In_81);
nor U379 (N_379,In_632,In_662);
nand U380 (N_380,In_154,In_871);
xnor U381 (N_381,In_116,In_831);
or U382 (N_382,In_1203,In_832);
nor U383 (N_383,N_280,N_83);
xnor U384 (N_384,In_1281,N_111);
or U385 (N_385,In_989,In_726);
and U386 (N_386,In_869,In_1235);
and U387 (N_387,In_739,In_148);
xor U388 (N_388,In_1497,In_1091);
nor U389 (N_389,In_1057,N_152);
nor U390 (N_390,In_0,In_1393);
or U391 (N_391,In_98,In_1166);
or U392 (N_392,N_283,In_129);
or U393 (N_393,In_1363,In_1456);
nand U394 (N_394,In_1095,In_906);
nand U395 (N_395,In_503,In_702);
nor U396 (N_396,N_189,N_222);
nor U397 (N_397,In_302,In_1401);
nor U398 (N_398,In_724,In_1180);
xnor U399 (N_399,N_35,In_972);
nand U400 (N_400,In_941,In_574);
xnor U401 (N_401,In_230,In_1040);
and U402 (N_402,N_278,In_365);
and U403 (N_403,N_295,In_1076);
or U404 (N_404,In_1120,N_166);
xnor U405 (N_405,In_395,In_1390);
xnor U406 (N_406,In_1135,In_610);
and U407 (N_407,In_240,In_1138);
or U408 (N_408,N_63,In_1340);
nand U409 (N_409,In_995,In_1109);
and U410 (N_410,In_304,In_615);
nand U411 (N_411,In_1215,In_1375);
and U412 (N_412,In_149,In_922);
nor U413 (N_413,In_1011,In_86);
nor U414 (N_414,N_109,In_834);
and U415 (N_415,In_644,N_151);
or U416 (N_416,In_676,N_45);
or U417 (N_417,N_155,In_592);
nand U418 (N_418,In_1395,In_99);
nor U419 (N_419,In_401,In_1322);
or U420 (N_420,In_156,N_267);
and U421 (N_421,N_266,N_233);
or U422 (N_422,N_159,In_126);
nand U423 (N_423,In_1037,N_293);
and U424 (N_424,N_5,In_829);
or U425 (N_425,In_913,N_86);
nand U426 (N_426,N_284,In_425);
nor U427 (N_427,In_133,In_60);
or U428 (N_428,In_199,In_138);
or U429 (N_429,N_220,N_297);
or U430 (N_430,N_239,In_1226);
or U431 (N_431,In_44,In_597);
or U432 (N_432,In_1458,In_704);
nor U433 (N_433,In_900,N_235);
xor U434 (N_434,In_41,N_104);
nand U435 (N_435,In_758,N_251);
xnor U436 (N_436,In_661,In_567);
nand U437 (N_437,In_225,In_842);
nor U438 (N_438,In_1140,N_149);
nor U439 (N_439,In_119,N_182);
xor U440 (N_440,In_936,N_240);
or U441 (N_441,In_1496,In_916);
nand U442 (N_442,N_22,In_877);
nand U443 (N_443,N_187,In_651);
nor U444 (N_444,In_1106,In_1345);
and U445 (N_445,In_561,In_607);
xor U446 (N_446,In_880,In_759);
nand U447 (N_447,In_889,In_1378);
xnor U448 (N_448,N_36,In_899);
nor U449 (N_449,In_741,In_789);
nand U450 (N_450,In_202,In_807);
nand U451 (N_451,In_801,In_1184);
and U452 (N_452,In_806,N_428);
xnor U453 (N_453,N_378,N_401);
nor U454 (N_454,In_1268,In_152);
xnor U455 (N_455,In_1186,N_440);
nor U456 (N_456,In_1348,In_13);
nor U457 (N_457,In_1016,N_92);
nor U458 (N_458,In_805,In_1391);
and U459 (N_459,In_1346,In_1370);
xnor U460 (N_460,N_225,In_1277);
and U461 (N_461,N_188,In_1010);
xor U462 (N_462,N_259,N_402);
xor U463 (N_463,N_360,N_186);
xor U464 (N_464,In_9,In_1332);
nor U465 (N_465,N_81,N_371);
nand U466 (N_466,In_997,N_201);
nor U467 (N_467,In_883,In_11);
nor U468 (N_468,In_1450,In_301);
and U469 (N_469,In_1243,In_1230);
nand U470 (N_470,In_1321,N_412);
nand U471 (N_471,In_1233,In_506);
xnor U472 (N_472,N_19,In_295);
nor U473 (N_473,In_874,In_328);
xnor U474 (N_474,In_43,In_155);
or U475 (N_475,N_393,In_1179);
xor U476 (N_476,In_1354,N_100);
and U477 (N_477,N_291,In_1400);
xor U478 (N_478,N_18,In_923);
nand U479 (N_479,In_952,In_542);
nor U480 (N_480,In_299,In_1077);
xnor U481 (N_481,In_1388,N_382);
or U482 (N_482,In_1110,In_1478);
and U483 (N_483,In_307,N_141);
nor U484 (N_484,In_573,N_139);
or U485 (N_485,N_230,N_179);
xor U486 (N_486,In_937,In_1134);
nor U487 (N_487,N_229,N_91);
xnor U488 (N_488,In_918,N_404);
nor U489 (N_489,N_30,In_445);
nand U490 (N_490,N_391,In_287);
and U491 (N_491,In_1020,In_1300);
or U492 (N_492,N_12,In_1334);
or U493 (N_493,N_136,In_885);
and U494 (N_494,In_263,N_127);
nand U495 (N_495,N_416,In_1358);
nor U496 (N_496,In_1052,In_1199);
nor U497 (N_497,In_1065,N_362);
xnor U498 (N_498,In_691,In_621);
xor U499 (N_499,In_879,In_1432);
nand U500 (N_500,In_811,In_967);
nand U501 (N_501,In_999,In_1023);
or U502 (N_502,In_920,In_207);
and U503 (N_503,In_914,In_1494);
or U504 (N_504,In_1436,N_84);
xor U505 (N_505,N_417,In_121);
and U506 (N_506,In_434,N_53);
or U507 (N_507,In_1159,N_292);
and U508 (N_508,N_262,N_185);
and U509 (N_509,N_173,N_118);
nand U510 (N_510,In_1101,In_746);
and U511 (N_511,In_281,In_1498);
xor U512 (N_512,N_95,N_305);
nor U513 (N_513,N_331,In_478);
or U514 (N_514,In_402,In_217);
and U515 (N_515,In_1073,N_385);
nand U516 (N_516,In_1350,In_828);
nand U517 (N_517,N_181,In_1265);
and U518 (N_518,In_284,In_373);
xor U519 (N_519,In_1376,N_328);
nor U520 (N_520,In_103,In_1158);
nor U521 (N_521,N_28,N_303);
and U522 (N_522,In_876,N_316);
nand U523 (N_523,N_1,N_348);
or U524 (N_524,N_405,N_64);
or U525 (N_525,In_76,In_1169);
nand U526 (N_526,In_1021,In_1266);
or U527 (N_527,N_314,In_703);
or U528 (N_528,In_1248,In_745);
nor U529 (N_529,In_1044,N_304);
nor U530 (N_530,In_1258,In_1058);
nand U531 (N_531,In_271,N_433);
and U532 (N_532,In_5,N_205);
nand U533 (N_533,N_359,In_730);
or U534 (N_534,In_1411,In_714);
and U535 (N_535,N_275,In_231);
nor U536 (N_536,In_964,In_564);
nor U537 (N_537,In_83,In_165);
and U538 (N_538,In_1163,N_11);
and U539 (N_539,In_769,In_310);
nand U540 (N_540,N_312,N_211);
and U541 (N_541,In_845,In_1419);
or U542 (N_542,N_287,In_720);
and U543 (N_543,N_327,In_820);
and U544 (N_544,In_150,N_103);
xor U545 (N_545,N_344,N_156);
and U546 (N_546,In_1161,In_897);
xor U547 (N_547,N_50,N_408);
or U548 (N_548,N_379,In_511);
nand U549 (N_549,In_137,In_1152);
nor U550 (N_550,N_323,In_992);
xnor U551 (N_551,In_678,N_298);
nand U552 (N_552,In_872,N_336);
xnor U553 (N_553,In_1392,In_412);
nor U554 (N_554,N_6,N_33);
and U555 (N_555,N_218,In_498);
nand U556 (N_556,In_112,In_1397);
nor U557 (N_557,In_545,In_1211);
or U558 (N_558,N_129,In_95);
and U559 (N_559,In_732,N_432);
xnor U560 (N_560,In_826,In_84);
and U561 (N_561,In_692,In_915);
nor U562 (N_562,N_167,In_333);
nand U563 (N_563,N_164,In_1338);
xnor U564 (N_564,In_1127,In_1459);
nand U565 (N_565,In_1492,N_3);
and U566 (N_566,N_367,N_135);
nor U567 (N_567,In_269,In_151);
nand U568 (N_568,N_330,In_1351);
and U569 (N_569,In_787,In_583);
or U570 (N_570,In_1142,N_352);
and U571 (N_571,In_189,In_427);
xor U572 (N_572,N_231,In_351);
nor U573 (N_573,N_426,In_1042);
xnor U574 (N_574,N_228,In_110);
nand U575 (N_575,In_943,N_268);
nor U576 (N_576,In_300,In_396);
nor U577 (N_577,In_1075,N_142);
nor U578 (N_578,In_107,In_1027);
and U579 (N_579,N_301,In_529);
xor U580 (N_580,N_398,In_157);
or U581 (N_581,N_439,In_1319);
nand U582 (N_582,In_1029,In_1324);
nand U583 (N_583,In_1371,In_979);
and U584 (N_584,N_363,In_286);
or U585 (N_585,N_313,In_146);
nand U586 (N_586,In_1050,In_326);
nor U587 (N_587,N_158,N_44);
or U588 (N_588,In_668,In_141);
xnor U589 (N_589,N_52,In_1162);
nor U590 (N_590,In_1293,In_802);
nor U591 (N_591,N_438,N_320);
nor U592 (N_592,N_203,N_209);
nand U593 (N_593,In_1254,In_114);
nor U594 (N_594,In_1194,In_1402);
xnor U595 (N_595,In_579,In_123);
nand U596 (N_596,In_1433,In_584);
or U597 (N_597,N_29,N_341);
xor U598 (N_598,In_1201,In_253);
or U599 (N_599,In_1317,In_791);
and U600 (N_600,N_131,N_134);
xnor U601 (N_601,N_517,N_552);
nand U602 (N_602,N_480,N_546);
nand U603 (N_603,N_146,In_340);
nor U604 (N_604,N_347,In_436);
and U605 (N_605,N_163,In_788);
xor U606 (N_606,In_1316,In_214);
or U607 (N_607,N_446,In_349);
and U608 (N_608,In_1413,In_945);
xnor U609 (N_609,In_200,N_522);
nor U610 (N_610,In_1282,N_554);
nand U611 (N_611,In_1160,In_660);
nand U612 (N_612,In_450,In_1024);
or U613 (N_613,In_85,In_344);
nand U614 (N_614,In_1191,N_102);
nand U615 (N_615,N_58,N_177);
xor U616 (N_616,In_707,N_421);
nand U617 (N_617,N_270,N_194);
or U618 (N_618,N_192,In_594);
nor U619 (N_619,N_411,In_1205);
and U620 (N_620,N_538,N_241);
and U621 (N_621,In_465,In_203);
nand U622 (N_622,N_541,N_108);
and U623 (N_623,N_273,In_667);
nor U624 (N_624,N_381,N_257);
nor U625 (N_625,N_471,In_715);
nor U626 (N_626,N_162,N_528);
and U627 (N_627,N_326,In_693);
nor U628 (N_628,N_306,In_1031);
and U629 (N_629,In_686,N_434);
and U630 (N_630,N_236,In_297);
nor U631 (N_631,N_559,N_390);
nand U632 (N_632,In_1287,In_1431);
nor U633 (N_633,In_1311,N_290);
nor U634 (N_634,In_237,N_176);
and U635 (N_635,In_495,In_1080);
nor U636 (N_636,In_613,In_631);
nand U637 (N_637,N_200,In_1068);
or U638 (N_638,In_770,N_445);
xnor U639 (N_639,In_1484,In_388);
and U640 (N_640,In_30,In_54);
nand U641 (N_641,N_365,N_99);
or U642 (N_642,In_369,N_450);
and U643 (N_643,N_504,N_544);
or U644 (N_644,In_982,In_451);
and U645 (N_645,N_513,In_907);
nand U646 (N_646,N_473,In_56);
nand U647 (N_647,N_322,N_286);
nor U648 (N_648,In_1437,N_551);
or U649 (N_649,In_187,N_456);
and U650 (N_650,N_126,In_799);
xor U651 (N_651,In_1439,N_383);
nand U652 (N_652,In_785,In_1093);
xor U653 (N_653,N_520,N_343);
nand U654 (N_654,In_1013,In_1487);
or U655 (N_655,In_1070,In_479);
nor U656 (N_656,N_452,N_310);
nor U657 (N_657,N_370,In_711);
nor U658 (N_658,In_14,In_118);
nor U659 (N_659,In_461,N_356);
or U660 (N_660,N_342,N_477);
nor U661 (N_661,In_382,In_520);
nor U662 (N_662,N_478,N_543);
and U663 (N_663,In_196,In_17);
nand U664 (N_664,N_249,In_1447);
xor U665 (N_665,In_996,In_1256);
nor U666 (N_666,N_444,In_1468);
or U667 (N_667,In_1481,N_319);
nor U668 (N_668,In_442,N_437);
xor U669 (N_669,N_55,In_1028);
nand U670 (N_670,N_96,In_1451);
or U671 (N_671,In_1089,N_540);
nor U672 (N_672,N_508,In_66);
and U673 (N_673,In_303,N_415);
or U674 (N_674,N_269,N_208);
nand U675 (N_675,N_539,N_154);
nor U676 (N_676,N_531,In_640);
and U677 (N_677,In_755,In_556);
and U678 (N_678,N_483,In_211);
nand U679 (N_679,N_107,N_198);
nand U680 (N_680,In_6,N_566);
or U681 (N_681,In_36,N_89);
nor U682 (N_682,N_418,In_1355);
nand U683 (N_683,N_376,In_898);
xor U684 (N_684,In_1228,N_193);
nand U685 (N_685,N_587,N_247);
nor U686 (N_686,In_234,N_373);
nand U687 (N_687,In_162,N_424);
or U688 (N_688,In_509,In_233);
and U689 (N_689,In_267,In_1380);
and U690 (N_690,In_786,In_51);
nand U691 (N_691,In_1104,In_935);
nand U692 (N_692,N_307,N_157);
nor U693 (N_693,In_350,In_904);
nor U694 (N_694,In_1475,N_474);
xnor U695 (N_695,N_219,N_423);
nand U696 (N_696,In_1472,N_550);
xnor U697 (N_697,In_82,In_886);
or U698 (N_698,In_169,N_16);
nand U699 (N_699,In_470,N_431);
xor U700 (N_700,In_1360,In_1012);
and U701 (N_701,In_1047,N_395);
and U702 (N_702,In_1435,In_153);
nand U703 (N_703,N_578,In_1007);
and U704 (N_704,In_973,N_582);
xor U705 (N_705,N_105,N_80);
and U706 (N_706,N_358,In_367);
nor U707 (N_707,In_537,In_452);
or U708 (N_708,In_276,N_0);
or U709 (N_709,N_87,N_355);
nor U710 (N_710,In_938,N_542);
or U711 (N_711,N_500,N_145);
or U712 (N_712,In_652,In_174);
nor U713 (N_713,In_314,In_751);
and U714 (N_714,N_32,N_377);
and U715 (N_715,In_247,N_243);
and U716 (N_716,In_67,In_844);
nor U717 (N_717,N_386,N_463);
or U718 (N_718,In_1398,In_1298);
or U719 (N_719,In_980,N_481);
or U720 (N_720,N_574,N_277);
and U721 (N_721,N_460,N_594);
or U722 (N_722,N_372,In_222);
and U723 (N_723,N_334,N_339);
or U724 (N_724,N_274,In_780);
nand U725 (N_725,N_132,In_1164);
and U726 (N_726,N_165,N_558);
or U727 (N_727,N_17,In_735);
xnor U728 (N_728,In_1061,N_160);
xnor U729 (N_729,In_507,N_97);
and U730 (N_730,N_143,In_1313);
or U731 (N_731,N_529,In_721);
nor U732 (N_732,In_1292,N_180);
and U733 (N_733,In_10,N_317);
and U734 (N_734,In_87,In_172);
and U735 (N_735,N_562,N_533);
or U736 (N_736,N_494,N_374);
nor U737 (N_737,In_474,N_467);
nand U738 (N_738,In_1183,N_548);
and U739 (N_739,N_576,N_488);
nand U740 (N_740,N_217,In_1389);
or U741 (N_741,N_147,In_218);
and U742 (N_742,N_285,In_255);
and U743 (N_743,In_1097,N_588);
nor U744 (N_744,In_1326,In_1102);
or U745 (N_745,N_125,In_1275);
nor U746 (N_746,In_1060,In_308);
nand U747 (N_747,In_616,In_1188);
or U748 (N_748,N_221,N_340);
nand U749 (N_749,In_729,In_376);
nand U750 (N_750,N_625,N_183);
nand U751 (N_751,In_500,N_557);
and U752 (N_752,N_724,In_1385);
nand U753 (N_753,N_638,N_687);
nand U754 (N_754,In_184,N_665);
and U755 (N_755,In_59,In_840);
and U756 (N_756,N_660,In_563);
and U757 (N_757,N_530,In_370);
nor U758 (N_758,N_455,In_1270);
xnor U759 (N_759,N_697,N_575);
or U760 (N_760,N_425,N_746);
nor U761 (N_761,In_418,In_185);
and U762 (N_762,N_555,In_524);
xor U763 (N_763,In_142,N_740);
or U764 (N_764,N_138,N_250);
and U765 (N_765,N_357,In_246);
xor U766 (N_766,In_90,N_565);
and U767 (N_767,N_244,N_375);
or U768 (N_768,N_527,N_721);
or U769 (N_769,In_128,In_372);
nor U770 (N_770,In_970,N_79);
or U771 (N_771,N_168,N_281);
or U772 (N_772,In_1206,N_353);
or U773 (N_773,N_674,N_675);
xnor U774 (N_774,N_429,In_1301);
nor U775 (N_775,N_475,N_617);
nor U776 (N_776,In_101,In_1408);
nor U777 (N_777,N_394,N_288);
xor U778 (N_778,N_389,In_321);
and U779 (N_779,N_388,N_503);
nand U780 (N_780,In_311,N_325);
xor U781 (N_781,In_338,N_294);
nand U782 (N_782,N_308,N_714);
nand U783 (N_783,N_302,In_1418);
xnor U784 (N_784,In_1086,In_1139);
or U785 (N_785,N_672,N_506);
nand U786 (N_786,In_341,In_530);
nor U787 (N_787,In_346,N_627);
xnor U788 (N_788,N_461,N_387);
nor U789 (N_789,N_430,In_1442);
xnor U790 (N_790,In_958,In_688);
and U791 (N_791,In_219,In_639);
and U792 (N_792,In_924,N_466);
nor U793 (N_793,In_220,N_512);
xor U794 (N_794,N_252,In_850);
nand U795 (N_795,In_236,In_1361);
nor U796 (N_796,N_485,N_636);
nor U797 (N_797,In_1083,N_26);
nor U798 (N_798,In_405,In_569);
or U799 (N_799,In_1464,In_42);
or U800 (N_800,N_604,N_616);
nor U801 (N_801,In_681,In_539);
and U802 (N_802,In_37,In_764);
or U803 (N_803,N_400,N_479);
or U804 (N_804,N_441,N_689);
nor U805 (N_805,N_414,N_21);
or U806 (N_806,In_893,N_628);
nor U807 (N_807,In_319,N_169);
and U808 (N_808,In_1255,N_191);
xnor U809 (N_809,In_180,In_238);
nor U810 (N_810,N_612,N_271);
nor U811 (N_811,N_368,N_639);
xor U812 (N_812,N_197,N_719);
or U813 (N_813,N_215,N_88);
or U814 (N_814,In_951,N_729);
nand U815 (N_815,N_454,N_101);
or U816 (N_816,In_423,In_1252);
nor U817 (N_817,In_487,N_472);
nor U818 (N_818,N_492,N_410);
xor U819 (N_819,N_276,In_1244);
and U820 (N_820,N_652,N_677);
xnor U821 (N_821,In_779,In_363);
xor U822 (N_822,In_1485,N_610);
xnor U823 (N_823,In_68,In_277);
nor U824 (N_824,In_435,N_703);
xor U825 (N_825,N_735,N_514);
nand U826 (N_826,N_650,In_293);
xor U827 (N_827,N_666,N_692);
xnor U828 (N_828,In_696,N_491);
xnor U829 (N_829,N_642,N_585);
nor U830 (N_830,In_259,N_122);
nand U831 (N_831,N_338,N_246);
xor U832 (N_832,N_662,In_1335);
xnor U833 (N_833,N_690,In_1434);
or U834 (N_834,N_621,N_153);
nand U835 (N_835,N_647,In_235);
nor U836 (N_836,N_204,N_623);
and U837 (N_837,In_361,In_1112);
nor U838 (N_838,In_1274,In_737);
and U839 (N_839,N_510,In_1359);
nor U840 (N_840,In_1202,N_300);
and U841 (N_841,In_510,In_315);
and U842 (N_842,N_172,In_232);
xor U843 (N_843,N_384,In_1273);
or U844 (N_844,N_603,N_289);
nand U845 (N_845,N_42,In_7);
nand U846 (N_846,In_1035,N_495);
and U847 (N_847,In_409,N_170);
xor U848 (N_848,In_576,In_968);
xor U849 (N_849,N_547,N_442);
nor U850 (N_850,In_768,N_556);
xor U851 (N_851,N_214,N_447);
or U852 (N_852,In_855,N_676);
nand U853 (N_853,In_1033,N_570);
nor U854 (N_854,In_1107,N_671);
nor U855 (N_855,N_515,In_1330);
and U856 (N_856,N_366,N_630);
or U857 (N_857,N_354,In_1039);
xnor U858 (N_858,In_127,N_739);
and U859 (N_859,N_599,N_648);
xor U860 (N_860,In_551,In_1290);
nor U861 (N_861,In_242,N_272);
xor U862 (N_862,In_178,In_1078);
nand U863 (N_863,In_298,N_651);
nor U864 (N_864,In_71,N_248);
or U865 (N_865,N_580,In_270);
or U866 (N_866,N_174,N_72);
or U867 (N_867,In_1115,N_511);
nor U868 (N_868,In_448,N_321);
nand U869 (N_869,In_586,N_620);
nor U870 (N_870,In_245,In_1124);
and U871 (N_871,In_48,N_256);
nor U872 (N_872,N_279,N_324);
xnor U873 (N_873,In_993,In_1297);
nand U874 (N_874,N_4,N_668);
or U875 (N_875,In_305,N_493);
nor U876 (N_876,In_853,In_431);
nor U877 (N_877,In_441,In_722);
nor U878 (N_878,In_617,In_1315);
xor U879 (N_879,N_712,N_59);
nand U880 (N_880,N_486,N_245);
nand U881 (N_881,N_581,In_954);
and U882 (N_882,In_862,In_1189);
and U883 (N_883,N_490,In_19);
nand U884 (N_884,N_663,N_69);
or U885 (N_885,In_1116,In_1382);
nor U886 (N_886,N_597,N_571);
xnor U887 (N_887,In_170,In_120);
and U888 (N_888,N_178,N_745);
xnor U889 (N_889,N_315,In_424);
nor U890 (N_890,N_661,In_598);
and U891 (N_891,In_397,N_7);
nand U892 (N_892,N_723,N_629);
and U893 (N_893,In_484,In_1131);
nand U894 (N_894,In_23,N_406);
and U895 (N_895,In_1197,In_447);
and U896 (N_896,In_1099,N_701);
nor U897 (N_897,N_563,In_216);
nand U898 (N_898,In_1242,N_744);
xor U899 (N_899,N_489,In_648);
and U900 (N_900,In_749,N_90);
and U901 (N_901,N_784,N_397);
and U902 (N_902,In_927,N_772);
and U903 (N_903,N_876,N_841);
nor U904 (N_904,N_175,N_584);
xor U905 (N_905,N_459,In_1440);
nand U906 (N_906,N_263,N_878);
xor U907 (N_907,N_679,N_545);
nor U908 (N_908,N_106,N_577);
or U909 (N_909,N_664,In_280);
or U910 (N_910,N_659,In_1414);
nor U911 (N_911,In_1064,N_568);
and U912 (N_912,N_759,In_1056);
or U913 (N_913,In_473,N_776);
or U914 (N_914,In_1214,N_762);
nor U915 (N_915,In_164,N_632);
nor U916 (N_916,N_823,N_282);
xnor U917 (N_917,N_443,N_656);
or U918 (N_918,N_706,N_896);
xor U919 (N_919,In_830,N_299);
and U920 (N_920,N_820,N_750);
and U921 (N_921,N_448,In_1001);
xnor U922 (N_922,In_80,N_863);
nor U923 (N_923,N_85,N_837);
and U924 (N_924,N_202,N_808);
nand U925 (N_925,In_895,In_356);
and U926 (N_926,In_191,In_248);
nor U927 (N_927,N_518,In_163);
and U928 (N_928,N_694,In_1424);
or U929 (N_929,In_1054,N_688);
or U930 (N_930,N_560,In_399);
xor U931 (N_931,In_173,N_653);
and U932 (N_932,In_132,N_351);
and U933 (N_933,N_611,N_778);
xnor U934 (N_934,In_981,In_1126);
xor U935 (N_935,N_757,N_715);
or U936 (N_936,N_507,N_741);
nand U937 (N_937,In_440,In_516);
xnor U938 (N_938,N_524,N_732);
and U939 (N_939,N_332,N_806);
nor U940 (N_940,N_794,N_685);
or U941 (N_941,N_822,N_756);
nor U942 (N_942,N_796,N_469);
or U943 (N_943,In_1302,In_695);
and U944 (N_944,In_1246,N_71);
xor U945 (N_945,In_334,In_1443);
xor U946 (N_946,In_278,In_540);
xor U947 (N_947,In_1495,In_1193);
xor U948 (N_948,In_700,N_764);
nor U949 (N_949,N_634,N_691);
and U950 (N_950,N_846,N_889);
and U951 (N_951,In_212,N_509);
xnor U952 (N_952,N_804,N_549);
and U953 (N_953,N_465,N_824);
and U954 (N_954,In_1404,N_699);
or U955 (N_955,N_258,N_56);
nand U956 (N_956,N_335,N_895);
and U957 (N_957,In_1247,N_553);
or U958 (N_958,N_502,In_1002);
or U959 (N_959,In_903,N_737);
or U960 (N_960,In_712,N_850);
nor U961 (N_961,N_836,N_70);
or U962 (N_962,In_733,N_708);
nor U963 (N_963,N_743,N_854);
nor U964 (N_964,N_525,N_851);
nor U965 (N_965,N_532,In_890);
xor U966 (N_966,In_623,In_1461);
nor U967 (N_967,N_613,In_26);
xor U968 (N_968,N_805,N_484);
or U969 (N_969,In_309,In_549);
nor U970 (N_970,In_1428,N_618);
xnor U971 (N_971,N_482,In_61);
or U972 (N_972,N_579,In_1174);
and U973 (N_973,N_615,In_1460);
nor U974 (N_974,N_874,N_897);
or U975 (N_975,N_898,N_887);
nor U976 (N_976,N_839,N_821);
xor U977 (N_977,N_844,In_213);
xnor U978 (N_978,In_761,N_780);
xor U979 (N_979,N_852,N_94);
or U980 (N_980,N_829,N_626);
xnor U981 (N_981,N_726,In_438);
xor U982 (N_982,N_601,In_1499);
nand U983 (N_983,N_774,N_700);
xnor U984 (N_984,N_885,In_1453);
xor U985 (N_985,N_644,N_840);
nand U986 (N_986,In_609,In_1153);
nand U987 (N_987,N_769,N_435);
nand U988 (N_988,N_871,N_797);
nand U989 (N_989,N_853,N_253);
nand U990 (N_990,In_619,In_38);
and U991 (N_991,N_396,N_65);
nand U992 (N_992,N_857,N_869);
nor U993 (N_993,N_150,N_583);
and U994 (N_994,In_956,N_890);
nand U995 (N_995,N_860,In_835);
xor U996 (N_996,In_571,N_501);
or U997 (N_997,In_1295,In_134);
xor U998 (N_998,In_73,N_171);
xor U999 (N_999,In_822,In_718);
or U1000 (N_1000,N_212,In_482);
nand U1001 (N_1001,In_1279,N_346);
or U1002 (N_1002,N_795,N_893);
nand U1003 (N_1003,N_206,N_875);
nand U1004 (N_1004,N_195,In_753);
nand U1005 (N_1005,In_736,N_831);
nor U1006 (N_1006,N_112,In_1213);
nor U1007 (N_1007,N_858,N_573);
xor U1008 (N_1008,N_802,In_790);
or U1009 (N_1009,In_677,N_864);
nand U1010 (N_1010,N_649,N_631);
nor U1011 (N_1011,N_861,N_686);
or U1012 (N_1012,N_877,N_350);
nand U1013 (N_1013,N_770,N_654);
nor U1014 (N_1014,In_444,N_196);
nand U1015 (N_1015,N_51,N_862);
nand U1016 (N_1016,In_272,N_684);
xnor U1017 (N_1017,N_819,N_807);
nor U1018 (N_1018,In_612,N_476);
xor U1019 (N_1019,N_590,N_606);
or U1020 (N_1020,In_1049,N_607);
nand U1021 (N_1021,N_536,N_399);
or U1022 (N_1022,N_788,In_1381);
xor U1023 (N_1023,In_1111,In_228);
and U1024 (N_1024,N_789,N_311);
xor U1025 (N_1025,N_468,N_57);
nand U1026 (N_1026,In_710,In_1216);
nor U1027 (N_1027,N_793,N_888);
nand U1028 (N_1028,In_224,N_47);
xnor U1029 (N_1029,N_364,N_419);
nand U1030 (N_1030,In_45,N_487);
nand U1031 (N_1031,N_718,N_695);
nor U1032 (N_1032,In_1403,In_97);
or U1033 (N_1033,N_835,In_966);
and U1034 (N_1034,N_727,In_505);
nor U1035 (N_1035,In_727,In_1379);
or U1036 (N_1036,N_9,N_790);
nand U1037 (N_1037,N_93,N_470);
nor U1038 (N_1038,In_1349,N_899);
xor U1039 (N_1039,N_255,N_717);
xnor U1040 (N_1040,N_891,In_525);
and U1041 (N_1041,N_894,N_883);
xor U1042 (N_1042,N_505,N_799);
xnor U1043 (N_1043,N_680,N_775);
and U1044 (N_1044,In_1147,N_519);
or U1045 (N_1045,N_755,In_176);
xnor U1046 (N_1046,In_111,N_749);
xnor U1047 (N_1047,N_673,N_569);
nor U1048 (N_1048,N_589,N_564);
nor U1049 (N_1049,N_881,N_667);
xnor U1050 (N_1050,N_761,N_1038);
xnor U1051 (N_1051,N_847,In_261);
xnor U1052 (N_1052,In_687,In_942);
xor U1053 (N_1053,N_237,N_633);
or U1054 (N_1054,N_462,N_830);
nor U1055 (N_1055,N_870,In_1480);
and U1056 (N_1056,N_963,N_773);
or U1057 (N_1057,N_1010,N_922);
xor U1058 (N_1058,N_595,In_773);
or U1059 (N_1059,N_133,In_353);
and U1060 (N_1060,In_1133,In_521);
nor U1061 (N_1061,N_921,N_994);
nor U1062 (N_1062,In_398,N_655);
nor U1063 (N_1063,In_161,N_913);
nor U1064 (N_1064,N_521,N_848);
or U1065 (N_1065,N_537,N_849);
nor U1066 (N_1066,N_637,N_782);
xor U1067 (N_1067,In_685,N_98);
or U1068 (N_1068,N_318,N_1014);
or U1069 (N_1069,In_766,In_1067);
nand U1070 (N_1070,In_1157,N_868);
and U1071 (N_1071,N_608,N_995);
nand U1072 (N_1072,N_670,In_888);
nor U1073 (N_1073,In_374,In_560);
nor U1074 (N_1074,N_865,In_863);
xnor U1075 (N_1075,N_1028,N_392);
nor U1076 (N_1076,N_925,N_991);
nand U1077 (N_1077,N_572,In_1429);
xnor U1078 (N_1078,N_935,N_1040);
nor U1079 (N_1079,N_1011,In_63);
nor U1080 (N_1080,N_380,N_705);
xnor U1081 (N_1081,N_962,N_2);
nor U1082 (N_1082,N_927,N_845);
or U1083 (N_1083,In_605,N_1042);
and U1084 (N_1084,N_602,N_622);
nand U1085 (N_1085,N_534,N_939);
xor U1086 (N_1086,N_1037,In_458);
xor U1087 (N_1087,N_681,N_978);
or U1088 (N_1088,N_1044,N_996);
nor U1089 (N_1089,N_27,N_949);
nor U1090 (N_1090,N_643,N_453);
and U1091 (N_1091,In_783,N_716);
nor U1092 (N_1092,N_369,In_1347);
xnor U1093 (N_1093,N_901,N_337);
or U1094 (N_1094,N_972,N_993);
and U1095 (N_1095,In_1337,N_526);
or U1096 (N_1096,N_856,In_437);
or U1097 (N_1097,In_1261,N_940);
and U1098 (N_1098,N_955,In_587);
nand U1099 (N_1099,N_702,N_834);
and U1100 (N_1100,N_753,N_722);
xnor U1101 (N_1101,In_1493,N_765);
nand U1102 (N_1102,In_256,In_336);
nor U1103 (N_1103,N_309,N_950);
nand U1104 (N_1104,N_951,N_976);
and U1105 (N_1105,N_37,N_329);
and U1106 (N_1106,N_728,N_1017);
nor U1107 (N_1107,N_954,N_242);
nand U1108 (N_1108,N_965,N_768);
or U1109 (N_1109,In_411,N_711);
xor U1110 (N_1110,N_1004,N_832);
xor U1111 (N_1111,N_641,In_1288);
nand U1112 (N_1112,N_814,N_786);
and U1113 (N_1113,N_966,N_683);
nand U1114 (N_1114,N_137,N_792);
nand U1115 (N_1115,N_945,N_457);
nand U1116 (N_1116,N_720,N_838);
and U1117 (N_1117,N_1024,N_956);
and U1118 (N_1118,N_731,N_682);
nand U1119 (N_1119,In_1372,N_911);
xnor U1120 (N_1120,N_953,N_345);
and U1121 (N_1121,N_1039,N_760);
nand U1122 (N_1122,N_781,N_25);
or U1123 (N_1123,N_1025,In_139);
nand U1124 (N_1124,N_983,N_975);
or U1125 (N_1125,N_496,N_986);
and U1126 (N_1126,N_1000,N_1015);
or U1127 (N_1127,N_586,N_825);
xnor U1128 (N_1128,In_1448,In_846);
or U1129 (N_1129,N_516,In_1260);
and U1130 (N_1130,N_499,N_420);
xnor U1131 (N_1131,N_61,N_910);
and U1132 (N_1132,N_707,In_984);
nand U1133 (N_1133,In_366,N_1013);
xor U1134 (N_1134,N_970,N_227);
or U1135 (N_1135,N_884,N_931);
and U1136 (N_1136,N_114,N_816);
and U1137 (N_1137,N_997,N_600);
nor U1138 (N_1138,In_477,N_886);
nor U1139 (N_1139,N_261,N_842);
xor U1140 (N_1140,In_653,N_464);
and U1141 (N_1141,N_917,N_941);
nor U1142 (N_1142,N_909,N_905);
or U1143 (N_1143,N_843,In_526);
xnor U1144 (N_1144,N_937,N_535);
or U1145 (N_1145,In_864,In_963);
or U1146 (N_1146,In_513,N_403);
nor U1147 (N_1147,N_763,In_756);
or U1148 (N_1148,N_973,In_868);
or U1149 (N_1149,N_1033,N_999);
nor U1150 (N_1150,N_811,In_408);
and U1151 (N_1151,In_198,N_906);
xnor U1152 (N_1152,N_1002,N_449);
nand U1153 (N_1153,N_1029,N_916);
nor U1154 (N_1154,N_1008,N_1023);
xnor U1155 (N_1155,N_1031,In_385);
nand U1156 (N_1156,N_880,In_1071);
nor U1157 (N_1157,N_964,N_990);
nor U1158 (N_1158,N_238,In_49);
nor U1159 (N_1159,N_912,In_102);
nand U1160 (N_1160,N_734,N_923);
and U1161 (N_1161,N_800,N_696);
nor U1162 (N_1162,In_1245,N_977);
or U1163 (N_1163,N_791,N_361);
and U1164 (N_1164,N_226,N_41);
xor U1165 (N_1165,N_1020,In_856);
nor U1166 (N_1166,N_738,N_932);
xnor U1167 (N_1167,N_713,N_859);
xor U1168 (N_1168,N_1034,N_982);
nand U1169 (N_1169,In_194,N_592);
xnor U1170 (N_1170,N_1016,In_1143);
and U1171 (N_1171,N_998,N_946);
and U1172 (N_1172,N_605,N_1009);
and U1173 (N_1173,In_562,N_733);
nor U1174 (N_1174,N_709,N_985);
xor U1175 (N_1175,N_930,N_812);
xor U1176 (N_1176,N_815,N_915);
and U1177 (N_1177,In_239,N_640);
xor U1178 (N_1178,N_785,N_903);
nor U1179 (N_1179,In_689,N_751);
xor U1180 (N_1180,N_1012,N_1006);
nor U1181 (N_1181,N_693,N_567);
or U1182 (N_1182,N_904,N_704);
xnor U1183 (N_1183,N_1005,N_929);
xor U1184 (N_1184,In_682,In_1396);
nand U1185 (N_1185,N_593,N_296);
and U1186 (N_1186,N_758,N_1032);
or U1187 (N_1187,N_1046,N_959);
or U1188 (N_1188,In_614,N_882);
nor U1189 (N_1189,In_249,N_1022);
and U1190 (N_1190,N_635,In_70);
nand U1191 (N_1191,N_974,N_422);
and U1192 (N_1192,N_771,N_752);
and U1193 (N_1193,N_952,In_518);
xor U1194 (N_1194,In_8,N_161);
nor U1195 (N_1195,In_375,N_813);
nor U1196 (N_1196,In_843,N_669);
nor U1197 (N_1197,N_614,In_538);
or U1198 (N_1198,N_818,N_958);
nand U1199 (N_1199,N_988,In_206);
and U1200 (N_1200,N_497,N_710);
nor U1201 (N_1201,N_1099,N_598);
nor U1202 (N_1202,N_803,N_1131);
or U1203 (N_1203,N_987,N_1075);
nor U1204 (N_1204,N_826,N_798);
xnor U1205 (N_1205,N_1068,N_828);
and U1206 (N_1206,N_1019,N_1198);
nor U1207 (N_1207,N_1151,N_1062);
xnor U1208 (N_1208,N_1045,In_767);
nor U1209 (N_1209,In_852,N_1184);
nand U1210 (N_1210,In_953,N_1160);
nor U1211 (N_1211,N_678,In_796);
or U1212 (N_1212,N_1110,N_409);
nand U1213 (N_1213,N_413,N_1041);
xnor U1214 (N_1214,N_1088,N_1093);
and U1215 (N_1215,N_1105,N_1137);
or U1216 (N_1216,N_920,N_1187);
xnor U1217 (N_1217,N_1108,N_596);
nand U1218 (N_1218,N_1081,N_928);
and U1219 (N_1219,N_1084,In_25);
nand U1220 (N_1220,N_1123,N_407);
xor U1221 (N_1221,N_333,In_1294);
nand U1222 (N_1222,N_879,N_1167);
nand U1223 (N_1223,N_748,N_1116);
xnor U1224 (N_1224,In_16,N_1118);
xor U1225 (N_1225,N_523,N_1018);
nor U1226 (N_1226,N_742,N_646);
and U1227 (N_1227,N_1049,N_10);
xnor U1228 (N_1228,N_957,N_971);
nor U1229 (N_1229,In_404,N_902);
nand U1230 (N_1230,N_1078,N_1141);
or U1231 (N_1231,In_1217,N_1182);
and U1232 (N_1232,N_936,N_779);
nor U1233 (N_1233,N_892,N_736);
nand U1234 (N_1234,N_1197,N_1190);
nand U1235 (N_1235,N_1001,N_1098);
and U1236 (N_1236,N_1095,N_645);
xor U1237 (N_1237,N_827,In_1476);
nand U1238 (N_1238,N_1007,N_1097);
or U1239 (N_1239,N_947,N_498);
nand U1240 (N_1240,N_1067,N_967);
and U1241 (N_1241,N_1174,N_1134);
nor U1242 (N_1242,N_960,N_754);
nand U1243 (N_1243,N_948,N_427);
and U1244 (N_1244,N_1127,N_1194);
nand U1245 (N_1245,N_1180,N_1152);
nor U1246 (N_1246,N_1047,N_1079);
xor U1247 (N_1247,N_919,In_420);
xor U1248 (N_1248,In_31,N_1103);
or U1249 (N_1249,N_1063,N_1087);
or U1250 (N_1250,In_986,N_436);
or U1251 (N_1251,N_968,N_1129);
nor U1252 (N_1252,N_1113,N_1094);
nor U1253 (N_1253,N_914,N_944);
xnor U1254 (N_1254,N_1163,N_1133);
nand U1255 (N_1255,N_1050,N_1173);
and U1256 (N_1256,N_1156,N_624);
nand U1257 (N_1257,N_1119,N_1193);
and U1258 (N_1258,N_1043,N_1125);
nor U1259 (N_1259,In_1046,N_766);
or U1260 (N_1260,N_1052,N_1145);
nor U1261 (N_1261,N_1055,N_867);
and U1262 (N_1262,In_1384,N_349);
nand U1263 (N_1263,N_1148,N_725);
or U1264 (N_1264,In_192,N_1195);
nand U1265 (N_1265,N_873,N_1053);
nor U1266 (N_1266,N_1083,N_924);
or U1267 (N_1267,N_1117,N_1085);
nor U1268 (N_1268,N_777,N_458);
or U1269 (N_1269,N_591,In_771);
xnor U1270 (N_1270,N_918,N_1090);
xnor U1271 (N_1271,N_1082,In_4);
and U1272 (N_1272,N_1107,N_1128);
xor U1273 (N_1273,N_1056,In_1386);
xnor U1274 (N_1274,N_1092,N_1199);
and U1275 (N_1275,N_1153,In_96);
or U1276 (N_1276,N_1070,N_1142);
xnor U1277 (N_1277,In_359,N_1166);
nand U1278 (N_1278,N_984,N_1077);
nand U1279 (N_1279,N_1066,N_1178);
and U1280 (N_1280,N_730,N_1136);
nor U1281 (N_1281,N_907,N_1074);
and U1282 (N_1282,In_1430,N_1189);
or U1283 (N_1283,N_1030,N_1181);
and U1284 (N_1284,N_1072,In_1123);
nand U1285 (N_1285,N_1191,N_767);
or U1286 (N_1286,N_1158,N_1057);
and U1287 (N_1287,In_1082,In_1454);
or U1288 (N_1288,N_980,N_1112);
xor U1289 (N_1289,N_1149,N_855);
nand U1290 (N_1290,In_1173,N_801);
nor U1291 (N_1291,In_390,N_1144);
and U1292 (N_1292,N_934,N_872);
nor U1293 (N_1293,N_1157,N_1138);
xnor U1294 (N_1294,N_619,In_656);
xnor U1295 (N_1295,N_900,N_1101);
nor U1296 (N_1296,N_969,N_1104);
and U1297 (N_1297,N_1143,N_1132);
or U1298 (N_1298,N_1135,N_1076);
or U1299 (N_1299,N_1080,N_981);
nand U1300 (N_1300,N_938,N_1051);
xnor U1301 (N_1301,N_451,N_1027);
and U1302 (N_1302,N_908,N_1086);
nand U1303 (N_1303,N_657,N_1186);
nand U1304 (N_1304,N_1188,N_1124);
nor U1305 (N_1305,N_1121,N_1171);
xor U1306 (N_1306,N_1089,N_1176);
nand U1307 (N_1307,N_1146,N_1073);
or U1308 (N_1308,N_1003,In_47);
xnor U1309 (N_1309,N_1061,N_1120);
nand U1310 (N_1310,In_1283,N_1026);
nand U1311 (N_1311,N_1036,N_1159);
nor U1312 (N_1312,N_1164,N_989);
and U1313 (N_1313,N_1059,N_1058);
xor U1314 (N_1314,In_1069,N_1155);
nor U1315 (N_1315,N_1165,N_1069);
nor U1316 (N_1316,N_1175,N_810);
or U1317 (N_1317,N_1048,N_1071);
nor U1318 (N_1318,N_609,N_264);
and U1319 (N_1319,N_1179,N_1021);
nand U1320 (N_1320,N_1147,N_1106);
nand U1321 (N_1321,N_1115,N_942);
nor U1322 (N_1322,N_1064,N_1169);
and U1323 (N_1323,N_1196,N_817);
nand U1324 (N_1324,N_783,N_1172);
and U1325 (N_1325,N_809,N_787);
or U1326 (N_1326,N_1114,N_992);
or U1327 (N_1327,In_577,N_1150);
nand U1328 (N_1328,N_1109,N_1170);
nand U1329 (N_1329,N_1139,N_1111);
or U1330 (N_1330,In_1000,N_833);
xnor U1331 (N_1331,N_1091,In_3);
nand U1332 (N_1332,N_1183,N_1122);
nor U1333 (N_1333,N_1126,N_747);
nand U1334 (N_1334,N_926,In_1128);
nand U1335 (N_1335,In_1466,N_1054);
nand U1336 (N_1336,N_1192,N_1154);
nor U1337 (N_1337,N_1130,In_572);
and U1338 (N_1338,N_961,N_77);
and U1339 (N_1339,N_698,N_1100);
nor U1340 (N_1340,N_1168,N_1185);
nand U1341 (N_1341,N_1102,N_1177);
xnor U1342 (N_1342,N_979,N_1162);
xnor U1343 (N_1343,N_1140,In_1471);
and U1344 (N_1344,In_627,N_866);
nand U1345 (N_1345,N_1035,N_943);
or U1346 (N_1346,N_1161,N_933);
nand U1347 (N_1347,N_1096,N_561);
and U1348 (N_1348,N_1060,N_117);
xnor U1349 (N_1349,N_658,N_1065);
xor U1350 (N_1350,N_1205,N_1342);
nor U1351 (N_1351,N_1287,N_1224);
and U1352 (N_1352,N_1264,N_1311);
and U1353 (N_1353,N_1253,N_1320);
nand U1354 (N_1354,N_1252,N_1209);
xor U1355 (N_1355,N_1312,N_1307);
nand U1356 (N_1356,N_1297,N_1200);
and U1357 (N_1357,N_1304,N_1243);
xor U1358 (N_1358,N_1267,N_1282);
xnor U1359 (N_1359,N_1214,N_1201);
or U1360 (N_1360,N_1303,N_1309);
nand U1361 (N_1361,N_1268,N_1315);
or U1362 (N_1362,N_1285,N_1278);
nor U1363 (N_1363,N_1247,N_1223);
nor U1364 (N_1364,N_1263,N_1251);
nand U1365 (N_1365,N_1241,N_1272);
and U1366 (N_1366,N_1301,N_1299);
nor U1367 (N_1367,N_1244,N_1273);
nand U1368 (N_1368,N_1237,N_1305);
and U1369 (N_1369,N_1226,N_1219);
or U1370 (N_1370,N_1333,N_1227);
and U1371 (N_1371,N_1292,N_1330);
nor U1372 (N_1372,N_1298,N_1323);
or U1373 (N_1373,N_1275,N_1274);
nor U1374 (N_1374,N_1348,N_1215);
and U1375 (N_1375,N_1208,N_1239);
nand U1376 (N_1376,N_1283,N_1341);
xnor U1377 (N_1377,N_1344,N_1257);
and U1378 (N_1378,N_1313,N_1216);
nand U1379 (N_1379,N_1322,N_1347);
nor U1380 (N_1380,N_1321,N_1254);
nor U1381 (N_1381,N_1334,N_1220);
nor U1382 (N_1382,N_1221,N_1233);
or U1383 (N_1383,N_1345,N_1336);
nand U1384 (N_1384,N_1255,N_1302);
xnor U1385 (N_1385,N_1249,N_1256);
nand U1386 (N_1386,N_1248,N_1235);
xor U1387 (N_1387,N_1225,N_1232);
or U1388 (N_1388,N_1324,N_1335);
and U1389 (N_1389,N_1266,N_1250);
and U1390 (N_1390,N_1259,N_1217);
or U1391 (N_1391,N_1337,N_1206);
nor U1392 (N_1392,N_1218,N_1343);
and U1393 (N_1393,N_1294,N_1242);
nor U1394 (N_1394,N_1314,N_1271);
or U1395 (N_1395,N_1318,N_1207);
and U1396 (N_1396,N_1306,N_1291);
or U1397 (N_1397,N_1210,N_1293);
and U1398 (N_1398,N_1325,N_1261);
or U1399 (N_1399,N_1228,N_1319);
nand U1400 (N_1400,N_1203,N_1234);
and U1401 (N_1401,N_1308,N_1331);
and U1402 (N_1402,N_1310,N_1276);
and U1403 (N_1403,N_1260,N_1346);
nor U1404 (N_1404,N_1230,N_1280);
and U1405 (N_1405,N_1326,N_1349);
and U1406 (N_1406,N_1258,N_1317);
nor U1407 (N_1407,N_1213,N_1202);
xor U1408 (N_1408,N_1240,N_1245);
or U1409 (N_1409,N_1269,N_1231);
nor U1410 (N_1410,N_1238,N_1300);
xor U1411 (N_1411,N_1288,N_1327);
and U1412 (N_1412,N_1329,N_1246);
or U1413 (N_1413,N_1279,N_1290);
and U1414 (N_1414,N_1265,N_1340);
nand U1415 (N_1415,N_1339,N_1204);
and U1416 (N_1416,N_1270,N_1296);
nand U1417 (N_1417,N_1328,N_1229);
or U1418 (N_1418,N_1289,N_1236);
or U1419 (N_1419,N_1316,N_1284);
nor U1420 (N_1420,N_1281,N_1211);
nand U1421 (N_1421,N_1295,N_1277);
or U1422 (N_1422,N_1262,N_1222);
nor U1423 (N_1423,N_1212,N_1286);
and U1424 (N_1424,N_1332,N_1338);
xnor U1425 (N_1425,N_1259,N_1219);
or U1426 (N_1426,N_1210,N_1213);
nand U1427 (N_1427,N_1325,N_1203);
and U1428 (N_1428,N_1236,N_1201);
xor U1429 (N_1429,N_1284,N_1334);
or U1430 (N_1430,N_1270,N_1339);
and U1431 (N_1431,N_1340,N_1243);
xor U1432 (N_1432,N_1302,N_1287);
nand U1433 (N_1433,N_1317,N_1334);
or U1434 (N_1434,N_1345,N_1301);
nand U1435 (N_1435,N_1265,N_1257);
or U1436 (N_1436,N_1237,N_1205);
xor U1437 (N_1437,N_1232,N_1256);
xnor U1438 (N_1438,N_1262,N_1231);
xor U1439 (N_1439,N_1226,N_1248);
and U1440 (N_1440,N_1265,N_1234);
and U1441 (N_1441,N_1309,N_1347);
nand U1442 (N_1442,N_1282,N_1258);
nor U1443 (N_1443,N_1297,N_1305);
and U1444 (N_1444,N_1204,N_1270);
nand U1445 (N_1445,N_1265,N_1301);
nor U1446 (N_1446,N_1255,N_1339);
nor U1447 (N_1447,N_1324,N_1329);
and U1448 (N_1448,N_1278,N_1206);
and U1449 (N_1449,N_1291,N_1283);
nor U1450 (N_1450,N_1326,N_1308);
nand U1451 (N_1451,N_1306,N_1261);
xnor U1452 (N_1452,N_1213,N_1263);
or U1453 (N_1453,N_1262,N_1239);
and U1454 (N_1454,N_1321,N_1337);
and U1455 (N_1455,N_1308,N_1311);
xor U1456 (N_1456,N_1238,N_1266);
and U1457 (N_1457,N_1237,N_1214);
nand U1458 (N_1458,N_1264,N_1334);
or U1459 (N_1459,N_1341,N_1247);
or U1460 (N_1460,N_1323,N_1243);
nor U1461 (N_1461,N_1332,N_1315);
or U1462 (N_1462,N_1213,N_1297);
nand U1463 (N_1463,N_1228,N_1303);
nor U1464 (N_1464,N_1206,N_1313);
nand U1465 (N_1465,N_1204,N_1206);
nand U1466 (N_1466,N_1321,N_1219);
nand U1467 (N_1467,N_1229,N_1212);
or U1468 (N_1468,N_1223,N_1231);
or U1469 (N_1469,N_1304,N_1276);
or U1470 (N_1470,N_1334,N_1214);
nor U1471 (N_1471,N_1215,N_1319);
nand U1472 (N_1472,N_1307,N_1203);
and U1473 (N_1473,N_1300,N_1306);
or U1474 (N_1474,N_1248,N_1218);
nand U1475 (N_1475,N_1202,N_1272);
or U1476 (N_1476,N_1263,N_1290);
nand U1477 (N_1477,N_1222,N_1307);
nor U1478 (N_1478,N_1312,N_1349);
and U1479 (N_1479,N_1283,N_1244);
or U1480 (N_1480,N_1266,N_1331);
nor U1481 (N_1481,N_1236,N_1337);
and U1482 (N_1482,N_1338,N_1236);
nand U1483 (N_1483,N_1214,N_1257);
nor U1484 (N_1484,N_1212,N_1221);
and U1485 (N_1485,N_1298,N_1292);
and U1486 (N_1486,N_1253,N_1274);
and U1487 (N_1487,N_1286,N_1304);
nand U1488 (N_1488,N_1250,N_1212);
nand U1489 (N_1489,N_1337,N_1318);
or U1490 (N_1490,N_1283,N_1267);
xor U1491 (N_1491,N_1280,N_1210);
and U1492 (N_1492,N_1281,N_1324);
nor U1493 (N_1493,N_1308,N_1280);
and U1494 (N_1494,N_1310,N_1339);
or U1495 (N_1495,N_1240,N_1258);
and U1496 (N_1496,N_1272,N_1286);
or U1497 (N_1497,N_1341,N_1216);
or U1498 (N_1498,N_1213,N_1209);
nand U1499 (N_1499,N_1304,N_1310);
or U1500 (N_1500,N_1401,N_1448);
or U1501 (N_1501,N_1412,N_1354);
nand U1502 (N_1502,N_1389,N_1431);
nor U1503 (N_1503,N_1423,N_1413);
nand U1504 (N_1504,N_1368,N_1387);
xnor U1505 (N_1505,N_1445,N_1472);
xnor U1506 (N_1506,N_1393,N_1470);
nand U1507 (N_1507,N_1432,N_1415);
xnor U1508 (N_1508,N_1436,N_1484);
nor U1509 (N_1509,N_1363,N_1366);
nand U1510 (N_1510,N_1396,N_1481);
nand U1511 (N_1511,N_1360,N_1455);
or U1512 (N_1512,N_1380,N_1407);
xor U1513 (N_1513,N_1422,N_1438);
and U1514 (N_1514,N_1483,N_1365);
xnor U1515 (N_1515,N_1398,N_1495);
xnor U1516 (N_1516,N_1410,N_1493);
or U1517 (N_1517,N_1482,N_1463);
nand U1518 (N_1518,N_1477,N_1358);
nand U1519 (N_1519,N_1459,N_1461);
xor U1520 (N_1520,N_1375,N_1454);
xor U1521 (N_1521,N_1476,N_1384);
nor U1522 (N_1522,N_1429,N_1467);
and U1523 (N_1523,N_1386,N_1462);
nor U1524 (N_1524,N_1373,N_1428);
xor U1525 (N_1525,N_1486,N_1499);
xor U1526 (N_1526,N_1468,N_1390);
nor U1527 (N_1527,N_1394,N_1383);
and U1528 (N_1528,N_1460,N_1439);
xor U1529 (N_1529,N_1487,N_1426);
xnor U1530 (N_1530,N_1367,N_1496);
nor U1531 (N_1531,N_1492,N_1403);
and U1532 (N_1532,N_1414,N_1427);
and U1533 (N_1533,N_1433,N_1453);
nor U1534 (N_1534,N_1471,N_1379);
or U1535 (N_1535,N_1377,N_1374);
nand U1536 (N_1536,N_1489,N_1498);
nor U1537 (N_1537,N_1444,N_1408);
nand U1538 (N_1538,N_1469,N_1392);
xnor U1539 (N_1539,N_1376,N_1385);
and U1540 (N_1540,N_1418,N_1442);
nand U1541 (N_1541,N_1359,N_1355);
and U1542 (N_1542,N_1494,N_1420);
nor U1543 (N_1543,N_1399,N_1424);
or U1544 (N_1544,N_1443,N_1425);
or U1545 (N_1545,N_1441,N_1406);
and U1546 (N_1546,N_1488,N_1421);
or U1547 (N_1547,N_1369,N_1361);
nand U1548 (N_1548,N_1364,N_1362);
and U1549 (N_1549,N_1430,N_1464);
and U1550 (N_1550,N_1475,N_1419);
or U1551 (N_1551,N_1447,N_1409);
nand U1552 (N_1552,N_1457,N_1485);
and U1553 (N_1553,N_1350,N_1497);
nand U1554 (N_1554,N_1395,N_1351);
or U1555 (N_1555,N_1402,N_1440);
and U1556 (N_1556,N_1473,N_1490);
and U1557 (N_1557,N_1382,N_1491);
nor U1558 (N_1558,N_1411,N_1352);
or U1559 (N_1559,N_1356,N_1446);
or U1560 (N_1560,N_1397,N_1434);
and U1561 (N_1561,N_1474,N_1405);
and U1562 (N_1562,N_1435,N_1449);
or U1563 (N_1563,N_1357,N_1381);
xnor U1564 (N_1564,N_1451,N_1458);
or U1565 (N_1565,N_1456,N_1372);
or U1566 (N_1566,N_1388,N_1353);
nand U1567 (N_1567,N_1400,N_1404);
and U1568 (N_1568,N_1378,N_1452);
xnor U1569 (N_1569,N_1417,N_1478);
nor U1570 (N_1570,N_1370,N_1371);
or U1571 (N_1571,N_1465,N_1437);
nand U1572 (N_1572,N_1480,N_1416);
xnor U1573 (N_1573,N_1466,N_1479);
or U1574 (N_1574,N_1391,N_1450);
nand U1575 (N_1575,N_1429,N_1409);
and U1576 (N_1576,N_1390,N_1430);
nand U1577 (N_1577,N_1364,N_1404);
xor U1578 (N_1578,N_1381,N_1403);
xor U1579 (N_1579,N_1355,N_1471);
nand U1580 (N_1580,N_1419,N_1397);
or U1581 (N_1581,N_1373,N_1417);
xor U1582 (N_1582,N_1416,N_1490);
or U1583 (N_1583,N_1473,N_1453);
or U1584 (N_1584,N_1464,N_1411);
or U1585 (N_1585,N_1424,N_1395);
nor U1586 (N_1586,N_1485,N_1380);
xor U1587 (N_1587,N_1416,N_1411);
nor U1588 (N_1588,N_1483,N_1429);
and U1589 (N_1589,N_1491,N_1481);
xor U1590 (N_1590,N_1432,N_1355);
or U1591 (N_1591,N_1490,N_1427);
and U1592 (N_1592,N_1442,N_1455);
nand U1593 (N_1593,N_1367,N_1493);
nor U1594 (N_1594,N_1386,N_1468);
or U1595 (N_1595,N_1483,N_1455);
and U1596 (N_1596,N_1412,N_1400);
nor U1597 (N_1597,N_1383,N_1371);
nand U1598 (N_1598,N_1465,N_1452);
or U1599 (N_1599,N_1493,N_1421);
xnor U1600 (N_1600,N_1402,N_1387);
xnor U1601 (N_1601,N_1389,N_1416);
or U1602 (N_1602,N_1499,N_1419);
and U1603 (N_1603,N_1363,N_1447);
nor U1604 (N_1604,N_1400,N_1480);
xnor U1605 (N_1605,N_1402,N_1439);
or U1606 (N_1606,N_1376,N_1425);
or U1607 (N_1607,N_1467,N_1379);
nor U1608 (N_1608,N_1483,N_1396);
or U1609 (N_1609,N_1460,N_1466);
or U1610 (N_1610,N_1385,N_1487);
nor U1611 (N_1611,N_1487,N_1428);
xor U1612 (N_1612,N_1496,N_1406);
nand U1613 (N_1613,N_1481,N_1429);
or U1614 (N_1614,N_1454,N_1413);
nor U1615 (N_1615,N_1394,N_1453);
xnor U1616 (N_1616,N_1416,N_1405);
nand U1617 (N_1617,N_1361,N_1415);
xor U1618 (N_1618,N_1411,N_1442);
nor U1619 (N_1619,N_1406,N_1400);
nand U1620 (N_1620,N_1472,N_1385);
nor U1621 (N_1621,N_1414,N_1492);
and U1622 (N_1622,N_1353,N_1458);
xor U1623 (N_1623,N_1423,N_1440);
and U1624 (N_1624,N_1414,N_1499);
nand U1625 (N_1625,N_1485,N_1477);
xor U1626 (N_1626,N_1450,N_1492);
nand U1627 (N_1627,N_1462,N_1362);
and U1628 (N_1628,N_1426,N_1364);
nor U1629 (N_1629,N_1400,N_1362);
or U1630 (N_1630,N_1411,N_1365);
nor U1631 (N_1631,N_1421,N_1415);
xor U1632 (N_1632,N_1352,N_1381);
and U1633 (N_1633,N_1497,N_1487);
nand U1634 (N_1634,N_1492,N_1413);
or U1635 (N_1635,N_1387,N_1493);
nand U1636 (N_1636,N_1467,N_1394);
xnor U1637 (N_1637,N_1364,N_1480);
and U1638 (N_1638,N_1435,N_1425);
or U1639 (N_1639,N_1403,N_1475);
nand U1640 (N_1640,N_1473,N_1465);
and U1641 (N_1641,N_1466,N_1490);
nor U1642 (N_1642,N_1351,N_1418);
or U1643 (N_1643,N_1371,N_1491);
nor U1644 (N_1644,N_1399,N_1485);
xor U1645 (N_1645,N_1360,N_1363);
and U1646 (N_1646,N_1412,N_1451);
or U1647 (N_1647,N_1496,N_1364);
nand U1648 (N_1648,N_1441,N_1431);
and U1649 (N_1649,N_1464,N_1456);
nand U1650 (N_1650,N_1576,N_1561);
or U1651 (N_1651,N_1596,N_1524);
nor U1652 (N_1652,N_1566,N_1500);
nor U1653 (N_1653,N_1568,N_1646);
nor U1654 (N_1654,N_1599,N_1515);
nand U1655 (N_1655,N_1555,N_1570);
xnor U1656 (N_1656,N_1635,N_1548);
nand U1657 (N_1657,N_1569,N_1551);
nand U1658 (N_1658,N_1638,N_1534);
xor U1659 (N_1659,N_1542,N_1629);
xor U1660 (N_1660,N_1527,N_1601);
xor U1661 (N_1661,N_1628,N_1508);
xnor U1662 (N_1662,N_1545,N_1594);
nor U1663 (N_1663,N_1567,N_1642);
xnor U1664 (N_1664,N_1631,N_1510);
nand U1665 (N_1665,N_1640,N_1511);
and U1666 (N_1666,N_1528,N_1584);
xor U1667 (N_1667,N_1554,N_1507);
nand U1668 (N_1668,N_1615,N_1636);
nor U1669 (N_1669,N_1564,N_1532);
or U1670 (N_1670,N_1536,N_1563);
nand U1671 (N_1671,N_1603,N_1578);
and U1672 (N_1672,N_1505,N_1591);
or U1673 (N_1673,N_1553,N_1546);
nor U1674 (N_1674,N_1624,N_1621);
or U1675 (N_1675,N_1580,N_1643);
or U1676 (N_1676,N_1610,N_1611);
or U1677 (N_1677,N_1627,N_1588);
or U1678 (N_1678,N_1620,N_1618);
xnor U1679 (N_1679,N_1521,N_1535);
and U1680 (N_1680,N_1587,N_1647);
or U1681 (N_1681,N_1529,N_1623);
nand U1682 (N_1682,N_1523,N_1522);
xnor U1683 (N_1683,N_1600,N_1541);
nor U1684 (N_1684,N_1614,N_1619);
xor U1685 (N_1685,N_1537,N_1519);
nor U1686 (N_1686,N_1612,N_1562);
or U1687 (N_1687,N_1645,N_1609);
or U1688 (N_1688,N_1598,N_1582);
xor U1689 (N_1689,N_1649,N_1581);
nand U1690 (N_1690,N_1543,N_1616);
xnor U1691 (N_1691,N_1574,N_1533);
and U1692 (N_1692,N_1589,N_1547);
xnor U1693 (N_1693,N_1602,N_1625);
nand U1694 (N_1694,N_1632,N_1549);
nand U1695 (N_1695,N_1552,N_1595);
nand U1696 (N_1696,N_1622,N_1592);
nor U1697 (N_1697,N_1514,N_1590);
nor U1698 (N_1698,N_1613,N_1501);
nor U1699 (N_1699,N_1558,N_1509);
nand U1700 (N_1700,N_1641,N_1556);
xnor U1701 (N_1701,N_1637,N_1512);
nor U1702 (N_1702,N_1506,N_1586);
and U1703 (N_1703,N_1504,N_1513);
nor U1704 (N_1704,N_1626,N_1559);
xnor U1705 (N_1705,N_1585,N_1571);
or U1706 (N_1706,N_1560,N_1630);
nand U1707 (N_1707,N_1517,N_1540);
nand U1708 (N_1708,N_1577,N_1572);
or U1709 (N_1709,N_1579,N_1593);
or U1710 (N_1710,N_1633,N_1573);
or U1711 (N_1711,N_1538,N_1607);
and U1712 (N_1712,N_1516,N_1525);
nand U1713 (N_1713,N_1597,N_1606);
and U1714 (N_1714,N_1605,N_1550);
or U1715 (N_1715,N_1604,N_1530);
or U1716 (N_1716,N_1526,N_1608);
nand U1717 (N_1717,N_1583,N_1502);
or U1718 (N_1718,N_1648,N_1634);
xnor U1719 (N_1719,N_1617,N_1639);
or U1720 (N_1720,N_1539,N_1644);
nand U1721 (N_1721,N_1518,N_1557);
or U1722 (N_1722,N_1520,N_1575);
xnor U1723 (N_1723,N_1565,N_1503);
nor U1724 (N_1724,N_1531,N_1544);
nor U1725 (N_1725,N_1611,N_1642);
nand U1726 (N_1726,N_1622,N_1606);
nand U1727 (N_1727,N_1562,N_1619);
nor U1728 (N_1728,N_1516,N_1606);
xor U1729 (N_1729,N_1500,N_1561);
or U1730 (N_1730,N_1623,N_1537);
nand U1731 (N_1731,N_1562,N_1566);
or U1732 (N_1732,N_1647,N_1502);
xor U1733 (N_1733,N_1528,N_1581);
or U1734 (N_1734,N_1620,N_1595);
nand U1735 (N_1735,N_1540,N_1593);
nor U1736 (N_1736,N_1606,N_1571);
or U1737 (N_1737,N_1504,N_1550);
and U1738 (N_1738,N_1550,N_1587);
xor U1739 (N_1739,N_1574,N_1568);
nand U1740 (N_1740,N_1521,N_1607);
and U1741 (N_1741,N_1552,N_1553);
nand U1742 (N_1742,N_1643,N_1624);
or U1743 (N_1743,N_1617,N_1599);
and U1744 (N_1744,N_1522,N_1554);
xor U1745 (N_1745,N_1632,N_1595);
and U1746 (N_1746,N_1575,N_1564);
and U1747 (N_1747,N_1628,N_1566);
nand U1748 (N_1748,N_1547,N_1530);
xnor U1749 (N_1749,N_1582,N_1618);
nand U1750 (N_1750,N_1649,N_1576);
nor U1751 (N_1751,N_1556,N_1569);
and U1752 (N_1752,N_1568,N_1537);
nor U1753 (N_1753,N_1509,N_1541);
nand U1754 (N_1754,N_1582,N_1570);
nand U1755 (N_1755,N_1541,N_1531);
nand U1756 (N_1756,N_1520,N_1599);
or U1757 (N_1757,N_1634,N_1529);
nand U1758 (N_1758,N_1604,N_1540);
or U1759 (N_1759,N_1638,N_1574);
xnor U1760 (N_1760,N_1557,N_1551);
xor U1761 (N_1761,N_1526,N_1564);
nand U1762 (N_1762,N_1620,N_1633);
and U1763 (N_1763,N_1543,N_1591);
and U1764 (N_1764,N_1518,N_1561);
nor U1765 (N_1765,N_1508,N_1536);
and U1766 (N_1766,N_1511,N_1594);
nand U1767 (N_1767,N_1558,N_1548);
xor U1768 (N_1768,N_1570,N_1527);
nand U1769 (N_1769,N_1516,N_1563);
or U1770 (N_1770,N_1526,N_1558);
nor U1771 (N_1771,N_1634,N_1629);
or U1772 (N_1772,N_1574,N_1603);
nor U1773 (N_1773,N_1618,N_1571);
nor U1774 (N_1774,N_1513,N_1547);
nand U1775 (N_1775,N_1622,N_1604);
and U1776 (N_1776,N_1577,N_1637);
xnor U1777 (N_1777,N_1592,N_1516);
nand U1778 (N_1778,N_1580,N_1553);
and U1779 (N_1779,N_1579,N_1523);
and U1780 (N_1780,N_1632,N_1509);
xor U1781 (N_1781,N_1575,N_1587);
or U1782 (N_1782,N_1524,N_1545);
xor U1783 (N_1783,N_1638,N_1565);
nand U1784 (N_1784,N_1605,N_1616);
nand U1785 (N_1785,N_1642,N_1635);
nand U1786 (N_1786,N_1545,N_1519);
or U1787 (N_1787,N_1628,N_1607);
and U1788 (N_1788,N_1537,N_1631);
nor U1789 (N_1789,N_1562,N_1575);
nand U1790 (N_1790,N_1627,N_1622);
or U1791 (N_1791,N_1575,N_1648);
nand U1792 (N_1792,N_1592,N_1582);
nand U1793 (N_1793,N_1548,N_1514);
or U1794 (N_1794,N_1536,N_1522);
nor U1795 (N_1795,N_1594,N_1553);
xor U1796 (N_1796,N_1555,N_1575);
nor U1797 (N_1797,N_1636,N_1641);
and U1798 (N_1798,N_1533,N_1534);
xor U1799 (N_1799,N_1617,N_1528);
nand U1800 (N_1800,N_1773,N_1696);
and U1801 (N_1801,N_1677,N_1685);
nand U1802 (N_1802,N_1704,N_1799);
nand U1803 (N_1803,N_1774,N_1686);
xnor U1804 (N_1804,N_1695,N_1690);
or U1805 (N_1805,N_1721,N_1660);
nor U1806 (N_1806,N_1666,N_1675);
and U1807 (N_1807,N_1658,N_1765);
xor U1808 (N_1808,N_1767,N_1705);
nor U1809 (N_1809,N_1661,N_1698);
nand U1810 (N_1810,N_1668,N_1679);
and U1811 (N_1811,N_1688,N_1709);
nor U1812 (N_1812,N_1735,N_1795);
nand U1813 (N_1813,N_1700,N_1790);
nor U1814 (N_1814,N_1723,N_1726);
and U1815 (N_1815,N_1663,N_1716);
nand U1816 (N_1816,N_1650,N_1654);
and U1817 (N_1817,N_1741,N_1775);
and U1818 (N_1818,N_1737,N_1656);
xnor U1819 (N_1819,N_1719,N_1669);
nand U1820 (N_1820,N_1713,N_1699);
or U1821 (N_1821,N_1702,N_1733);
xor U1822 (N_1822,N_1672,N_1744);
nor U1823 (N_1823,N_1732,N_1693);
or U1824 (N_1824,N_1710,N_1760);
nand U1825 (N_1825,N_1667,N_1684);
and U1826 (N_1826,N_1791,N_1736);
nand U1827 (N_1827,N_1683,N_1752);
xor U1828 (N_1828,N_1780,N_1772);
xnor U1829 (N_1829,N_1758,N_1725);
xor U1830 (N_1830,N_1708,N_1793);
nor U1831 (N_1831,N_1764,N_1792);
nor U1832 (N_1832,N_1715,N_1755);
nor U1833 (N_1833,N_1787,N_1757);
nor U1834 (N_1834,N_1694,N_1697);
or U1835 (N_1835,N_1753,N_1712);
and U1836 (N_1836,N_1729,N_1680);
or U1837 (N_1837,N_1745,N_1771);
and U1838 (N_1838,N_1797,N_1794);
or U1839 (N_1839,N_1769,N_1749);
and U1840 (N_1840,N_1730,N_1671);
or U1841 (N_1841,N_1783,N_1662);
nand U1842 (N_1842,N_1653,N_1740);
or U1843 (N_1843,N_1651,N_1652);
and U1844 (N_1844,N_1766,N_1657);
xnor U1845 (N_1845,N_1786,N_1743);
xor U1846 (N_1846,N_1659,N_1748);
and U1847 (N_1847,N_1718,N_1689);
xor U1848 (N_1848,N_1701,N_1761);
and U1849 (N_1849,N_1776,N_1756);
and U1850 (N_1850,N_1687,N_1751);
nor U1851 (N_1851,N_1750,N_1739);
or U1852 (N_1852,N_1682,N_1763);
nand U1853 (N_1853,N_1691,N_1711);
or U1854 (N_1854,N_1728,N_1788);
nor U1855 (N_1855,N_1742,N_1717);
nor U1856 (N_1856,N_1678,N_1759);
xor U1857 (N_1857,N_1727,N_1768);
nor U1858 (N_1858,N_1778,N_1681);
and U1859 (N_1859,N_1714,N_1747);
or U1860 (N_1860,N_1785,N_1738);
xor U1861 (N_1861,N_1798,N_1777);
xor U1862 (N_1862,N_1731,N_1707);
or U1863 (N_1863,N_1796,N_1692);
nand U1864 (N_1864,N_1655,N_1703);
xnor U1865 (N_1865,N_1784,N_1781);
xnor U1866 (N_1866,N_1665,N_1724);
xnor U1867 (N_1867,N_1664,N_1779);
and U1868 (N_1868,N_1734,N_1770);
xnor U1869 (N_1869,N_1789,N_1670);
xor U1870 (N_1870,N_1754,N_1674);
or U1871 (N_1871,N_1762,N_1676);
xnor U1872 (N_1872,N_1673,N_1782);
xnor U1873 (N_1873,N_1720,N_1722);
nor U1874 (N_1874,N_1706,N_1746);
xnor U1875 (N_1875,N_1714,N_1796);
or U1876 (N_1876,N_1786,N_1674);
or U1877 (N_1877,N_1655,N_1666);
or U1878 (N_1878,N_1773,N_1714);
nor U1879 (N_1879,N_1777,N_1787);
nand U1880 (N_1880,N_1689,N_1668);
and U1881 (N_1881,N_1651,N_1791);
and U1882 (N_1882,N_1707,N_1706);
xor U1883 (N_1883,N_1667,N_1677);
or U1884 (N_1884,N_1798,N_1757);
nand U1885 (N_1885,N_1795,N_1759);
nor U1886 (N_1886,N_1701,N_1691);
nor U1887 (N_1887,N_1761,N_1756);
or U1888 (N_1888,N_1750,N_1765);
xor U1889 (N_1889,N_1701,N_1673);
or U1890 (N_1890,N_1656,N_1748);
or U1891 (N_1891,N_1689,N_1757);
and U1892 (N_1892,N_1743,N_1748);
or U1893 (N_1893,N_1692,N_1651);
or U1894 (N_1894,N_1714,N_1666);
or U1895 (N_1895,N_1792,N_1680);
nor U1896 (N_1896,N_1703,N_1671);
nor U1897 (N_1897,N_1762,N_1763);
xnor U1898 (N_1898,N_1784,N_1703);
xor U1899 (N_1899,N_1710,N_1731);
and U1900 (N_1900,N_1767,N_1656);
nand U1901 (N_1901,N_1776,N_1768);
nand U1902 (N_1902,N_1753,N_1673);
and U1903 (N_1903,N_1787,N_1756);
nand U1904 (N_1904,N_1714,N_1727);
and U1905 (N_1905,N_1711,N_1701);
xor U1906 (N_1906,N_1779,N_1773);
nand U1907 (N_1907,N_1797,N_1657);
xor U1908 (N_1908,N_1736,N_1707);
nor U1909 (N_1909,N_1693,N_1769);
xor U1910 (N_1910,N_1675,N_1700);
xor U1911 (N_1911,N_1748,N_1745);
xor U1912 (N_1912,N_1700,N_1667);
or U1913 (N_1913,N_1740,N_1680);
or U1914 (N_1914,N_1789,N_1701);
nor U1915 (N_1915,N_1737,N_1681);
xnor U1916 (N_1916,N_1774,N_1667);
and U1917 (N_1917,N_1745,N_1708);
or U1918 (N_1918,N_1748,N_1709);
xnor U1919 (N_1919,N_1660,N_1751);
xor U1920 (N_1920,N_1671,N_1775);
and U1921 (N_1921,N_1763,N_1681);
and U1922 (N_1922,N_1716,N_1667);
or U1923 (N_1923,N_1760,N_1762);
nand U1924 (N_1924,N_1725,N_1795);
nand U1925 (N_1925,N_1680,N_1783);
nand U1926 (N_1926,N_1651,N_1672);
or U1927 (N_1927,N_1651,N_1709);
xnor U1928 (N_1928,N_1767,N_1765);
and U1929 (N_1929,N_1737,N_1731);
nor U1930 (N_1930,N_1715,N_1690);
or U1931 (N_1931,N_1666,N_1783);
or U1932 (N_1932,N_1786,N_1741);
and U1933 (N_1933,N_1726,N_1768);
nor U1934 (N_1934,N_1708,N_1682);
and U1935 (N_1935,N_1689,N_1675);
and U1936 (N_1936,N_1672,N_1777);
xnor U1937 (N_1937,N_1653,N_1773);
xnor U1938 (N_1938,N_1703,N_1650);
and U1939 (N_1939,N_1673,N_1757);
nor U1940 (N_1940,N_1765,N_1715);
xnor U1941 (N_1941,N_1671,N_1738);
nand U1942 (N_1942,N_1792,N_1654);
nand U1943 (N_1943,N_1766,N_1737);
and U1944 (N_1944,N_1660,N_1681);
xor U1945 (N_1945,N_1653,N_1720);
xor U1946 (N_1946,N_1769,N_1735);
or U1947 (N_1947,N_1788,N_1767);
and U1948 (N_1948,N_1768,N_1787);
and U1949 (N_1949,N_1721,N_1675);
xor U1950 (N_1950,N_1843,N_1906);
xor U1951 (N_1951,N_1856,N_1886);
nor U1952 (N_1952,N_1804,N_1845);
xnor U1953 (N_1953,N_1897,N_1880);
xor U1954 (N_1954,N_1944,N_1914);
nor U1955 (N_1955,N_1803,N_1852);
or U1956 (N_1956,N_1817,N_1891);
nand U1957 (N_1957,N_1801,N_1899);
nand U1958 (N_1958,N_1908,N_1802);
nand U1959 (N_1959,N_1830,N_1858);
and U1960 (N_1960,N_1820,N_1828);
nor U1961 (N_1961,N_1869,N_1824);
or U1962 (N_1962,N_1805,N_1919);
or U1963 (N_1963,N_1943,N_1923);
nor U1964 (N_1964,N_1825,N_1933);
nor U1965 (N_1965,N_1862,N_1833);
nor U1966 (N_1966,N_1827,N_1829);
nand U1967 (N_1967,N_1903,N_1889);
nor U1968 (N_1968,N_1866,N_1922);
nand U1969 (N_1969,N_1909,N_1915);
xnor U1970 (N_1970,N_1859,N_1815);
nor U1971 (N_1971,N_1935,N_1940);
nand U1972 (N_1972,N_1882,N_1892);
or U1973 (N_1973,N_1912,N_1808);
and U1974 (N_1974,N_1870,N_1902);
nand U1975 (N_1975,N_1885,N_1879);
xor U1976 (N_1976,N_1871,N_1839);
xor U1977 (N_1977,N_1890,N_1835);
and U1978 (N_1978,N_1937,N_1800);
nand U1979 (N_1979,N_1894,N_1920);
or U1980 (N_1980,N_1924,N_1874);
xor U1981 (N_1981,N_1900,N_1818);
nor U1982 (N_1982,N_1934,N_1868);
and U1983 (N_1983,N_1887,N_1911);
and U1984 (N_1984,N_1893,N_1939);
nor U1985 (N_1985,N_1930,N_1842);
and U1986 (N_1986,N_1855,N_1905);
nand U1987 (N_1987,N_1901,N_1936);
xor U1988 (N_1988,N_1844,N_1819);
nor U1989 (N_1989,N_1896,N_1836);
and U1990 (N_1990,N_1875,N_1916);
or U1991 (N_1991,N_1929,N_1888);
xor U1992 (N_1992,N_1910,N_1898);
or U1993 (N_1993,N_1816,N_1895);
xnor U1994 (N_1994,N_1877,N_1913);
xnor U1995 (N_1995,N_1813,N_1851);
xor U1996 (N_1996,N_1942,N_1907);
or U1997 (N_1997,N_1904,N_1861);
nand U1998 (N_1998,N_1867,N_1947);
nor U1999 (N_1999,N_1812,N_1848);
or U2000 (N_2000,N_1850,N_1823);
and U2001 (N_2001,N_1883,N_1928);
nand U2002 (N_2002,N_1821,N_1873);
and U2003 (N_2003,N_1872,N_1921);
nor U2004 (N_2004,N_1837,N_1941);
nand U2005 (N_2005,N_1810,N_1925);
nand U2006 (N_2006,N_1949,N_1807);
nand U2007 (N_2007,N_1841,N_1945);
or U2008 (N_2008,N_1932,N_1857);
nor U2009 (N_2009,N_1865,N_1881);
xnor U2010 (N_2010,N_1948,N_1832);
xnor U2011 (N_2011,N_1926,N_1840);
or U2012 (N_2012,N_1864,N_1814);
or U2013 (N_2013,N_1938,N_1838);
nand U2014 (N_2014,N_1826,N_1917);
nor U2015 (N_2015,N_1809,N_1849);
nand U2016 (N_2016,N_1847,N_1854);
and U2017 (N_2017,N_1884,N_1927);
nor U2018 (N_2018,N_1946,N_1822);
nor U2019 (N_2019,N_1931,N_1834);
xnor U2020 (N_2020,N_1853,N_1811);
xnor U2021 (N_2021,N_1831,N_1846);
or U2022 (N_2022,N_1860,N_1878);
nand U2023 (N_2023,N_1918,N_1863);
xnor U2024 (N_2024,N_1806,N_1876);
xnor U2025 (N_2025,N_1948,N_1867);
nand U2026 (N_2026,N_1890,N_1945);
and U2027 (N_2027,N_1814,N_1836);
or U2028 (N_2028,N_1939,N_1936);
or U2029 (N_2029,N_1832,N_1919);
or U2030 (N_2030,N_1887,N_1843);
xor U2031 (N_2031,N_1855,N_1851);
and U2032 (N_2032,N_1940,N_1834);
nor U2033 (N_2033,N_1829,N_1816);
and U2034 (N_2034,N_1896,N_1807);
and U2035 (N_2035,N_1906,N_1949);
or U2036 (N_2036,N_1824,N_1840);
or U2037 (N_2037,N_1877,N_1892);
xor U2038 (N_2038,N_1898,N_1923);
and U2039 (N_2039,N_1921,N_1814);
nand U2040 (N_2040,N_1896,N_1820);
xnor U2041 (N_2041,N_1801,N_1834);
or U2042 (N_2042,N_1801,N_1937);
or U2043 (N_2043,N_1843,N_1872);
or U2044 (N_2044,N_1851,N_1904);
nor U2045 (N_2045,N_1946,N_1941);
nand U2046 (N_2046,N_1922,N_1876);
nor U2047 (N_2047,N_1912,N_1824);
nor U2048 (N_2048,N_1864,N_1803);
nor U2049 (N_2049,N_1937,N_1853);
xnor U2050 (N_2050,N_1884,N_1899);
or U2051 (N_2051,N_1932,N_1887);
or U2052 (N_2052,N_1890,N_1923);
nand U2053 (N_2053,N_1916,N_1870);
xnor U2054 (N_2054,N_1933,N_1920);
and U2055 (N_2055,N_1836,N_1850);
and U2056 (N_2056,N_1866,N_1872);
nor U2057 (N_2057,N_1898,N_1922);
nor U2058 (N_2058,N_1902,N_1909);
and U2059 (N_2059,N_1866,N_1804);
or U2060 (N_2060,N_1830,N_1883);
or U2061 (N_2061,N_1843,N_1925);
nand U2062 (N_2062,N_1940,N_1830);
xnor U2063 (N_2063,N_1927,N_1819);
and U2064 (N_2064,N_1938,N_1936);
nand U2065 (N_2065,N_1923,N_1828);
nor U2066 (N_2066,N_1866,N_1887);
nor U2067 (N_2067,N_1825,N_1808);
nor U2068 (N_2068,N_1856,N_1827);
nand U2069 (N_2069,N_1903,N_1850);
xnor U2070 (N_2070,N_1916,N_1905);
or U2071 (N_2071,N_1903,N_1852);
and U2072 (N_2072,N_1815,N_1818);
xor U2073 (N_2073,N_1856,N_1896);
xnor U2074 (N_2074,N_1908,N_1931);
nand U2075 (N_2075,N_1936,N_1909);
xnor U2076 (N_2076,N_1940,N_1929);
xor U2077 (N_2077,N_1931,N_1915);
or U2078 (N_2078,N_1830,N_1816);
xor U2079 (N_2079,N_1827,N_1931);
nor U2080 (N_2080,N_1866,N_1933);
and U2081 (N_2081,N_1894,N_1853);
nor U2082 (N_2082,N_1890,N_1858);
or U2083 (N_2083,N_1912,N_1904);
nand U2084 (N_2084,N_1812,N_1811);
or U2085 (N_2085,N_1824,N_1944);
xnor U2086 (N_2086,N_1844,N_1937);
nand U2087 (N_2087,N_1831,N_1840);
xnor U2088 (N_2088,N_1835,N_1898);
and U2089 (N_2089,N_1899,N_1889);
nand U2090 (N_2090,N_1847,N_1834);
xor U2091 (N_2091,N_1859,N_1841);
xor U2092 (N_2092,N_1834,N_1802);
and U2093 (N_2093,N_1805,N_1913);
or U2094 (N_2094,N_1886,N_1805);
nor U2095 (N_2095,N_1866,N_1856);
or U2096 (N_2096,N_1885,N_1821);
nor U2097 (N_2097,N_1930,N_1860);
or U2098 (N_2098,N_1874,N_1940);
xnor U2099 (N_2099,N_1864,N_1817);
and U2100 (N_2100,N_2071,N_2003);
or U2101 (N_2101,N_2074,N_1952);
xor U2102 (N_2102,N_1980,N_1999);
nor U2103 (N_2103,N_1993,N_2006);
nand U2104 (N_2104,N_2096,N_2000);
xor U2105 (N_2105,N_1979,N_1962);
xnor U2106 (N_2106,N_2017,N_2098);
xor U2107 (N_2107,N_1965,N_1958);
nor U2108 (N_2108,N_2030,N_2091);
nor U2109 (N_2109,N_2070,N_2060);
nor U2110 (N_2110,N_2029,N_2058);
nand U2111 (N_2111,N_2059,N_2021);
or U2112 (N_2112,N_2087,N_2081);
nor U2113 (N_2113,N_2072,N_2079);
nor U2114 (N_2114,N_2043,N_1973);
xor U2115 (N_2115,N_2051,N_2088);
xnor U2116 (N_2116,N_2036,N_2026);
xnor U2117 (N_2117,N_1997,N_1976);
nand U2118 (N_2118,N_2068,N_2042);
xor U2119 (N_2119,N_2039,N_2015);
nor U2120 (N_2120,N_1954,N_2078);
and U2121 (N_2121,N_2057,N_2046);
xor U2122 (N_2122,N_2086,N_2027);
or U2123 (N_2123,N_2012,N_1964);
or U2124 (N_2124,N_1968,N_2033);
xor U2125 (N_2125,N_2031,N_2093);
nor U2126 (N_2126,N_1984,N_2050);
or U2127 (N_2127,N_2077,N_1987);
xor U2128 (N_2128,N_1955,N_1989);
or U2129 (N_2129,N_2009,N_2061);
nor U2130 (N_2130,N_2099,N_2034);
xnor U2131 (N_2131,N_2023,N_1992);
nor U2132 (N_2132,N_1970,N_2094);
and U2133 (N_2133,N_1975,N_2024);
or U2134 (N_2134,N_1956,N_2095);
and U2135 (N_2135,N_1998,N_1950);
and U2136 (N_2136,N_2004,N_2038);
and U2137 (N_2137,N_2002,N_1988);
nand U2138 (N_2138,N_2007,N_2089);
nor U2139 (N_2139,N_2073,N_2016);
or U2140 (N_2140,N_1986,N_2056);
or U2141 (N_2141,N_1969,N_2010);
or U2142 (N_2142,N_2041,N_2097);
nor U2143 (N_2143,N_2075,N_2076);
nand U2144 (N_2144,N_1985,N_1994);
nor U2145 (N_2145,N_2069,N_2035);
and U2146 (N_2146,N_2052,N_2085);
nor U2147 (N_2147,N_2013,N_2045);
nand U2148 (N_2148,N_2055,N_2084);
and U2149 (N_2149,N_1974,N_1967);
or U2150 (N_2150,N_2001,N_1957);
xor U2151 (N_2151,N_2065,N_1972);
or U2152 (N_2152,N_2063,N_2090);
xnor U2153 (N_2153,N_1960,N_1981);
or U2154 (N_2154,N_1951,N_1990);
nor U2155 (N_2155,N_2048,N_2005);
and U2156 (N_2156,N_2080,N_1991);
nor U2157 (N_2157,N_1966,N_2044);
nor U2158 (N_2158,N_2011,N_2053);
xnor U2159 (N_2159,N_1982,N_2083);
nor U2160 (N_2160,N_1978,N_1983);
or U2161 (N_2161,N_2025,N_1995);
nor U2162 (N_2162,N_2064,N_2067);
and U2163 (N_2163,N_2020,N_2018);
and U2164 (N_2164,N_2008,N_2019);
xor U2165 (N_2165,N_1971,N_2092);
or U2166 (N_2166,N_2049,N_2037);
nand U2167 (N_2167,N_1996,N_2040);
xor U2168 (N_2168,N_1953,N_2066);
nor U2169 (N_2169,N_2062,N_1959);
nand U2170 (N_2170,N_2054,N_2082);
xnor U2171 (N_2171,N_1963,N_2014);
xor U2172 (N_2172,N_2022,N_1961);
nand U2173 (N_2173,N_1977,N_2028);
and U2174 (N_2174,N_2047,N_2032);
nand U2175 (N_2175,N_1964,N_2092);
nor U2176 (N_2176,N_2077,N_1954);
nand U2177 (N_2177,N_1997,N_2045);
and U2178 (N_2178,N_2059,N_2029);
and U2179 (N_2179,N_2061,N_1976);
nand U2180 (N_2180,N_2026,N_2037);
or U2181 (N_2181,N_2016,N_2030);
xor U2182 (N_2182,N_1980,N_2084);
xnor U2183 (N_2183,N_1962,N_1997);
or U2184 (N_2184,N_2085,N_2065);
xor U2185 (N_2185,N_1968,N_2095);
and U2186 (N_2186,N_2011,N_2015);
and U2187 (N_2187,N_1990,N_2066);
xor U2188 (N_2188,N_1979,N_2087);
and U2189 (N_2189,N_2000,N_2045);
xnor U2190 (N_2190,N_2014,N_1970);
or U2191 (N_2191,N_2052,N_1985);
or U2192 (N_2192,N_2040,N_1997);
xor U2193 (N_2193,N_2090,N_2013);
and U2194 (N_2194,N_2044,N_2072);
nand U2195 (N_2195,N_2052,N_2010);
nand U2196 (N_2196,N_2095,N_1965);
nor U2197 (N_2197,N_1978,N_2019);
and U2198 (N_2198,N_2059,N_2022);
nand U2199 (N_2199,N_1983,N_2043);
xnor U2200 (N_2200,N_1974,N_1979);
nor U2201 (N_2201,N_1979,N_1997);
nand U2202 (N_2202,N_2045,N_1960);
xor U2203 (N_2203,N_2045,N_2082);
or U2204 (N_2204,N_2097,N_1970);
and U2205 (N_2205,N_2024,N_1993);
and U2206 (N_2206,N_2099,N_2058);
nand U2207 (N_2207,N_2045,N_1993);
and U2208 (N_2208,N_2094,N_2050);
nor U2209 (N_2209,N_1980,N_1964);
nand U2210 (N_2210,N_2031,N_1959);
and U2211 (N_2211,N_1985,N_2080);
and U2212 (N_2212,N_2012,N_2008);
xor U2213 (N_2213,N_2069,N_2081);
xor U2214 (N_2214,N_2045,N_2047);
nand U2215 (N_2215,N_1999,N_2085);
nor U2216 (N_2216,N_2085,N_2075);
xnor U2217 (N_2217,N_1987,N_1971);
or U2218 (N_2218,N_1970,N_2051);
and U2219 (N_2219,N_1977,N_2000);
nand U2220 (N_2220,N_2081,N_2039);
or U2221 (N_2221,N_2030,N_2096);
and U2222 (N_2222,N_2018,N_2090);
or U2223 (N_2223,N_2081,N_2055);
xor U2224 (N_2224,N_1989,N_1999);
and U2225 (N_2225,N_2014,N_1995);
xor U2226 (N_2226,N_1966,N_2068);
nand U2227 (N_2227,N_2099,N_2029);
nor U2228 (N_2228,N_2028,N_2081);
nand U2229 (N_2229,N_2084,N_1968);
xnor U2230 (N_2230,N_2029,N_2003);
and U2231 (N_2231,N_2063,N_2004);
xnor U2232 (N_2232,N_2040,N_2095);
nand U2233 (N_2233,N_2097,N_2091);
nand U2234 (N_2234,N_2080,N_2090);
or U2235 (N_2235,N_2057,N_2072);
and U2236 (N_2236,N_2041,N_2086);
nor U2237 (N_2237,N_2042,N_1973);
xor U2238 (N_2238,N_2027,N_2063);
or U2239 (N_2239,N_1979,N_2060);
nand U2240 (N_2240,N_2039,N_2082);
nand U2241 (N_2241,N_2006,N_2091);
and U2242 (N_2242,N_2081,N_1958);
and U2243 (N_2243,N_1960,N_2049);
xnor U2244 (N_2244,N_2079,N_2030);
and U2245 (N_2245,N_2085,N_1950);
and U2246 (N_2246,N_2022,N_1953);
nand U2247 (N_2247,N_2077,N_2050);
and U2248 (N_2248,N_2030,N_2012);
nor U2249 (N_2249,N_1957,N_1997);
and U2250 (N_2250,N_2206,N_2129);
and U2251 (N_2251,N_2109,N_2170);
and U2252 (N_2252,N_2208,N_2145);
nor U2253 (N_2253,N_2149,N_2199);
nand U2254 (N_2254,N_2217,N_2173);
or U2255 (N_2255,N_2183,N_2125);
and U2256 (N_2256,N_2188,N_2119);
nand U2257 (N_2257,N_2174,N_2165);
xnor U2258 (N_2258,N_2142,N_2233);
nor U2259 (N_2259,N_2113,N_2246);
or U2260 (N_2260,N_2126,N_2240);
xor U2261 (N_2261,N_2229,N_2245);
or U2262 (N_2262,N_2242,N_2166);
nand U2263 (N_2263,N_2244,N_2127);
or U2264 (N_2264,N_2136,N_2191);
xor U2265 (N_2265,N_2107,N_2140);
nand U2266 (N_2266,N_2118,N_2168);
xor U2267 (N_2267,N_2111,N_2146);
nor U2268 (N_2268,N_2224,N_2100);
nor U2269 (N_2269,N_2185,N_2222);
nand U2270 (N_2270,N_2198,N_2161);
nor U2271 (N_2271,N_2101,N_2160);
xnor U2272 (N_2272,N_2235,N_2241);
and U2273 (N_2273,N_2175,N_2176);
nor U2274 (N_2274,N_2110,N_2139);
and U2275 (N_2275,N_2186,N_2141);
and U2276 (N_2276,N_2231,N_2122);
or U2277 (N_2277,N_2128,N_2152);
and U2278 (N_2278,N_2237,N_2212);
or U2279 (N_2279,N_2193,N_2226);
and U2280 (N_2280,N_2123,N_2158);
xor U2281 (N_2281,N_2156,N_2105);
or U2282 (N_2282,N_2223,N_2247);
and U2283 (N_2283,N_2210,N_2154);
xnor U2284 (N_2284,N_2187,N_2121);
xor U2285 (N_2285,N_2196,N_2232);
or U2286 (N_2286,N_2178,N_2159);
nor U2287 (N_2287,N_2230,N_2135);
or U2288 (N_2288,N_2115,N_2184);
or U2289 (N_2289,N_2124,N_2219);
or U2290 (N_2290,N_2108,N_2137);
xnor U2291 (N_2291,N_2227,N_2243);
nor U2292 (N_2292,N_2106,N_2138);
nand U2293 (N_2293,N_2164,N_2192);
and U2294 (N_2294,N_2203,N_2239);
nand U2295 (N_2295,N_2189,N_2150);
xor U2296 (N_2296,N_2163,N_2205);
xor U2297 (N_2297,N_2197,N_2228);
nor U2298 (N_2298,N_2153,N_2134);
and U2299 (N_2299,N_2216,N_2211);
and U2300 (N_2300,N_2234,N_2236);
and U2301 (N_2301,N_2130,N_2120);
xnor U2302 (N_2302,N_2132,N_2200);
and U2303 (N_2303,N_2220,N_2213);
or U2304 (N_2304,N_2249,N_2112);
xor U2305 (N_2305,N_2155,N_2204);
xor U2306 (N_2306,N_2194,N_2209);
xnor U2307 (N_2307,N_2177,N_2179);
nand U2308 (N_2308,N_2131,N_2180);
and U2309 (N_2309,N_2172,N_2143);
and U2310 (N_2310,N_2201,N_2116);
or U2311 (N_2311,N_2167,N_2238);
nor U2312 (N_2312,N_2214,N_2195);
nor U2313 (N_2313,N_2218,N_2207);
or U2314 (N_2314,N_2103,N_2147);
xor U2315 (N_2315,N_2221,N_2148);
or U2316 (N_2316,N_2102,N_2248);
xnor U2317 (N_2317,N_2181,N_2114);
and U2318 (N_2318,N_2171,N_2162);
or U2319 (N_2319,N_2225,N_2190);
or U2320 (N_2320,N_2182,N_2202);
nand U2321 (N_2321,N_2144,N_2215);
and U2322 (N_2322,N_2151,N_2104);
or U2323 (N_2323,N_2117,N_2157);
xor U2324 (N_2324,N_2169,N_2133);
or U2325 (N_2325,N_2162,N_2218);
xnor U2326 (N_2326,N_2111,N_2136);
and U2327 (N_2327,N_2223,N_2137);
or U2328 (N_2328,N_2156,N_2218);
nor U2329 (N_2329,N_2225,N_2115);
nor U2330 (N_2330,N_2112,N_2189);
nand U2331 (N_2331,N_2192,N_2144);
nand U2332 (N_2332,N_2137,N_2138);
or U2333 (N_2333,N_2220,N_2201);
nand U2334 (N_2334,N_2188,N_2201);
and U2335 (N_2335,N_2119,N_2145);
xor U2336 (N_2336,N_2161,N_2241);
or U2337 (N_2337,N_2208,N_2185);
nor U2338 (N_2338,N_2199,N_2113);
nor U2339 (N_2339,N_2192,N_2145);
or U2340 (N_2340,N_2248,N_2122);
xnor U2341 (N_2341,N_2234,N_2167);
nand U2342 (N_2342,N_2123,N_2151);
nand U2343 (N_2343,N_2189,N_2165);
xnor U2344 (N_2344,N_2224,N_2129);
and U2345 (N_2345,N_2104,N_2180);
nor U2346 (N_2346,N_2113,N_2167);
or U2347 (N_2347,N_2200,N_2125);
nor U2348 (N_2348,N_2120,N_2128);
nand U2349 (N_2349,N_2112,N_2153);
nand U2350 (N_2350,N_2222,N_2241);
nor U2351 (N_2351,N_2130,N_2150);
nor U2352 (N_2352,N_2147,N_2176);
nand U2353 (N_2353,N_2235,N_2146);
nor U2354 (N_2354,N_2205,N_2171);
xor U2355 (N_2355,N_2158,N_2155);
nand U2356 (N_2356,N_2221,N_2110);
and U2357 (N_2357,N_2208,N_2219);
or U2358 (N_2358,N_2238,N_2213);
nand U2359 (N_2359,N_2123,N_2114);
nor U2360 (N_2360,N_2189,N_2111);
nor U2361 (N_2361,N_2109,N_2221);
or U2362 (N_2362,N_2213,N_2158);
nor U2363 (N_2363,N_2222,N_2140);
and U2364 (N_2364,N_2145,N_2180);
xnor U2365 (N_2365,N_2110,N_2198);
nor U2366 (N_2366,N_2166,N_2183);
nor U2367 (N_2367,N_2209,N_2164);
or U2368 (N_2368,N_2119,N_2249);
and U2369 (N_2369,N_2235,N_2145);
and U2370 (N_2370,N_2105,N_2100);
or U2371 (N_2371,N_2218,N_2188);
nor U2372 (N_2372,N_2187,N_2143);
xor U2373 (N_2373,N_2109,N_2248);
xnor U2374 (N_2374,N_2108,N_2136);
nor U2375 (N_2375,N_2249,N_2224);
nor U2376 (N_2376,N_2155,N_2206);
and U2377 (N_2377,N_2192,N_2179);
and U2378 (N_2378,N_2141,N_2245);
nor U2379 (N_2379,N_2150,N_2146);
nor U2380 (N_2380,N_2208,N_2180);
and U2381 (N_2381,N_2173,N_2109);
and U2382 (N_2382,N_2228,N_2176);
nor U2383 (N_2383,N_2137,N_2170);
and U2384 (N_2384,N_2217,N_2222);
and U2385 (N_2385,N_2235,N_2207);
or U2386 (N_2386,N_2145,N_2172);
nor U2387 (N_2387,N_2153,N_2107);
and U2388 (N_2388,N_2168,N_2145);
nand U2389 (N_2389,N_2108,N_2146);
or U2390 (N_2390,N_2191,N_2174);
xor U2391 (N_2391,N_2213,N_2120);
xor U2392 (N_2392,N_2168,N_2128);
and U2393 (N_2393,N_2244,N_2126);
nand U2394 (N_2394,N_2238,N_2111);
xor U2395 (N_2395,N_2226,N_2222);
and U2396 (N_2396,N_2193,N_2206);
nor U2397 (N_2397,N_2216,N_2101);
or U2398 (N_2398,N_2132,N_2241);
nand U2399 (N_2399,N_2175,N_2138);
and U2400 (N_2400,N_2350,N_2305);
and U2401 (N_2401,N_2309,N_2372);
nor U2402 (N_2402,N_2302,N_2289);
nor U2403 (N_2403,N_2316,N_2314);
nor U2404 (N_2404,N_2349,N_2326);
or U2405 (N_2405,N_2318,N_2331);
or U2406 (N_2406,N_2363,N_2351);
and U2407 (N_2407,N_2262,N_2365);
and U2408 (N_2408,N_2285,N_2345);
or U2409 (N_2409,N_2384,N_2319);
and U2410 (N_2410,N_2303,N_2388);
and U2411 (N_2411,N_2361,N_2357);
nand U2412 (N_2412,N_2291,N_2389);
and U2413 (N_2413,N_2250,N_2281);
or U2414 (N_2414,N_2393,N_2396);
or U2415 (N_2415,N_2296,N_2324);
and U2416 (N_2416,N_2269,N_2275);
xor U2417 (N_2417,N_2399,N_2353);
or U2418 (N_2418,N_2317,N_2292);
or U2419 (N_2419,N_2323,N_2253);
nand U2420 (N_2420,N_2290,N_2272);
xnor U2421 (N_2421,N_2295,N_2348);
nor U2422 (N_2422,N_2397,N_2369);
xor U2423 (N_2423,N_2320,N_2368);
or U2424 (N_2424,N_2342,N_2287);
nor U2425 (N_2425,N_2313,N_2267);
or U2426 (N_2426,N_2286,N_2339);
and U2427 (N_2427,N_2328,N_2284);
and U2428 (N_2428,N_2352,N_2355);
xnor U2429 (N_2429,N_2346,N_2322);
xor U2430 (N_2430,N_2330,N_2338);
xnor U2431 (N_2431,N_2391,N_2276);
or U2432 (N_2432,N_2370,N_2255);
nor U2433 (N_2433,N_2367,N_2260);
nor U2434 (N_2434,N_2297,N_2298);
or U2435 (N_2435,N_2343,N_2383);
xnor U2436 (N_2436,N_2356,N_2288);
nor U2437 (N_2437,N_2283,N_2263);
or U2438 (N_2438,N_2266,N_2380);
and U2439 (N_2439,N_2307,N_2268);
and U2440 (N_2440,N_2334,N_2252);
and U2441 (N_2441,N_2315,N_2347);
or U2442 (N_2442,N_2277,N_2386);
or U2443 (N_2443,N_2394,N_2382);
and U2444 (N_2444,N_2273,N_2294);
or U2445 (N_2445,N_2374,N_2337);
nor U2446 (N_2446,N_2256,N_2310);
or U2447 (N_2447,N_2358,N_2395);
nor U2448 (N_2448,N_2254,N_2278);
nor U2449 (N_2449,N_2341,N_2311);
xnor U2450 (N_2450,N_2259,N_2371);
nor U2451 (N_2451,N_2306,N_2392);
and U2452 (N_2452,N_2321,N_2271);
nor U2453 (N_2453,N_2274,N_2360);
nand U2454 (N_2454,N_2354,N_2304);
xor U2455 (N_2455,N_2377,N_2362);
xnor U2456 (N_2456,N_2376,N_2264);
nand U2457 (N_2457,N_2300,N_2270);
xor U2458 (N_2458,N_2335,N_2340);
xnor U2459 (N_2459,N_2280,N_2398);
xnor U2460 (N_2460,N_2381,N_2279);
or U2461 (N_2461,N_2379,N_2373);
nand U2462 (N_2462,N_2387,N_2344);
nor U2463 (N_2463,N_2385,N_2282);
nor U2464 (N_2464,N_2325,N_2366);
or U2465 (N_2465,N_2308,N_2251);
nor U2466 (N_2466,N_2329,N_2390);
nand U2467 (N_2467,N_2265,N_2378);
xnor U2468 (N_2468,N_2261,N_2299);
nand U2469 (N_2469,N_2257,N_2333);
or U2470 (N_2470,N_2359,N_2327);
nor U2471 (N_2471,N_2375,N_2258);
nand U2472 (N_2472,N_2293,N_2336);
xnor U2473 (N_2473,N_2364,N_2332);
nand U2474 (N_2474,N_2301,N_2312);
nand U2475 (N_2475,N_2257,N_2302);
and U2476 (N_2476,N_2271,N_2383);
nor U2477 (N_2477,N_2255,N_2263);
or U2478 (N_2478,N_2339,N_2311);
xor U2479 (N_2479,N_2305,N_2346);
and U2480 (N_2480,N_2303,N_2370);
or U2481 (N_2481,N_2329,N_2330);
xor U2482 (N_2482,N_2261,N_2258);
nand U2483 (N_2483,N_2385,N_2360);
xor U2484 (N_2484,N_2363,N_2335);
xnor U2485 (N_2485,N_2362,N_2324);
nor U2486 (N_2486,N_2306,N_2333);
xnor U2487 (N_2487,N_2253,N_2397);
or U2488 (N_2488,N_2270,N_2318);
and U2489 (N_2489,N_2255,N_2315);
nor U2490 (N_2490,N_2327,N_2334);
nand U2491 (N_2491,N_2292,N_2307);
nand U2492 (N_2492,N_2357,N_2288);
xor U2493 (N_2493,N_2337,N_2289);
nand U2494 (N_2494,N_2256,N_2294);
or U2495 (N_2495,N_2361,N_2285);
xnor U2496 (N_2496,N_2359,N_2307);
xor U2497 (N_2497,N_2275,N_2397);
or U2498 (N_2498,N_2309,N_2392);
and U2499 (N_2499,N_2381,N_2367);
or U2500 (N_2500,N_2304,N_2356);
or U2501 (N_2501,N_2370,N_2399);
or U2502 (N_2502,N_2259,N_2275);
nor U2503 (N_2503,N_2286,N_2291);
nor U2504 (N_2504,N_2256,N_2369);
nor U2505 (N_2505,N_2357,N_2370);
nand U2506 (N_2506,N_2262,N_2299);
nor U2507 (N_2507,N_2322,N_2340);
and U2508 (N_2508,N_2268,N_2338);
and U2509 (N_2509,N_2269,N_2357);
or U2510 (N_2510,N_2267,N_2275);
xor U2511 (N_2511,N_2260,N_2352);
or U2512 (N_2512,N_2256,N_2381);
xnor U2513 (N_2513,N_2263,N_2326);
or U2514 (N_2514,N_2397,N_2352);
xor U2515 (N_2515,N_2295,N_2270);
and U2516 (N_2516,N_2374,N_2381);
nand U2517 (N_2517,N_2279,N_2284);
or U2518 (N_2518,N_2358,N_2329);
nor U2519 (N_2519,N_2297,N_2355);
nand U2520 (N_2520,N_2267,N_2256);
nand U2521 (N_2521,N_2393,N_2398);
or U2522 (N_2522,N_2394,N_2267);
and U2523 (N_2523,N_2353,N_2326);
xnor U2524 (N_2524,N_2349,N_2331);
xor U2525 (N_2525,N_2344,N_2314);
or U2526 (N_2526,N_2255,N_2293);
xor U2527 (N_2527,N_2294,N_2340);
nand U2528 (N_2528,N_2339,N_2278);
nand U2529 (N_2529,N_2292,N_2319);
nor U2530 (N_2530,N_2261,N_2284);
xor U2531 (N_2531,N_2340,N_2334);
nand U2532 (N_2532,N_2376,N_2292);
nor U2533 (N_2533,N_2345,N_2349);
nand U2534 (N_2534,N_2316,N_2282);
nor U2535 (N_2535,N_2310,N_2336);
xnor U2536 (N_2536,N_2318,N_2351);
nor U2537 (N_2537,N_2366,N_2294);
xnor U2538 (N_2538,N_2271,N_2268);
nor U2539 (N_2539,N_2349,N_2363);
nand U2540 (N_2540,N_2383,N_2286);
and U2541 (N_2541,N_2351,N_2332);
nor U2542 (N_2542,N_2262,N_2313);
and U2543 (N_2543,N_2299,N_2290);
xor U2544 (N_2544,N_2274,N_2380);
and U2545 (N_2545,N_2320,N_2287);
nor U2546 (N_2546,N_2374,N_2303);
xnor U2547 (N_2547,N_2348,N_2270);
and U2548 (N_2548,N_2268,N_2343);
xnor U2549 (N_2549,N_2286,N_2333);
nor U2550 (N_2550,N_2532,N_2448);
nand U2551 (N_2551,N_2435,N_2421);
and U2552 (N_2552,N_2504,N_2500);
nand U2553 (N_2553,N_2491,N_2422);
nand U2554 (N_2554,N_2471,N_2446);
nand U2555 (N_2555,N_2503,N_2492);
nand U2556 (N_2556,N_2400,N_2482);
and U2557 (N_2557,N_2493,N_2549);
xnor U2558 (N_2558,N_2476,N_2487);
nor U2559 (N_2559,N_2501,N_2461);
nand U2560 (N_2560,N_2402,N_2429);
nand U2561 (N_2561,N_2439,N_2425);
nand U2562 (N_2562,N_2447,N_2480);
and U2563 (N_2563,N_2510,N_2519);
nand U2564 (N_2564,N_2535,N_2415);
nor U2565 (N_2565,N_2521,N_2511);
or U2566 (N_2566,N_2543,N_2426);
xnor U2567 (N_2567,N_2484,N_2442);
xor U2568 (N_2568,N_2534,N_2508);
nor U2569 (N_2569,N_2479,N_2518);
nand U2570 (N_2570,N_2516,N_2536);
or U2571 (N_2571,N_2433,N_2514);
and U2572 (N_2572,N_2494,N_2526);
nand U2573 (N_2573,N_2485,N_2432);
nand U2574 (N_2574,N_2440,N_2405);
xor U2575 (N_2575,N_2423,N_2546);
xor U2576 (N_2576,N_2467,N_2455);
or U2577 (N_2577,N_2530,N_2541);
nor U2578 (N_2578,N_2488,N_2507);
or U2579 (N_2579,N_2473,N_2443);
nand U2580 (N_2580,N_2468,N_2437);
nand U2581 (N_2581,N_2542,N_2436);
nand U2582 (N_2582,N_2520,N_2403);
nand U2583 (N_2583,N_2481,N_2469);
nor U2584 (N_2584,N_2509,N_2407);
nor U2585 (N_2585,N_2472,N_2545);
xor U2586 (N_2586,N_2496,N_2527);
nand U2587 (N_2587,N_2529,N_2441);
nand U2588 (N_2588,N_2401,N_2457);
and U2589 (N_2589,N_2463,N_2466);
nor U2590 (N_2590,N_2548,N_2450);
or U2591 (N_2591,N_2462,N_2539);
or U2592 (N_2592,N_2547,N_2445);
or U2593 (N_2593,N_2489,N_2413);
nand U2594 (N_2594,N_2404,N_2506);
nor U2595 (N_2595,N_2419,N_2499);
or U2596 (N_2596,N_2428,N_2416);
nor U2597 (N_2597,N_2458,N_2524);
nand U2598 (N_2598,N_2451,N_2464);
nor U2599 (N_2599,N_2495,N_2417);
or U2600 (N_2600,N_2418,N_2474);
and U2601 (N_2601,N_2523,N_2411);
and U2602 (N_2602,N_2459,N_2460);
nor U2603 (N_2603,N_2408,N_2525);
nand U2604 (N_2604,N_2470,N_2456);
xor U2605 (N_2605,N_2477,N_2512);
xor U2606 (N_2606,N_2414,N_2537);
and U2607 (N_2607,N_2490,N_2424);
xnor U2608 (N_2608,N_2538,N_2533);
nand U2609 (N_2609,N_2431,N_2517);
or U2610 (N_2610,N_2454,N_2430);
and U2611 (N_2611,N_2540,N_2544);
or U2612 (N_2612,N_2444,N_2515);
and U2613 (N_2613,N_2452,N_2449);
nand U2614 (N_2614,N_2438,N_2513);
xor U2615 (N_2615,N_2505,N_2483);
nor U2616 (N_2616,N_2410,N_2522);
nor U2617 (N_2617,N_2409,N_2478);
and U2618 (N_2618,N_2412,N_2434);
nor U2619 (N_2619,N_2497,N_2453);
and U2620 (N_2620,N_2531,N_2427);
nand U2621 (N_2621,N_2502,N_2406);
and U2622 (N_2622,N_2420,N_2498);
nand U2623 (N_2623,N_2465,N_2528);
or U2624 (N_2624,N_2486,N_2475);
nand U2625 (N_2625,N_2408,N_2462);
and U2626 (N_2626,N_2445,N_2455);
or U2627 (N_2627,N_2502,N_2439);
or U2628 (N_2628,N_2444,N_2405);
nand U2629 (N_2629,N_2433,N_2475);
or U2630 (N_2630,N_2492,N_2539);
nand U2631 (N_2631,N_2423,N_2517);
and U2632 (N_2632,N_2490,N_2506);
or U2633 (N_2633,N_2543,N_2423);
xnor U2634 (N_2634,N_2457,N_2481);
nor U2635 (N_2635,N_2420,N_2484);
and U2636 (N_2636,N_2420,N_2427);
nand U2637 (N_2637,N_2460,N_2458);
xnor U2638 (N_2638,N_2437,N_2545);
xnor U2639 (N_2639,N_2467,N_2431);
xnor U2640 (N_2640,N_2427,N_2532);
xor U2641 (N_2641,N_2452,N_2436);
or U2642 (N_2642,N_2452,N_2466);
xor U2643 (N_2643,N_2545,N_2520);
xor U2644 (N_2644,N_2426,N_2548);
nand U2645 (N_2645,N_2475,N_2425);
nor U2646 (N_2646,N_2532,N_2409);
nor U2647 (N_2647,N_2456,N_2503);
nor U2648 (N_2648,N_2461,N_2443);
xor U2649 (N_2649,N_2403,N_2538);
and U2650 (N_2650,N_2504,N_2421);
or U2651 (N_2651,N_2544,N_2438);
or U2652 (N_2652,N_2408,N_2460);
and U2653 (N_2653,N_2470,N_2485);
or U2654 (N_2654,N_2520,N_2466);
or U2655 (N_2655,N_2492,N_2450);
and U2656 (N_2656,N_2439,N_2482);
nor U2657 (N_2657,N_2545,N_2465);
and U2658 (N_2658,N_2436,N_2426);
nand U2659 (N_2659,N_2468,N_2488);
and U2660 (N_2660,N_2467,N_2515);
nand U2661 (N_2661,N_2539,N_2442);
or U2662 (N_2662,N_2484,N_2489);
nor U2663 (N_2663,N_2496,N_2516);
and U2664 (N_2664,N_2526,N_2437);
xnor U2665 (N_2665,N_2505,N_2464);
xor U2666 (N_2666,N_2542,N_2452);
nand U2667 (N_2667,N_2484,N_2434);
nand U2668 (N_2668,N_2466,N_2449);
or U2669 (N_2669,N_2432,N_2501);
xor U2670 (N_2670,N_2516,N_2415);
nand U2671 (N_2671,N_2544,N_2434);
or U2672 (N_2672,N_2404,N_2435);
nor U2673 (N_2673,N_2421,N_2516);
or U2674 (N_2674,N_2535,N_2481);
or U2675 (N_2675,N_2537,N_2484);
nor U2676 (N_2676,N_2405,N_2402);
xnor U2677 (N_2677,N_2525,N_2507);
or U2678 (N_2678,N_2491,N_2521);
nor U2679 (N_2679,N_2459,N_2433);
nor U2680 (N_2680,N_2475,N_2470);
xnor U2681 (N_2681,N_2458,N_2401);
nand U2682 (N_2682,N_2542,N_2478);
or U2683 (N_2683,N_2464,N_2421);
xor U2684 (N_2684,N_2528,N_2420);
xor U2685 (N_2685,N_2527,N_2456);
xor U2686 (N_2686,N_2437,N_2458);
nand U2687 (N_2687,N_2497,N_2458);
nor U2688 (N_2688,N_2470,N_2501);
nand U2689 (N_2689,N_2476,N_2402);
nor U2690 (N_2690,N_2440,N_2406);
nand U2691 (N_2691,N_2407,N_2406);
nand U2692 (N_2692,N_2461,N_2538);
and U2693 (N_2693,N_2458,N_2517);
nor U2694 (N_2694,N_2498,N_2497);
nand U2695 (N_2695,N_2418,N_2468);
and U2696 (N_2696,N_2460,N_2451);
or U2697 (N_2697,N_2411,N_2486);
xor U2698 (N_2698,N_2493,N_2449);
nor U2699 (N_2699,N_2400,N_2439);
and U2700 (N_2700,N_2694,N_2588);
nor U2701 (N_2701,N_2607,N_2661);
nor U2702 (N_2702,N_2646,N_2682);
nand U2703 (N_2703,N_2554,N_2572);
xor U2704 (N_2704,N_2685,N_2672);
nor U2705 (N_2705,N_2575,N_2552);
nand U2706 (N_2706,N_2644,N_2555);
nand U2707 (N_2707,N_2616,N_2624);
nor U2708 (N_2708,N_2650,N_2623);
xor U2709 (N_2709,N_2684,N_2574);
or U2710 (N_2710,N_2641,N_2604);
nand U2711 (N_2711,N_2615,N_2573);
xnor U2712 (N_2712,N_2660,N_2556);
xor U2713 (N_2713,N_2611,N_2583);
xor U2714 (N_2714,N_2570,N_2638);
xnor U2715 (N_2715,N_2691,N_2675);
xnor U2716 (N_2716,N_2656,N_2643);
or U2717 (N_2717,N_2589,N_2612);
or U2718 (N_2718,N_2681,N_2560);
or U2719 (N_2719,N_2621,N_2582);
or U2720 (N_2720,N_2686,N_2629);
and U2721 (N_2721,N_2587,N_2618);
nor U2722 (N_2722,N_2576,N_2592);
or U2723 (N_2723,N_2596,N_2565);
nand U2724 (N_2724,N_2680,N_2567);
nand U2725 (N_2725,N_2601,N_2668);
and U2726 (N_2726,N_2627,N_2674);
xnor U2727 (N_2727,N_2630,N_2666);
xor U2728 (N_2728,N_2605,N_2563);
xor U2729 (N_2729,N_2632,N_2649);
nor U2730 (N_2730,N_2693,N_2593);
or U2731 (N_2731,N_2626,N_2688);
nand U2732 (N_2732,N_2559,N_2631);
xnor U2733 (N_2733,N_2595,N_2602);
nand U2734 (N_2734,N_2640,N_2571);
or U2735 (N_2735,N_2676,N_2608);
nand U2736 (N_2736,N_2653,N_2578);
nand U2737 (N_2737,N_2606,N_2622);
xor U2738 (N_2738,N_2667,N_2695);
xnor U2739 (N_2739,N_2581,N_2699);
or U2740 (N_2740,N_2619,N_2698);
nor U2741 (N_2741,N_2690,N_2642);
xor U2742 (N_2742,N_2586,N_2665);
nand U2743 (N_2743,N_2671,N_2663);
or U2744 (N_2744,N_2564,N_2633);
nand U2745 (N_2745,N_2591,N_2566);
nand U2746 (N_2746,N_2692,N_2678);
xnor U2747 (N_2747,N_2696,N_2620);
or U2748 (N_2748,N_2579,N_2677);
nor U2749 (N_2749,N_2628,N_2568);
nand U2750 (N_2750,N_2577,N_2657);
xnor U2751 (N_2751,N_2580,N_2664);
and U2752 (N_2752,N_2658,N_2600);
and U2753 (N_2753,N_2639,N_2617);
and U2754 (N_2754,N_2597,N_2648);
and U2755 (N_2755,N_2651,N_2697);
nor U2756 (N_2756,N_2614,N_2585);
or U2757 (N_2757,N_2599,N_2636);
or U2758 (N_2758,N_2669,N_2645);
nor U2759 (N_2759,N_2613,N_2647);
nor U2760 (N_2760,N_2553,N_2590);
or U2761 (N_2761,N_2683,N_2562);
or U2762 (N_2762,N_2689,N_2609);
and U2763 (N_2763,N_2558,N_2610);
nand U2764 (N_2764,N_2635,N_2662);
xnor U2765 (N_2765,N_2655,N_2584);
or U2766 (N_2766,N_2634,N_2670);
or U2767 (N_2767,N_2598,N_2550);
and U2768 (N_2768,N_2557,N_2659);
nor U2769 (N_2769,N_2561,N_2569);
and U2770 (N_2770,N_2687,N_2679);
and U2771 (N_2771,N_2673,N_2594);
xor U2772 (N_2772,N_2654,N_2652);
xor U2773 (N_2773,N_2603,N_2551);
nand U2774 (N_2774,N_2637,N_2625);
nor U2775 (N_2775,N_2669,N_2672);
or U2776 (N_2776,N_2590,N_2690);
xor U2777 (N_2777,N_2646,N_2583);
or U2778 (N_2778,N_2552,N_2677);
nor U2779 (N_2779,N_2685,N_2560);
nor U2780 (N_2780,N_2634,N_2570);
or U2781 (N_2781,N_2663,N_2581);
nor U2782 (N_2782,N_2616,N_2553);
xnor U2783 (N_2783,N_2571,N_2606);
nor U2784 (N_2784,N_2582,N_2638);
xnor U2785 (N_2785,N_2679,N_2675);
nand U2786 (N_2786,N_2612,N_2617);
or U2787 (N_2787,N_2624,N_2620);
or U2788 (N_2788,N_2639,N_2643);
and U2789 (N_2789,N_2682,N_2563);
nor U2790 (N_2790,N_2674,N_2575);
nand U2791 (N_2791,N_2686,N_2574);
nand U2792 (N_2792,N_2653,N_2654);
or U2793 (N_2793,N_2666,N_2628);
and U2794 (N_2794,N_2694,N_2673);
nand U2795 (N_2795,N_2575,N_2613);
nand U2796 (N_2796,N_2678,N_2688);
xnor U2797 (N_2797,N_2661,N_2649);
nand U2798 (N_2798,N_2563,N_2637);
or U2799 (N_2799,N_2657,N_2696);
nand U2800 (N_2800,N_2655,N_2637);
nor U2801 (N_2801,N_2610,N_2645);
nor U2802 (N_2802,N_2668,N_2574);
xnor U2803 (N_2803,N_2608,N_2675);
or U2804 (N_2804,N_2574,N_2681);
xnor U2805 (N_2805,N_2684,N_2672);
and U2806 (N_2806,N_2569,N_2555);
nand U2807 (N_2807,N_2689,N_2613);
and U2808 (N_2808,N_2667,N_2568);
or U2809 (N_2809,N_2691,N_2553);
nor U2810 (N_2810,N_2550,N_2679);
and U2811 (N_2811,N_2582,N_2623);
or U2812 (N_2812,N_2687,N_2596);
nand U2813 (N_2813,N_2618,N_2592);
or U2814 (N_2814,N_2577,N_2568);
or U2815 (N_2815,N_2580,N_2645);
nor U2816 (N_2816,N_2558,N_2587);
and U2817 (N_2817,N_2629,N_2609);
xor U2818 (N_2818,N_2650,N_2615);
nand U2819 (N_2819,N_2592,N_2560);
xnor U2820 (N_2820,N_2693,N_2590);
or U2821 (N_2821,N_2572,N_2588);
and U2822 (N_2822,N_2614,N_2602);
nor U2823 (N_2823,N_2621,N_2557);
xor U2824 (N_2824,N_2690,N_2555);
nor U2825 (N_2825,N_2584,N_2634);
xor U2826 (N_2826,N_2550,N_2699);
nand U2827 (N_2827,N_2655,N_2672);
xnor U2828 (N_2828,N_2684,N_2671);
nand U2829 (N_2829,N_2569,N_2654);
xnor U2830 (N_2830,N_2615,N_2631);
or U2831 (N_2831,N_2622,N_2695);
nand U2832 (N_2832,N_2587,N_2605);
or U2833 (N_2833,N_2653,N_2694);
nand U2834 (N_2834,N_2698,N_2552);
or U2835 (N_2835,N_2699,N_2594);
nor U2836 (N_2836,N_2682,N_2660);
nand U2837 (N_2837,N_2678,N_2593);
nand U2838 (N_2838,N_2589,N_2631);
or U2839 (N_2839,N_2626,N_2624);
nand U2840 (N_2840,N_2691,N_2670);
or U2841 (N_2841,N_2597,N_2697);
and U2842 (N_2842,N_2613,N_2588);
nor U2843 (N_2843,N_2677,N_2686);
nand U2844 (N_2844,N_2617,N_2646);
nand U2845 (N_2845,N_2566,N_2562);
nand U2846 (N_2846,N_2686,N_2643);
nand U2847 (N_2847,N_2601,N_2619);
and U2848 (N_2848,N_2657,N_2684);
or U2849 (N_2849,N_2667,N_2684);
xor U2850 (N_2850,N_2830,N_2734);
or U2851 (N_2851,N_2794,N_2848);
nand U2852 (N_2852,N_2829,N_2800);
and U2853 (N_2853,N_2725,N_2721);
nand U2854 (N_2854,N_2804,N_2729);
nand U2855 (N_2855,N_2724,N_2743);
nor U2856 (N_2856,N_2844,N_2700);
nor U2857 (N_2857,N_2774,N_2733);
nand U2858 (N_2858,N_2756,N_2835);
nand U2859 (N_2859,N_2790,N_2738);
nand U2860 (N_2860,N_2785,N_2788);
or U2861 (N_2861,N_2819,N_2707);
xnor U2862 (N_2862,N_2839,N_2717);
and U2863 (N_2863,N_2779,N_2757);
xor U2864 (N_2864,N_2816,N_2780);
xor U2865 (N_2865,N_2801,N_2842);
or U2866 (N_2866,N_2792,N_2755);
xnor U2867 (N_2867,N_2767,N_2846);
and U2868 (N_2868,N_2781,N_2766);
nand U2869 (N_2869,N_2748,N_2843);
nand U2870 (N_2870,N_2718,N_2798);
nor U2871 (N_2871,N_2726,N_2809);
and U2872 (N_2872,N_2732,N_2728);
nand U2873 (N_2873,N_2823,N_2831);
nor U2874 (N_2874,N_2838,N_2824);
or U2875 (N_2875,N_2768,N_2736);
and U2876 (N_2876,N_2713,N_2723);
or U2877 (N_2877,N_2793,N_2737);
and U2878 (N_2878,N_2849,N_2763);
or U2879 (N_2879,N_2761,N_2784);
or U2880 (N_2880,N_2741,N_2709);
nor U2881 (N_2881,N_2772,N_2778);
nor U2882 (N_2882,N_2840,N_2731);
and U2883 (N_2883,N_2777,N_2751);
xor U2884 (N_2884,N_2828,N_2716);
xnor U2885 (N_2885,N_2833,N_2811);
nor U2886 (N_2886,N_2834,N_2783);
or U2887 (N_2887,N_2727,N_2712);
and U2888 (N_2888,N_2703,N_2808);
nor U2889 (N_2889,N_2765,N_2771);
nand U2890 (N_2890,N_2752,N_2826);
nor U2891 (N_2891,N_2742,N_2847);
nand U2892 (N_2892,N_2730,N_2820);
or U2893 (N_2893,N_2735,N_2789);
or U2894 (N_2894,N_2837,N_2822);
nand U2895 (N_2895,N_2827,N_2787);
or U2896 (N_2896,N_2813,N_2720);
nand U2897 (N_2897,N_2799,N_2739);
and U2898 (N_2898,N_2758,N_2708);
nand U2899 (N_2899,N_2769,N_2762);
or U2900 (N_2900,N_2764,N_2796);
or U2901 (N_2901,N_2817,N_2719);
nand U2902 (N_2902,N_2802,N_2841);
and U2903 (N_2903,N_2749,N_2759);
nand U2904 (N_2904,N_2797,N_2704);
and U2905 (N_2905,N_2814,N_2806);
or U2906 (N_2906,N_2747,N_2750);
and U2907 (N_2907,N_2754,N_2702);
nand U2908 (N_2908,N_2705,N_2803);
nand U2909 (N_2909,N_2795,N_2715);
nand U2910 (N_2910,N_2740,N_2706);
nor U2911 (N_2911,N_2770,N_2810);
or U2912 (N_2912,N_2745,N_2782);
or U2913 (N_2913,N_2714,N_2845);
nor U2914 (N_2914,N_2832,N_2760);
xnor U2915 (N_2915,N_2815,N_2773);
nor U2916 (N_2916,N_2701,N_2711);
or U2917 (N_2917,N_2805,N_2825);
and U2918 (N_2918,N_2753,N_2836);
nor U2919 (N_2919,N_2812,N_2775);
or U2920 (N_2920,N_2710,N_2818);
nand U2921 (N_2921,N_2786,N_2746);
xor U2922 (N_2922,N_2744,N_2776);
xnor U2923 (N_2923,N_2722,N_2821);
nand U2924 (N_2924,N_2791,N_2807);
xor U2925 (N_2925,N_2812,N_2727);
and U2926 (N_2926,N_2834,N_2847);
or U2927 (N_2927,N_2782,N_2817);
nor U2928 (N_2928,N_2832,N_2843);
xor U2929 (N_2929,N_2839,N_2846);
or U2930 (N_2930,N_2827,N_2790);
nand U2931 (N_2931,N_2814,N_2758);
nand U2932 (N_2932,N_2721,N_2753);
nor U2933 (N_2933,N_2724,N_2755);
nand U2934 (N_2934,N_2782,N_2739);
nand U2935 (N_2935,N_2801,N_2841);
nand U2936 (N_2936,N_2753,N_2710);
xor U2937 (N_2937,N_2702,N_2773);
or U2938 (N_2938,N_2792,N_2765);
or U2939 (N_2939,N_2778,N_2798);
nor U2940 (N_2940,N_2701,N_2714);
xor U2941 (N_2941,N_2789,N_2787);
nand U2942 (N_2942,N_2761,N_2724);
or U2943 (N_2943,N_2720,N_2705);
and U2944 (N_2944,N_2839,N_2749);
xor U2945 (N_2945,N_2746,N_2800);
nand U2946 (N_2946,N_2768,N_2756);
or U2947 (N_2947,N_2844,N_2728);
nor U2948 (N_2948,N_2706,N_2765);
and U2949 (N_2949,N_2775,N_2810);
nand U2950 (N_2950,N_2820,N_2817);
and U2951 (N_2951,N_2791,N_2729);
or U2952 (N_2952,N_2799,N_2824);
xor U2953 (N_2953,N_2739,N_2829);
and U2954 (N_2954,N_2732,N_2718);
and U2955 (N_2955,N_2792,N_2820);
nand U2956 (N_2956,N_2807,N_2779);
nand U2957 (N_2957,N_2849,N_2755);
or U2958 (N_2958,N_2805,N_2793);
and U2959 (N_2959,N_2774,N_2723);
nor U2960 (N_2960,N_2837,N_2770);
nor U2961 (N_2961,N_2849,N_2811);
nand U2962 (N_2962,N_2758,N_2788);
and U2963 (N_2963,N_2740,N_2791);
nor U2964 (N_2964,N_2807,N_2776);
or U2965 (N_2965,N_2825,N_2739);
or U2966 (N_2966,N_2702,N_2772);
nor U2967 (N_2967,N_2741,N_2745);
nand U2968 (N_2968,N_2761,N_2732);
and U2969 (N_2969,N_2751,N_2826);
nand U2970 (N_2970,N_2740,N_2750);
xor U2971 (N_2971,N_2830,N_2766);
and U2972 (N_2972,N_2833,N_2733);
or U2973 (N_2973,N_2791,N_2805);
and U2974 (N_2974,N_2772,N_2836);
nor U2975 (N_2975,N_2745,N_2848);
or U2976 (N_2976,N_2749,N_2740);
or U2977 (N_2977,N_2729,N_2781);
nor U2978 (N_2978,N_2849,N_2707);
and U2979 (N_2979,N_2781,N_2755);
or U2980 (N_2980,N_2783,N_2732);
xnor U2981 (N_2981,N_2768,N_2843);
xor U2982 (N_2982,N_2725,N_2773);
or U2983 (N_2983,N_2831,N_2754);
nand U2984 (N_2984,N_2780,N_2726);
nor U2985 (N_2985,N_2833,N_2813);
and U2986 (N_2986,N_2777,N_2730);
xnor U2987 (N_2987,N_2796,N_2843);
xor U2988 (N_2988,N_2782,N_2822);
or U2989 (N_2989,N_2777,N_2794);
and U2990 (N_2990,N_2841,N_2707);
nor U2991 (N_2991,N_2842,N_2786);
or U2992 (N_2992,N_2817,N_2720);
and U2993 (N_2993,N_2789,N_2830);
xnor U2994 (N_2994,N_2782,N_2823);
nand U2995 (N_2995,N_2824,N_2744);
or U2996 (N_2996,N_2783,N_2752);
xor U2997 (N_2997,N_2792,N_2783);
xor U2998 (N_2998,N_2825,N_2709);
and U2999 (N_2999,N_2823,N_2806);
or U3000 (N_3000,N_2969,N_2857);
nand U3001 (N_3001,N_2988,N_2856);
and U3002 (N_3002,N_2995,N_2903);
nor U3003 (N_3003,N_2927,N_2886);
xor U3004 (N_3004,N_2949,N_2944);
xnor U3005 (N_3005,N_2968,N_2972);
and U3006 (N_3006,N_2885,N_2983);
xnor U3007 (N_3007,N_2924,N_2992);
nand U3008 (N_3008,N_2905,N_2858);
or U3009 (N_3009,N_2855,N_2881);
nor U3010 (N_3010,N_2975,N_2953);
nand U3011 (N_3011,N_2893,N_2880);
and U3012 (N_3012,N_2882,N_2911);
nor U3013 (N_3013,N_2922,N_2962);
xor U3014 (N_3014,N_2956,N_2850);
and U3015 (N_3015,N_2965,N_2851);
xnor U3016 (N_3016,N_2930,N_2947);
xnor U3017 (N_3017,N_2966,N_2990);
and U3018 (N_3018,N_2912,N_2928);
and U3019 (N_3019,N_2877,N_2909);
xor U3020 (N_3020,N_2868,N_2984);
nand U3021 (N_3021,N_2957,N_2982);
and U3022 (N_3022,N_2959,N_2871);
and U3023 (N_3023,N_2998,N_2925);
nand U3024 (N_3024,N_2894,N_2952);
or U3025 (N_3025,N_2865,N_2904);
nor U3026 (N_3026,N_2933,N_2940);
nand U3027 (N_3027,N_2964,N_2993);
xnor U3028 (N_3028,N_2948,N_2853);
xor U3029 (N_3029,N_2986,N_2914);
nand U3030 (N_3030,N_2864,N_2951);
or U3031 (N_3031,N_2931,N_2961);
or U3032 (N_3032,N_2985,N_2870);
nor U3033 (N_3033,N_2997,N_2888);
or U3034 (N_3034,N_2884,N_2854);
xnor U3035 (N_3035,N_2921,N_2967);
and U3036 (N_3036,N_2963,N_2867);
nand U3037 (N_3037,N_2869,N_2994);
and U3038 (N_3038,N_2936,N_2879);
or U3039 (N_3039,N_2906,N_2898);
nor U3040 (N_3040,N_2973,N_2980);
nor U3041 (N_3041,N_2938,N_2883);
and U3042 (N_3042,N_2939,N_2878);
and U3043 (N_3043,N_2971,N_2974);
nor U3044 (N_3044,N_2977,N_2875);
nor U3045 (N_3045,N_2874,N_2908);
or U3046 (N_3046,N_2918,N_2916);
nor U3047 (N_3047,N_2873,N_2900);
or U3048 (N_3048,N_2902,N_2946);
and U3049 (N_3049,N_2862,N_2976);
nor U3050 (N_3050,N_2901,N_2934);
and U3051 (N_3051,N_2932,N_2899);
xnor U3052 (N_3052,N_2910,N_2917);
or U3053 (N_3053,N_2923,N_2979);
xor U3054 (N_3054,N_2915,N_2890);
and U3055 (N_3055,N_2860,N_2852);
and U3056 (N_3056,N_2919,N_2981);
nand U3057 (N_3057,N_2991,N_2897);
or U3058 (N_3058,N_2987,N_2970);
nor U3059 (N_3059,N_2929,N_2896);
nor U3060 (N_3060,N_2937,N_2891);
nor U3061 (N_3061,N_2920,N_2887);
or U3062 (N_3062,N_2989,N_2960);
xor U3063 (N_3063,N_2945,N_2943);
and U3064 (N_3064,N_2955,N_2941);
nor U3065 (N_3065,N_2978,N_2950);
and U3066 (N_3066,N_2872,N_2926);
nand U3067 (N_3067,N_2892,N_2859);
nand U3068 (N_3068,N_2958,N_2889);
xor U3069 (N_3069,N_2942,N_2999);
nand U3070 (N_3070,N_2907,N_2935);
and U3071 (N_3071,N_2996,N_2913);
and U3072 (N_3072,N_2895,N_2863);
nand U3073 (N_3073,N_2866,N_2861);
nand U3074 (N_3074,N_2954,N_2876);
or U3075 (N_3075,N_2896,N_2980);
and U3076 (N_3076,N_2920,N_2894);
xnor U3077 (N_3077,N_2922,N_2978);
nand U3078 (N_3078,N_2870,N_2913);
or U3079 (N_3079,N_2968,N_2992);
xor U3080 (N_3080,N_2977,N_2945);
xnor U3081 (N_3081,N_2903,N_2863);
nand U3082 (N_3082,N_2864,N_2990);
xor U3083 (N_3083,N_2971,N_2953);
nor U3084 (N_3084,N_2906,N_2964);
nand U3085 (N_3085,N_2891,N_2867);
or U3086 (N_3086,N_2939,N_2886);
xnor U3087 (N_3087,N_2974,N_2890);
and U3088 (N_3088,N_2884,N_2970);
or U3089 (N_3089,N_2897,N_2988);
nand U3090 (N_3090,N_2969,N_2949);
and U3091 (N_3091,N_2992,N_2994);
or U3092 (N_3092,N_2988,N_2901);
and U3093 (N_3093,N_2855,N_2871);
or U3094 (N_3094,N_2932,N_2873);
nor U3095 (N_3095,N_2938,N_2893);
nand U3096 (N_3096,N_2972,N_2986);
and U3097 (N_3097,N_2919,N_2937);
and U3098 (N_3098,N_2865,N_2920);
nor U3099 (N_3099,N_2918,N_2887);
and U3100 (N_3100,N_2992,N_2888);
nand U3101 (N_3101,N_2999,N_2936);
xor U3102 (N_3102,N_2934,N_2931);
nor U3103 (N_3103,N_2859,N_2952);
or U3104 (N_3104,N_2922,N_2882);
xnor U3105 (N_3105,N_2949,N_2878);
nand U3106 (N_3106,N_2930,N_2985);
nor U3107 (N_3107,N_2922,N_2852);
xor U3108 (N_3108,N_2908,N_2896);
and U3109 (N_3109,N_2914,N_2867);
nand U3110 (N_3110,N_2857,N_2942);
and U3111 (N_3111,N_2907,N_2868);
and U3112 (N_3112,N_2919,N_2893);
or U3113 (N_3113,N_2936,N_2909);
nor U3114 (N_3114,N_2900,N_2865);
xnor U3115 (N_3115,N_2860,N_2998);
nand U3116 (N_3116,N_2891,N_2882);
nor U3117 (N_3117,N_2890,N_2943);
xnor U3118 (N_3118,N_2924,N_2958);
xor U3119 (N_3119,N_2909,N_2987);
nand U3120 (N_3120,N_2872,N_2917);
or U3121 (N_3121,N_2993,N_2970);
and U3122 (N_3122,N_2934,N_2998);
xnor U3123 (N_3123,N_2904,N_2998);
and U3124 (N_3124,N_2978,N_2999);
xor U3125 (N_3125,N_2945,N_2881);
nand U3126 (N_3126,N_2950,N_2941);
or U3127 (N_3127,N_2946,N_2939);
and U3128 (N_3128,N_2935,N_2868);
xnor U3129 (N_3129,N_2991,N_2996);
xor U3130 (N_3130,N_2996,N_2902);
nor U3131 (N_3131,N_2974,N_2931);
xnor U3132 (N_3132,N_2949,N_2923);
and U3133 (N_3133,N_2869,N_2938);
nand U3134 (N_3134,N_2938,N_2937);
xor U3135 (N_3135,N_2935,N_2881);
nand U3136 (N_3136,N_2984,N_2854);
nor U3137 (N_3137,N_2935,N_2884);
nand U3138 (N_3138,N_2929,N_2901);
or U3139 (N_3139,N_2922,N_2903);
and U3140 (N_3140,N_2863,N_2964);
nor U3141 (N_3141,N_2873,N_2944);
xnor U3142 (N_3142,N_2871,N_2969);
xor U3143 (N_3143,N_2896,N_2887);
nand U3144 (N_3144,N_2924,N_2852);
nor U3145 (N_3145,N_2965,N_2896);
xnor U3146 (N_3146,N_2938,N_2878);
nor U3147 (N_3147,N_2934,N_2994);
nand U3148 (N_3148,N_2961,N_2894);
nand U3149 (N_3149,N_2919,N_2989);
or U3150 (N_3150,N_3050,N_3110);
xnor U3151 (N_3151,N_3122,N_3101);
nor U3152 (N_3152,N_3053,N_3045);
and U3153 (N_3153,N_3082,N_3123);
or U3154 (N_3154,N_3097,N_3070);
nand U3155 (N_3155,N_3112,N_3061);
xnor U3156 (N_3156,N_3039,N_3056);
nand U3157 (N_3157,N_3148,N_3079);
and U3158 (N_3158,N_3012,N_3098);
or U3159 (N_3159,N_3114,N_3144);
nand U3160 (N_3160,N_3067,N_3095);
and U3161 (N_3161,N_3049,N_3085);
xor U3162 (N_3162,N_3010,N_3076);
and U3163 (N_3163,N_3033,N_3024);
xor U3164 (N_3164,N_3038,N_3134);
nor U3165 (N_3165,N_3022,N_3060);
nand U3166 (N_3166,N_3058,N_3140);
nor U3167 (N_3167,N_3073,N_3020);
and U3168 (N_3168,N_3002,N_3102);
xnor U3169 (N_3169,N_3072,N_3126);
nor U3170 (N_3170,N_3115,N_3054);
nor U3171 (N_3171,N_3104,N_3078);
nand U3172 (N_3172,N_3041,N_3121);
nor U3173 (N_3173,N_3088,N_3129);
nand U3174 (N_3174,N_3145,N_3003);
nor U3175 (N_3175,N_3040,N_3127);
or U3176 (N_3176,N_3028,N_3089);
or U3177 (N_3177,N_3015,N_3023);
and U3178 (N_3178,N_3069,N_3000);
xnor U3179 (N_3179,N_3030,N_3025);
xnor U3180 (N_3180,N_3014,N_3139);
nor U3181 (N_3181,N_3027,N_3042);
or U3182 (N_3182,N_3086,N_3111);
and U3183 (N_3183,N_3108,N_3064);
or U3184 (N_3184,N_3035,N_3034);
nor U3185 (N_3185,N_3131,N_3135);
and U3186 (N_3186,N_3081,N_3109);
or U3187 (N_3187,N_3092,N_3103);
and U3188 (N_3188,N_3013,N_3055);
and U3189 (N_3189,N_3004,N_3087);
or U3190 (N_3190,N_3063,N_3071);
nor U3191 (N_3191,N_3066,N_3105);
xnor U3192 (N_3192,N_3133,N_3062);
nor U3193 (N_3193,N_3100,N_3051);
or U3194 (N_3194,N_3107,N_3009);
xor U3195 (N_3195,N_3117,N_3119);
nor U3196 (N_3196,N_3147,N_3093);
nor U3197 (N_3197,N_3143,N_3007);
nor U3198 (N_3198,N_3017,N_3080);
xnor U3199 (N_3199,N_3090,N_3057);
and U3200 (N_3200,N_3074,N_3036);
or U3201 (N_3201,N_3021,N_3130);
or U3202 (N_3202,N_3083,N_3096);
nand U3203 (N_3203,N_3068,N_3113);
nand U3204 (N_3204,N_3032,N_3137);
nand U3205 (N_3205,N_3124,N_3142);
or U3206 (N_3206,N_3016,N_3006);
nand U3207 (N_3207,N_3008,N_3059);
and U3208 (N_3208,N_3094,N_3044);
and U3209 (N_3209,N_3011,N_3128);
xnor U3210 (N_3210,N_3149,N_3075);
nor U3211 (N_3211,N_3120,N_3019);
or U3212 (N_3212,N_3138,N_3047);
nand U3213 (N_3213,N_3106,N_3132);
xnor U3214 (N_3214,N_3125,N_3136);
nand U3215 (N_3215,N_3048,N_3077);
or U3216 (N_3216,N_3046,N_3118);
nor U3217 (N_3217,N_3116,N_3031);
nor U3218 (N_3218,N_3037,N_3026);
or U3219 (N_3219,N_3084,N_3029);
nor U3220 (N_3220,N_3005,N_3001);
nor U3221 (N_3221,N_3099,N_3018);
and U3222 (N_3222,N_3065,N_3141);
and U3223 (N_3223,N_3043,N_3091);
xnor U3224 (N_3224,N_3052,N_3146);
nor U3225 (N_3225,N_3003,N_3034);
xnor U3226 (N_3226,N_3117,N_3148);
or U3227 (N_3227,N_3071,N_3119);
xnor U3228 (N_3228,N_3068,N_3087);
nor U3229 (N_3229,N_3111,N_3050);
and U3230 (N_3230,N_3117,N_3141);
and U3231 (N_3231,N_3127,N_3132);
or U3232 (N_3232,N_3002,N_3084);
and U3233 (N_3233,N_3065,N_3006);
or U3234 (N_3234,N_3132,N_3039);
xor U3235 (N_3235,N_3024,N_3015);
or U3236 (N_3236,N_3099,N_3116);
and U3237 (N_3237,N_3132,N_3019);
or U3238 (N_3238,N_3035,N_3006);
nand U3239 (N_3239,N_3020,N_3043);
nand U3240 (N_3240,N_3138,N_3087);
nand U3241 (N_3241,N_3145,N_3058);
and U3242 (N_3242,N_3114,N_3079);
xor U3243 (N_3243,N_3072,N_3100);
or U3244 (N_3244,N_3037,N_3070);
xor U3245 (N_3245,N_3146,N_3065);
nor U3246 (N_3246,N_3052,N_3119);
and U3247 (N_3247,N_3131,N_3099);
and U3248 (N_3248,N_3054,N_3037);
and U3249 (N_3249,N_3140,N_3044);
and U3250 (N_3250,N_3035,N_3007);
xor U3251 (N_3251,N_3089,N_3108);
nand U3252 (N_3252,N_3139,N_3130);
nand U3253 (N_3253,N_3027,N_3108);
and U3254 (N_3254,N_3096,N_3065);
nor U3255 (N_3255,N_3140,N_3082);
xor U3256 (N_3256,N_3095,N_3029);
or U3257 (N_3257,N_3072,N_3067);
nand U3258 (N_3258,N_3070,N_3129);
and U3259 (N_3259,N_3101,N_3013);
nor U3260 (N_3260,N_3096,N_3122);
and U3261 (N_3261,N_3081,N_3049);
nand U3262 (N_3262,N_3065,N_3127);
nor U3263 (N_3263,N_3038,N_3050);
and U3264 (N_3264,N_3056,N_3005);
nand U3265 (N_3265,N_3065,N_3074);
xor U3266 (N_3266,N_3129,N_3120);
xnor U3267 (N_3267,N_3059,N_3029);
nand U3268 (N_3268,N_3078,N_3071);
and U3269 (N_3269,N_3084,N_3062);
nand U3270 (N_3270,N_3034,N_3121);
nor U3271 (N_3271,N_3133,N_3025);
or U3272 (N_3272,N_3025,N_3116);
nor U3273 (N_3273,N_3148,N_3027);
nand U3274 (N_3274,N_3100,N_3111);
nor U3275 (N_3275,N_3051,N_3075);
xor U3276 (N_3276,N_3114,N_3149);
or U3277 (N_3277,N_3044,N_3100);
nand U3278 (N_3278,N_3142,N_3079);
nor U3279 (N_3279,N_3072,N_3053);
and U3280 (N_3280,N_3148,N_3093);
or U3281 (N_3281,N_3076,N_3052);
or U3282 (N_3282,N_3104,N_3109);
and U3283 (N_3283,N_3085,N_3073);
xor U3284 (N_3284,N_3039,N_3116);
nor U3285 (N_3285,N_3132,N_3097);
or U3286 (N_3286,N_3053,N_3126);
nand U3287 (N_3287,N_3032,N_3133);
nor U3288 (N_3288,N_3028,N_3054);
nor U3289 (N_3289,N_3131,N_3026);
nor U3290 (N_3290,N_3130,N_3069);
xnor U3291 (N_3291,N_3137,N_3017);
xor U3292 (N_3292,N_3120,N_3115);
and U3293 (N_3293,N_3048,N_3001);
and U3294 (N_3294,N_3104,N_3086);
or U3295 (N_3295,N_3137,N_3105);
nor U3296 (N_3296,N_3095,N_3017);
xnor U3297 (N_3297,N_3104,N_3120);
nand U3298 (N_3298,N_3096,N_3070);
xor U3299 (N_3299,N_3141,N_3097);
nand U3300 (N_3300,N_3265,N_3259);
xnor U3301 (N_3301,N_3178,N_3220);
xnor U3302 (N_3302,N_3217,N_3266);
nand U3303 (N_3303,N_3272,N_3224);
and U3304 (N_3304,N_3226,N_3237);
xnor U3305 (N_3305,N_3181,N_3164);
and U3306 (N_3306,N_3299,N_3157);
or U3307 (N_3307,N_3161,N_3222);
nand U3308 (N_3308,N_3187,N_3212);
or U3309 (N_3309,N_3227,N_3241);
xor U3310 (N_3310,N_3193,N_3273);
nor U3311 (N_3311,N_3208,N_3160);
nand U3312 (N_3312,N_3196,N_3159);
nand U3313 (N_3313,N_3150,N_3213);
and U3314 (N_3314,N_3173,N_3278);
xor U3315 (N_3315,N_3295,N_3236);
or U3316 (N_3316,N_3205,N_3185);
and U3317 (N_3317,N_3169,N_3177);
or U3318 (N_3318,N_3297,N_3257);
and U3319 (N_3319,N_3230,N_3274);
nor U3320 (N_3320,N_3183,N_3249);
nor U3321 (N_3321,N_3240,N_3168);
and U3322 (N_3322,N_3290,N_3292);
or U3323 (N_3323,N_3293,N_3242);
nor U3324 (N_3324,N_3268,N_3235);
nand U3325 (N_3325,N_3234,N_3288);
nor U3326 (N_3326,N_3190,N_3247);
and U3327 (N_3327,N_3166,N_3206);
nor U3328 (N_3328,N_3195,N_3232);
nand U3329 (N_3329,N_3223,N_3194);
and U3330 (N_3330,N_3270,N_3152);
nand U3331 (N_3331,N_3219,N_3280);
nor U3332 (N_3332,N_3192,N_3228);
xor U3333 (N_3333,N_3244,N_3210);
xnor U3334 (N_3334,N_3170,N_3281);
nand U3335 (N_3335,N_3251,N_3179);
nand U3336 (N_3336,N_3277,N_3229);
nand U3337 (N_3337,N_3167,N_3260);
xnor U3338 (N_3338,N_3291,N_3180);
nand U3339 (N_3339,N_3182,N_3258);
nand U3340 (N_3340,N_3207,N_3162);
and U3341 (N_3341,N_3198,N_3191);
or U3342 (N_3342,N_3248,N_3282);
nor U3343 (N_3343,N_3284,N_3254);
nor U3344 (N_3344,N_3252,N_3209);
and U3345 (N_3345,N_3184,N_3188);
nand U3346 (N_3346,N_3174,N_3239);
nor U3347 (N_3347,N_3151,N_3250);
xor U3348 (N_3348,N_3154,N_3201);
and U3349 (N_3349,N_3218,N_3221);
nand U3350 (N_3350,N_3298,N_3216);
nor U3351 (N_3351,N_3264,N_3286);
nor U3352 (N_3352,N_3225,N_3199);
xnor U3353 (N_3353,N_3172,N_3163);
and U3354 (N_3354,N_3246,N_3289);
or U3355 (N_3355,N_3267,N_3271);
nand U3356 (N_3356,N_3283,N_3186);
xnor U3357 (N_3357,N_3287,N_3197);
xnor U3358 (N_3358,N_3263,N_3175);
nand U3359 (N_3359,N_3171,N_3262);
and U3360 (N_3360,N_3215,N_3231);
xnor U3361 (N_3361,N_3165,N_3200);
xor U3362 (N_3362,N_3158,N_3189);
nor U3363 (N_3363,N_3256,N_3176);
nand U3364 (N_3364,N_3214,N_3155);
xnor U3365 (N_3365,N_3285,N_3204);
xor U3366 (N_3366,N_3245,N_3156);
nor U3367 (N_3367,N_3203,N_3233);
nor U3368 (N_3368,N_3294,N_3253);
xnor U3369 (N_3369,N_3261,N_3153);
xnor U3370 (N_3370,N_3255,N_3296);
xnor U3371 (N_3371,N_3243,N_3269);
nand U3372 (N_3372,N_3276,N_3238);
nor U3373 (N_3373,N_3275,N_3279);
nor U3374 (N_3374,N_3202,N_3211);
or U3375 (N_3375,N_3240,N_3251);
xnor U3376 (N_3376,N_3187,N_3280);
xnor U3377 (N_3377,N_3197,N_3224);
nor U3378 (N_3378,N_3279,N_3292);
and U3379 (N_3379,N_3164,N_3294);
nand U3380 (N_3380,N_3170,N_3242);
nand U3381 (N_3381,N_3213,N_3172);
nand U3382 (N_3382,N_3268,N_3270);
and U3383 (N_3383,N_3218,N_3165);
nand U3384 (N_3384,N_3189,N_3234);
or U3385 (N_3385,N_3154,N_3236);
nor U3386 (N_3386,N_3263,N_3199);
nand U3387 (N_3387,N_3277,N_3153);
and U3388 (N_3388,N_3191,N_3274);
or U3389 (N_3389,N_3229,N_3248);
nand U3390 (N_3390,N_3154,N_3186);
xor U3391 (N_3391,N_3153,N_3193);
and U3392 (N_3392,N_3222,N_3169);
and U3393 (N_3393,N_3221,N_3161);
and U3394 (N_3394,N_3203,N_3283);
and U3395 (N_3395,N_3275,N_3210);
nor U3396 (N_3396,N_3210,N_3160);
xnor U3397 (N_3397,N_3226,N_3227);
nor U3398 (N_3398,N_3172,N_3205);
xnor U3399 (N_3399,N_3272,N_3218);
and U3400 (N_3400,N_3183,N_3244);
and U3401 (N_3401,N_3282,N_3168);
nand U3402 (N_3402,N_3189,N_3297);
nand U3403 (N_3403,N_3156,N_3213);
xor U3404 (N_3404,N_3163,N_3294);
and U3405 (N_3405,N_3289,N_3208);
or U3406 (N_3406,N_3241,N_3181);
xor U3407 (N_3407,N_3294,N_3268);
and U3408 (N_3408,N_3152,N_3298);
xor U3409 (N_3409,N_3177,N_3165);
nor U3410 (N_3410,N_3254,N_3155);
and U3411 (N_3411,N_3228,N_3213);
nor U3412 (N_3412,N_3168,N_3267);
and U3413 (N_3413,N_3202,N_3168);
nand U3414 (N_3414,N_3248,N_3222);
xnor U3415 (N_3415,N_3190,N_3150);
xor U3416 (N_3416,N_3212,N_3257);
and U3417 (N_3417,N_3286,N_3269);
nor U3418 (N_3418,N_3219,N_3226);
xnor U3419 (N_3419,N_3166,N_3247);
xor U3420 (N_3420,N_3259,N_3296);
nor U3421 (N_3421,N_3233,N_3256);
nor U3422 (N_3422,N_3170,N_3217);
and U3423 (N_3423,N_3162,N_3173);
nor U3424 (N_3424,N_3262,N_3196);
and U3425 (N_3425,N_3216,N_3209);
nand U3426 (N_3426,N_3247,N_3200);
xor U3427 (N_3427,N_3257,N_3221);
and U3428 (N_3428,N_3248,N_3263);
and U3429 (N_3429,N_3175,N_3221);
nor U3430 (N_3430,N_3269,N_3234);
nor U3431 (N_3431,N_3291,N_3235);
xor U3432 (N_3432,N_3200,N_3216);
xnor U3433 (N_3433,N_3240,N_3213);
nor U3434 (N_3434,N_3168,N_3157);
nor U3435 (N_3435,N_3150,N_3204);
and U3436 (N_3436,N_3253,N_3251);
and U3437 (N_3437,N_3280,N_3252);
xor U3438 (N_3438,N_3199,N_3179);
or U3439 (N_3439,N_3219,N_3218);
or U3440 (N_3440,N_3224,N_3288);
or U3441 (N_3441,N_3197,N_3158);
and U3442 (N_3442,N_3161,N_3244);
nor U3443 (N_3443,N_3196,N_3171);
nor U3444 (N_3444,N_3263,N_3189);
xnor U3445 (N_3445,N_3166,N_3230);
nand U3446 (N_3446,N_3204,N_3254);
xnor U3447 (N_3447,N_3150,N_3272);
or U3448 (N_3448,N_3240,N_3211);
or U3449 (N_3449,N_3169,N_3227);
nor U3450 (N_3450,N_3324,N_3415);
nor U3451 (N_3451,N_3395,N_3339);
xnor U3452 (N_3452,N_3365,N_3425);
xnor U3453 (N_3453,N_3333,N_3427);
nand U3454 (N_3454,N_3449,N_3306);
nand U3455 (N_3455,N_3404,N_3420);
and U3456 (N_3456,N_3335,N_3341);
nand U3457 (N_3457,N_3414,N_3399);
xor U3458 (N_3458,N_3442,N_3349);
nand U3459 (N_3459,N_3325,N_3434);
nand U3460 (N_3460,N_3428,N_3383);
xnor U3461 (N_3461,N_3374,N_3366);
and U3462 (N_3462,N_3326,N_3437);
or U3463 (N_3463,N_3301,N_3387);
nand U3464 (N_3464,N_3440,N_3444);
nand U3465 (N_3465,N_3358,N_3413);
nor U3466 (N_3466,N_3400,N_3369);
and U3467 (N_3467,N_3309,N_3344);
or U3468 (N_3468,N_3328,N_3410);
or U3469 (N_3469,N_3323,N_3360);
or U3470 (N_3470,N_3407,N_3350);
or U3471 (N_3471,N_3313,N_3429);
xnor U3472 (N_3472,N_3443,N_3319);
nand U3473 (N_3473,N_3375,N_3391);
or U3474 (N_3474,N_3378,N_3353);
and U3475 (N_3475,N_3435,N_3331);
xor U3476 (N_3476,N_3439,N_3438);
nand U3477 (N_3477,N_3364,N_3403);
nand U3478 (N_3478,N_3447,N_3385);
nand U3479 (N_3479,N_3408,N_3384);
and U3480 (N_3480,N_3315,N_3363);
xnor U3481 (N_3481,N_3307,N_3320);
and U3482 (N_3482,N_3377,N_3412);
and U3483 (N_3483,N_3343,N_3419);
nand U3484 (N_3484,N_3336,N_3340);
nand U3485 (N_3485,N_3421,N_3359);
or U3486 (N_3486,N_3386,N_3396);
or U3487 (N_3487,N_3357,N_3322);
nor U3488 (N_3488,N_3373,N_3446);
and U3489 (N_3489,N_3436,N_3372);
xnor U3490 (N_3490,N_3423,N_3448);
xnor U3491 (N_3491,N_3382,N_3345);
xor U3492 (N_3492,N_3416,N_3394);
and U3493 (N_3493,N_3371,N_3445);
and U3494 (N_3494,N_3332,N_3308);
nor U3495 (N_3495,N_3411,N_3389);
and U3496 (N_3496,N_3351,N_3418);
nand U3497 (N_3497,N_3424,N_3300);
nand U3498 (N_3498,N_3390,N_3314);
or U3499 (N_3499,N_3417,N_3338);
nand U3500 (N_3500,N_3330,N_3381);
xor U3501 (N_3501,N_3304,N_3342);
nand U3502 (N_3502,N_3370,N_3352);
nand U3503 (N_3503,N_3367,N_3327);
nor U3504 (N_3504,N_3441,N_3376);
or U3505 (N_3505,N_3406,N_3398);
nor U3506 (N_3506,N_3310,N_3317);
and U3507 (N_3507,N_3355,N_3432);
nor U3508 (N_3508,N_3393,N_3433);
nand U3509 (N_3509,N_3354,N_3405);
or U3510 (N_3510,N_3392,N_3379);
xnor U3511 (N_3511,N_3401,N_3426);
xnor U3512 (N_3512,N_3430,N_3329);
xnor U3513 (N_3513,N_3316,N_3337);
xnor U3514 (N_3514,N_3318,N_3321);
xnor U3515 (N_3515,N_3348,N_3422);
xnor U3516 (N_3516,N_3409,N_3346);
nand U3517 (N_3517,N_3302,N_3305);
or U3518 (N_3518,N_3361,N_3334);
nor U3519 (N_3519,N_3311,N_3347);
nor U3520 (N_3520,N_3303,N_3397);
nor U3521 (N_3521,N_3380,N_3388);
nor U3522 (N_3522,N_3402,N_3356);
xnor U3523 (N_3523,N_3312,N_3362);
xor U3524 (N_3524,N_3431,N_3368);
or U3525 (N_3525,N_3311,N_3433);
nor U3526 (N_3526,N_3340,N_3301);
nor U3527 (N_3527,N_3433,N_3310);
nand U3528 (N_3528,N_3351,N_3354);
xnor U3529 (N_3529,N_3361,N_3368);
nor U3530 (N_3530,N_3413,N_3417);
or U3531 (N_3531,N_3385,N_3404);
xor U3532 (N_3532,N_3367,N_3439);
nand U3533 (N_3533,N_3447,N_3327);
and U3534 (N_3534,N_3324,N_3444);
and U3535 (N_3535,N_3426,N_3335);
or U3536 (N_3536,N_3383,N_3361);
or U3537 (N_3537,N_3421,N_3420);
xnor U3538 (N_3538,N_3382,N_3359);
nor U3539 (N_3539,N_3381,N_3448);
and U3540 (N_3540,N_3394,N_3408);
and U3541 (N_3541,N_3306,N_3355);
and U3542 (N_3542,N_3378,N_3314);
and U3543 (N_3543,N_3307,N_3393);
nand U3544 (N_3544,N_3378,N_3409);
and U3545 (N_3545,N_3342,N_3364);
xnor U3546 (N_3546,N_3442,N_3432);
nand U3547 (N_3547,N_3300,N_3329);
and U3548 (N_3548,N_3409,N_3305);
xor U3549 (N_3549,N_3408,N_3347);
nor U3550 (N_3550,N_3331,N_3354);
and U3551 (N_3551,N_3423,N_3429);
or U3552 (N_3552,N_3302,N_3370);
nor U3553 (N_3553,N_3404,N_3358);
nand U3554 (N_3554,N_3419,N_3350);
nand U3555 (N_3555,N_3315,N_3417);
or U3556 (N_3556,N_3309,N_3444);
nand U3557 (N_3557,N_3412,N_3347);
and U3558 (N_3558,N_3368,N_3369);
xor U3559 (N_3559,N_3373,N_3404);
nand U3560 (N_3560,N_3443,N_3402);
nor U3561 (N_3561,N_3402,N_3395);
xnor U3562 (N_3562,N_3321,N_3394);
nor U3563 (N_3563,N_3375,N_3359);
nor U3564 (N_3564,N_3362,N_3300);
or U3565 (N_3565,N_3420,N_3386);
nand U3566 (N_3566,N_3405,N_3356);
xnor U3567 (N_3567,N_3330,N_3366);
and U3568 (N_3568,N_3368,N_3342);
nor U3569 (N_3569,N_3320,N_3336);
nand U3570 (N_3570,N_3360,N_3405);
nand U3571 (N_3571,N_3407,N_3372);
and U3572 (N_3572,N_3300,N_3395);
nor U3573 (N_3573,N_3401,N_3318);
and U3574 (N_3574,N_3440,N_3398);
xor U3575 (N_3575,N_3309,N_3312);
and U3576 (N_3576,N_3361,N_3371);
xor U3577 (N_3577,N_3408,N_3428);
nand U3578 (N_3578,N_3310,N_3350);
and U3579 (N_3579,N_3314,N_3446);
xor U3580 (N_3580,N_3339,N_3301);
nand U3581 (N_3581,N_3432,N_3383);
xnor U3582 (N_3582,N_3338,N_3334);
nand U3583 (N_3583,N_3444,N_3379);
nand U3584 (N_3584,N_3400,N_3389);
or U3585 (N_3585,N_3432,N_3352);
or U3586 (N_3586,N_3447,N_3407);
xnor U3587 (N_3587,N_3441,N_3448);
nand U3588 (N_3588,N_3368,N_3378);
nor U3589 (N_3589,N_3310,N_3323);
nor U3590 (N_3590,N_3338,N_3336);
xnor U3591 (N_3591,N_3318,N_3341);
and U3592 (N_3592,N_3307,N_3314);
xnor U3593 (N_3593,N_3371,N_3342);
and U3594 (N_3594,N_3346,N_3324);
or U3595 (N_3595,N_3327,N_3446);
and U3596 (N_3596,N_3423,N_3444);
xnor U3597 (N_3597,N_3354,N_3427);
xnor U3598 (N_3598,N_3433,N_3446);
nand U3599 (N_3599,N_3409,N_3357);
xnor U3600 (N_3600,N_3529,N_3585);
xnor U3601 (N_3601,N_3514,N_3521);
nor U3602 (N_3602,N_3583,N_3554);
nand U3603 (N_3603,N_3573,N_3473);
or U3604 (N_3604,N_3456,N_3475);
and U3605 (N_3605,N_3485,N_3450);
nor U3606 (N_3606,N_3541,N_3537);
nand U3607 (N_3607,N_3518,N_3566);
and U3608 (N_3608,N_3551,N_3539);
or U3609 (N_3609,N_3580,N_3451);
and U3610 (N_3610,N_3477,N_3463);
nand U3611 (N_3611,N_3496,N_3457);
nor U3612 (N_3612,N_3474,N_3568);
nand U3613 (N_3613,N_3587,N_3593);
xnor U3614 (N_3614,N_3507,N_3502);
xor U3615 (N_3615,N_3506,N_3527);
nor U3616 (N_3616,N_3552,N_3523);
and U3617 (N_3617,N_3486,N_3516);
nand U3618 (N_3618,N_3536,N_3522);
and U3619 (N_3619,N_3520,N_3563);
nand U3620 (N_3620,N_3581,N_3543);
nor U3621 (N_3621,N_3578,N_3510);
xor U3622 (N_3622,N_3576,N_3598);
nand U3623 (N_3623,N_3482,N_3586);
nor U3624 (N_3624,N_3567,N_3530);
and U3625 (N_3625,N_3540,N_3542);
nor U3626 (N_3626,N_3517,N_3584);
and U3627 (N_3627,N_3558,N_3575);
and U3628 (N_3628,N_3579,N_3546);
nor U3629 (N_3629,N_3462,N_3511);
nor U3630 (N_3630,N_3533,N_3508);
nand U3631 (N_3631,N_3478,N_3498);
and U3632 (N_3632,N_3479,N_3549);
xnor U3633 (N_3633,N_3505,N_3509);
and U3634 (N_3634,N_3548,N_3545);
xor U3635 (N_3635,N_3562,N_3513);
xnor U3636 (N_3636,N_3515,N_3564);
and U3637 (N_3637,N_3531,N_3495);
and U3638 (N_3638,N_3492,N_3550);
or U3639 (N_3639,N_3499,N_3544);
nor U3640 (N_3640,N_3465,N_3582);
xnor U3641 (N_3641,N_3455,N_3452);
nor U3642 (N_3642,N_3488,N_3487);
xor U3643 (N_3643,N_3472,N_3476);
nor U3644 (N_3644,N_3553,N_3469);
nand U3645 (N_3645,N_3577,N_3560);
nor U3646 (N_3646,N_3572,N_3466);
or U3647 (N_3647,N_3570,N_3458);
nand U3648 (N_3648,N_3524,N_3459);
or U3649 (N_3649,N_3519,N_3470);
or U3650 (N_3650,N_3483,N_3561);
xor U3651 (N_3651,N_3526,N_3569);
xor U3652 (N_3652,N_3512,N_3591);
nand U3653 (N_3653,N_3501,N_3594);
xnor U3654 (N_3654,N_3504,N_3491);
xnor U3655 (N_3655,N_3493,N_3480);
nor U3656 (N_3656,N_3464,N_3532);
and U3657 (N_3657,N_3590,N_3565);
nand U3658 (N_3658,N_3497,N_3571);
or U3659 (N_3659,N_3468,N_3471);
nand U3660 (N_3660,N_3589,N_3453);
xor U3661 (N_3661,N_3461,N_3489);
xnor U3662 (N_3662,N_3547,N_3595);
nor U3663 (N_3663,N_3460,N_3559);
and U3664 (N_3664,N_3525,N_3503);
xor U3665 (N_3665,N_3535,N_3494);
and U3666 (N_3666,N_3597,N_3467);
nand U3667 (N_3667,N_3556,N_3484);
and U3668 (N_3668,N_3596,N_3599);
nor U3669 (N_3669,N_3528,N_3588);
or U3670 (N_3670,N_3574,N_3557);
xnor U3671 (N_3671,N_3555,N_3592);
and U3672 (N_3672,N_3538,N_3490);
nor U3673 (N_3673,N_3534,N_3500);
nor U3674 (N_3674,N_3481,N_3454);
or U3675 (N_3675,N_3588,N_3592);
and U3676 (N_3676,N_3548,N_3525);
or U3677 (N_3677,N_3476,N_3590);
or U3678 (N_3678,N_3588,N_3586);
xor U3679 (N_3679,N_3548,N_3451);
xor U3680 (N_3680,N_3494,N_3477);
and U3681 (N_3681,N_3470,N_3527);
xnor U3682 (N_3682,N_3545,N_3482);
and U3683 (N_3683,N_3566,N_3459);
or U3684 (N_3684,N_3479,N_3462);
nand U3685 (N_3685,N_3582,N_3553);
nor U3686 (N_3686,N_3549,N_3582);
nand U3687 (N_3687,N_3538,N_3542);
or U3688 (N_3688,N_3560,N_3591);
nand U3689 (N_3689,N_3491,N_3526);
nor U3690 (N_3690,N_3577,N_3584);
or U3691 (N_3691,N_3513,N_3570);
xor U3692 (N_3692,N_3452,N_3556);
and U3693 (N_3693,N_3560,N_3464);
xnor U3694 (N_3694,N_3469,N_3549);
xor U3695 (N_3695,N_3538,N_3594);
or U3696 (N_3696,N_3459,N_3539);
or U3697 (N_3697,N_3507,N_3538);
nand U3698 (N_3698,N_3559,N_3557);
nor U3699 (N_3699,N_3503,N_3526);
and U3700 (N_3700,N_3495,N_3525);
xnor U3701 (N_3701,N_3533,N_3599);
xnor U3702 (N_3702,N_3450,N_3507);
nand U3703 (N_3703,N_3566,N_3488);
nor U3704 (N_3704,N_3483,N_3540);
nand U3705 (N_3705,N_3461,N_3522);
xor U3706 (N_3706,N_3513,N_3597);
xor U3707 (N_3707,N_3511,N_3528);
or U3708 (N_3708,N_3464,N_3556);
or U3709 (N_3709,N_3535,N_3462);
xor U3710 (N_3710,N_3493,N_3478);
and U3711 (N_3711,N_3492,N_3456);
or U3712 (N_3712,N_3544,N_3568);
nand U3713 (N_3713,N_3479,N_3569);
or U3714 (N_3714,N_3486,N_3483);
xnor U3715 (N_3715,N_3514,N_3574);
nor U3716 (N_3716,N_3503,N_3516);
or U3717 (N_3717,N_3576,N_3484);
and U3718 (N_3718,N_3453,N_3521);
nand U3719 (N_3719,N_3526,N_3473);
xor U3720 (N_3720,N_3553,N_3593);
xor U3721 (N_3721,N_3487,N_3500);
nor U3722 (N_3722,N_3526,N_3570);
nand U3723 (N_3723,N_3455,N_3530);
nand U3724 (N_3724,N_3456,N_3485);
xnor U3725 (N_3725,N_3471,N_3460);
xnor U3726 (N_3726,N_3591,N_3485);
and U3727 (N_3727,N_3476,N_3585);
and U3728 (N_3728,N_3530,N_3597);
and U3729 (N_3729,N_3594,N_3473);
nand U3730 (N_3730,N_3598,N_3461);
nand U3731 (N_3731,N_3470,N_3557);
xnor U3732 (N_3732,N_3575,N_3490);
and U3733 (N_3733,N_3467,N_3460);
xnor U3734 (N_3734,N_3453,N_3459);
and U3735 (N_3735,N_3536,N_3491);
or U3736 (N_3736,N_3567,N_3571);
and U3737 (N_3737,N_3572,N_3499);
xor U3738 (N_3738,N_3566,N_3477);
and U3739 (N_3739,N_3454,N_3589);
and U3740 (N_3740,N_3532,N_3545);
or U3741 (N_3741,N_3571,N_3475);
nor U3742 (N_3742,N_3584,N_3513);
xor U3743 (N_3743,N_3507,N_3569);
nand U3744 (N_3744,N_3493,N_3565);
xor U3745 (N_3745,N_3489,N_3594);
nor U3746 (N_3746,N_3473,N_3596);
nand U3747 (N_3747,N_3541,N_3451);
and U3748 (N_3748,N_3568,N_3463);
xor U3749 (N_3749,N_3545,N_3565);
or U3750 (N_3750,N_3686,N_3687);
and U3751 (N_3751,N_3679,N_3601);
or U3752 (N_3752,N_3658,N_3627);
nand U3753 (N_3753,N_3656,N_3628);
and U3754 (N_3754,N_3654,N_3659);
xnor U3755 (N_3755,N_3700,N_3634);
and U3756 (N_3756,N_3643,N_3640);
nand U3757 (N_3757,N_3690,N_3729);
or U3758 (N_3758,N_3615,N_3709);
nor U3759 (N_3759,N_3630,N_3617);
nor U3760 (N_3760,N_3607,N_3741);
and U3761 (N_3761,N_3663,N_3653);
or U3762 (N_3762,N_3684,N_3675);
nand U3763 (N_3763,N_3667,N_3747);
or U3764 (N_3764,N_3662,N_3676);
and U3765 (N_3765,N_3665,N_3735);
or U3766 (N_3766,N_3714,N_3603);
nand U3767 (N_3767,N_3613,N_3704);
nand U3768 (N_3768,N_3695,N_3638);
or U3769 (N_3769,N_3621,N_3723);
nand U3770 (N_3770,N_3652,N_3733);
nand U3771 (N_3771,N_3701,N_3651);
nor U3772 (N_3772,N_3710,N_3673);
xor U3773 (N_3773,N_3713,N_3619);
nand U3774 (N_3774,N_3722,N_3718);
nor U3775 (N_3775,N_3626,N_3728);
and U3776 (N_3776,N_3648,N_3683);
nor U3777 (N_3777,N_3711,N_3748);
or U3778 (N_3778,N_3641,N_3719);
nand U3779 (N_3779,N_3698,N_3660);
or U3780 (N_3780,N_3730,N_3670);
or U3781 (N_3781,N_3632,N_3642);
nand U3782 (N_3782,N_3602,N_3604);
nor U3783 (N_3783,N_3623,N_3639);
nand U3784 (N_3784,N_3631,N_3649);
nor U3785 (N_3785,N_3629,N_3666);
and U3786 (N_3786,N_3600,N_3669);
nand U3787 (N_3787,N_3678,N_3739);
or U3788 (N_3788,N_3744,N_3740);
and U3789 (N_3789,N_3696,N_3635);
or U3790 (N_3790,N_3726,N_3693);
xor U3791 (N_3791,N_3672,N_3708);
xnor U3792 (N_3792,N_3720,N_3655);
nand U3793 (N_3793,N_3705,N_3688);
nand U3794 (N_3794,N_3717,N_3738);
or U3795 (N_3795,N_3606,N_3707);
nand U3796 (N_3796,N_3681,N_3732);
and U3797 (N_3797,N_3742,N_3682);
nand U3798 (N_3798,N_3625,N_3745);
nand U3799 (N_3799,N_3605,N_3715);
nor U3800 (N_3800,N_3612,N_3661);
xor U3801 (N_3801,N_3637,N_3685);
nor U3802 (N_3802,N_3724,N_3614);
nor U3803 (N_3803,N_3680,N_3727);
nor U3804 (N_3804,N_3636,N_3706);
nand U3805 (N_3805,N_3725,N_3610);
and U3806 (N_3806,N_3734,N_3749);
xnor U3807 (N_3807,N_3674,N_3691);
and U3808 (N_3808,N_3699,N_3677);
xor U3809 (N_3809,N_3743,N_3712);
nor U3810 (N_3810,N_3620,N_3616);
nand U3811 (N_3811,N_3608,N_3611);
xnor U3812 (N_3812,N_3689,N_3731);
and U3813 (N_3813,N_3657,N_3721);
nor U3814 (N_3814,N_3737,N_3668);
nor U3815 (N_3815,N_3702,N_3716);
or U3816 (N_3816,N_3622,N_3646);
nor U3817 (N_3817,N_3694,N_3647);
xor U3818 (N_3818,N_3609,N_3618);
nand U3819 (N_3819,N_3633,N_3671);
xnor U3820 (N_3820,N_3697,N_3650);
and U3821 (N_3821,N_3692,N_3644);
and U3822 (N_3822,N_3736,N_3746);
nor U3823 (N_3823,N_3624,N_3645);
nand U3824 (N_3824,N_3664,N_3703);
nor U3825 (N_3825,N_3655,N_3642);
nor U3826 (N_3826,N_3659,N_3653);
xnor U3827 (N_3827,N_3737,N_3676);
nor U3828 (N_3828,N_3616,N_3615);
nand U3829 (N_3829,N_3621,N_3707);
nand U3830 (N_3830,N_3699,N_3602);
nand U3831 (N_3831,N_3667,N_3660);
nand U3832 (N_3832,N_3632,N_3707);
xor U3833 (N_3833,N_3621,N_3652);
nand U3834 (N_3834,N_3733,N_3663);
or U3835 (N_3835,N_3658,N_3735);
and U3836 (N_3836,N_3610,N_3603);
xnor U3837 (N_3837,N_3687,N_3619);
xor U3838 (N_3838,N_3641,N_3738);
xnor U3839 (N_3839,N_3738,N_3733);
xor U3840 (N_3840,N_3606,N_3616);
nand U3841 (N_3841,N_3727,N_3691);
and U3842 (N_3842,N_3633,N_3730);
or U3843 (N_3843,N_3726,N_3707);
nor U3844 (N_3844,N_3604,N_3663);
xnor U3845 (N_3845,N_3732,N_3736);
or U3846 (N_3846,N_3656,N_3633);
xor U3847 (N_3847,N_3692,N_3614);
nand U3848 (N_3848,N_3696,N_3737);
and U3849 (N_3849,N_3707,N_3627);
nor U3850 (N_3850,N_3643,N_3664);
and U3851 (N_3851,N_3698,N_3702);
and U3852 (N_3852,N_3663,N_3714);
nand U3853 (N_3853,N_3616,N_3669);
xor U3854 (N_3854,N_3684,N_3623);
nor U3855 (N_3855,N_3723,N_3689);
and U3856 (N_3856,N_3659,N_3687);
nand U3857 (N_3857,N_3661,N_3633);
nor U3858 (N_3858,N_3641,N_3657);
nor U3859 (N_3859,N_3637,N_3649);
xnor U3860 (N_3860,N_3737,N_3692);
or U3861 (N_3861,N_3615,N_3622);
nand U3862 (N_3862,N_3706,N_3661);
xor U3863 (N_3863,N_3652,N_3628);
nor U3864 (N_3864,N_3680,N_3600);
and U3865 (N_3865,N_3684,N_3605);
or U3866 (N_3866,N_3622,N_3634);
nor U3867 (N_3867,N_3688,N_3624);
or U3868 (N_3868,N_3660,N_3716);
nand U3869 (N_3869,N_3671,N_3699);
and U3870 (N_3870,N_3623,N_3601);
nor U3871 (N_3871,N_3668,N_3632);
xor U3872 (N_3872,N_3644,N_3668);
and U3873 (N_3873,N_3663,N_3606);
or U3874 (N_3874,N_3612,N_3687);
xor U3875 (N_3875,N_3613,N_3605);
or U3876 (N_3876,N_3746,N_3743);
or U3877 (N_3877,N_3700,N_3710);
xor U3878 (N_3878,N_3708,N_3700);
nor U3879 (N_3879,N_3607,N_3701);
nand U3880 (N_3880,N_3637,N_3667);
and U3881 (N_3881,N_3715,N_3683);
or U3882 (N_3882,N_3642,N_3639);
nor U3883 (N_3883,N_3625,N_3679);
nand U3884 (N_3884,N_3652,N_3661);
xor U3885 (N_3885,N_3711,N_3641);
xor U3886 (N_3886,N_3651,N_3671);
and U3887 (N_3887,N_3691,N_3728);
and U3888 (N_3888,N_3659,N_3663);
xnor U3889 (N_3889,N_3695,N_3735);
nand U3890 (N_3890,N_3649,N_3688);
nor U3891 (N_3891,N_3715,N_3712);
nor U3892 (N_3892,N_3747,N_3638);
nor U3893 (N_3893,N_3693,N_3663);
nor U3894 (N_3894,N_3741,N_3620);
xnor U3895 (N_3895,N_3711,N_3701);
and U3896 (N_3896,N_3689,N_3684);
and U3897 (N_3897,N_3676,N_3645);
nand U3898 (N_3898,N_3603,N_3685);
and U3899 (N_3899,N_3634,N_3626);
nor U3900 (N_3900,N_3835,N_3796);
and U3901 (N_3901,N_3899,N_3889);
nand U3902 (N_3902,N_3789,N_3836);
nor U3903 (N_3903,N_3882,N_3773);
xor U3904 (N_3904,N_3777,N_3751);
nor U3905 (N_3905,N_3775,N_3764);
nor U3906 (N_3906,N_3793,N_3772);
nand U3907 (N_3907,N_3890,N_3824);
or U3908 (N_3908,N_3876,N_3818);
or U3909 (N_3909,N_3897,N_3830);
xor U3910 (N_3910,N_3837,N_3754);
nor U3911 (N_3911,N_3786,N_3875);
and U3912 (N_3912,N_3812,N_3866);
nand U3913 (N_3913,N_3771,N_3766);
or U3914 (N_3914,N_3828,N_3842);
and U3915 (N_3915,N_3778,N_3803);
or U3916 (N_3916,N_3829,N_3848);
or U3917 (N_3917,N_3809,N_3768);
and U3918 (N_3918,N_3854,N_3834);
nand U3919 (N_3919,N_3785,N_3805);
nand U3920 (N_3920,N_3867,N_3756);
nor U3921 (N_3921,N_3753,N_3801);
xor U3922 (N_3922,N_3826,N_3863);
nand U3923 (N_3923,N_3795,N_3841);
nor U3924 (N_3924,N_3877,N_3861);
and U3925 (N_3925,N_3891,N_3781);
or U3926 (N_3926,N_3847,N_3868);
nand U3927 (N_3927,N_3831,N_3816);
nand U3928 (N_3928,N_3871,N_3849);
or U3929 (N_3929,N_3758,N_3760);
or U3930 (N_3930,N_3878,N_3864);
or U3931 (N_3931,N_3832,N_3892);
nand U3932 (N_3932,N_3880,N_3791);
nor U3933 (N_3933,N_3757,N_3774);
or U3934 (N_3934,N_3788,N_3838);
and U3935 (N_3935,N_3762,N_3843);
nand U3936 (N_3936,N_3853,N_3845);
and U3937 (N_3937,N_3782,N_3800);
nor U3938 (N_3938,N_3894,N_3893);
nand U3939 (N_3939,N_3815,N_3851);
nor U3940 (N_3940,N_3783,N_3784);
nor U3941 (N_3941,N_3761,N_3833);
and U3942 (N_3942,N_3865,N_3879);
or U3943 (N_3943,N_3857,N_3881);
and U3944 (N_3944,N_3770,N_3898);
nor U3945 (N_3945,N_3817,N_3822);
and U3946 (N_3946,N_3895,N_3827);
nor U3947 (N_3947,N_3792,N_3872);
nor U3948 (N_3948,N_3811,N_3810);
and U3949 (N_3949,N_3763,N_3844);
and U3950 (N_3950,N_3797,N_3790);
or U3951 (N_3951,N_3856,N_3821);
or U3952 (N_3952,N_3769,N_3873);
and U3953 (N_3953,N_3886,N_3870);
nand U3954 (N_3954,N_3855,N_3806);
nor U3955 (N_3955,N_3823,N_3896);
nand U3956 (N_3956,N_3808,N_3825);
nor U3957 (N_3957,N_3814,N_3819);
xnor U3958 (N_3958,N_3862,N_3888);
nand U3959 (N_3959,N_3776,N_3852);
xor U3960 (N_3960,N_3850,N_3885);
or U3961 (N_3961,N_3807,N_3813);
or U3962 (N_3962,N_3869,N_3755);
nor U3963 (N_3963,N_3846,N_3883);
xnor U3964 (N_3964,N_3884,N_3820);
nor U3965 (N_3965,N_3887,N_3859);
xor U3966 (N_3966,N_3759,N_3780);
and U3967 (N_3967,N_3767,N_3798);
and U3968 (N_3968,N_3752,N_3794);
xor U3969 (N_3969,N_3804,N_3787);
and U3970 (N_3970,N_3839,N_3840);
or U3971 (N_3971,N_3799,N_3779);
and U3972 (N_3972,N_3858,N_3750);
nor U3973 (N_3973,N_3765,N_3802);
or U3974 (N_3974,N_3874,N_3860);
xnor U3975 (N_3975,N_3884,N_3828);
nand U3976 (N_3976,N_3874,N_3865);
nand U3977 (N_3977,N_3816,N_3780);
and U3978 (N_3978,N_3793,N_3849);
nand U3979 (N_3979,N_3790,N_3814);
xnor U3980 (N_3980,N_3771,N_3820);
nand U3981 (N_3981,N_3784,N_3767);
or U3982 (N_3982,N_3834,N_3813);
nand U3983 (N_3983,N_3891,N_3834);
and U3984 (N_3984,N_3769,N_3759);
or U3985 (N_3985,N_3831,N_3835);
nor U3986 (N_3986,N_3759,N_3854);
and U3987 (N_3987,N_3771,N_3872);
xor U3988 (N_3988,N_3883,N_3779);
or U3989 (N_3989,N_3832,N_3802);
nand U3990 (N_3990,N_3814,N_3876);
xor U3991 (N_3991,N_3816,N_3820);
xnor U3992 (N_3992,N_3816,N_3773);
xor U3993 (N_3993,N_3864,N_3826);
and U3994 (N_3994,N_3750,N_3753);
nor U3995 (N_3995,N_3837,N_3876);
nand U3996 (N_3996,N_3866,N_3750);
nand U3997 (N_3997,N_3803,N_3750);
nand U3998 (N_3998,N_3809,N_3808);
and U3999 (N_3999,N_3836,N_3790);
nor U4000 (N_4000,N_3890,N_3862);
or U4001 (N_4001,N_3884,N_3812);
nor U4002 (N_4002,N_3884,N_3853);
nand U4003 (N_4003,N_3769,N_3768);
and U4004 (N_4004,N_3892,N_3781);
or U4005 (N_4005,N_3750,N_3827);
nand U4006 (N_4006,N_3884,N_3872);
nand U4007 (N_4007,N_3806,N_3823);
nor U4008 (N_4008,N_3883,N_3758);
and U4009 (N_4009,N_3786,N_3886);
or U4010 (N_4010,N_3895,N_3824);
xor U4011 (N_4011,N_3772,N_3833);
nor U4012 (N_4012,N_3821,N_3899);
xor U4013 (N_4013,N_3766,N_3805);
nor U4014 (N_4014,N_3767,N_3799);
or U4015 (N_4015,N_3788,N_3860);
xor U4016 (N_4016,N_3810,N_3768);
or U4017 (N_4017,N_3810,N_3783);
nor U4018 (N_4018,N_3809,N_3830);
and U4019 (N_4019,N_3892,N_3877);
and U4020 (N_4020,N_3833,N_3786);
nor U4021 (N_4021,N_3842,N_3790);
nor U4022 (N_4022,N_3765,N_3883);
nand U4023 (N_4023,N_3795,N_3783);
nor U4024 (N_4024,N_3851,N_3800);
xnor U4025 (N_4025,N_3835,N_3785);
xnor U4026 (N_4026,N_3823,N_3837);
or U4027 (N_4027,N_3890,N_3816);
and U4028 (N_4028,N_3786,N_3795);
nor U4029 (N_4029,N_3801,N_3835);
nand U4030 (N_4030,N_3858,N_3777);
nand U4031 (N_4031,N_3809,N_3850);
nand U4032 (N_4032,N_3857,N_3757);
nor U4033 (N_4033,N_3758,N_3824);
nand U4034 (N_4034,N_3753,N_3854);
nand U4035 (N_4035,N_3839,N_3820);
or U4036 (N_4036,N_3894,N_3871);
and U4037 (N_4037,N_3846,N_3836);
nor U4038 (N_4038,N_3864,N_3758);
or U4039 (N_4039,N_3834,N_3847);
nor U4040 (N_4040,N_3804,N_3755);
or U4041 (N_4041,N_3794,N_3891);
and U4042 (N_4042,N_3829,N_3795);
nor U4043 (N_4043,N_3818,N_3770);
nand U4044 (N_4044,N_3888,N_3833);
or U4045 (N_4045,N_3833,N_3777);
nand U4046 (N_4046,N_3781,N_3834);
and U4047 (N_4047,N_3868,N_3885);
nand U4048 (N_4048,N_3890,N_3893);
xnor U4049 (N_4049,N_3807,N_3801);
and U4050 (N_4050,N_4044,N_4038);
or U4051 (N_4051,N_4008,N_4004);
or U4052 (N_4052,N_4022,N_3950);
nand U4053 (N_4053,N_3932,N_4026);
and U4054 (N_4054,N_3929,N_3973);
nand U4055 (N_4055,N_4002,N_3983);
and U4056 (N_4056,N_3905,N_3934);
nand U4057 (N_4057,N_3977,N_4041);
xnor U4058 (N_4058,N_3994,N_3923);
and U4059 (N_4059,N_4048,N_3976);
and U4060 (N_4060,N_3996,N_3967);
and U4061 (N_4061,N_4046,N_4015);
and U4062 (N_4062,N_3936,N_4030);
nand U4063 (N_4063,N_3908,N_4011);
xnor U4064 (N_4064,N_3988,N_3972);
xor U4065 (N_4065,N_4024,N_3942);
nand U4066 (N_4066,N_3917,N_3933);
or U4067 (N_4067,N_3904,N_3910);
and U4068 (N_4068,N_4023,N_3978);
nand U4069 (N_4069,N_4043,N_3963);
nor U4070 (N_4070,N_3943,N_4034);
nor U4071 (N_4071,N_3926,N_3939);
and U4072 (N_4072,N_3906,N_3991);
and U4073 (N_4073,N_3944,N_4027);
nand U4074 (N_4074,N_4017,N_3900);
or U4075 (N_4075,N_3916,N_3951);
and U4076 (N_4076,N_3907,N_4014);
nand U4077 (N_4077,N_3958,N_3953);
nand U4078 (N_4078,N_3989,N_3985);
xor U4079 (N_4079,N_4025,N_4020);
nor U4080 (N_4080,N_3961,N_3938);
nor U4081 (N_4081,N_3965,N_4031);
nand U4082 (N_4082,N_4007,N_3968);
xor U4083 (N_4083,N_3981,N_3971);
and U4084 (N_4084,N_3928,N_3992);
or U4085 (N_4085,N_3979,N_3964);
xor U4086 (N_4086,N_3935,N_3986);
nand U4087 (N_4087,N_4029,N_3921);
or U4088 (N_4088,N_3995,N_3975);
and U4089 (N_4089,N_3966,N_4032);
nand U4090 (N_4090,N_3980,N_4003);
xor U4091 (N_4091,N_3945,N_3997);
xor U4092 (N_4092,N_4021,N_4000);
nand U4093 (N_4093,N_3940,N_3999);
nand U4094 (N_4094,N_3937,N_3913);
nor U4095 (N_4095,N_4047,N_3962);
or U4096 (N_4096,N_4012,N_3915);
nor U4097 (N_4097,N_3924,N_3998);
or U4098 (N_4098,N_4045,N_3948);
nand U4099 (N_4099,N_3969,N_4016);
and U4100 (N_4100,N_3912,N_3909);
nand U4101 (N_4101,N_3987,N_4010);
nor U4102 (N_4102,N_3925,N_4028);
nor U4103 (N_4103,N_3927,N_3922);
xnor U4104 (N_4104,N_4013,N_3902);
and U4105 (N_4105,N_3974,N_4001);
and U4106 (N_4106,N_3959,N_4042);
nor U4107 (N_4107,N_4036,N_3914);
or U4108 (N_4108,N_3930,N_3984);
or U4109 (N_4109,N_4049,N_3982);
or U4110 (N_4110,N_3901,N_3949);
nand U4111 (N_4111,N_3903,N_3956);
or U4112 (N_4112,N_3931,N_3919);
nand U4113 (N_4113,N_4019,N_4018);
or U4114 (N_4114,N_3918,N_3970);
or U4115 (N_4115,N_3993,N_3957);
or U4116 (N_4116,N_3954,N_3960);
nor U4117 (N_4117,N_3947,N_4039);
or U4118 (N_4118,N_4040,N_3990);
or U4119 (N_4119,N_3920,N_4006);
and U4120 (N_4120,N_4037,N_3941);
and U4121 (N_4121,N_3955,N_4033);
nand U4122 (N_4122,N_4035,N_4009);
and U4123 (N_4123,N_3946,N_3952);
nor U4124 (N_4124,N_4005,N_3911);
xnor U4125 (N_4125,N_4040,N_4000);
xor U4126 (N_4126,N_4038,N_3978);
nor U4127 (N_4127,N_3940,N_3915);
nand U4128 (N_4128,N_3901,N_3917);
nand U4129 (N_4129,N_4049,N_3964);
or U4130 (N_4130,N_3939,N_3936);
nor U4131 (N_4131,N_3918,N_4041);
and U4132 (N_4132,N_4000,N_3998);
nor U4133 (N_4133,N_3924,N_3962);
nor U4134 (N_4134,N_3915,N_3952);
and U4135 (N_4135,N_3938,N_3916);
nand U4136 (N_4136,N_3954,N_3986);
nand U4137 (N_4137,N_3952,N_4025);
and U4138 (N_4138,N_4027,N_3987);
nand U4139 (N_4139,N_4003,N_3912);
nor U4140 (N_4140,N_3903,N_3931);
or U4141 (N_4141,N_3933,N_4042);
xor U4142 (N_4142,N_3916,N_3922);
or U4143 (N_4143,N_3906,N_3965);
and U4144 (N_4144,N_4039,N_3919);
or U4145 (N_4145,N_4035,N_3970);
nand U4146 (N_4146,N_3986,N_3998);
nor U4147 (N_4147,N_4030,N_4003);
or U4148 (N_4148,N_3912,N_3910);
and U4149 (N_4149,N_4011,N_3972);
and U4150 (N_4150,N_4041,N_3949);
and U4151 (N_4151,N_4047,N_3960);
and U4152 (N_4152,N_3915,N_3966);
and U4153 (N_4153,N_4012,N_3911);
and U4154 (N_4154,N_4010,N_3917);
and U4155 (N_4155,N_4011,N_3910);
nand U4156 (N_4156,N_4041,N_4023);
or U4157 (N_4157,N_3994,N_3978);
nand U4158 (N_4158,N_3988,N_4019);
and U4159 (N_4159,N_3933,N_3928);
nor U4160 (N_4160,N_4000,N_3958);
xor U4161 (N_4161,N_4019,N_3922);
nor U4162 (N_4162,N_3956,N_3955);
nor U4163 (N_4163,N_3923,N_4031);
xnor U4164 (N_4164,N_4039,N_4003);
nand U4165 (N_4165,N_3971,N_3923);
and U4166 (N_4166,N_3967,N_4015);
or U4167 (N_4167,N_4016,N_3932);
and U4168 (N_4168,N_3906,N_3908);
or U4169 (N_4169,N_3942,N_4047);
and U4170 (N_4170,N_3981,N_3967);
and U4171 (N_4171,N_4045,N_3956);
and U4172 (N_4172,N_4015,N_3908);
nor U4173 (N_4173,N_3929,N_3960);
or U4174 (N_4174,N_3963,N_3903);
nor U4175 (N_4175,N_3973,N_4045);
nand U4176 (N_4176,N_3986,N_3993);
nor U4177 (N_4177,N_3944,N_4039);
and U4178 (N_4178,N_3950,N_4036);
or U4179 (N_4179,N_3934,N_3943);
or U4180 (N_4180,N_3922,N_3972);
and U4181 (N_4181,N_3989,N_3956);
and U4182 (N_4182,N_4011,N_3953);
nand U4183 (N_4183,N_3936,N_3934);
or U4184 (N_4184,N_3963,N_4018);
nand U4185 (N_4185,N_3980,N_4031);
or U4186 (N_4186,N_3953,N_3940);
and U4187 (N_4187,N_3942,N_4002);
and U4188 (N_4188,N_3961,N_4009);
nor U4189 (N_4189,N_3976,N_3914);
and U4190 (N_4190,N_3918,N_3967);
nand U4191 (N_4191,N_3924,N_3979);
and U4192 (N_4192,N_3942,N_3935);
xor U4193 (N_4193,N_3912,N_3934);
nor U4194 (N_4194,N_3943,N_4011);
nand U4195 (N_4195,N_3969,N_3974);
xor U4196 (N_4196,N_4034,N_3902);
nor U4197 (N_4197,N_4011,N_3981);
nand U4198 (N_4198,N_3991,N_4039);
nand U4199 (N_4199,N_4015,N_3930);
nor U4200 (N_4200,N_4140,N_4159);
and U4201 (N_4201,N_4131,N_4085);
xnor U4202 (N_4202,N_4165,N_4100);
and U4203 (N_4203,N_4168,N_4145);
nand U4204 (N_4204,N_4171,N_4169);
or U4205 (N_4205,N_4080,N_4107);
and U4206 (N_4206,N_4097,N_4146);
nand U4207 (N_4207,N_4185,N_4110);
and U4208 (N_4208,N_4178,N_4139);
or U4209 (N_4209,N_4108,N_4106);
and U4210 (N_4210,N_4063,N_4102);
and U4211 (N_4211,N_4091,N_4114);
nor U4212 (N_4212,N_4153,N_4193);
nor U4213 (N_4213,N_4198,N_4104);
nor U4214 (N_4214,N_4088,N_4156);
nor U4215 (N_4215,N_4172,N_4113);
nor U4216 (N_4216,N_4116,N_4115);
xnor U4217 (N_4217,N_4136,N_4109);
nor U4218 (N_4218,N_4078,N_4167);
nand U4219 (N_4219,N_4187,N_4180);
xnor U4220 (N_4220,N_4074,N_4083);
and U4221 (N_4221,N_4123,N_4189);
nand U4222 (N_4222,N_4134,N_4150);
and U4223 (N_4223,N_4073,N_4191);
and U4224 (N_4224,N_4112,N_4059);
nor U4225 (N_4225,N_4164,N_4160);
xnor U4226 (N_4226,N_4166,N_4090);
and U4227 (N_4227,N_4183,N_4062);
xnor U4228 (N_4228,N_4119,N_4053);
and U4229 (N_4229,N_4126,N_4154);
nand U4230 (N_4230,N_4143,N_4184);
and U4231 (N_4231,N_4081,N_4196);
xnor U4232 (N_4232,N_4174,N_4130);
nand U4233 (N_4233,N_4142,N_4157);
nor U4234 (N_4234,N_4148,N_4067);
nor U4235 (N_4235,N_4163,N_4069);
xor U4236 (N_4236,N_4175,N_4176);
nor U4237 (N_4237,N_4066,N_4056);
and U4238 (N_4238,N_4132,N_4181);
and U4239 (N_4239,N_4095,N_4192);
and U4240 (N_4240,N_4099,N_4087);
nor U4241 (N_4241,N_4190,N_4161);
nor U4242 (N_4242,N_4179,N_4072);
nor U4243 (N_4243,N_4127,N_4060);
or U4244 (N_4244,N_4122,N_4151);
xor U4245 (N_4245,N_4050,N_4089);
or U4246 (N_4246,N_4186,N_4182);
nor U4247 (N_4247,N_4082,N_4077);
and U4248 (N_4248,N_4125,N_4135);
xor U4249 (N_4249,N_4057,N_4155);
and U4250 (N_4250,N_4118,N_4177);
xnor U4251 (N_4251,N_4117,N_4064);
nor U4252 (N_4252,N_4144,N_4197);
or U4253 (N_4253,N_4199,N_4068);
or U4254 (N_4254,N_4101,N_4075);
or U4255 (N_4255,N_4129,N_4070);
nand U4256 (N_4256,N_4188,N_4103);
or U4257 (N_4257,N_4141,N_4058);
or U4258 (N_4258,N_4111,N_4147);
nand U4259 (N_4259,N_4194,N_4137);
or U4260 (N_4260,N_4121,N_4124);
xnor U4261 (N_4261,N_4079,N_4054);
nand U4262 (N_4262,N_4133,N_4138);
or U4263 (N_4263,N_4061,N_4086);
xnor U4264 (N_4264,N_4071,N_4120);
and U4265 (N_4265,N_4162,N_4152);
or U4266 (N_4266,N_4092,N_4105);
xor U4267 (N_4267,N_4052,N_4170);
xnor U4268 (N_4268,N_4076,N_4093);
nand U4269 (N_4269,N_4065,N_4094);
and U4270 (N_4270,N_4128,N_4195);
or U4271 (N_4271,N_4098,N_4158);
xnor U4272 (N_4272,N_4173,N_4051);
nor U4273 (N_4273,N_4055,N_4096);
and U4274 (N_4274,N_4084,N_4149);
and U4275 (N_4275,N_4154,N_4087);
nor U4276 (N_4276,N_4192,N_4070);
nand U4277 (N_4277,N_4180,N_4152);
nor U4278 (N_4278,N_4192,N_4088);
xor U4279 (N_4279,N_4130,N_4094);
and U4280 (N_4280,N_4152,N_4125);
and U4281 (N_4281,N_4158,N_4126);
or U4282 (N_4282,N_4158,N_4167);
or U4283 (N_4283,N_4104,N_4116);
nand U4284 (N_4284,N_4169,N_4069);
nor U4285 (N_4285,N_4052,N_4051);
or U4286 (N_4286,N_4053,N_4194);
nor U4287 (N_4287,N_4059,N_4144);
nor U4288 (N_4288,N_4056,N_4110);
or U4289 (N_4289,N_4131,N_4125);
nor U4290 (N_4290,N_4058,N_4088);
nand U4291 (N_4291,N_4100,N_4166);
nor U4292 (N_4292,N_4139,N_4074);
or U4293 (N_4293,N_4112,N_4146);
and U4294 (N_4294,N_4074,N_4174);
or U4295 (N_4295,N_4073,N_4062);
and U4296 (N_4296,N_4063,N_4052);
nand U4297 (N_4297,N_4069,N_4056);
or U4298 (N_4298,N_4187,N_4175);
xor U4299 (N_4299,N_4133,N_4197);
nor U4300 (N_4300,N_4156,N_4050);
or U4301 (N_4301,N_4063,N_4058);
nor U4302 (N_4302,N_4149,N_4085);
and U4303 (N_4303,N_4138,N_4131);
nor U4304 (N_4304,N_4149,N_4117);
or U4305 (N_4305,N_4056,N_4053);
nand U4306 (N_4306,N_4192,N_4132);
nor U4307 (N_4307,N_4189,N_4137);
xor U4308 (N_4308,N_4151,N_4147);
nand U4309 (N_4309,N_4106,N_4061);
and U4310 (N_4310,N_4075,N_4185);
xor U4311 (N_4311,N_4162,N_4118);
xnor U4312 (N_4312,N_4107,N_4106);
or U4313 (N_4313,N_4107,N_4185);
xnor U4314 (N_4314,N_4085,N_4125);
or U4315 (N_4315,N_4131,N_4070);
nand U4316 (N_4316,N_4127,N_4059);
xor U4317 (N_4317,N_4107,N_4130);
and U4318 (N_4318,N_4101,N_4070);
and U4319 (N_4319,N_4111,N_4150);
and U4320 (N_4320,N_4105,N_4170);
and U4321 (N_4321,N_4102,N_4052);
xnor U4322 (N_4322,N_4069,N_4132);
nor U4323 (N_4323,N_4091,N_4110);
or U4324 (N_4324,N_4163,N_4128);
or U4325 (N_4325,N_4119,N_4152);
and U4326 (N_4326,N_4158,N_4123);
nand U4327 (N_4327,N_4151,N_4102);
xnor U4328 (N_4328,N_4121,N_4051);
nor U4329 (N_4329,N_4134,N_4153);
nand U4330 (N_4330,N_4090,N_4111);
nor U4331 (N_4331,N_4090,N_4164);
nand U4332 (N_4332,N_4087,N_4093);
nor U4333 (N_4333,N_4102,N_4154);
or U4334 (N_4334,N_4149,N_4186);
nand U4335 (N_4335,N_4107,N_4100);
and U4336 (N_4336,N_4147,N_4079);
nor U4337 (N_4337,N_4142,N_4069);
xnor U4338 (N_4338,N_4128,N_4091);
and U4339 (N_4339,N_4052,N_4140);
and U4340 (N_4340,N_4152,N_4106);
nor U4341 (N_4341,N_4098,N_4080);
nor U4342 (N_4342,N_4142,N_4088);
or U4343 (N_4343,N_4186,N_4116);
xnor U4344 (N_4344,N_4159,N_4128);
and U4345 (N_4345,N_4168,N_4151);
or U4346 (N_4346,N_4180,N_4178);
or U4347 (N_4347,N_4180,N_4087);
nand U4348 (N_4348,N_4136,N_4070);
nand U4349 (N_4349,N_4105,N_4123);
and U4350 (N_4350,N_4297,N_4241);
nor U4351 (N_4351,N_4205,N_4215);
or U4352 (N_4352,N_4289,N_4299);
xor U4353 (N_4353,N_4308,N_4275);
nor U4354 (N_4354,N_4228,N_4235);
xor U4355 (N_4355,N_4218,N_4283);
nor U4356 (N_4356,N_4236,N_4233);
nand U4357 (N_4357,N_4277,N_4312);
and U4358 (N_4358,N_4206,N_4260);
and U4359 (N_4359,N_4246,N_4325);
nor U4360 (N_4360,N_4295,N_4272);
xnor U4361 (N_4361,N_4225,N_4292);
xor U4362 (N_4362,N_4268,N_4224);
or U4363 (N_4363,N_4300,N_4262);
nand U4364 (N_4364,N_4238,N_4333);
or U4365 (N_4365,N_4222,N_4247);
xor U4366 (N_4366,N_4264,N_4254);
nand U4367 (N_4367,N_4344,N_4212);
xor U4368 (N_4368,N_4261,N_4230);
and U4369 (N_4369,N_4267,N_4332);
xnor U4370 (N_4370,N_4273,N_4282);
nand U4371 (N_4371,N_4338,N_4217);
nor U4372 (N_4372,N_4310,N_4326);
xor U4373 (N_4373,N_4263,N_4330);
nor U4374 (N_4374,N_4340,N_4303);
or U4375 (N_4375,N_4204,N_4278);
nand U4376 (N_4376,N_4324,N_4328);
and U4377 (N_4377,N_4223,N_4309);
or U4378 (N_4378,N_4311,N_4293);
nor U4379 (N_4379,N_4207,N_4280);
nand U4380 (N_4380,N_4231,N_4208);
or U4381 (N_4381,N_4347,N_4316);
xnor U4382 (N_4382,N_4251,N_4243);
nor U4383 (N_4383,N_4253,N_4334);
nand U4384 (N_4384,N_4346,N_4329);
and U4385 (N_4385,N_4276,N_4256);
nand U4386 (N_4386,N_4284,N_4302);
xor U4387 (N_4387,N_4336,N_4327);
nor U4388 (N_4388,N_4341,N_4318);
nand U4389 (N_4389,N_4305,N_4258);
and U4390 (N_4390,N_4287,N_4249);
or U4391 (N_4391,N_4210,N_4239);
or U4392 (N_4392,N_4322,N_4257);
or U4393 (N_4393,N_4245,N_4286);
nor U4394 (N_4394,N_4211,N_4294);
and U4395 (N_4395,N_4266,N_4234);
nor U4396 (N_4396,N_4342,N_4209);
and U4397 (N_4397,N_4214,N_4255);
or U4398 (N_4398,N_4242,N_4288);
and U4399 (N_4399,N_4269,N_4213);
nand U4400 (N_4400,N_4221,N_4271);
nand U4401 (N_4401,N_4219,N_4229);
and U4402 (N_4402,N_4343,N_4265);
and U4403 (N_4403,N_4270,N_4259);
or U4404 (N_4404,N_4307,N_4227);
xnor U4405 (N_4405,N_4290,N_4331);
nor U4406 (N_4406,N_4345,N_4248);
or U4407 (N_4407,N_4200,N_4244);
xor U4408 (N_4408,N_4320,N_4313);
and U4409 (N_4409,N_4232,N_4202);
nand U4410 (N_4410,N_4298,N_4201);
or U4411 (N_4411,N_4216,N_4291);
nand U4412 (N_4412,N_4348,N_4323);
nor U4413 (N_4413,N_4240,N_4321);
or U4414 (N_4414,N_4304,N_4317);
nor U4415 (N_4415,N_4349,N_4274);
or U4416 (N_4416,N_4279,N_4315);
and U4417 (N_4417,N_4203,N_4319);
nand U4418 (N_4418,N_4337,N_4226);
nor U4419 (N_4419,N_4335,N_4301);
nor U4420 (N_4420,N_4314,N_4281);
nor U4421 (N_4421,N_4306,N_4339);
xor U4422 (N_4422,N_4296,N_4250);
or U4423 (N_4423,N_4252,N_4285);
nand U4424 (N_4424,N_4237,N_4220);
or U4425 (N_4425,N_4269,N_4229);
xor U4426 (N_4426,N_4345,N_4281);
xor U4427 (N_4427,N_4301,N_4309);
and U4428 (N_4428,N_4230,N_4270);
nand U4429 (N_4429,N_4300,N_4264);
or U4430 (N_4430,N_4305,N_4247);
nand U4431 (N_4431,N_4309,N_4344);
xor U4432 (N_4432,N_4348,N_4246);
and U4433 (N_4433,N_4295,N_4342);
nor U4434 (N_4434,N_4269,N_4345);
xor U4435 (N_4435,N_4300,N_4344);
nand U4436 (N_4436,N_4284,N_4339);
or U4437 (N_4437,N_4306,N_4322);
or U4438 (N_4438,N_4211,N_4246);
nor U4439 (N_4439,N_4290,N_4243);
nand U4440 (N_4440,N_4202,N_4203);
nand U4441 (N_4441,N_4348,N_4347);
nand U4442 (N_4442,N_4265,N_4315);
nand U4443 (N_4443,N_4227,N_4264);
or U4444 (N_4444,N_4332,N_4281);
nand U4445 (N_4445,N_4215,N_4234);
nor U4446 (N_4446,N_4327,N_4328);
nand U4447 (N_4447,N_4283,N_4214);
or U4448 (N_4448,N_4318,N_4346);
xnor U4449 (N_4449,N_4205,N_4311);
nand U4450 (N_4450,N_4208,N_4200);
nand U4451 (N_4451,N_4264,N_4274);
or U4452 (N_4452,N_4334,N_4344);
xor U4453 (N_4453,N_4202,N_4218);
and U4454 (N_4454,N_4245,N_4225);
or U4455 (N_4455,N_4313,N_4338);
nor U4456 (N_4456,N_4296,N_4219);
or U4457 (N_4457,N_4280,N_4262);
nand U4458 (N_4458,N_4268,N_4339);
and U4459 (N_4459,N_4291,N_4234);
xnor U4460 (N_4460,N_4341,N_4269);
and U4461 (N_4461,N_4233,N_4330);
nand U4462 (N_4462,N_4330,N_4346);
nand U4463 (N_4463,N_4254,N_4249);
or U4464 (N_4464,N_4277,N_4337);
nand U4465 (N_4465,N_4310,N_4277);
nor U4466 (N_4466,N_4204,N_4295);
and U4467 (N_4467,N_4244,N_4304);
xnor U4468 (N_4468,N_4228,N_4332);
nor U4469 (N_4469,N_4251,N_4315);
and U4470 (N_4470,N_4340,N_4265);
or U4471 (N_4471,N_4265,N_4236);
xor U4472 (N_4472,N_4206,N_4332);
xor U4473 (N_4473,N_4219,N_4325);
or U4474 (N_4474,N_4216,N_4218);
nand U4475 (N_4475,N_4274,N_4260);
nand U4476 (N_4476,N_4227,N_4267);
and U4477 (N_4477,N_4256,N_4299);
nand U4478 (N_4478,N_4225,N_4229);
xor U4479 (N_4479,N_4220,N_4292);
and U4480 (N_4480,N_4278,N_4337);
or U4481 (N_4481,N_4227,N_4226);
and U4482 (N_4482,N_4203,N_4236);
nand U4483 (N_4483,N_4226,N_4210);
xnor U4484 (N_4484,N_4306,N_4219);
nor U4485 (N_4485,N_4298,N_4204);
and U4486 (N_4486,N_4213,N_4283);
and U4487 (N_4487,N_4303,N_4257);
nand U4488 (N_4488,N_4211,N_4345);
nand U4489 (N_4489,N_4304,N_4340);
nor U4490 (N_4490,N_4273,N_4290);
xor U4491 (N_4491,N_4339,N_4239);
nor U4492 (N_4492,N_4212,N_4207);
and U4493 (N_4493,N_4215,N_4200);
or U4494 (N_4494,N_4206,N_4281);
and U4495 (N_4495,N_4321,N_4344);
or U4496 (N_4496,N_4321,N_4268);
xor U4497 (N_4497,N_4219,N_4281);
or U4498 (N_4498,N_4262,N_4249);
or U4499 (N_4499,N_4213,N_4343);
nand U4500 (N_4500,N_4416,N_4350);
xor U4501 (N_4501,N_4428,N_4383);
and U4502 (N_4502,N_4358,N_4377);
nand U4503 (N_4503,N_4449,N_4393);
nand U4504 (N_4504,N_4414,N_4390);
and U4505 (N_4505,N_4433,N_4370);
xnor U4506 (N_4506,N_4485,N_4352);
nor U4507 (N_4507,N_4482,N_4472);
and U4508 (N_4508,N_4404,N_4469);
nor U4509 (N_4509,N_4395,N_4464);
nor U4510 (N_4510,N_4354,N_4412);
or U4511 (N_4511,N_4399,N_4458);
or U4512 (N_4512,N_4442,N_4415);
nand U4513 (N_4513,N_4438,N_4367);
xor U4514 (N_4514,N_4364,N_4391);
or U4515 (N_4515,N_4487,N_4479);
xnor U4516 (N_4516,N_4476,N_4398);
nor U4517 (N_4517,N_4466,N_4448);
nand U4518 (N_4518,N_4493,N_4489);
or U4519 (N_4519,N_4477,N_4436);
xor U4520 (N_4520,N_4380,N_4402);
and U4521 (N_4521,N_4351,N_4403);
nand U4522 (N_4522,N_4440,N_4473);
nor U4523 (N_4523,N_4446,N_4460);
or U4524 (N_4524,N_4392,N_4411);
nand U4525 (N_4525,N_4420,N_4407);
nor U4526 (N_4526,N_4375,N_4389);
and U4527 (N_4527,N_4397,N_4445);
or U4528 (N_4528,N_4447,N_4454);
or U4529 (N_4529,N_4491,N_4483);
nand U4530 (N_4530,N_4356,N_4456);
and U4531 (N_4531,N_4372,N_4429);
and U4532 (N_4532,N_4441,N_4388);
nor U4533 (N_4533,N_4384,N_4425);
and U4534 (N_4534,N_4386,N_4359);
and U4535 (N_4535,N_4462,N_4465);
and U4536 (N_4536,N_4421,N_4362);
xnor U4537 (N_4537,N_4451,N_4379);
or U4538 (N_4538,N_4475,N_4486);
and U4539 (N_4539,N_4490,N_4478);
xnor U4540 (N_4540,N_4357,N_4387);
nor U4541 (N_4541,N_4405,N_4366);
and U4542 (N_4542,N_4468,N_4385);
and U4543 (N_4543,N_4484,N_4426);
xor U4544 (N_4544,N_4492,N_4471);
nand U4545 (N_4545,N_4439,N_4363);
nand U4546 (N_4546,N_4400,N_4431);
xor U4547 (N_4547,N_4443,N_4396);
nor U4548 (N_4548,N_4408,N_4394);
nor U4549 (N_4549,N_4488,N_4437);
and U4550 (N_4550,N_4481,N_4498);
and U4551 (N_4551,N_4406,N_4453);
or U4552 (N_4552,N_4470,N_4463);
nand U4553 (N_4553,N_4474,N_4369);
nand U4554 (N_4554,N_4381,N_4424);
and U4555 (N_4555,N_4378,N_4419);
nor U4556 (N_4556,N_4376,N_4444);
xor U4557 (N_4557,N_4373,N_4360);
and U4558 (N_4558,N_4417,N_4361);
or U4559 (N_4559,N_4423,N_4459);
xor U4560 (N_4560,N_4382,N_4413);
nand U4561 (N_4561,N_4461,N_4499);
nor U4562 (N_4562,N_4457,N_4422);
or U4563 (N_4563,N_4432,N_4410);
nand U4564 (N_4564,N_4374,N_4365);
nor U4565 (N_4565,N_4368,N_4497);
xor U4566 (N_4566,N_4494,N_4467);
or U4567 (N_4567,N_4401,N_4418);
and U4568 (N_4568,N_4495,N_4353);
and U4569 (N_4569,N_4430,N_4496);
and U4570 (N_4570,N_4435,N_4427);
and U4571 (N_4571,N_4455,N_4452);
or U4572 (N_4572,N_4434,N_4371);
xor U4573 (N_4573,N_4480,N_4409);
and U4574 (N_4574,N_4355,N_4450);
and U4575 (N_4575,N_4368,N_4374);
or U4576 (N_4576,N_4472,N_4477);
or U4577 (N_4577,N_4384,N_4450);
nand U4578 (N_4578,N_4452,N_4441);
xor U4579 (N_4579,N_4491,N_4391);
nor U4580 (N_4580,N_4383,N_4490);
xor U4581 (N_4581,N_4486,N_4411);
xor U4582 (N_4582,N_4481,N_4419);
and U4583 (N_4583,N_4390,N_4392);
and U4584 (N_4584,N_4450,N_4439);
nor U4585 (N_4585,N_4361,N_4391);
or U4586 (N_4586,N_4463,N_4472);
nand U4587 (N_4587,N_4486,N_4493);
nand U4588 (N_4588,N_4428,N_4399);
nand U4589 (N_4589,N_4472,N_4439);
or U4590 (N_4590,N_4468,N_4421);
nor U4591 (N_4591,N_4387,N_4394);
xor U4592 (N_4592,N_4493,N_4445);
xnor U4593 (N_4593,N_4368,N_4489);
or U4594 (N_4594,N_4359,N_4351);
nand U4595 (N_4595,N_4404,N_4411);
or U4596 (N_4596,N_4430,N_4494);
xor U4597 (N_4597,N_4365,N_4401);
nor U4598 (N_4598,N_4482,N_4450);
xnor U4599 (N_4599,N_4477,N_4374);
or U4600 (N_4600,N_4392,N_4374);
nor U4601 (N_4601,N_4428,N_4445);
nor U4602 (N_4602,N_4468,N_4451);
nand U4603 (N_4603,N_4384,N_4364);
and U4604 (N_4604,N_4474,N_4366);
xor U4605 (N_4605,N_4474,N_4389);
and U4606 (N_4606,N_4451,N_4476);
nor U4607 (N_4607,N_4364,N_4400);
nand U4608 (N_4608,N_4453,N_4480);
or U4609 (N_4609,N_4490,N_4499);
or U4610 (N_4610,N_4406,N_4481);
and U4611 (N_4611,N_4364,N_4447);
or U4612 (N_4612,N_4457,N_4481);
nor U4613 (N_4613,N_4477,N_4362);
nor U4614 (N_4614,N_4425,N_4361);
xnor U4615 (N_4615,N_4393,N_4397);
nor U4616 (N_4616,N_4439,N_4486);
xor U4617 (N_4617,N_4391,N_4484);
nand U4618 (N_4618,N_4477,N_4370);
or U4619 (N_4619,N_4471,N_4366);
nor U4620 (N_4620,N_4472,N_4416);
xnor U4621 (N_4621,N_4366,N_4463);
and U4622 (N_4622,N_4369,N_4376);
nand U4623 (N_4623,N_4467,N_4458);
and U4624 (N_4624,N_4424,N_4390);
nand U4625 (N_4625,N_4388,N_4393);
nand U4626 (N_4626,N_4363,N_4366);
nor U4627 (N_4627,N_4498,N_4464);
xor U4628 (N_4628,N_4409,N_4377);
nand U4629 (N_4629,N_4457,N_4449);
xnor U4630 (N_4630,N_4416,N_4471);
xor U4631 (N_4631,N_4440,N_4452);
nor U4632 (N_4632,N_4474,N_4360);
xnor U4633 (N_4633,N_4491,N_4404);
xor U4634 (N_4634,N_4484,N_4480);
or U4635 (N_4635,N_4475,N_4487);
xnor U4636 (N_4636,N_4395,N_4424);
and U4637 (N_4637,N_4418,N_4483);
nand U4638 (N_4638,N_4416,N_4391);
nor U4639 (N_4639,N_4360,N_4450);
xnor U4640 (N_4640,N_4464,N_4459);
xor U4641 (N_4641,N_4408,N_4456);
nand U4642 (N_4642,N_4415,N_4401);
nand U4643 (N_4643,N_4361,N_4499);
nand U4644 (N_4644,N_4413,N_4427);
or U4645 (N_4645,N_4498,N_4405);
xor U4646 (N_4646,N_4358,N_4456);
nand U4647 (N_4647,N_4387,N_4396);
xnor U4648 (N_4648,N_4458,N_4406);
xnor U4649 (N_4649,N_4479,N_4356);
nor U4650 (N_4650,N_4578,N_4569);
nand U4651 (N_4651,N_4614,N_4504);
xnor U4652 (N_4652,N_4630,N_4620);
or U4653 (N_4653,N_4519,N_4585);
and U4654 (N_4654,N_4598,N_4517);
and U4655 (N_4655,N_4548,N_4524);
or U4656 (N_4656,N_4514,N_4576);
xor U4657 (N_4657,N_4538,N_4512);
xor U4658 (N_4658,N_4570,N_4513);
or U4659 (N_4659,N_4619,N_4587);
and U4660 (N_4660,N_4539,N_4574);
nor U4661 (N_4661,N_4594,N_4520);
or U4662 (N_4662,N_4638,N_4528);
nor U4663 (N_4663,N_4532,N_4625);
or U4664 (N_4664,N_4612,N_4617);
or U4665 (N_4665,N_4613,N_4571);
or U4666 (N_4666,N_4525,N_4597);
xnor U4667 (N_4667,N_4611,N_4502);
nor U4668 (N_4668,N_4564,N_4503);
or U4669 (N_4669,N_4534,N_4561);
or U4670 (N_4670,N_4508,N_4608);
or U4671 (N_4671,N_4515,N_4631);
or U4672 (N_4672,N_4510,N_4544);
nor U4673 (N_4673,N_4545,N_4639);
nand U4674 (N_4674,N_4605,N_4560);
nor U4675 (N_4675,N_4540,N_4500);
xnor U4676 (N_4676,N_4599,N_4579);
nand U4677 (N_4677,N_4588,N_4527);
or U4678 (N_4678,N_4553,N_4629);
nand U4679 (N_4679,N_4600,N_4603);
nand U4680 (N_4680,N_4550,N_4501);
and U4681 (N_4681,N_4535,N_4645);
or U4682 (N_4682,N_4511,N_4556);
or U4683 (N_4683,N_4648,N_4521);
xor U4684 (N_4684,N_4559,N_4552);
and U4685 (N_4685,N_4529,N_4551);
nor U4686 (N_4686,N_4547,N_4644);
xnor U4687 (N_4687,N_4546,N_4640);
nand U4688 (N_4688,N_4628,N_4622);
nor U4689 (N_4689,N_4568,N_4609);
nor U4690 (N_4690,N_4506,N_4643);
and U4691 (N_4691,N_4649,N_4582);
nand U4692 (N_4692,N_4526,N_4610);
xnor U4693 (N_4693,N_4566,N_4567);
and U4694 (N_4694,N_4618,N_4621);
nand U4695 (N_4695,N_4616,N_4575);
nand U4696 (N_4696,N_4607,N_4615);
or U4697 (N_4697,N_4531,N_4536);
nor U4698 (N_4698,N_4522,N_4509);
nor U4699 (N_4699,N_4518,N_4516);
and U4700 (N_4700,N_4633,N_4601);
or U4701 (N_4701,N_4634,N_4543);
nor U4702 (N_4702,N_4592,N_4623);
or U4703 (N_4703,N_4573,N_4557);
xor U4704 (N_4704,N_4646,N_4589);
or U4705 (N_4705,N_4523,N_4596);
nand U4706 (N_4706,N_4505,N_4586);
or U4707 (N_4707,N_4635,N_4604);
nand U4708 (N_4708,N_4606,N_4580);
or U4709 (N_4709,N_4602,N_4590);
and U4710 (N_4710,N_4637,N_4541);
or U4711 (N_4711,N_4647,N_4572);
or U4712 (N_4712,N_4537,N_4642);
or U4713 (N_4713,N_4549,N_4584);
nor U4714 (N_4714,N_4577,N_4530);
nor U4715 (N_4715,N_4565,N_4641);
xor U4716 (N_4716,N_4593,N_4581);
nor U4717 (N_4717,N_4533,N_4542);
nor U4718 (N_4718,N_4624,N_4632);
or U4719 (N_4719,N_4627,N_4583);
nor U4720 (N_4720,N_4626,N_4636);
and U4721 (N_4721,N_4555,N_4507);
xor U4722 (N_4722,N_4591,N_4554);
and U4723 (N_4723,N_4562,N_4558);
nand U4724 (N_4724,N_4595,N_4563);
and U4725 (N_4725,N_4535,N_4611);
and U4726 (N_4726,N_4547,N_4586);
or U4727 (N_4727,N_4535,N_4609);
nand U4728 (N_4728,N_4614,N_4585);
and U4729 (N_4729,N_4619,N_4584);
nor U4730 (N_4730,N_4504,N_4618);
and U4731 (N_4731,N_4623,N_4572);
or U4732 (N_4732,N_4524,N_4578);
and U4733 (N_4733,N_4603,N_4532);
xor U4734 (N_4734,N_4506,N_4515);
nor U4735 (N_4735,N_4546,N_4600);
and U4736 (N_4736,N_4612,N_4647);
nand U4737 (N_4737,N_4593,N_4523);
nand U4738 (N_4738,N_4548,N_4628);
xnor U4739 (N_4739,N_4551,N_4619);
or U4740 (N_4740,N_4587,N_4596);
nor U4741 (N_4741,N_4636,N_4535);
or U4742 (N_4742,N_4584,N_4573);
and U4743 (N_4743,N_4639,N_4546);
or U4744 (N_4744,N_4641,N_4515);
xnor U4745 (N_4745,N_4523,N_4501);
nor U4746 (N_4746,N_4513,N_4603);
or U4747 (N_4747,N_4614,N_4558);
or U4748 (N_4748,N_4578,N_4625);
nand U4749 (N_4749,N_4556,N_4522);
nand U4750 (N_4750,N_4600,N_4620);
or U4751 (N_4751,N_4609,N_4580);
or U4752 (N_4752,N_4597,N_4590);
or U4753 (N_4753,N_4549,N_4513);
or U4754 (N_4754,N_4605,N_4594);
xnor U4755 (N_4755,N_4608,N_4610);
and U4756 (N_4756,N_4556,N_4519);
or U4757 (N_4757,N_4644,N_4506);
xnor U4758 (N_4758,N_4648,N_4528);
or U4759 (N_4759,N_4618,N_4570);
and U4760 (N_4760,N_4571,N_4601);
or U4761 (N_4761,N_4564,N_4571);
and U4762 (N_4762,N_4554,N_4542);
nor U4763 (N_4763,N_4519,N_4573);
or U4764 (N_4764,N_4511,N_4526);
nor U4765 (N_4765,N_4642,N_4584);
xor U4766 (N_4766,N_4527,N_4600);
or U4767 (N_4767,N_4649,N_4597);
nand U4768 (N_4768,N_4599,N_4501);
or U4769 (N_4769,N_4631,N_4527);
nand U4770 (N_4770,N_4516,N_4584);
or U4771 (N_4771,N_4612,N_4591);
xor U4772 (N_4772,N_4628,N_4551);
nand U4773 (N_4773,N_4555,N_4580);
or U4774 (N_4774,N_4639,N_4631);
or U4775 (N_4775,N_4590,N_4558);
nand U4776 (N_4776,N_4623,N_4585);
nand U4777 (N_4777,N_4637,N_4514);
and U4778 (N_4778,N_4550,N_4609);
nand U4779 (N_4779,N_4505,N_4530);
and U4780 (N_4780,N_4505,N_4637);
and U4781 (N_4781,N_4501,N_4593);
nand U4782 (N_4782,N_4606,N_4592);
nand U4783 (N_4783,N_4612,N_4649);
nand U4784 (N_4784,N_4541,N_4564);
nand U4785 (N_4785,N_4539,N_4648);
and U4786 (N_4786,N_4587,N_4581);
or U4787 (N_4787,N_4504,N_4564);
xnor U4788 (N_4788,N_4599,N_4536);
nand U4789 (N_4789,N_4594,N_4607);
xnor U4790 (N_4790,N_4603,N_4568);
or U4791 (N_4791,N_4598,N_4648);
nor U4792 (N_4792,N_4530,N_4555);
xor U4793 (N_4793,N_4641,N_4618);
xnor U4794 (N_4794,N_4628,N_4507);
xor U4795 (N_4795,N_4643,N_4630);
nand U4796 (N_4796,N_4539,N_4640);
nand U4797 (N_4797,N_4528,N_4639);
nor U4798 (N_4798,N_4539,N_4556);
and U4799 (N_4799,N_4642,N_4626);
or U4800 (N_4800,N_4797,N_4715);
nand U4801 (N_4801,N_4663,N_4710);
or U4802 (N_4802,N_4745,N_4757);
xor U4803 (N_4803,N_4732,N_4682);
nand U4804 (N_4804,N_4792,N_4665);
or U4805 (N_4805,N_4719,N_4695);
and U4806 (N_4806,N_4703,N_4664);
or U4807 (N_4807,N_4752,N_4786);
nor U4808 (N_4808,N_4736,N_4662);
nand U4809 (N_4809,N_4699,N_4653);
nand U4810 (N_4810,N_4650,N_4658);
nor U4811 (N_4811,N_4668,N_4731);
nor U4812 (N_4812,N_4756,N_4796);
nor U4813 (N_4813,N_4783,N_4689);
xor U4814 (N_4814,N_4744,N_4739);
xnor U4815 (N_4815,N_4669,N_4680);
nand U4816 (N_4816,N_4696,N_4656);
nand U4817 (N_4817,N_4743,N_4694);
or U4818 (N_4818,N_4780,N_4782);
and U4819 (N_4819,N_4759,N_4708);
xnor U4820 (N_4820,N_4767,N_4730);
xnor U4821 (N_4821,N_4725,N_4654);
nor U4822 (N_4822,N_4749,N_4765);
xnor U4823 (N_4823,N_4798,N_4709);
xnor U4824 (N_4824,N_4762,N_4723);
and U4825 (N_4825,N_4671,N_4761);
and U4826 (N_4826,N_4779,N_4661);
nand U4827 (N_4827,N_4758,N_4793);
nor U4828 (N_4828,N_4746,N_4660);
nor U4829 (N_4829,N_4673,N_4707);
xnor U4830 (N_4830,N_4712,N_4705);
nand U4831 (N_4831,N_4713,N_4681);
and U4832 (N_4832,N_4716,N_4706);
and U4833 (N_4833,N_4733,N_4776);
xnor U4834 (N_4834,N_4720,N_4691);
nand U4835 (N_4835,N_4678,N_4679);
and U4836 (N_4836,N_4795,N_4741);
or U4837 (N_4837,N_4772,N_4675);
nor U4838 (N_4838,N_4688,N_4676);
xnor U4839 (N_4839,N_4714,N_4687);
or U4840 (N_4840,N_4750,N_4734);
xnor U4841 (N_4841,N_4726,N_4657);
nor U4842 (N_4842,N_4701,N_4789);
xor U4843 (N_4843,N_4718,N_4727);
or U4844 (N_4844,N_4685,N_4677);
xnor U4845 (N_4845,N_4700,N_4670);
xor U4846 (N_4846,N_4771,N_4799);
or U4847 (N_4847,N_4740,N_4704);
xnor U4848 (N_4848,N_4770,N_4785);
or U4849 (N_4849,N_4652,N_4764);
or U4850 (N_4850,N_4692,N_4672);
xor U4851 (N_4851,N_4753,N_4755);
xor U4852 (N_4852,N_4735,N_4717);
and U4853 (N_4853,N_4683,N_4666);
xnor U4854 (N_4854,N_4674,N_4777);
xnor U4855 (N_4855,N_4768,N_4698);
nand U4856 (N_4856,N_4737,N_4791);
nand U4857 (N_4857,N_4781,N_4787);
or U4858 (N_4858,N_4655,N_4697);
or U4859 (N_4859,N_4693,N_4686);
and U4860 (N_4860,N_4775,N_4769);
xor U4861 (N_4861,N_4760,N_4738);
and U4862 (N_4862,N_4651,N_4721);
nand U4863 (N_4863,N_4748,N_4724);
xnor U4864 (N_4864,N_4763,N_4722);
and U4865 (N_4865,N_4711,N_4729);
nor U4866 (N_4866,N_4728,N_4788);
or U4867 (N_4867,N_4684,N_4667);
or U4868 (N_4868,N_4742,N_4690);
and U4869 (N_4869,N_4773,N_4702);
or U4870 (N_4870,N_4659,N_4794);
nand U4871 (N_4871,N_4778,N_4747);
or U4872 (N_4872,N_4751,N_4790);
or U4873 (N_4873,N_4766,N_4774);
xor U4874 (N_4874,N_4754,N_4784);
xor U4875 (N_4875,N_4722,N_4785);
or U4876 (N_4876,N_4681,N_4770);
xor U4877 (N_4877,N_4712,N_4741);
or U4878 (N_4878,N_4784,N_4658);
or U4879 (N_4879,N_4778,N_4736);
or U4880 (N_4880,N_4659,N_4756);
xnor U4881 (N_4881,N_4668,N_4782);
and U4882 (N_4882,N_4765,N_4769);
nor U4883 (N_4883,N_4675,N_4751);
xor U4884 (N_4884,N_4782,N_4698);
xor U4885 (N_4885,N_4673,N_4659);
xnor U4886 (N_4886,N_4676,N_4726);
and U4887 (N_4887,N_4694,N_4720);
nand U4888 (N_4888,N_4774,N_4735);
or U4889 (N_4889,N_4777,N_4798);
nor U4890 (N_4890,N_4772,N_4733);
xor U4891 (N_4891,N_4756,N_4729);
nor U4892 (N_4892,N_4704,N_4746);
or U4893 (N_4893,N_4790,N_4715);
nand U4894 (N_4894,N_4671,N_4697);
and U4895 (N_4895,N_4671,N_4692);
nand U4896 (N_4896,N_4798,N_4702);
nand U4897 (N_4897,N_4729,N_4793);
or U4898 (N_4898,N_4713,N_4787);
and U4899 (N_4899,N_4787,N_4679);
xor U4900 (N_4900,N_4722,N_4748);
or U4901 (N_4901,N_4714,N_4701);
and U4902 (N_4902,N_4722,N_4703);
xnor U4903 (N_4903,N_4793,N_4696);
and U4904 (N_4904,N_4774,N_4730);
and U4905 (N_4905,N_4683,N_4792);
and U4906 (N_4906,N_4772,N_4652);
xor U4907 (N_4907,N_4675,N_4735);
nor U4908 (N_4908,N_4665,N_4730);
and U4909 (N_4909,N_4688,N_4651);
nor U4910 (N_4910,N_4716,N_4702);
or U4911 (N_4911,N_4778,N_4675);
or U4912 (N_4912,N_4675,N_4719);
nor U4913 (N_4913,N_4723,N_4703);
and U4914 (N_4914,N_4764,N_4659);
or U4915 (N_4915,N_4754,N_4796);
nor U4916 (N_4916,N_4734,N_4688);
and U4917 (N_4917,N_4656,N_4679);
nand U4918 (N_4918,N_4755,N_4793);
xnor U4919 (N_4919,N_4766,N_4740);
and U4920 (N_4920,N_4719,N_4714);
xor U4921 (N_4921,N_4678,N_4756);
nand U4922 (N_4922,N_4731,N_4650);
nand U4923 (N_4923,N_4794,N_4708);
nor U4924 (N_4924,N_4792,N_4697);
or U4925 (N_4925,N_4753,N_4776);
nor U4926 (N_4926,N_4786,N_4676);
and U4927 (N_4927,N_4659,N_4654);
nand U4928 (N_4928,N_4655,N_4761);
nor U4929 (N_4929,N_4679,N_4788);
and U4930 (N_4930,N_4677,N_4652);
nand U4931 (N_4931,N_4671,N_4652);
and U4932 (N_4932,N_4794,N_4715);
nor U4933 (N_4933,N_4799,N_4651);
nand U4934 (N_4934,N_4708,N_4689);
and U4935 (N_4935,N_4730,N_4707);
or U4936 (N_4936,N_4702,N_4772);
nor U4937 (N_4937,N_4759,N_4740);
and U4938 (N_4938,N_4680,N_4715);
or U4939 (N_4939,N_4693,N_4799);
xor U4940 (N_4940,N_4770,N_4771);
or U4941 (N_4941,N_4742,N_4716);
or U4942 (N_4942,N_4666,N_4662);
or U4943 (N_4943,N_4717,N_4779);
and U4944 (N_4944,N_4760,N_4708);
nor U4945 (N_4945,N_4661,N_4732);
nor U4946 (N_4946,N_4701,N_4685);
nand U4947 (N_4947,N_4798,N_4706);
xnor U4948 (N_4948,N_4722,N_4670);
nand U4949 (N_4949,N_4719,N_4750);
nor U4950 (N_4950,N_4882,N_4808);
xnor U4951 (N_4951,N_4849,N_4875);
xor U4952 (N_4952,N_4909,N_4802);
xnor U4953 (N_4953,N_4830,N_4861);
nor U4954 (N_4954,N_4879,N_4869);
nor U4955 (N_4955,N_4844,N_4938);
and U4956 (N_4956,N_4835,N_4846);
xnor U4957 (N_4957,N_4922,N_4949);
nand U4958 (N_4958,N_4945,N_4921);
nand U4959 (N_4959,N_4890,N_4944);
and U4960 (N_4960,N_4824,N_4812);
and U4961 (N_4961,N_4816,N_4943);
and U4962 (N_4962,N_4877,N_4946);
xor U4963 (N_4963,N_4941,N_4857);
xnor U4964 (N_4964,N_4819,N_4845);
xor U4965 (N_4965,N_4817,N_4923);
or U4966 (N_4966,N_4896,N_4929);
nor U4967 (N_4967,N_4833,N_4881);
nor U4968 (N_4968,N_4806,N_4820);
nand U4969 (N_4969,N_4935,N_4892);
or U4970 (N_4970,N_4856,N_4828);
nor U4971 (N_4971,N_4918,N_4880);
and U4972 (N_4972,N_4851,N_4889);
xor U4973 (N_4973,N_4810,N_4910);
xnor U4974 (N_4974,N_4897,N_4899);
xnor U4975 (N_4975,N_4940,N_4873);
or U4976 (N_4976,N_4859,N_4904);
or U4977 (N_4977,N_4840,N_4903);
xor U4978 (N_4978,N_4804,N_4927);
xnor U4979 (N_4979,N_4908,N_4843);
xor U4980 (N_4980,N_4866,N_4936);
or U4981 (N_4981,N_4809,N_4807);
nor U4982 (N_4982,N_4905,N_4919);
xnor U4983 (N_4983,N_4831,N_4838);
and U4984 (N_4984,N_4860,N_4818);
nor U4985 (N_4985,N_4811,N_4834);
xor U4986 (N_4986,N_4884,N_4878);
xor U4987 (N_4987,N_4850,N_4822);
or U4988 (N_4988,N_4823,N_4914);
and U4989 (N_4989,N_4931,N_4867);
and U4990 (N_4990,N_4911,N_4948);
nor U4991 (N_4991,N_4815,N_4915);
or U4992 (N_4992,N_4900,N_4864);
nor U4993 (N_4993,N_4803,N_4805);
or U4994 (N_4994,N_4893,N_4853);
xnor U4995 (N_4995,N_4801,N_4891);
xor U4996 (N_4996,N_4836,N_4847);
nand U4997 (N_4997,N_4932,N_4855);
and U4998 (N_4998,N_4895,N_4876);
or U4999 (N_4999,N_4930,N_4800);
xnor U5000 (N_5000,N_4924,N_4814);
or U5001 (N_5001,N_4813,N_4858);
or U5002 (N_5002,N_4874,N_4829);
xor U5003 (N_5003,N_4939,N_4942);
and U5004 (N_5004,N_4862,N_4934);
and U5005 (N_5005,N_4871,N_4826);
nor U5006 (N_5006,N_4865,N_4821);
nor U5007 (N_5007,N_4870,N_4933);
or U5008 (N_5008,N_4898,N_4827);
or U5009 (N_5009,N_4868,N_4848);
nor U5010 (N_5010,N_4885,N_4907);
xor U5011 (N_5011,N_4906,N_4852);
or U5012 (N_5012,N_4894,N_4917);
or U5013 (N_5013,N_4925,N_4872);
nor U5014 (N_5014,N_4928,N_4863);
nand U5015 (N_5015,N_4842,N_4886);
nand U5016 (N_5016,N_4901,N_4920);
nand U5017 (N_5017,N_4912,N_4837);
xor U5018 (N_5018,N_4888,N_4916);
nand U5019 (N_5019,N_4902,N_4887);
nand U5020 (N_5020,N_4883,N_4825);
xor U5021 (N_5021,N_4841,N_4937);
and U5022 (N_5022,N_4839,N_4947);
xnor U5023 (N_5023,N_4913,N_4926);
nand U5024 (N_5024,N_4832,N_4854);
or U5025 (N_5025,N_4801,N_4941);
nand U5026 (N_5026,N_4925,N_4896);
nor U5027 (N_5027,N_4887,N_4856);
nor U5028 (N_5028,N_4808,N_4809);
or U5029 (N_5029,N_4853,N_4918);
nor U5030 (N_5030,N_4882,N_4835);
nand U5031 (N_5031,N_4915,N_4937);
or U5032 (N_5032,N_4913,N_4811);
nand U5033 (N_5033,N_4832,N_4891);
and U5034 (N_5034,N_4857,N_4864);
or U5035 (N_5035,N_4909,N_4817);
xor U5036 (N_5036,N_4875,N_4845);
and U5037 (N_5037,N_4874,N_4898);
and U5038 (N_5038,N_4826,N_4869);
nor U5039 (N_5039,N_4920,N_4867);
nor U5040 (N_5040,N_4947,N_4891);
and U5041 (N_5041,N_4804,N_4912);
nand U5042 (N_5042,N_4840,N_4910);
and U5043 (N_5043,N_4944,N_4896);
xor U5044 (N_5044,N_4867,N_4904);
nand U5045 (N_5045,N_4874,N_4909);
nand U5046 (N_5046,N_4817,N_4818);
or U5047 (N_5047,N_4939,N_4872);
or U5048 (N_5048,N_4940,N_4862);
or U5049 (N_5049,N_4893,N_4921);
or U5050 (N_5050,N_4914,N_4893);
xor U5051 (N_5051,N_4859,N_4926);
or U5052 (N_5052,N_4803,N_4838);
xnor U5053 (N_5053,N_4843,N_4841);
and U5054 (N_5054,N_4882,N_4933);
nor U5055 (N_5055,N_4857,N_4899);
or U5056 (N_5056,N_4884,N_4862);
nor U5057 (N_5057,N_4832,N_4886);
and U5058 (N_5058,N_4902,N_4949);
nand U5059 (N_5059,N_4880,N_4874);
nor U5060 (N_5060,N_4880,N_4855);
nor U5061 (N_5061,N_4927,N_4863);
nand U5062 (N_5062,N_4887,N_4823);
and U5063 (N_5063,N_4813,N_4864);
nor U5064 (N_5064,N_4857,N_4845);
and U5065 (N_5065,N_4921,N_4838);
xnor U5066 (N_5066,N_4845,N_4904);
nor U5067 (N_5067,N_4866,N_4830);
nand U5068 (N_5068,N_4899,N_4910);
nand U5069 (N_5069,N_4886,N_4884);
nor U5070 (N_5070,N_4817,N_4821);
nor U5071 (N_5071,N_4856,N_4816);
nand U5072 (N_5072,N_4806,N_4883);
xnor U5073 (N_5073,N_4832,N_4918);
xnor U5074 (N_5074,N_4805,N_4905);
xnor U5075 (N_5075,N_4893,N_4877);
or U5076 (N_5076,N_4810,N_4890);
nor U5077 (N_5077,N_4833,N_4883);
or U5078 (N_5078,N_4895,N_4837);
xnor U5079 (N_5079,N_4910,N_4916);
xnor U5080 (N_5080,N_4913,N_4863);
nor U5081 (N_5081,N_4934,N_4864);
nor U5082 (N_5082,N_4876,N_4848);
nand U5083 (N_5083,N_4869,N_4926);
nor U5084 (N_5084,N_4900,N_4851);
xnor U5085 (N_5085,N_4861,N_4887);
or U5086 (N_5086,N_4931,N_4808);
xnor U5087 (N_5087,N_4805,N_4906);
xor U5088 (N_5088,N_4907,N_4902);
xnor U5089 (N_5089,N_4885,N_4890);
nand U5090 (N_5090,N_4825,N_4891);
xnor U5091 (N_5091,N_4861,N_4913);
and U5092 (N_5092,N_4849,N_4927);
and U5093 (N_5093,N_4850,N_4892);
or U5094 (N_5094,N_4941,N_4815);
nand U5095 (N_5095,N_4938,N_4890);
or U5096 (N_5096,N_4949,N_4905);
nand U5097 (N_5097,N_4810,N_4863);
nor U5098 (N_5098,N_4825,N_4923);
and U5099 (N_5099,N_4900,N_4930);
xnor U5100 (N_5100,N_5008,N_4954);
and U5101 (N_5101,N_5019,N_5044);
nand U5102 (N_5102,N_5042,N_5028);
or U5103 (N_5103,N_4971,N_5065);
nand U5104 (N_5104,N_5041,N_5046);
nor U5105 (N_5105,N_5062,N_5024);
or U5106 (N_5106,N_5078,N_5029);
nor U5107 (N_5107,N_5098,N_5088);
nand U5108 (N_5108,N_4976,N_4950);
or U5109 (N_5109,N_4983,N_4998);
xor U5110 (N_5110,N_4958,N_4952);
nor U5111 (N_5111,N_5031,N_5045);
and U5112 (N_5112,N_5059,N_5094);
nand U5113 (N_5113,N_4977,N_5081);
xnor U5114 (N_5114,N_4988,N_4984);
xnor U5115 (N_5115,N_5055,N_4974);
xor U5116 (N_5116,N_4996,N_5010);
xor U5117 (N_5117,N_5034,N_5097);
or U5118 (N_5118,N_5001,N_5083);
or U5119 (N_5119,N_5014,N_5035);
or U5120 (N_5120,N_5032,N_5086);
and U5121 (N_5121,N_4969,N_5057);
and U5122 (N_5122,N_5043,N_5068);
and U5123 (N_5123,N_4961,N_5033);
nand U5124 (N_5124,N_5089,N_5037);
or U5125 (N_5125,N_5016,N_5072);
xor U5126 (N_5126,N_5036,N_5079);
nor U5127 (N_5127,N_5069,N_5002);
xnor U5128 (N_5128,N_5077,N_5027);
or U5129 (N_5129,N_4972,N_5020);
nand U5130 (N_5130,N_4989,N_4981);
or U5131 (N_5131,N_5054,N_5006);
nand U5132 (N_5132,N_4956,N_5026);
and U5133 (N_5133,N_5073,N_5013);
xnor U5134 (N_5134,N_5048,N_5018);
xor U5135 (N_5135,N_4960,N_4999);
nor U5136 (N_5136,N_5052,N_4962);
xor U5137 (N_5137,N_4966,N_5056);
or U5138 (N_5138,N_5047,N_4995);
xnor U5139 (N_5139,N_5095,N_5003);
nand U5140 (N_5140,N_4991,N_5000);
nor U5141 (N_5141,N_5096,N_5093);
and U5142 (N_5142,N_5017,N_5050);
nand U5143 (N_5143,N_5009,N_4993);
or U5144 (N_5144,N_4985,N_5012);
nor U5145 (N_5145,N_5007,N_4963);
and U5146 (N_5146,N_5066,N_4994);
nor U5147 (N_5147,N_5053,N_5030);
xor U5148 (N_5148,N_5011,N_4953);
or U5149 (N_5149,N_5076,N_5061);
xnor U5150 (N_5150,N_5085,N_4982);
xnor U5151 (N_5151,N_4965,N_4987);
or U5152 (N_5152,N_4964,N_4979);
xnor U5153 (N_5153,N_5082,N_4986);
nor U5154 (N_5154,N_5005,N_4951);
nand U5155 (N_5155,N_5021,N_5075);
and U5156 (N_5156,N_5090,N_5051);
xor U5157 (N_5157,N_4968,N_5023);
or U5158 (N_5158,N_4957,N_5038);
or U5159 (N_5159,N_5087,N_5040);
nand U5160 (N_5160,N_5084,N_4992);
or U5161 (N_5161,N_5099,N_4973);
and U5162 (N_5162,N_5091,N_4975);
or U5163 (N_5163,N_5060,N_5049);
xor U5164 (N_5164,N_4980,N_5074);
and U5165 (N_5165,N_5080,N_5004);
or U5166 (N_5166,N_5067,N_5071);
or U5167 (N_5167,N_5092,N_4970);
nand U5168 (N_5168,N_4990,N_5015);
nand U5169 (N_5169,N_4978,N_5070);
nand U5170 (N_5170,N_5025,N_5039);
nand U5171 (N_5171,N_4959,N_5058);
xor U5172 (N_5172,N_5063,N_4955);
and U5173 (N_5173,N_5022,N_5064);
nor U5174 (N_5174,N_4967,N_4997);
nor U5175 (N_5175,N_5000,N_5042);
or U5176 (N_5176,N_5016,N_5007);
xor U5177 (N_5177,N_4969,N_5072);
xor U5178 (N_5178,N_5053,N_4993);
nor U5179 (N_5179,N_5030,N_5027);
and U5180 (N_5180,N_4969,N_4974);
nor U5181 (N_5181,N_5054,N_4963);
nand U5182 (N_5182,N_5044,N_4968);
or U5183 (N_5183,N_5074,N_5082);
and U5184 (N_5184,N_5047,N_5054);
xor U5185 (N_5185,N_5036,N_5049);
xnor U5186 (N_5186,N_4997,N_4982);
and U5187 (N_5187,N_4982,N_5031);
or U5188 (N_5188,N_5011,N_5059);
or U5189 (N_5189,N_5082,N_4978);
xnor U5190 (N_5190,N_5090,N_4983);
nand U5191 (N_5191,N_5087,N_4967);
xor U5192 (N_5192,N_5009,N_5022);
and U5193 (N_5193,N_5065,N_5084);
nand U5194 (N_5194,N_4972,N_4954);
and U5195 (N_5195,N_5063,N_5049);
or U5196 (N_5196,N_5074,N_5097);
or U5197 (N_5197,N_4959,N_4951);
nand U5198 (N_5198,N_5021,N_5082);
nor U5199 (N_5199,N_5045,N_4955);
and U5200 (N_5200,N_5025,N_4975);
nand U5201 (N_5201,N_5068,N_5058);
xor U5202 (N_5202,N_4975,N_5068);
xor U5203 (N_5203,N_5056,N_5025);
nor U5204 (N_5204,N_5027,N_4975);
xnor U5205 (N_5205,N_5073,N_5089);
xnor U5206 (N_5206,N_5023,N_4971);
nand U5207 (N_5207,N_4987,N_4971);
xor U5208 (N_5208,N_5025,N_5034);
and U5209 (N_5209,N_5018,N_5033);
nor U5210 (N_5210,N_4989,N_5027);
nand U5211 (N_5211,N_5012,N_5037);
xor U5212 (N_5212,N_5056,N_5089);
nor U5213 (N_5213,N_5056,N_5024);
and U5214 (N_5214,N_5055,N_5008);
or U5215 (N_5215,N_4995,N_5075);
or U5216 (N_5216,N_5025,N_5021);
and U5217 (N_5217,N_5055,N_4978);
xor U5218 (N_5218,N_5069,N_4991);
and U5219 (N_5219,N_5000,N_5098);
xor U5220 (N_5220,N_5029,N_5033);
nor U5221 (N_5221,N_5060,N_5036);
and U5222 (N_5222,N_5023,N_5082);
nand U5223 (N_5223,N_5048,N_4972);
xnor U5224 (N_5224,N_4996,N_4998);
or U5225 (N_5225,N_4956,N_5083);
or U5226 (N_5226,N_5036,N_5059);
xnor U5227 (N_5227,N_4958,N_4967);
and U5228 (N_5228,N_5091,N_5085);
or U5229 (N_5229,N_4971,N_5059);
nand U5230 (N_5230,N_4984,N_5019);
nor U5231 (N_5231,N_5087,N_5077);
xnor U5232 (N_5232,N_5069,N_5012);
and U5233 (N_5233,N_5071,N_4995);
or U5234 (N_5234,N_5042,N_5027);
nand U5235 (N_5235,N_5012,N_5028);
nor U5236 (N_5236,N_5022,N_5042);
xnor U5237 (N_5237,N_5030,N_5086);
nand U5238 (N_5238,N_4983,N_4971);
xnor U5239 (N_5239,N_5030,N_5000);
nand U5240 (N_5240,N_5000,N_5037);
xnor U5241 (N_5241,N_5091,N_4973);
xor U5242 (N_5242,N_5059,N_5018);
nor U5243 (N_5243,N_5046,N_5053);
and U5244 (N_5244,N_5074,N_5099);
nor U5245 (N_5245,N_5087,N_4995);
and U5246 (N_5246,N_4952,N_5052);
or U5247 (N_5247,N_5099,N_5044);
nor U5248 (N_5248,N_4989,N_4988);
or U5249 (N_5249,N_4994,N_5098);
nor U5250 (N_5250,N_5131,N_5235);
or U5251 (N_5251,N_5130,N_5248);
and U5252 (N_5252,N_5102,N_5236);
or U5253 (N_5253,N_5245,N_5241);
or U5254 (N_5254,N_5157,N_5113);
or U5255 (N_5255,N_5233,N_5192);
nor U5256 (N_5256,N_5112,N_5207);
nor U5257 (N_5257,N_5204,N_5211);
or U5258 (N_5258,N_5119,N_5159);
nand U5259 (N_5259,N_5124,N_5189);
nor U5260 (N_5260,N_5190,N_5132);
nand U5261 (N_5261,N_5203,N_5155);
xnor U5262 (N_5262,N_5120,N_5225);
xor U5263 (N_5263,N_5175,N_5101);
nand U5264 (N_5264,N_5185,N_5135);
nand U5265 (N_5265,N_5249,N_5178);
nand U5266 (N_5266,N_5221,N_5141);
nand U5267 (N_5267,N_5126,N_5147);
nor U5268 (N_5268,N_5195,N_5144);
xnor U5269 (N_5269,N_5109,N_5143);
nor U5270 (N_5270,N_5186,N_5129);
xnor U5271 (N_5271,N_5172,N_5156);
nor U5272 (N_5272,N_5164,N_5152);
or U5273 (N_5273,N_5244,N_5219);
nand U5274 (N_5274,N_5179,N_5217);
nand U5275 (N_5275,N_5138,N_5163);
or U5276 (N_5276,N_5196,N_5121);
or U5277 (N_5277,N_5194,N_5208);
nand U5278 (N_5278,N_5148,N_5160);
xor U5279 (N_5279,N_5213,N_5134);
nor U5280 (N_5280,N_5218,N_5215);
nor U5281 (N_5281,N_5223,N_5122);
or U5282 (N_5282,N_5238,N_5107);
and U5283 (N_5283,N_5154,N_5222);
nand U5284 (N_5284,N_5182,N_5198);
or U5285 (N_5285,N_5242,N_5111);
nand U5286 (N_5286,N_5193,N_5116);
or U5287 (N_5287,N_5243,N_5180);
nand U5288 (N_5288,N_5158,N_5184);
xor U5289 (N_5289,N_5240,N_5214);
nor U5290 (N_5290,N_5128,N_5183);
xor U5291 (N_5291,N_5165,N_5200);
xnor U5292 (N_5292,N_5133,N_5103);
and U5293 (N_5293,N_5229,N_5212);
nand U5294 (N_5294,N_5171,N_5227);
nand U5295 (N_5295,N_5210,N_5123);
nand U5296 (N_5296,N_5216,N_5118);
nor U5297 (N_5297,N_5205,N_5191);
nand U5298 (N_5298,N_5127,N_5246);
xor U5299 (N_5299,N_5177,N_5199);
and U5300 (N_5300,N_5106,N_5140);
and U5301 (N_5301,N_5170,N_5150);
and U5302 (N_5302,N_5104,N_5187);
nand U5303 (N_5303,N_5149,N_5176);
xor U5304 (N_5304,N_5188,N_5226);
or U5305 (N_5305,N_5239,N_5168);
nor U5306 (N_5306,N_5174,N_5197);
and U5307 (N_5307,N_5202,N_5224);
xor U5308 (N_5308,N_5247,N_5105);
xor U5309 (N_5309,N_5181,N_5145);
xnor U5310 (N_5310,N_5115,N_5146);
or U5311 (N_5311,N_5231,N_5206);
or U5312 (N_5312,N_5167,N_5234);
or U5313 (N_5313,N_5220,N_5137);
nand U5314 (N_5314,N_5139,N_5169);
xnor U5315 (N_5315,N_5110,N_5100);
xnor U5316 (N_5316,N_5209,N_5142);
or U5317 (N_5317,N_5162,N_5114);
and U5318 (N_5318,N_5228,N_5125);
and U5319 (N_5319,N_5161,N_5108);
xnor U5320 (N_5320,N_5151,N_5166);
nor U5321 (N_5321,N_5136,N_5201);
nor U5322 (N_5322,N_5153,N_5230);
nand U5323 (N_5323,N_5173,N_5232);
nor U5324 (N_5324,N_5237,N_5117);
nor U5325 (N_5325,N_5189,N_5207);
xnor U5326 (N_5326,N_5117,N_5114);
and U5327 (N_5327,N_5234,N_5222);
or U5328 (N_5328,N_5183,N_5205);
and U5329 (N_5329,N_5189,N_5143);
or U5330 (N_5330,N_5114,N_5213);
and U5331 (N_5331,N_5222,N_5127);
or U5332 (N_5332,N_5146,N_5242);
and U5333 (N_5333,N_5159,N_5237);
nor U5334 (N_5334,N_5113,N_5122);
or U5335 (N_5335,N_5201,N_5132);
and U5336 (N_5336,N_5246,N_5183);
xor U5337 (N_5337,N_5198,N_5233);
nor U5338 (N_5338,N_5187,N_5101);
nand U5339 (N_5339,N_5104,N_5182);
xor U5340 (N_5340,N_5120,N_5238);
and U5341 (N_5341,N_5238,N_5100);
and U5342 (N_5342,N_5232,N_5220);
or U5343 (N_5343,N_5222,N_5114);
and U5344 (N_5344,N_5114,N_5146);
xor U5345 (N_5345,N_5173,N_5128);
nor U5346 (N_5346,N_5244,N_5150);
xnor U5347 (N_5347,N_5206,N_5180);
nand U5348 (N_5348,N_5242,N_5186);
or U5349 (N_5349,N_5139,N_5108);
or U5350 (N_5350,N_5156,N_5166);
or U5351 (N_5351,N_5224,N_5146);
or U5352 (N_5352,N_5204,N_5180);
xnor U5353 (N_5353,N_5248,N_5104);
or U5354 (N_5354,N_5244,N_5140);
nor U5355 (N_5355,N_5127,N_5128);
and U5356 (N_5356,N_5152,N_5219);
xor U5357 (N_5357,N_5192,N_5242);
nor U5358 (N_5358,N_5182,N_5240);
and U5359 (N_5359,N_5147,N_5245);
nand U5360 (N_5360,N_5230,N_5112);
nand U5361 (N_5361,N_5111,N_5116);
nand U5362 (N_5362,N_5143,N_5172);
and U5363 (N_5363,N_5158,N_5247);
or U5364 (N_5364,N_5121,N_5148);
and U5365 (N_5365,N_5220,N_5116);
nand U5366 (N_5366,N_5249,N_5144);
or U5367 (N_5367,N_5241,N_5242);
and U5368 (N_5368,N_5180,N_5226);
and U5369 (N_5369,N_5235,N_5163);
nand U5370 (N_5370,N_5214,N_5129);
or U5371 (N_5371,N_5152,N_5246);
or U5372 (N_5372,N_5242,N_5239);
nor U5373 (N_5373,N_5188,N_5113);
and U5374 (N_5374,N_5141,N_5228);
nand U5375 (N_5375,N_5238,N_5196);
or U5376 (N_5376,N_5246,N_5124);
nor U5377 (N_5377,N_5117,N_5159);
xor U5378 (N_5378,N_5228,N_5226);
nor U5379 (N_5379,N_5123,N_5179);
xor U5380 (N_5380,N_5213,N_5233);
or U5381 (N_5381,N_5209,N_5222);
xor U5382 (N_5382,N_5131,N_5168);
xnor U5383 (N_5383,N_5172,N_5115);
xor U5384 (N_5384,N_5200,N_5194);
xor U5385 (N_5385,N_5195,N_5135);
xnor U5386 (N_5386,N_5156,N_5143);
and U5387 (N_5387,N_5107,N_5218);
nand U5388 (N_5388,N_5202,N_5148);
nor U5389 (N_5389,N_5216,N_5180);
nand U5390 (N_5390,N_5226,N_5136);
xor U5391 (N_5391,N_5130,N_5152);
nand U5392 (N_5392,N_5133,N_5223);
nand U5393 (N_5393,N_5246,N_5136);
or U5394 (N_5394,N_5181,N_5237);
nand U5395 (N_5395,N_5202,N_5167);
nand U5396 (N_5396,N_5237,N_5216);
xor U5397 (N_5397,N_5159,N_5158);
xor U5398 (N_5398,N_5211,N_5184);
and U5399 (N_5399,N_5123,N_5196);
xor U5400 (N_5400,N_5383,N_5256);
or U5401 (N_5401,N_5306,N_5265);
xnor U5402 (N_5402,N_5291,N_5390);
nor U5403 (N_5403,N_5375,N_5333);
or U5404 (N_5404,N_5299,N_5318);
or U5405 (N_5405,N_5281,N_5272);
nor U5406 (N_5406,N_5371,N_5374);
and U5407 (N_5407,N_5268,N_5297);
and U5408 (N_5408,N_5336,N_5398);
nand U5409 (N_5409,N_5385,N_5278);
and U5410 (N_5410,N_5293,N_5305);
nor U5411 (N_5411,N_5275,N_5391);
nand U5412 (N_5412,N_5253,N_5370);
or U5413 (N_5413,N_5289,N_5315);
nor U5414 (N_5414,N_5277,N_5252);
and U5415 (N_5415,N_5368,N_5324);
nor U5416 (N_5416,N_5396,N_5377);
xnor U5417 (N_5417,N_5307,N_5397);
nor U5418 (N_5418,N_5351,N_5271);
nor U5419 (N_5419,N_5261,N_5382);
and U5420 (N_5420,N_5355,N_5258);
nor U5421 (N_5421,N_5376,N_5316);
or U5422 (N_5422,N_5269,N_5326);
nor U5423 (N_5423,N_5266,N_5313);
and U5424 (N_5424,N_5274,N_5394);
or U5425 (N_5425,N_5262,N_5331);
nor U5426 (N_5426,N_5317,N_5386);
and U5427 (N_5427,N_5392,N_5300);
xnor U5428 (N_5428,N_5358,N_5367);
and U5429 (N_5429,N_5290,N_5310);
xnor U5430 (N_5430,N_5294,N_5314);
nand U5431 (N_5431,N_5288,N_5381);
xor U5432 (N_5432,N_5325,N_5276);
nand U5433 (N_5433,N_5321,N_5395);
xor U5434 (N_5434,N_5347,N_5279);
nand U5435 (N_5435,N_5399,N_5339);
xnor U5436 (N_5436,N_5360,N_5267);
nand U5437 (N_5437,N_5364,N_5337);
xor U5438 (N_5438,N_5263,N_5303);
nor U5439 (N_5439,N_5328,N_5349);
nand U5440 (N_5440,N_5250,N_5362);
and U5441 (N_5441,N_5257,N_5379);
nand U5442 (N_5442,N_5342,N_5330);
nand U5443 (N_5443,N_5283,N_5372);
nor U5444 (N_5444,N_5366,N_5359);
nor U5445 (N_5445,N_5319,N_5340);
nand U5446 (N_5446,N_5345,N_5344);
or U5447 (N_5447,N_5348,N_5387);
or U5448 (N_5448,N_5323,N_5311);
and U5449 (N_5449,N_5341,N_5329);
xnor U5450 (N_5450,N_5365,N_5363);
and U5451 (N_5451,N_5335,N_5302);
nand U5452 (N_5452,N_5361,N_5312);
nor U5453 (N_5453,N_5334,N_5284);
nor U5454 (N_5454,N_5389,N_5388);
or U5455 (N_5455,N_5254,N_5295);
nand U5456 (N_5456,N_5384,N_5343);
nand U5457 (N_5457,N_5327,N_5369);
xor U5458 (N_5458,N_5356,N_5292);
nand U5459 (N_5459,N_5282,N_5260);
and U5460 (N_5460,N_5346,N_5308);
nor U5461 (N_5461,N_5353,N_5380);
or U5462 (N_5462,N_5301,N_5350);
nand U5463 (N_5463,N_5304,N_5285);
nor U5464 (N_5464,N_5338,N_5251);
nor U5465 (N_5465,N_5332,N_5270);
xnor U5466 (N_5466,N_5273,N_5354);
or U5467 (N_5467,N_5255,N_5373);
xnor U5468 (N_5468,N_5298,N_5259);
nor U5469 (N_5469,N_5393,N_5357);
xnor U5470 (N_5470,N_5286,N_5280);
nand U5471 (N_5471,N_5378,N_5309);
nor U5472 (N_5472,N_5264,N_5296);
and U5473 (N_5473,N_5287,N_5322);
nand U5474 (N_5474,N_5352,N_5320);
or U5475 (N_5475,N_5388,N_5256);
nand U5476 (N_5476,N_5301,N_5340);
and U5477 (N_5477,N_5334,N_5341);
xnor U5478 (N_5478,N_5327,N_5340);
nor U5479 (N_5479,N_5263,N_5342);
or U5480 (N_5480,N_5386,N_5332);
or U5481 (N_5481,N_5312,N_5397);
nor U5482 (N_5482,N_5305,N_5258);
or U5483 (N_5483,N_5326,N_5392);
xor U5484 (N_5484,N_5327,N_5364);
xor U5485 (N_5485,N_5352,N_5323);
nor U5486 (N_5486,N_5264,N_5381);
nand U5487 (N_5487,N_5396,N_5268);
nand U5488 (N_5488,N_5341,N_5374);
or U5489 (N_5489,N_5394,N_5254);
xor U5490 (N_5490,N_5328,N_5290);
nand U5491 (N_5491,N_5370,N_5332);
nor U5492 (N_5492,N_5385,N_5260);
nand U5493 (N_5493,N_5392,N_5372);
and U5494 (N_5494,N_5347,N_5297);
nand U5495 (N_5495,N_5270,N_5268);
nand U5496 (N_5496,N_5381,N_5364);
and U5497 (N_5497,N_5288,N_5277);
nand U5498 (N_5498,N_5321,N_5317);
and U5499 (N_5499,N_5265,N_5365);
and U5500 (N_5500,N_5321,N_5296);
nor U5501 (N_5501,N_5296,N_5355);
nand U5502 (N_5502,N_5362,N_5351);
nor U5503 (N_5503,N_5345,N_5256);
nand U5504 (N_5504,N_5386,N_5352);
nand U5505 (N_5505,N_5396,N_5301);
or U5506 (N_5506,N_5324,N_5313);
and U5507 (N_5507,N_5250,N_5378);
nand U5508 (N_5508,N_5371,N_5292);
and U5509 (N_5509,N_5390,N_5387);
xnor U5510 (N_5510,N_5287,N_5388);
and U5511 (N_5511,N_5331,N_5324);
or U5512 (N_5512,N_5347,N_5373);
nand U5513 (N_5513,N_5336,N_5399);
xor U5514 (N_5514,N_5303,N_5304);
nand U5515 (N_5515,N_5366,N_5331);
or U5516 (N_5516,N_5342,N_5368);
and U5517 (N_5517,N_5385,N_5364);
or U5518 (N_5518,N_5356,N_5388);
nand U5519 (N_5519,N_5384,N_5256);
nor U5520 (N_5520,N_5329,N_5359);
nor U5521 (N_5521,N_5288,N_5301);
or U5522 (N_5522,N_5354,N_5318);
xnor U5523 (N_5523,N_5286,N_5391);
xnor U5524 (N_5524,N_5314,N_5361);
or U5525 (N_5525,N_5373,N_5289);
and U5526 (N_5526,N_5300,N_5325);
nand U5527 (N_5527,N_5272,N_5250);
and U5528 (N_5528,N_5304,N_5399);
nor U5529 (N_5529,N_5316,N_5295);
nand U5530 (N_5530,N_5281,N_5257);
nor U5531 (N_5531,N_5363,N_5324);
or U5532 (N_5532,N_5315,N_5381);
or U5533 (N_5533,N_5252,N_5347);
and U5534 (N_5534,N_5300,N_5391);
xor U5535 (N_5535,N_5258,N_5344);
and U5536 (N_5536,N_5285,N_5305);
nand U5537 (N_5537,N_5398,N_5353);
or U5538 (N_5538,N_5338,N_5299);
nor U5539 (N_5539,N_5275,N_5388);
and U5540 (N_5540,N_5284,N_5369);
xnor U5541 (N_5541,N_5263,N_5385);
or U5542 (N_5542,N_5287,N_5378);
nand U5543 (N_5543,N_5334,N_5346);
and U5544 (N_5544,N_5334,N_5365);
and U5545 (N_5545,N_5276,N_5278);
nor U5546 (N_5546,N_5264,N_5356);
xnor U5547 (N_5547,N_5332,N_5363);
xor U5548 (N_5548,N_5303,N_5393);
xnor U5549 (N_5549,N_5375,N_5346);
or U5550 (N_5550,N_5543,N_5441);
nand U5551 (N_5551,N_5407,N_5425);
xnor U5552 (N_5552,N_5502,N_5546);
nor U5553 (N_5553,N_5438,N_5405);
and U5554 (N_5554,N_5529,N_5413);
nor U5555 (N_5555,N_5533,N_5421);
and U5556 (N_5556,N_5445,N_5453);
nand U5557 (N_5557,N_5408,N_5536);
nor U5558 (N_5558,N_5459,N_5464);
nand U5559 (N_5559,N_5468,N_5479);
nor U5560 (N_5560,N_5481,N_5488);
nand U5561 (N_5561,N_5508,N_5507);
and U5562 (N_5562,N_5495,N_5420);
and U5563 (N_5563,N_5540,N_5548);
or U5564 (N_5564,N_5415,N_5527);
or U5565 (N_5565,N_5449,N_5513);
or U5566 (N_5566,N_5492,N_5443);
and U5567 (N_5567,N_5410,N_5418);
or U5568 (N_5568,N_5520,N_5444);
xnor U5569 (N_5569,N_5528,N_5439);
and U5570 (N_5570,N_5491,N_5432);
and U5571 (N_5571,N_5470,N_5514);
and U5572 (N_5572,N_5482,N_5496);
nor U5573 (N_5573,N_5480,N_5451);
nor U5574 (N_5574,N_5426,N_5467);
or U5575 (N_5575,N_5519,N_5431);
and U5576 (N_5576,N_5458,N_5537);
and U5577 (N_5577,N_5474,N_5517);
and U5578 (N_5578,N_5430,N_5503);
and U5579 (N_5579,N_5484,N_5494);
xnor U5580 (N_5580,N_5518,N_5462);
nand U5581 (N_5581,N_5455,N_5423);
or U5582 (N_5582,N_5416,N_5506);
xnor U5583 (N_5583,N_5487,N_5489);
or U5584 (N_5584,N_5505,N_5476);
xor U5585 (N_5585,N_5547,N_5549);
and U5586 (N_5586,N_5523,N_5406);
xor U5587 (N_5587,N_5526,N_5469);
xor U5588 (N_5588,N_5404,N_5436);
xnor U5589 (N_5589,N_5531,N_5499);
and U5590 (N_5590,N_5440,N_5448);
nor U5591 (N_5591,N_5498,N_5500);
or U5592 (N_5592,N_5539,N_5411);
or U5593 (N_5593,N_5545,N_5477);
xnor U5594 (N_5594,N_5501,N_5437);
nor U5595 (N_5595,N_5486,N_5428);
nand U5596 (N_5596,N_5433,N_5454);
nor U5597 (N_5597,N_5417,N_5532);
nor U5598 (N_5598,N_5475,N_5419);
xor U5599 (N_5599,N_5461,N_5402);
xnor U5600 (N_5600,N_5521,N_5400);
or U5601 (N_5601,N_5512,N_5457);
and U5602 (N_5602,N_5465,N_5460);
and U5603 (N_5603,N_5534,N_5434);
xnor U5604 (N_5604,N_5493,N_5497);
or U5605 (N_5605,N_5463,N_5483);
or U5606 (N_5606,N_5530,N_5424);
nand U5607 (N_5607,N_5524,N_5511);
nand U5608 (N_5608,N_5442,N_5525);
nor U5609 (N_5609,N_5427,N_5429);
nand U5610 (N_5610,N_5412,N_5504);
nand U5611 (N_5611,N_5472,N_5538);
nor U5612 (N_5612,N_5542,N_5447);
or U5613 (N_5613,N_5452,N_5473);
or U5614 (N_5614,N_5535,N_5435);
nor U5615 (N_5615,N_5478,N_5510);
or U5616 (N_5616,N_5515,N_5541);
nor U5617 (N_5617,N_5414,N_5516);
nand U5618 (N_5618,N_5485,N_5409);
nand U5619 (N_5619,N_5446,N_5466);
nand U5620 (N_5620,N_5522,N_5509);
and U5621 (N_5621,N_5422,N_5401);
nand U5622 (N_5622,N_5450,N_5490);
and U5623 (N_5623,N_5456,N_5471);
xnor U5624 (N_5624,N_5403,N_5544);
nand U5625 (N_5625,N_5430,N_5548);
or U5626 (N_5626,N_5407,N_5423);
nand U5627 (N_5627,N_5411,N_5513);
nand U5628 (N_5628,N_5465,N_5466);
xnor U5629 (N_5629,N_5415,N_5466);
nand U5630 (N_5630,N_5442,N_5505);
nand U5631 (N_5631,N_5443,N_5497);
or U5632 (N_5632,N_5529,N_5416);
nor U5633 (N_5633,N_5417,N_5514);
xor U5634 (N_5634,N_5454,N_5468);
and U5635 (N_5635,N_5488,N_5461);
nand U5636 (N_5636,N_5500,N_5508);
xor U5637 (N_5637,N_5459,N_5537);
and U5638 (N_5638,N_5438,N_5431);
nor U5639 (N_5639,N_5512,N_5456);
or U5640 (N_5640,N_5401,N_5418);
xor U5641 (N_5641,N_5499,N_5509);
or U5642 (N_5642,N_5495,N_5488);
xnor U5643 (N_5643,N_5457,N_5531);
nor U5644 (N_5644,N_5509,N_5473);
xnor U5645 (N_5645,N_5536,N_5437);
nand U5646 (N_5646,N_5455,N_5422);
nor U5647 (N_5647,N_5443,N_5511);
and U5648 (N_5648,N_5413,N_5505);
xnor U5649 (N_5649,N_5532,N_5538);
nand U5650 (N_5650,N_5428,N_5543);
and U5651 (N_5651,N_5449,N_5538);
nor U5652 (N_5652,N_5469,N_5509);
and U5653 (N_5653,N_5482,N_5497);
nand U5654 (N_5654,N_5541,N_5537);
or U5655 (N_5655,N_5533,N_5486);
nor U5656 (N_5656,N_5406,N_5546);
or U5657 (N_5657,N_5409,N_5428);
xnor U5658 (N_5658,N_5421,N_5453);
xnor U5659 (N_5659,N_5527,N_5409);
nor U5660 (N_5660,N_5500,N_5506);
or U5661 (N_5661,N_5407,N_5529);
or U5662 (N_5662,N_5444,N_5532);
and U5663 (N_5663,N_5492,N_5526);
nor U5664 (N_5664,N_5420,N_5438);
nand U5665 (N_5665,N_5502,N_5435);
xor U5666 (N_5666,N_5505,N_5420);
nor U5667 (N_5667,N_5448,N_5458);
nor U5668 (N_5668,N_5527,N_5521);
or U5669 (N_5669,N_5423,N_5513);
xor U5670 (N_5670,N_5453,N_5526);
or U5671 (N_5671,N_5474,N_5428);
nor U5672 (N_5672,N_5409,N_5548);
or U5673 (N_5673,N_5411,N_5493);
xnor U5674 (N_5674,N_5526,N_5503);
nand U5675 (N_5675,N_5467,N_5414);
and U5676 (N_5676,N_5443,N_5440);
or U5677 (N_5677,N_5491,N_5452);
xor U5678 (N_5678,N_5526,N_5509);
nor U5679 (N_5679,N_5518,N_5455);
or U5680 (N_5680,N_5514,N_5402);
nor U5681 (N_5681,N_5529,N_5496);
nor U5682 (N_5682,N_5430,N_5533);
xnor U5683 (N_5683,N_5454,N_5461);
nor U5684 (N_5684,N_5473,N_5418);
and U5685 (N_5685,N_5404,N_5461);
nor U5686 (N_5686,N_5443,N_5480);
nor U5687 (N_5687,N_5415,N_5444);
nand U5688 (N_5688,N_5501,N_5433);
nor U5689 (N_5689,N_5452,N_5533);
nand U5690 (N_5690,N_5491,N_5527);
nor U5691 (N_5691,N_5485,N_5426);
and U5692 (N_5692,N_5439,N_5526);
xnor U5693 (N_5693,N_5508,N_5488);
xnor U5694 (N_5694,N_5536,N_5489);
and U5695 (N_5695,N_5446,N_5473);
nand U5696 (N_5696,N_5517,N_5449);
or U5697 (N_5697,N_5544,N_5414);
and U5698 (N_5698,N_5420,N_5461);
or U5699 (N_5699,N_5498,N_5485);
and U5700 (N_5700,N_5595,N_5699);
and U5701 (N_5701,N_5684,N_5593);
nor U5702 (N_5702,N_5666,N_5698);
nor U5703 (N_5703,N_5675,N_5609);
xor U5704 (N_5704,N_5578,N_5563);
nand U5705 (N_5705,N_5587,N_5581);
nand U5706 (N_5706,N_5617,N_5667);
xnor U5707 (N_5707,N_5682,N_5550);
nand U5708 (N_5708,N_5697,N_5692);
nor U5709 (N_5709,N_5688,N_5621);
and U5710 (N_5710,N_5600,N_5589);
and U5711 (N_5711,N_5637,N_5565);
nor U5712 (N_5712,N_5645,N_5566);
or U5713 (N_5713,N_5661,N_5570);
or U5714 (N_5714,N_5574,N_5653);
nor U5715 (N_5715,N_5572,N_5611);
nand U5716 (N_5716,N_5649,N_5628);
nor U5717 (N_5717,N_5654,N_5632);
and U5718 (N_5718,N_5559,N_5672);
nor U5719 (N_5719,N_5660,N_5644);
and U5720 (N_5720,N_5608,N_5612);
nand U5721 (N_5721,N_5561,N_5659);
nand U5722 (N_5722,N_5626,N_5596);
nor U5723 (N_5723,N_5629,N_5582);
or U5724 (N_5724,N_5691,N_5634);
nand U5725 (N_5725,N_5671,N_5552);
nor U5726 (N_5726,N_5681,N_5610);
xnor U5727 (N_5727,N_5686,N_5562);
nand U5728 (N_5728,N_5607,N_5594);
nor U5729 (N_5729,N_5657,N_5683);
or U5730 (N_5730,N_5603,N_5636);
or U5731 (N_5731,N_5604,N_5590);
and U5732 (N_5732,N_5579,N_5555);
or U5733 (N_5733,N_5655,N_5668);
or U5734 (N_5734,N_5598,N_5631);
nor U5735 (N_5735,N_5568,N_5597);
or U5736 (N_5736,N_5647,N_5618);
and U5737 (N_5737,N_5576,N_5696);
nand U5738 (N_5738,N_5588,N_5642);
xnor U5739 (N_5739,N_5687,N_5680);
or U5740 (N_5740,N_5665,N_5586);
xor U5741 (N_5741,N_5567,N_5619);
and U5742 (N_5742,N_5616,N_5551);
xor U5743 (N_5743,N_5557,N_5569);
and U5744 (N_5744,N_5592,N_5679);
xnor U5745 (N_5745,N_5571,N_5658);
xnor U5746 (N_5746,N_5613,N_5640);
nor U5747 (N_5747,N_5630,N_5663);
or U5748 (N_5748,N_5620,N_5677);
nand U5749 (N_5749,N_5662,N_5556);
xnor U5750 (N_5750,N_5577,N_5639);
or U5751 (N_5751,N_5633,N_5615);
xnor U5752 (N_5752,N_5650,N_5606);
nor U5753 (N_5753,N_5689,N_5635);
or U5754 (N_5754,N_5673,N_5685);
xnor U5755 (N_5755,N_5584,N_5641);
and U5756 (N_5756,N_5646,N_5614);
or U5757 (N_5757,N_5638,N_5669);
nand U5758 (N_5758,N_5622,N_5580);
or U5759 (N_5759,N_5605,N_5585);
or U5760 (N_5760,N_5695,N_5678);
nor U5761 (N_5761,N_5624,N_5625);
or U5762 (N_5762,N_5656,N_5648);
or U5763 (N_5763,N_5599,N_5560);
nor U5764 (N_5764,N_5690,N_5573);
and U5765 (N_5765,N_5651,N_5693);
nand U5766 (N_5766,N_5575,N_5602);
and U5767 (N_5767,N_5591,N_5676);
xor U5768 (N_5768,N_5583,N_5670);
or U5769 (N_5769,N_5652,N_5674);
nor U5770 (N_5770,N_5554,N_5627);
nor U5771 (N_5771,N_5564,N_5643);
or U5772 (N_5772,N_5664,N_5553);
nor U5773 (N_5773,N_5558,N_5694);
and U5774 (N_5774,N_5601,N_5623);
xnor U5775 (N_5775,N_5594,N_5595);
or U5776 (N_5776,N_5599,N_5569);
and U5777 (N_5777,N_5627,N_5577);
xnor U5778 (N_5778,N_5577,N_5656);
or U5779 (N_5779,N_5553,N_5559);
and U5780 (N_5780,N_5668,N_5671);
nand U5781 (N_5781,N_5627,N_5696);
and U5782 (N_5782,N_5586,N_5675);
nor U5783 (N_5783,N_5638,N_5570);
nand U5784 (N_5784,N_5602,N_5588);
nand U5785 (N_5785,N_5696,N_5646);
and U5786 (N_5786,N_5637,N_5575);
and U5787 (N_5787,N_5599,N_5606);
xor U5788 (N_5788,N_5691,N_5621);
nand U5789 (N_5789,N_5584,N_5637);
nor U5790 (N_5790,N_5688,N_5565);
and U5791 (N_5791,N_5617,N_5683);
or U5792 (N_5792,N_5555,N_5696);
xnor U5793 (N_5793,N_5584,N_5668);
and U5794 (N_5794,N_5673,N_5602);
nor U5795 (N_5795,N_5595,N_5564);
nand U5796 (N_5796,N_5668,N_5562);
or U5797 (N_5797,N_5553,N_5569);
nand U5798 (N_5798,N_5658,N_5662);
nand U5799 (N_5799,N_5673,N_5659);
xor U5800 (N_5800,N_5636,N_5560);
and U5801 (N_5801,N_5580,N_5679);
nand U5802 (N_5802,N_5688,N_5695);
or U5803 (N_5803,N_5554,N_5686);
nand U5804 (N_5804,N_5688,N_5646);
and U5805 (N_5805,N_5654,N_5606);
nor U5806 (N_5806,N_5671,N_5653);
nand U5807 (N_5807,N_5661,N_5557);
and U5808 (N_5808,N_5637,N_5570);
nand U5809 (N_5809,N_5574,N_5554);
and U5810 (N_5810,N_5560,N_5639);
xor U5811 (N_5811,N_5660,N_5650);
nand U5812 (N_5812,N_5581,N_5676);
xor U5813 (N_5813,N_5660,N_5569);
xor U5814 (N_5814,N_5612,N_5688);
nor U5815 (N_5815,N_5608,N_5607);
nor U5816 (N_5816,N_5677,N_5678);
or U5817 (N_5817,N_5600,N_5679);
xnor U5818 (N_5818,N_5570,N_5590);
nand U5819 (N_5819,N_5620,N_5623);
xor U5820 (N_5820,N_5674,N_5585);
xnor U5821 (N_5821,N_5590,N_5666);
nand U5822 (N_5822,N_5650,N_5629);
xnor U5823 (N_5823,N_5673,N_5660);
and U5824 (N_5824,N_5582,N_5655);
nor U5825 (N_5825,N_5693,N_5563);
or U5826 (N_5826,N_5680,N_5562);
nor U5827 (N_5827,N_5616,N_5618);
nand U5828 (N_5828,N_5651,N_5580);
xnor U5829 (N_5829,N_5660,N_5600);
nand U5830 (N_5830,N_5578,N_5650);
xnor U5831 (N_5831,N_5597,N_5606);
nor U5832 (N_5832,N_5618,N_5641);
and U5833 (N_5833,N_5590,N_5643);
or U5834 (N_5834,N_5552,N_5690);
and U5835 (N_5835,N_5656,N_5583);
and U5836 (N_5836,N_5642,N_5585);
and U5837 (N_5837,N_5597,N_5659);
nor U5838 (N_5838,N_5656,N_5559);
or U5839 (N_5839,N_5582,N_5607);
nand U5840 (N_5840,N_5608,N_5603);
nand U5841 (N_5841,N_5601,N_5614);
xnor U5842 (N_5842,N_5570,N_5609);
or U5843 (N_5843,N_5583,N_5595);
nor U5844 (N_5844,N_5562,N_5678);
xnor U5845 (N_5845,N_5619,N_5659);
and U5846 (N_5846,N_5696,N_5679);
nor U5847 (N_5847,N_5557,N_5596);
and U5848 (N_5848,N_5696,N_5633);
and U5849 (N_5849,N_5616,N_5629);
nand U5850 (N_5850,N_5790,N_5728);
nor U5851 (N_5851,N_5782,N_5748);
and U5852 (N_5852,N_5796,N_5750);
and U5853 (N_5853,N_5822,N_5737);
nor U5854 (N_5854,N_5705,N_5788);
and U5855 (N_5855,N_5834,N_5771);
and U5856 (N_5856,N_5800,N_5746);
xor U5857 (N_5857,N_5846,N_5801);
nand U5858 (N_5858,N_5726,N_5794);
and U5859 (N_5859,N_5773,N_5747);
or U5860 (N_5860,N_5762,N_5751);
or U5861 (N_5861,N_5845,N_5824);
or U5862 (N_5862,N_5701,N_5725);
or U5863 (N_5863,N_5811,N_5786);
nor U5864 (N_5864,N_5848,N_5849);
xor U5865 (N_5865,N_5793,N_5778);
or U5866 (N_5866,N_5819,N_5755);
nor U5867 (N_5867,N_5807,N_5787);
nor U5868 (N_5868,N_5767,N_5826);
xnor U5869 (N_5869,N_5769,N_5843);
or U5870 (N_5870,N_5831,N_5772);
or U5871 (N_5871,N_5710,N_5765);
nor U5872 (N_5872,N_5842,N_5820);
nand U5873 (N_5873,N_5736,N_5797);
nor U5874 (N_5874,N_5722,N_5829);
or U5875 (N_5875,N_5818,N_5799);
xor U5876 (N_5876,N_5832,N_5830);
or U5877 (N_5877,N_5789,N_5717);
or U5878 (N_5878,N_5744,N_5702);
xor U5879 (N_5879,N_5735,N_5720);
or U5880 (N_5880,N_5847,N_5732);
or U5881 (N_5881,N_5753,N_5809);
xnor U5882 (N_5882,N_5740,N_5752);
nor U5883 (N_5883,N_5730,N_5835);
nor U5884 (N_5884,N_5731,N_5741);
or U5885 (N_5885,N_5754,N_5723);
nand U5886 (N_5886,N_5704,N_5758);
or U5887 (N_5887,N_5768,N_5838);
xnor U5888 (N_5888,N_5714,N_5745);
and U5889 (N_5889,N_5763,N_5810);
or U5890 (N_5890,N_5700,N_5775);
and U5891 (N_5891,N_5776,N_5805);
nand U5892 (N_5892,N_5711,N_5839);
xor U5893 (N_5893,N_5783,N_5708);
nor U5894 (N_5894,N_5812,N_5749);
xnor U5895 (N_5895,N_5804,N_5825);
and U5896 (N_5896,N_5817,N_5823);
and U5897 (N_5897,N_5709,N_5779);
nor U5898 (N_5898,N_5792,N_5733);
nand U5899 (N_5899,N_5815,N_5734);
nor U5900 (N_5900,N_5781,N_5713);
and U5901 (N_5901,N_5724,N_5759);
nor U5902 (N_5902,N_5739,N_5816);
and U5903 (N_5903,N_5795,N_5774);
nor U5904 (N_5904,N_5721,N_5770);
xor U5905 (N_5905,N_5707,N_5837);
xor U5906 (N_5906,N_5780,N_5764);
or U5907 (N_5907,N_5756,N_5738);
nand U5908 (N_5908,N_5791,N_5798);
nor U5909 (N_5909,N_5743,N_5706);
nor U5910 (N_5910,N_5827,N_5729);
nand U5911 (N_5911,N_5712,N_5833);
or U5912 (N_5912,N_5802,N_5840);
or U5913 (N_5913,N_5841,N_5766);
nand U5914 (N_5914,N_5784,N_5742);
nor U5915 (N_5915,N_5836,N_5806);
nor U5916 (N_5916,N_5808,N_5844);
or U5917 (N_5917,N_5785,N_5757);
and U5918 (N_5918,N_5761,N_5821);
and U5919 (N_5919,N_5703,N_5760);
nor U5920 (N_5920,N_5814,N_5718);
nand U5921 (N_5921,N_5813,N_5828);
or U5922 (N_5922,N_5777,N_5727);
nand U5923 (N_5923,N_5716,N_5719);
nand U5924 (N_5924,N_5715,N_5803);
or U5925 (N_5925,N_5757,N_5817);
xor U5926 (N_5926,N_5800,N_5712);
and U5927 (N_5927,N_5776,N_5768);
and U5928 (N_5928,N_5742,N_5777);
nand U5929 (N_5929,N_5811,N_5740);
nand U5930 (N_5930,N_5746,N_5788);
and U5931 (N_5931,N_5832,N_5750);
xor U5932 (N_5932,N_5733,N_5737);
xnor U5933 (N_5933,N_5712,N_5782);
xnor U5934 (N_5934,N_5741,N_5705);
and U5935 (N_5935,N_5752,N_5700);
or U5936 (N_5936,N_5837,N_5773);
xnor U5937 (N_5937,N_5724,N_5780);
nor U5938 (N_5938,N_5844,N_5756);
nand U5939 (N_5939,N_5764,N_5849);
nand U5940 (N_5940,N_5795,N_5828);
and U5941 (N_5941,N_5728,N_5808);
nor U5942 (N_5942,N_5829,N_5723);
nor U5943 (N_5943,N_5772,N_5702);
nand U5944 (N_5944,N_5714,N_5736);
xnor U5945 (N_5945,N_5807,N_5725);
or U5946 (N_5946,N_5807,N_5712);
and U5947 (N_5947,N_5744,N_5773);
nand U5948 (N_5948,N_5738,N_5744);
or U5949 (N_5949,N_5825,N_5755);
nand U5950 (N_5950,N_5793,N_5764);
xnor U5951 (N_5951,N_5781,N_5767);
nor U5952 (N_5952,N_5841,N_5716);
xnor U5953 (N_5953,N_5829,N_5728);
nand U5954 (N_5954,N_5732,N_5800);
or U5955 (N_5955,N_5703,N_5711);
nor U5956 (N_5956,N_5768,N_5791);
and U5957 (N_5957,N_5732,N_5844);
xor U5958 (N_5958,N_5767,N_5768);
or U5959 (N_5959,N_5835,N_5736);
xnor U5960 (N_5960,N_5727,N_5793);
xor U5961 (N_5961,N_5828,N_5796);
xor U5962 (N_5962,N_5843,N_5808);
nor U5963 (N_5963,N_5791,N_5749);
or U5964 (N_5964,N_5784,N_5753);
nand U5965 (N_5965,N_5811,N_5799);
nor U5966 (N_5966,N_5741,N_5739);
and U5967 (N_5967,N_5834,N_5701);
nand U5968 (N_5968,N_5823,N_5720);
nand U5969 (N_5969,N_5744,N_5750);
and U5970 (N_5970,N_5841,N_5754);
and U5971 (N_5971,N_5716,N_5806);
and U5972 (N_5972,N_5832,N_5833);
and U5973 (N_5973,N_5825,N_5738);
or U5974 (N_5974,N_5705,N_5762);
or U5975 (N_5975,N_5839,N_5778);
and U5976 (N_5976,N_5709,N_5730);
xnor U5977 (N_5977,N_5836,N_5735);
or U5978 (N_5978,N_5754,N_5733);
or U5979 (N_5979,N_5822,N_5828);
nor U5980 (N_5980,N_5720,N_5814);
nor U5981 (N_5981,N_5766,N_5847);
and U5982 (N_5982,N_5742,N_5736);
nor U5983 (N_5983,N_5742,N_5760);
nor U5984 (N_5984,N_5847,N_5765);
xnor U5985 (N_5985,N_5825,N_5813);
or U5986 (N_5986,N_5747,N_5816);
xor U5987 (N_5987,N_5795,N_5701);
nand U5988 (N_5988,N_5771,N_5753);
xnor U5989 (N_5989,N_5705,N_5763);
and U5990 (N_5990,N_5773,N_5785);
xnor U5991 (N_5991,N_5762,N_5756);
nand U5992 (N_5992,N_5700,N_5795);
and U5993 (N_5993,N_5830,N_5729);
and U5994 (N_5994,N_5732,N_5787);
nor U5995 (N_5995,N_5716,N_5753);
xor U5996 (N_5996,N_5780,N_5849);
or U5997 (N_5997,N_5731,N_5778);
and U5998 (N_5998,N_5704,N_5796);
xnor U5999 (N_5999,N_5796,N_5705);
xor U6000 (N_6000,N_5898,N_5854);
and U6001 (N_6001,N_5856,N_5955);
nand U6002 (N_6002,N_5954,N_5864);
or U6003 (N_6003,N_5937,N_5980);
and U6004 (N_6004,N_5858,N_5901);
nand U6005 (N_6005,N_5890,N_5940);
and U6006 (N_6006,N_5884,N_5870);
nor U6007 (N_6007,N_5969,N_5982);
xor U6008 (N_6008,N_5880,N_5956);
or U6009 (N_6009,N_5906,N_5863);
nand U6010 (N_6010,N_5896,N_5876);
nand U6011 (N_6011,N_5857,N_5914);
nand U6012 (N_6012,N_5855,N_5936);
and U6013 (N_6013,N_5965,N_5889);
xnor U6014 (N_6014,N_5860,N_5939);
xnor U6015 (N_6015,N_5902,N_5910);
xor U6016 (N_6016,N_5873,N_5948);
nand U6017 (N_6017,N_5951,N_5960);
nor U6018 (N_6018,N_5952,N_5893);
and U6019 (N_6019,N_5924,N_5975);
nand U6020 (N_6020,N_5859,N_5881);
xnor U6021 (N_6021,N_5989,N_5976);
nand U6022 (N_6022,N_5932,N_5851);
and U6023 (N_6023,N_5934,N_5981);
or U6024 (N_6024,N_5900,N_5929);
xnor U6025 (N_6025,N_5922,N_5915);
xor U6026 (N_6026,N_5899,N_5966);
and U6027 (N_6027,N_5988,N_5996);
nand U6028 (N_6028,N_5962,N_5938);
or U6029 (N_6029,N_5923,N_5943);
nand U6030 (N_6030,N_5973,N_5882);
nor U6031 (N_6031,N_5909,N_5968);
xnor U6032 (N_6032,N_5861,N_5986);
nor U6033 (N_6033,N_5897,N_5891);
or U6034 (N_6034,N_5983,N_5868);
and U6035 (N_6035,N_5925,N_5871);
or U6036 (N_6036,N_5978,N_5886);
nand U6037 (N_6037,N_5991,N_5994);
nand U6038 (N_6038,N_5892,N_5904);
nand U6039 (N_6039,N_5974,N_5958);
xor U6040 (N_6040,N_5850,N_5967);
nand U6041 (N_6041,N_5927,N_5919);
nor U6042 (N_6042,N_5885,N_5878);
nand U6043 (N_6043,N_5947,N_5874);
or U6044 (N_6044,N_5930,N_5963);
and U6045 (N_6045,N_5977,N_5888);
and U6046 (N_6046,N_5979,N_5877);
xnor U6047 (N_6047,N_5933,N_5872);
and U6048 (N_6048,N_5972,N_5964);
xnor U6049 (N_6049,N_5852,N_5853);
or U6050 (N_6050,N_5970,N_5944);
nor U6051 (N_6051,N_5931,N_5928);
and U6052 (N_6052,N_5905,N_5935);
nor U6053 (N_6053,N_5942,N_5887);
and U6054 (N_6054,N_5926,N_5879);
and U6055 (N_6055,N_5895,N_5971);
xnor U6056 (N_6056,N_5987,N_5992);
nor U6057 (N_6057,N_5990,N_5869);
and U6058 (N_6058,N_5993,N_5961);
or U6059 (N_6059,N_5946,N_5917);
or U6060 (N_6060,N_5867,N_5949);
xnor U6061 (N_6061,N_5865,N_5903);
or U6062 (N_6062,N_5883,N_5912);
or U6063 (N_6063,N_5953,N_5875);
nor U6064 (N_6064,N_5950,N_5913);
or U6065 (N_6065,N_5984,N_5957);
and U6066 (N_6066,N_5997,N_5998);
xnor U6067 (N_6067,N_5916,N_5920);
or U6068 (N_6068,N_5921,N_5894);
xor U6069 (N_6069,N_5911,N_5941);
and U6070 (N_6070,N_5862,N_5959);
nand U6071 (N_6071,N_5945,N_5918);
nand U6072 (N_6072,N_5999,N_5985);
nor U6073 (N_6073,N_5907,N_5995);
nor U6074 (N_6074,N_5908,N_5866);
and U6075 (N_6075,N_5920,N_5939);
xor U6076 (N_6076,N_5951,N_5957);
xor U6077 (N_6077,N_5957,N_5906);
or U6078 (N_6078,N_5877,N_5859);
xor U6079 (N_6079,N_5923,N_5985);
or U6080 (N_6080,N_5976,N_5938);
nor U6081 (N_6081,N_5946,N_5918);
and U6082 (N_6082,N_5886,N_5995);
and U6083 (N_6083,N_5899,N_5922);
nor U6084 (N_6084,N_5949,N_5970);
and U6085 (N_6085,N_5996,N_5859);
or U6086 (N_6086,N_5915,N_5918);
or U6087 (N_6087,N_5971,N_5951);
xor U6088 (N_6088,N_5860,N_5941);
nand U6089 (N_6089,N_5936,N_5884);
and U6090 (N_6090,N_5942,N_5967);
nand U6091 (N_6091,N_5989,N_5913);
nor U6092 (N_6092,N_5960,N_5976);
nand U6093 (N_6093,N_5860,N_5985);
xor U6094 (N_6094,N_5928,N_5968);
and U6095 (N_6095,N_5906,N_5995);
or U6096 (N_6096,N_5899,N_5987);
or U6097 (N_6097,N_5936,N_5893);
xor U6098 (N_6098,N_5900,N_5990);
nor U6099 (N_6099,N_5921,N_5916);
nor U6100 (N_6100,N_5942,N_5908);
nor U6101 (N_6101,N_5879,N_5918);
nand U6102 (N_6102,N_5885,N_5874);
or U6103 (N_6103,N_5958,N_5989);
or U6104 (N_6104,N_5991,N_5962);
nand U6105 (N_6105,N_5890,N_5856);
and U6106 (N_6106,N_5934,N_5968);
or U6107 (N_6107,N_5990,N_5930);
or U6108 (N_6108,N_5911,N_5907);
xor U6109 (N_6109,N_5979,N_5950);
and U6110 (N_6110,N_5890,N_5967);
and U6111 (N_6111,N_5975,N_5884);
xor U6112 (N_6112,N_5923,N_5859);
and U6113 (N_6113,N_5852,N_5910);
nor U6114 (N_6114,N_5883,N_5886);
nand U6115 (N_6115,N_5866,N_5971);
xor U6116 (N_6116,N_5958,N_5953);
nor U6117 (N_6117,N_5969,N_5892);
nand U6118 (N_6118,N_5882,N_5974);
and U6119 (N_6119,N_5869,N_5998);
nor U6120 (N_6120,N_5858,N_5863);
or U6121 (N_6121,N_5923,N_5924);
and U6122 (N_6122,N_5967,N_5889);
nand U6123 (N_6123,N_5902,N_5877);
or U6124 (N_6124,N_5989,N_5956);
nand U6125 (N_6125,N_5948,N_5872);
and U6126 (N_6126,N_5936,N_5850);
or U6127 (N_6127,N_5963,N_5927);
xor U6128 (N_6128,N_5971,N_5873);
nand U6129 (N_6129,N_5861,N_5999);
nor U6130 (N_6130,N_5973,N_5910);
nand U6131 (N_6131,N_5990,N_5884);
and U6132 (N_6132,N_5866,N_5876);
and U6133 (N_6133,N_5975,N_5949);
or U6134 (N_6134,N_5863,N_5953);
or U6135 (N_6135,N_5905,N_5874);
xor U6136 (N_6136,N_5974,N_5993);
and U6137 (N_6137,N_5911,N_5960);
and U6138 (N_6138,N_5908,N_5996);
and U6139 (N_6139,N_5904,N_5861);
or U6140 (N_6140,N_5898,N_5989);
nand U6141 (N_6141,N_5903,N_5967);
or U6142 (N_6142,N_5853,N_5982);
xnor U6143 (N_6143,N_5942,N_5866);
xor U6144 (N_6144,N_5966,N_5863);
and U6145 (N_6145,N_5985,N_5886);
and U6146 (N_6146,N_5939,N_5970);
and U6147 (N_6147,N_5907,N_5937);
xnor U6148 (N_6148,N_5997,N_5946);
or U6149 (N_6149,N_5964,N_5930);
and U6150 (N_6150,N_6140,N_6138);
nand U6151 (N_6151,N_6020,N_6133);
or U6152 (N_6152,N_6003,N_6129);
nand U6153 (N_6153,N_6013,N_6086);
and U6154 (N_6154,N_6096,N_6097);
or U6155 (N_6155,N_6027,N_6076);
nand U6156 (N_6156,N_6098,N_6116);
and U6157 (N_6157,N_6145,N_6068);
nand U6158 (N_6158,N_6092,N_6002);
nand U6159 (N_6159,N_6106,N_6095);
nor U6160 (N_6160,N_6084,N_6114);
or U6161 (N_6161,N_6072,N_6037);
nand U6162 (N_6162,N_6078,N_6118);
or U6163 (N_6163,N_6107,N_6099);
nor U6164 (N_6164,N_6043,N_6074);
xnor U6165 (N_6165,N_6119,N_6058);
or U6166 (N_6166,N_6124,N_6066);
xor U6167 (N_6167,N_6050,N_6073);
and U6168 (N_6168,N_6070,N_6014);
and U6169 (N_6169,N_6012,N_6089);
nand U6170 (N_6170,N_6031,N_6018);
nand U6171 (N_6171,N_6141,N_6046);
nand U6172 (N_6172,N_6139,N_6069);
and U6173 (N_6173,N_6094,N_6060);
xnor U6174 (N_6174,N_6065,N_6000);
xnor U6175 (N_6175,N_6144,N_6064);
xor U6176 (N_6176,N_6022,N_6080);
xor U6177 (N_6177,N_6075,N_6104);
nor U6178 (N_6178,N_6128,N_6059);
and U6179 (N_6179,N_6047,N_6103);
nand U6180 (N_6180,N_6035,N_6038);
nand U6181 (N_6181,N_6004,N_6036);
nor U6182 (N_6182,N_6148,N_6083);
nor U6183 (N_6183,N_6082,N_6123);
xnor U6184 (N_6184,N_6121,N_6052);
or U6185 (N_6185,N_6053,N_6111);
and U6186 (N_6186,N_6125,N_6093);
nand U6187 (N_6187,N_6044,N_6010);
nor U6188 (N_6188,N_6005,N_6011);
nand U6189 (N_6189,N_6113,N_6131);
xor U6190 (N_6190,N_6102,N_6019);
or U6191 (N_6191,N_6147,N_6120);
nor U6192 (N_6192,N_6023,N_6026);
nor U6193 (N_6193,N_6045,N_6100);
nand U6194 (N_6194,N_6146,N_6067);
xnor U6195 (N_6195,N_6142,N_6017);
and U6196 (N_6196,N_6015,N_6049);
and U6197 (N_6197,N_6122,N_6112);
or U6198 (N_6198,N_6127,N_6115);
or U6199 (N_6199,N_6087,N_6051);
or U6200 (N_6200,N_6024,N_6101);
xnor U6201 (N_6201,N_6117,N_6054);
nand U6202 (N_6202,N_6032,N_6149);
nand U6203 (N_6203,N_6137,N_6016);
nor U6204 (N_6204,N_6057,N_6091);
nor U6205 (N_6205,N_6132,N_6021);
or U6206 (N_6206,N_6001,N_6105);
xor U6207 (N_6207,N_6028,N_6025);
or U6208 (N_6208,N_6048,N_6056);
nor U6209 (N_6209,N_6063,N_6061);
or U6210 (N_6210,N_6136,N_6135);
or U6211 (N_6211,N_6126,N_6090);
and U6212 (N_6212,N_6108,N_6030);
or U6213 (N_6213,N_6041,N_6040);
and U6214 (N_6214,N_6143,N_6034);
or U6215 (N_6215,N_6081,N_6134);
or U6216 (N_6216,N_6085,N_6007);
and U6217 (N_6217,N_6088,N_6062);
or U6218 (N_6218,N_6077,N_6110);
nor U6219 (N_6219,N_6042,N_6009);
or U6220 (N_6220,N_6006,N_6033);
and U6221 (N_6221,N_6008,N_6055);
and U6222 (N_6222,N_6071,N_6130);
and U6223 (N_6223,N_6109,N_6029);
and U6224 (N_6224,N_6079,N_6039);
nor U6225 (N_6225,N_6051,N_6146);
xor U6226 (N_6226,N_6090,N_6093);
xnor U6227 (N_6227,N_6135,N_6049);
xnor U6228 (N_6228,N_6034,N_6024);
and U6229 (N_6229,N_6014,N_6135);
nor U6230 (N_6230,N_6072,N_6137);
or U6231 (N_6231,N_6121,N_6147);
or U6232 (N_6232,N_6105,N_6088);
nand U6233 (N_6233,N_6101,N_6019);
xor U6234 (N_6234,N_6078,N_6039);
and U6235 (N_6235,N_6139,N_6117);
xnor U6236 (N_6236,N_6083,N_6053);
nand U6237 (N_6237,N_6057,N_6038);
xor U6238 (N_6238,N_6092,N_6036);
nand U6239 (N_6239,N_6018,N_6111);
and U6240 (N_6240,N_6079,N_6075);
nor U6241 (N_6241,N_6086,N_6068);
and U6242 (N_6242,N_6143,N_6125);
nand U6243 (N_6243,N_6138,N_6059);
or U6244 (N_6244,N_6142,N_6065);
or U6245 (N_6245,N_6128,N_6138);
nor U6246 (N_6246,N_6060,N_6124);
nor U6247 (N_6247,N_6026,N_6073);
nor U6248 (N_6248,N_6060,N_6001);
nand U6249 (N_6249,N_6127,N_6126);
xor U6250 (N_6250,N_6059,N_6149);
nor U6251 (N_6251,N_6027,N_6006);
xor U6252 (N_6252,N_6136,N_6043);
nor U6253 (N_6253,N_6074,N_6011);
nor U6254 (N_6254,N_6009,N_6065);
nor U6255 (N_6255,N_6057,N_6145);
xor U6256 (N_6256,N_6033,N_6129);
and U6257 (N_6257,N_6109,N_6145);
nor U6258 (N_6258,N_6133,N_6118);
and U6259 (N_6259,N_6096,N_6141);
xnor U6260 (N_6260,N_6094,N_6047);
or U6261 (N_6261,N_6033,N_6121);
nor U6262 (N_6262,N_6029,N_6073);
nand U6263 (N_6263,N_6081,N_6102);
xor U6264 (N_6264,N_6043,N_6037);
or U6265 (N_6265,N_6012,N_6045);
and U6266 (N_6266,N_6093,N_6094);
nor U6267 (N_6267,N_6097,N_6131);
xor U6268 (N_6268,N_6086,N_6044);
nor U6269 (N_6269,N_6052,N_6014);
xnor U6270 (N_6270,N_6056,N_6043);
and U6271 (N_6271,N_6038,N_6098);
nor U6272 (N_6272,N_6082,N_6015);
nor U6273 (N_6273,N_6121,N_6036);
nor U6274 (N_6274,N_6030,N_6098);
or U6275 (N_6275,N_6050,N_6115);
xor U6276 (N_6276,N_6010,N_6032);
nor U6277 (N_6277,N_6052,N_6107);
xor U6278 (N_6278,N_6030,N_6083);
and U6279 (N_6279,N_6046,N_6131);
and U6280 (N_6280,N_6120,N_6009);
and U6281 (N_6281,N_6002,N_6100);
and U6282 (N_6282,N_6016,N_6067);
nor U6283 (N_6283,N_6034,N_6086);
xor U6284 (N_6284,N_6107,N_6104);
nor U6285 (N_6285,N_6141,N_6147);
xor U6286 (N_6286,N_6079,N_6049);
or U6287 (N_6287,N_6060,N_6086);
or U6288 (N_6288,N_6109,N_6139);
or U6289 (N_6289,N_6107,N_6011);
nor U6290 (N_6290,N_6079,N_6015);
xor U6291 (N_6291,N_6090,N_6147);
and U6292 (N_6292,N_6052,N_6129);
nand U6293 (N_6293,N_6003,N_6000);
nor U6294 (N_6294,N_6124,N_6039);
nand U6295 (N_6295,N_6019,N_6052);
nor U6296 (N_6296,N_6038,N_6107);
xnor U6297 (N_6297,N_6142,N_6092);
xor U6298 (N_6298,N_6090,N_6076);
nand U6299 (N_6299,N_6131,N_6115);
nor U6300 (N_6300,N_6155,N_6275);
nand U6301 (N_6301,N_6299,N_6263);
nand U6302 (N_6302,N_6161,N_6195);
and U6303 (N_6303,N_6237,N_6276);
and U6304 (N_6304,N_6264,N_6217);
nand U6305 (N_6305,N_6215,N_6178);
and U6306 (N_6306,N_6278,N_6203);
nor U6307 (N_6307,N_6223,N_6289);
or U6308 (N_6308,N_6251,N_6230);
nor U6309 (N_6309,N_6216,N_6265);
nor U6310 (N_6310,N_6181,N_6282);
xor U6311 (N_6311,N_6200,N_6254);
or U6312 (N_6312,N_6210,N_6151);
and U6313 (N_6313,N_6248,N_6219);
xor U6314 (N_6314,N_6287,N_6288);
or U6315 (N_6315,N_6165,N_6245);
or U6316 (N_6316,N_6191,N_6175);
nand U6317 (N_6317,N_6221,N_6247);
nand U6318 (N_6318,N_6242,N_6296);
xor U6319 (N_6319,N_6182,N_6295);
xor U6320 (N_6320,N_6260,N_6224);
and U6321 (N_6321,N_6189,N_6229);
or U6322 (N_6322,N_6177,N_6255);
nand U6323 (N_6323,N_6272,N_6298);
and U6324 (N_6324,N_6198,N_6171);
and U6325 (N_6325,N_6257,N_6158);
nor U6326 (N_6326,N_6222,N_6180);
nand U6327 (N_6327,N_6205,N_6162);
xnor U6328 (N_6328,N_6252,N_6283);
and U6329 (N_6329,N_6253,N_6174);
and U6330 (N_6330,N_6207,N_6235);
and U6331 (N_6331,N_6160,N_6281);
nand U6332 (N_6332,N_6268,N_6190);
nand U6333 (N_6333,N_6167,N_6294);
xor U6334 (N_6334,N_6150,N_6246);
xnor U6335 (N_6335,N_6183,N_6233);
and U6336 (N_6336,N_6184,N_6225);
and U6337 (N_6337,N_6214,N_6193);
and U6338 (N_6338,N_6166,N_6258);
xor U6339 (N_6339,N_6293,N_6292);
or U6340 (N_6340,N_6226,N_6279);
xnor U6341 (N_6341,N_6290,N_6164);
or U6342 (N_6342,N_6250,N_6199);
nand U6343 (N_6343,N_6176,N_6249);
nor U6344 (N_6344,N_6194,N_6243);
or U6345 (N_6345,N_6153,N_6234);
or U6346 (N_6346,N_6154,N_6280);
nor U6347 (N_6347,N_6269,N_6266);
xor U6348 (N_6348,N_6172,N_6170);
nand U6349 (N_6349,N_6188,N_6156);
nor U6350 (N_6350,N_6208,N_6274);
and U6351 (N_6351,N_6297,N_6227);
xor U6352 (N_6352,N_6192,N_6185);
or U6353 (N_6353,N_6197,N_6204);
and U6354 (N_6354,N_6201,N_6179);
nand U6355 (N_6355,N_6277,N_6218);
and U6356 (N_6356,N_6267,N_6261);
and U6357 (N_6357,N_6239,N_6163);
or U6358 (N_6358,N_6271,N_6236);
or U6359 (N_6359,N_6173,N_6259);
or U6360 (N_6360,N_6284,N_6256);
or U6361 (N_6361,N_6270,N_6169);
or U6362 (N_6362,N_6212,N_6206);
nor U6363 (N_6363,N_6244,N_6291);
nand U6364 (N_6364,N_6285,N_6157);
nor U6365 (N_6365,N_6187,N_6202);
and U6366 (N_6366,N_6241,N_6209);
and U6367 (N_6367,N_6168,N_6220);
or U6368 (N_6368,N_6238,N_6273);
and U6369 (N_6369,N_6228,N_6231);
xor U6370 (N_6370,N_6240,N_6213);
or U6371 (N_6371,N_6186,N_6211);
or U6372 (N_6372,N_6286,N_6232);
nand U6373 (N_6373,N_6262,N_6159);
xnor U6374 (N_6374,N_6196,N_6152);
xnor U6375 (N_6375,N_6201,N_6206);
nand U6376 (N_6376,N_6211,N_6168);
xnor U6377 (N_6377,N_6264,N_6261);
xnor U6378 (N_6378,N_6170,N_6292);
or U6379 (N_6379,N_6174,N_6194);
xnor U6380 (N_6380,N_6230,N_6202);
nor U6381 (N_6381,N_6204,N_6209);
nand U6382 (N_6382,N_6248,N_6268);
nor U6383 (N_6383,N_6261,N_6215);
and U6384 (N_6384,N_6218,N_6187);
xor U6385 (N_6385,N_6189,N_6243);
nor U6386 (N_6386,N_6236,N_6293);
and U6387 (N_6387,N_6213,N_6214);
nor U6388 (N_6388,N_6242,N_6194);
and U6389 (N_6389,N_6293,N_6275);
or U6390 (N_6390,N_6208,N_6267);
nor U6391 (N_6391,N_6289,N_6229);
xnor U6392 (N_6392,N_6222,N_6231);
nand U6393 (N_6393,N_6191,N_6163);
nor U6394 (N_6394,N_6284,N_6233);
and U6395 (N_6395,N_6253,N_6165);
xnor U6396 (N_6396,N_6150,N_6280);
or U6397 (N_6397,N_6245,N_6281);
nor U6398 (N_6398,N_6178,N_6234);
xor U6399 (N_6399,N_6256,N_6282);
nor U6400 (N_6400,N_6181,N_6212);
or U6401 (N_6401,N_6279,N_6218);
xnor U6402 (N_6402,N_6171,N_6234);
nor U6403 (N_6403,N_6232,N_6158);
xnor U6404 (N_6404,N_6247,N_6266);
xnor U6405 (N_6405,N_6258,N_6230);
xor U6406 (N_6406,N_6153,N_6178);
nor U6407 (N_6407,N_6178,N_6202);
and U6408 (N_6408,N_6179,N_6211);
or U6409 (N_6409,N_6188,N_6214);
nor U6410 (N_6410,N_6182,N_6208);
nand U6411 (N_6411,N_6172,N_6246);
xnor U6412 (N_6412,N_6291,N_6151);
xnor U6413 (N_6413,N_6205,N_6257);
and U6414 (N_6414,N_6270,N_6241);
xor U6415 (N_6415,N_6237,N_6266);
or U6416 (N_6416,N_6261,N_6276);
nor U6417 (N_6417,N_6151,N_6270);
nand U6418 (N_6418,N_6252,N_6282);
xnor U6419 (N_6419,N_6235,N_6201);
nor U6420 (N_6420,N_6299,N_6168);
or U6421 (N_6421,N_6249,N_6203);
nand U6422 (N_6422,N_6213,N_6290);
or U6423 (N_6423,N_6278,N_6181);
nor U6424 (N_6424,N_6268,N_6159);
or U6425 (N_6425,N_6182,N_6245);
nor U6426 (N_6426,N_6158,N_6295);
nand U6427 (N_6427,N_6289,N_6267);
or U6428 (N_6428,N_6274,N_6283);
or U6429 (N_6429,N_6204,N_6287);
or U6430 (N_6430,N_6256,N_6153);
nand U6431 (N_6431,N_6298,N_6257);
nand U6432 (N_6432,N_6273,N_6192);
xor U6433 (N_6433,N_6183,N_6216);
nand U6434 (N_6434,N_6284,N_6189);
or U6435 (N_6435,N_6216,N_6163);
nor U6436 (N_6436,N_6204,N_6265);
nor U6437 (N_6437,N_6157,N_6155);
nor U6438 (N_6438,N_6298,N_6299);
or U6439 (N_6439,N_6243,N_6207);
and U6440 (N_6440,N_6162,N_6161);
xor U6441 (N_6441,N_6252,N_6299);
and U6442 (N_6442,N_6253,N_6242);
xnor U6443 (N_6443,N_6163,N_6211);
or U6444 (N_6444,N_6282,N_6247);
nor U6445 (N_6445,N_6220,N_6196);
xnor U6446 (N_6446,N_6214,N_6170);
xor U6447 (N_6447,N_6205,N_6291);
nor U6448 (N_6448,N_6182,N_6210);
or U6449 (N_6449,N_6296,N_6245);
nor U6450 (N_6450,N_6308,N_6375);
nand U6451 (N_6451,N_6422,N_6377);
nor U6452 (N_6452,N_6382,N_6318);
nand U6453 (N_6453,N_6418,N_6345);
xnor U6454 (N_6454,N_6338,N_6307);
xor U6455 (N_6455,N_6446,N_6328);
and U6456 (N_6456,N_6416,N_6432);
nor U6457 (N_6457,N_6369,N_6306);
and U6458 (N_6458,N_6309,N_6447);
nor U6459 (N_6459,N_6439,N_6372);
and U6460 (N_6460,N_6426,N_6398);
nor U6461 (N_6461,N_6431,N_6429);
nor U6462 (N_6462,N_6441,N_6317);
xor U6463 (N_6463,N_6443,N_6344);
nand U6464 (N_6464,N_6384,N_6341);
nand U6465 (N_6465,N_6348,N_6379);
or U6466 (N_6466,N_6406,N_6410);
or U6467 (N_6467,N_6436,N_6365);
or U6468 (N_6468,N_6347,N_6411);
nand U6469 (N_6469,N_6364,N_6357);
nand U6470 (N_6470,N_6373,N_6337);
or U6471 (N_6471,N_6305,N_6424);
or U6472 (N_6472,N_6423,N_6433);
or U6473 (N_6473,N_6339,N_6437);
and U6474 (N_6474,N_6427,N_6430);
nor U6475 (N_6475,N_6445,N_6312);
nor U6476 (N_6476,N_6351,N_6353);
or U6477 (N_6477,N_6381,N_6335);
xnor U6478 (N_6478,N_6327,N_6334);
nor U6479 (N_6479,N_6371,N_6326);
and U6480 (N_6480,N_6301,N_6389);
or U6481 (N_6481,N_6388,N_6378);
and U6482 (N_6482,N_6444,N_6362);
and U6483 (N_6483,N_6354,N_6387);
nor U6484 (N_6484,N_6415,N_6329);
nor U6485 (N_6485,N_6409,N_6325);
or U6486 (N_6486,N_6352,N_6303);
or U6487 (N_6487,N_6385,N_6396);
nor U6488 (N_6488,N_6333,N_6331);
or U6489 (N_6489,N_6425,N_6340);
or U6490 (N_6490,N_6408,N_6413);
and U6491 (N_6491,N_6394,N_6403);
nand U6492 (N_6492,N_6435,N_6405);
and U6493 (N_6493,N_6342,N_6304);
or U6494 (N_6494,N_6361,N_6370);
and U6495 (N_6495,N_6376,N_6434);
nor U6496 (N_6496,N_6383,N_6402);
nor U6497 (N_6497,N_6336,N_6324);
nor U6498 (N_6498,N_6392,N_6400);
or U6499 (N_6499,N_6358,N_6314);
xor U6500 (N_6500,N_6440,N_6419);
xor U6501 (N_6501,N_6420,N_6428);
xnor U6502 (N_6502,N_6349,N_6380);
nor U6503 (N_6503,N_6442,N_6356);
and U6504 (N_6504,N_6368,N_6311);
nor U6505 (N_6505,N_6401,N_6449);
or U6506 (N_6506,N_6448,N_6395);
nand U6507 (N_6507,N_6315,N_6320);
xor U6508 (N_6508,N_6321,N_6300);
nor U6509 (N_6509,N_6316,N_6397);
or U6510 (N_6510,N_6346,N_6355);
nor U6511 (N_6511,N_6374,N_6386);
nand U6512 (N_6512,N_6391,N_6438);
nand U6513 (N_6513,N_6390,N_6412);
nand U6514 (N_6514,N_6302,N_6363);
nor U6515 (N_6515,N_6313,N_6404);
nor U6516 (N_6516,N_6323,N_6310);
or U6517 (N_6517,N_6399,N_6322);
nand U6518 (N_6518,N_6332,N_6407);
or U6519 (N_6519,N_6343,N_6330);
or U6520 (N_6520,N_6393,N_6359);
or U6521 (N_6521,N_6350,N_6360);
nor U6522 (N_6522,N_6414,N_6421);
and U6523 (N_6523,N_6417,N_6366);
nor U6524 (N_6524,N_6367,N_6319);
nand U6525 (N_6525,N_6356,N_6320);
nor U6526 (N_6526,N_6431,N_6347);
nand U6527 (N_6527,N_6324,N_6351);
xnor U6528 (N_6528,N_6438,N_6385);
xnor U6529 (N_6529,N_6376,N_6384);
nand U6530 (N_6530,N_6377,N_6427);
nor U6531 (N_6531,N_6368,N_6399);
nor U6532 (N_6532,N_6388,N_6379);
nand U6533 (N_6533,N_6371,N_6383);
or U6534 (N_6534,N_6317,N_6449);
nor U6535 (N_6535,N_6373,N_6384);
xor U6536 (N_6536,N_6408,N_6418);
nor U6537 (N_6537,N_6360,N_6380);
or U6538 (N_6538,N_6411,N_6384);
nor U6539 (N_6539,N_6328,N_6394);
and U6540 (N_6540,N_6317,N_6374);
or U6541 (N_6541,N_6385,N_6388);
nor U6542 (N_6542,N_6396,N_6314);
nor U6543 (N_6543,N_6379,N_6374);
and U6544 (N_6544,N_6416,N_6372);
nor U6545 (N_6545,N_6425,N_6347);
or U6546 (N_6546,N_6335,N_6397);
or U6547 (N_6547,N_6325,N_6417);
nor U6548 (N_6548,N_6391,N_6340);
nand U6549 (N_6549,N_6355,N_6425);
and U6550 (N_6550,N_6436,N_6405);
xor U6551 (N_6551,N_6396,N_6449);
and U6552 (N_6552,N_6339,N_6436);
or U6553 (N_6553,N_6356,N_6359);
nor U6554 (N_6554,N_6410,N_6333);
or U6555 (N_6555,N_6418,N_6327);
or U6556 (N_6556,N_6302,N_6341);
nand U6557 (N_6557,N_6441,N_6435);
nand U6558 (N_6558,N_6397,N_6343);
nand U6559 (N_6559,N_6400,N_6390);
nor U6560 (N_6560,N_6422,N_6394);
nand U6561 (N_6561,N_6384,N_6413);
or U6562 (N_6562,N_6335,N_6448);
nand U6563 (N_6563,N_6327,N_6393);
xor U6564 (N_6564,N_6348,N_6409);
and U6565 (N_6565,N_6317,N_6322);
xnor U6566 (N_6566,N_6370,N_6324);
and U6567 (N_6567,N_6383,N_6398);
nand U6568 (N_6568,N_6421,N_6392);
or U6569 (N_6569,N_6307,N_6368);
and U6570 (N_6570,N_6438,N_6426);
nand U6571 (N_6571,N_6380,N_6432);
or U6572 (N_6572,N_6393,N_6397);
and U6573 (N_6573,N_6429,N_6442);
and U6574 (N_6574,N_6330,N_6421);
nand U6575 (N_6575,N_6429,N_6438);
nand U6576 (N_6576,N_6426,N_6417);
and U6577 (N_6577,N_6328,N_6338);
nand U6578 (N_6578,N_6434,N_6379);
and U6579 (N_6579,N_6413,N_6439);
xor U6580 (N_6580,N_6343,N_6358);
nor U6581 (N_6581,N_6303,N_6429);
nor U6582 (N_6582,N_6448,N_6424);
and U6583 (N_6583,N_6367,N_6336);
or U6584 (N_6584,N_6338,N_6329);
and U6585 (N_6585,N_6436,N_6414);
nand U6586 (N_6586,N_6378,N_6411);
xnor U6587 (N_6587,N_6386,N_6304);
xor U6588 (N_6588,N_6316,N_6441);
nor U6589 (N_6589,N_6433,N_6406);
nand U6590 (N_6590,N_6436,N_6442);
nand U6591 (N_6591,N_6319,N_6393);
and U6592 (N_6592,N_6302,N_6334);
or U6593 (N_6593,N_6430,N_6404);
nor U6594 (N_6594,N_6415,N_6416);
nand U6595 (N_6595,N_6392,N_6317);
nor U6596 (N_6596,N_6348,N_6335);
and U6597 (N_6597,N_6390,N_6303);
nand U6598 (N_6598,N_6328,N_6418);
or U6599 (N_6599,N_6315,N_6353);
xnor U6600 (N_6600,N_6546,N_6486);
nor U6601 (N_6601,N_6516,N_6489);
and U6602 (N_6602,N_6588,N_6577);
nand U6603 (N_6603,N_6578,N_6551);
nor U6604 (N_6604,N_6460,N_6527);
or U6605 (N_6605,N_6572,N_6511);
xor U6606 (N_6606,N_6476,N_6548);
xnor U6607 (N_6607,N_6462,N_6458);
nand U6608 (N_6608,N_6478,N_6568);
xnor U6609 (N_6609,N_6512,N_6484);
nand U6610 (N_6610,N_6480,N_6494);
and U6611 (N_6611,N_6581,N_6554);
and U6612 (N_6612,N_6457,N_6450);
xnor U6613 (N_6613,N_6495,N_6563);
or U6614 (N_6614,N_6580,N_6515);
nand U6615 (N_6615,N_6540,N_6467);
or U6616 (N_6616,N_6465,N_6526);
or U6617 (N_6617,N_6496,N_6452);
and U6618 (N_6618,N_6524,N_6505);
xor U6619 (N_6619,N_6575,N_6593);
or U6620 (N_6620,N_6453,N_6522);
xor U6621 (N_6621,N_6487,N_6541);
nand U6622 (N_6622,N_6592,N_6594);
xnor U6623 (N_6623,N_6565,N_6474);
or U6624 (N_6624,N_6557,N_6523);
and U6625 (N_6625,N_6454,N_6517);
nor U6626 (N_6626,N_6477,N_6596);
xnor U6627 (N_6627,N_6525,N_6536);
nor U6628 (N_6628,N_6520,N_6573);
xnor U6629 (N_6629,N_6564,N_6552);
or U6630 (N_6630,N_6485,N_6451);
and U6631 (N_6631,N_6555,N_6514);
or U6632 (N_6632,N_6459,N_6483);
and U6633 (N_6633,N_6519,N_6499);
xnor U6634 (N_6634,N_6497,N_6531);
or U6635 (N_6635,N_6510,N_6533);
or U6636 (N_6636,N_6542,N_6561);
or U6637 (N_6637,N_6560,N_6455);
nand U6638 (N_6638,N_6583,N_6569);
xor U6639 (N_6639,N_6598,N_6558);
or U6640 (N_6640,N_6549,N_6509);
or U6641 (N_6641,N_6585,N_6481);
or U6642 (N_6642,N_6534,N_6539);
and U6643 (N_6643,N_6550,N_6518);
xnor U6644 (N_6644,N_6456,N_6466);
or U6645 (N_6645,N_6538,N_6503);
and U6646 (N_6646,N_6579,N_6591);
nand U6647 (N_6647,N_6587,N_6513);
nor U6648 (N_6648,N_6464,N_6472);
or U6649 (N_6649,N_6491,N_6500);
nand U6650 (N_6650,N_6566,N_6488);
nand U6651 (N_6651,N_6553,N_6586);
nand U6652 (N_6652,N_6532,N_6528);
nor U6653 (N_6653,N_6475,N_6556);
and U6654 (N_6654,N_6521,N_6463);
xnor U6655 (N_6655,N_6576,N_6493);
or U6656 (N_6656,N_6461,N_6570);
and U6657 (N_6657,N_6530,N_6562);
or U6658 (N_6658,N_6589,N_6470);
nand U6659 (N_6659,N_6469,N_6544);
or U6660 (N_6660,N_6545,N_6473);
xor U6661 (N_6661,N_6597,N_6507);
or U6662 (N_6662,N_6492,N_6547);
and U6663 (N_6663,N_6498,N_6502);
and U6664 (N_6664,N_6590,N_6506);
nand U6665 (N_6665,N_6535,N_6529);
or U6666 (N_6666,N_6501,N_6468);
nor U6667 (N_6667,N_6537,N_6508);
nand U6668 (N_6668,N_6582,N_6490);
and U6669 (N_6669,N_6559,N_6574);
or U6670 (N_6670,N_6567,N_6571);
or U6671 (N_6671,N_6599,N_6543);
nand U6672 (N_6672,N_6482,N_6471);
nor U6673 (N_6673,N_6584,N_6595);
xnor U6674 (N_6674,N_6479,N_6504);
and U6675 (N_6675,N_6479,N_6547);
nand U6676 (N_6676,N_6470,N_6592);
nor U6677 (N_6677,N_6455,N_6467);
xnor U6678 (N_6678,N_6587,N_6555);
and U6679 (N_6679,N_6471,N_6521);
and U6680 (N_6680,N_6598,N_6581);
nand U6681 (N_6681,N_6504,N_6564);
nor U6682 (N_6682,N_6547,N_6507);
or U6683 (N_6683,N_6506,N_6502);
nand U6684 (N_6684,N_6482,N_6541);
nand U6685 (N_6685,N_6568,N_6457);
nor U6686 (N_6686,N_6521,N_6530);
nor U6687 (N_6687,N_6477,N_6470);
or U6688 (N_6688,N_6579,N_6515);
xnor U6689 (N_6689,N_6553,N_6518);
xor U6690 (N_6690,N_6531,N_6454);
or U6691 (N_6691,N_6542,N_6544);
xor U6692 (N_6692,N_6544,N_6541);
and U6693 (N_6693,N_6454,N_6472);
nand U6694 (N_6694,N_6545,N_6544);
or U6695 (N_6695,N_6477,N_6452);
or U6696 (N_6696,N_6599,N_6451);
nor U6697 (N_6697,N_6522,N_6598);
nor U6698 (N_6698,N_6559,N_6549);
nor U6699 (N_6699,N_6559,N_6477);
nor U6700 (N_6700,N_6474,N_6536);
and U6701 (N_6701,N_6453,N_6598);
or U6702 (N_6702,N_6526,N_6587);
nor U6703 (N_6703,N_6522,N_6491);
nand U6704 (N_6704,N_6452,N_6585);
nor U6705 (N_6705,N_6517,N_6537);
or U6706 (N_6706,N_6507,N_6538);
nand U6707 (N_6707,N_6453,N_6599);
xor U6708 (N_6708,N_6538,N_6568);
and U6709 (N_6709,N_6548,N_6585);
nor U6710 (N_6710,N_6540,N_6553);
nand U6711 (N_6711,N_6547,N_6595);
or U6712 (N_6712,N_6519,N_6545);
and U6713 (N_6713,N_6511,N_6519);
or U6714 (N_6714,N_6453,N_6568);
nand U6715 (N_6715,N_6490,N_6528);
and U6716 (N_6716,N_6487,N_6521);
and U6717 (N_6717,N_6547,N_6537);
xor U6718 (N_6718,N_6570,N_6550);
nand U6719 (N_6719,N_6560,N_6527);
nand U6720 (N_6720,N_6527,N_6483);
nand U6721 (N_6721,N_6554,N_6573);
xor U6722 (N_6722,N_6545,N_6581);
and U6723 (N_6723,N_6519,N_6488);
and U6724 (N_6724,N_6578,N_6475);
nand U6725 (N_6725,N_6561,N_6589);
nand U6726 (N_6726,N_6512,N_6594);
or U6727 (N_6727,N_6595,N_6554);
xor U6728 (N_6728,N_6588,N_6519);
nor U6729 (N_6729,N_6598,N_6534);
nand U6730 (N_6730,N_6507,N_6568);
and U6731 (N_6731,N_6588,N_6571);
xor U6732 (N_6732,N_6467,N_6594);
nand U6733 (N_6733,N_6542,N_6464);
or U6734 (N_6734,N_6456,N_6458);
xor U6735 (N_6735,N_6484,N_6526);
nand U6736 (N_6736,N_6530,N_6597);
nor U6737 (N_6737,N_6571,N_6521);
and U6738 (N_6738,N_6549,N_6470);
or U6739 (N_6739,N_6495,N_6579);
and U6740 (N_6740,N_6575,N_6523);
nor U6741 (N_6741,N_6541,N_6525);
nand U6742 (N_6742,N_6549,N_6497);
nand U6743 (N_6743,N_6562,N_6531);
nand U6744 (N_6744,N_6584,N_6483);
and U6745 (N_6745,N_6541,N_6460);
xor U6746 (N_6746,N_6564,N_6464);
nand U6747 (N_6747,N_6458,N_6597);
nor U6748 (N_6748,N_6546,N_6587);
or U6749 (N_6749,N_6594,N_6596);
xor U6750 (N_6750,N_6648,N_6633);
nand U6751 (N_6751,N_6665,N_6725);
and U6752 (N_6752,N_6638,N_6676);
nor U6753 (N_6753,N_6670,N_6685);
and U6754 (N_6754,N_6611,N_6631);
nor U6755 (N_6755,N_6720,N_6733);
xor U6756 (N_6756,N_6716,N_6622);
or U6757 (N_6757,N_6635,N_6726);
and U6758 (N_6758,N_6601,N_6683);
xor U6759 (N_6759,N_6603,N_6744);
or U6760 (N_6760,N_6653,N_6710);
and U6761 (N_6761,N_6686,N_6620);
nor U6762 (N_6762,N_6694,N_6660);
xor U6763 (N_6763,N_6732,N_6628);
and U6764 (N_6764,N_6719,N_6636);
or U6765 (N_6765,N_6667,N_6619);
and U6766 (N_6766,N_6618,N_6668);
nor U6767 (N_6767,N_6637,N_6708);
or U6768 (N_6768,N_6729,N_6730);
and U6769 (N_6769,N_6711,N_6658);
and U6770 (N_6770,N_6738,N_6727);
nand U6771 (N_6771,N_6604,N_6680);
nor U6772 (N_6772,N_6722,N_6627);
and U6773 (N_6773,N_6659,N_6650);
nand U6774 (N_6774,N_6689,N_6723);
nand U6775 (N_6775,N_6697,N_6712);
nand U6776 (N_6776,N_6735,N_6656);
nor U6777 (N_6777,N_6669,N_6613);
and U6778 (N_6778,N_6693,N_6605);
nor U6779 (N_6779,N_6600,N_6609);
nand U6780 (N_6780,N_6645,N_6614);
and U6781 (N_6781,N_6649,N_6629);
or U6782 (N_6782,N_6717,N_6625);
nor U6783 (N_6783,N_6646,N_6715);
or U6784 (N_6784,N_6703,N_6639);
xnor U6785 (N_6785,N_6731,N_6734);
or U6786 (N_6786,N_6664,N_6675);
nor U6787 (N_6787,N_6632,N_6654);
and U6788 (N_6788,N_6663,N_6709);
xor U6789 (N_6789,N_6721,N_6749);
or U6790 (N_6790,N_6748,N_6747);
or U6791 (N_6791,N_6692,N_6674);
nor U6792 (N_6792,N_6702,N_6700);
nor U6793 (N_6793,N_6671,N_6696);
nor U6794 (N_6794,N_6606,N_6737);
nor U6795 (N_6795,N_6607,N_6678);
and U6796 (N_6796,N_6673,N_6666);
or U6797 (N_6797,N_6657,N_6699);
nor U6798 (N_6798,N_6704,N_6736);
nor U6799 (N_6799,N_6679,N_6621);
and U6800 (N_6800,N_6691,N_6707);
or U6801 (N_6801,N_6740,N_6724);
nor U6802 (N_6802,N_6718,N_6623);
xnor U6803 (N_6803,N_6651,N_6610);
nand U6804 (N_6804,N_6687,N_6612);
xnor U6805 (N_6805,N_6617,N_6662);
and U6806 (N_6806,N_6742,N_6655);
xor U6807 (N_6807,N_6642,N_6713);
and U6808 (N_6808,N_6684,N_6634);
or U6809 (N_6809,N_6652,N_6743);
nand U6810 (N_6810,N_6644,N_6641);
xor U6811 (N_6811,N_6745,N_6682);
or U6812 (N_6812,N_6688,N_6602);
nor U6813 (N_6813,N_6640,N_6608);
and U6814 (N_6814,N_6672,N_6705);
or U6815 (N_6815,N_6630,N_6728);
and U6816 (N_6816,N_6661,N_6624);
xor U6817 (N_6817,N_6698,N_6643);
nor U6818 (N_6818,N_6739,N_6626);
nand U6819 (N_6819,N_6677,N_6615);
xor U6820 (N_6820,N_6695,N_6681);
or U6821 (N_6821,N_6616,N_6690);
xnor U6822 (N_6822,N_6746,N_6741);
xor U6823 (N_6823,N_6647,N_6706);
nor U6824 (N_6824,N_6714,N_6701);
nor U6825 (N_6825,N_6646,N_6706);
and U6826 (N_6826,N_6742,N_6738);
xnor U6827 (N_6827,N_6668,N_6731);
xnor U6828 (N_6828,N_6714,N_6744);
nand U6829 (N_6829,N_6627,N_6709);
and U6830 (N_6830,N_6601,N_6705);
nand U6831 (N_6831,N_6693,N_6637);
nor U6832 (N_6832,N_6624,N_6738);
xnor U6833 (N_6833,N_6621,N_6712);
or U6834 (N_6834,N_6687,N_6675);
nor U6835 (N_6835,N_6662,N_6623);
or U6836 (N_6836,N_6666,N_6602);
or U6837 (N_6837,N_6708,N_6738);
nor U6838 (N_6838,N_6708,N_6743);
nor U6839 (N_6839,N_6617,N_6716);
and U6840 (N_6840,N_6671,N_6738);
or U6841 (N_6841,N_6640,N_6600);
or U6842 (N_6842,N_6662,N_6739);
nor U6843 (N_6843,N_6664,N_6683);
nor U6844 (N_6844,N_6689,N_6730);
nor U6845 (N_6845,N_6666,N_6710);
xnor U6846 (N_6846,N_6616,N_6601);
xor U6847 (N_6847,N_6693,N_6611);
nand U6848 (N_6848,N_6618,N_6627);
nor U6849 (N_6849,N_6640,N_6698);
nor U6850 (N_6850,N_6628,N_6655);
and U6851 (N_6851,N_6620,N_6740);
nor U6852 (N_6852,N_6649,N_6654);
nor U6853 (N_6853,N_6743,N_6695);
nand U6854 (N_6854,N_6712,N_6636);
or U6855 (N_6855,N_6666,N_6676);
and U6856 (N_6856,N_6653,N_6737);
nor U6857 (N_6857,N_6623,N_6673);
or U6858 (N_6858,N_6677,N_6657);
nand U6859 (N_6859,N_6702,N_6625);
nor U6860 (N_6860,N_6626,N_6710);
nand U6861 (N_6861,N_6741,N_6629);
and U6862 (N_6862,N_6727,N_6650);
and U6863 (N_6863,N_6609,N_6740);
and U6864 (N_6864,N_6615,N_6716);
xnor U6865 (N_6865,N_6695,N_6732);
nand U6866 (N_6866,N_6653,N_6643);
xnor U6867 (N_6867,N_6638,N_6685);
or U6868 (N_6868,N_6641,N_6664);
nand U6869 (N_6869,N_6630,N_6668);
nand U6870 (N_6870,N_6714,N_6683);
xor U6871 (N_6871,N_6730,N_6618);
or U6872 (N_6872,N_6626,N_6666);
nor U6873 (N_6873,N_6647,N_6633);
and U6874 (N_6874,N_6664,N_6687);
or U6875 (N_6875,N_6649,N_6615);
and U6876 (N_6876,N_6605,N_6663);
nand U6877 (N_6877,N_6617,N_6664);
xnor U6878 (N_6878,N_6702,N_6668);
or U6879 (N_6879,N_6640,N_6615);
or U6880 (N_6880,N_6624,N_6697);
nor U6881 (N_6881,N_6619,N_6702);
or U6882 (N_6882,N_6726,N_6716);
and U6883 (N_6883,N_6618,N_6696);
and U6884 (N_6884,N_6623,N_6672);
nor U6885 (N_6885,N_6679,N_6662);
xnor U6886 (N_6886,N_6672,N_6691);
xnor U6887 (N_6887,N_6735,N_6627);
xnor U6888 (N_6888,N_6622,N_6695);
or U6889 (N_6889,N_6622,N_6661);
and U6890 (N_6890,N_6634,N_6705);
and U6891 (N_6891,N_6738,N_6635);
and U6892 (N_6892,N_6643,N_6743);
xnor U6893 (N_6893,N_6748,N_6671);
and U6894 (N_6894,N_6652,N_6629);
and U6895 (N_6895,N_6619,N_6656);
xnor U6896 (N_6896,N_6679,N_6685);
xor U6897 (N_6897,N_6625,N_6675);
and U6898 (N_6898,N_6695,N_6636);
and U6899 (N_6899,N_6706,N_6654);
and U6900 (N_6900,N_6813,N_6877);
nand U6901 (N_6901,N_6875,N_6852);
nand U6902 (N_6902,N_6887,N_6899);
and U6903 (N_6903,N_6823,N_6896);
or U6904 (N_6904,N_6751,N_6800);
or U6905 (N_6905,N_6857,N_6859);
or U6906 (N_6906,N_6882,N_6809);
xor U6907 (N_6907,N_6866,N_6829);
xor U6908 (N_6908,N_6753,N_6895);
or U6909 (N_6909,N_6861,N_6805);
xor U6910 (N_6910,N_6892,N_6757);
nor U6911 (N_6911,N_6837,N_6826);
nor U6912 (N_6912,N_6885,N_6860);
nor U6913 (N_6913,N_6867,N_6771);
xnor U6914 (N_6914,N_6766,N_6858);
nor U6915 (N_6915,N_6818,N_6897);
and U6916 (N_6916,N_6756,N_6844);
and U6917 (N_6917,N_6789,N_6865);
nor U6918 (N_6918,N_6776,N_6898);
nor U6919 (N_6919,N_6817,N_6886);
nor U6920 (N_6920,N_6758,N_6839);
or U6921 (N_6921,N_6773,N_6786);
or U6922 (N_6922,N_6827,N_6798);
or U6923 (N_6923,N_6750,N_6814);
or U6924 (N_6924,N_6787,N_6799);
and U6925 (N_6925,N_6774,N_6838);
nor U6926 (N_6926,N_6815,N_6890);
nor U6927 (N_6927,N_6894,N_6797);
or U6928 (N_6928,N_6816,N_6862);
or U6929 (N_6929,N_6811,N_6770);
xnor U6930 (N_6930,N_6795,N_6788);
or U6931 (N_6931,N_6842,N_6768);
or U6932 (N_6932,N_6848,N_6845);
nand U6933 (N_6933,N_6775,N_6840);
xor U6934 (N_6934,N_6828,N_6764);
nand U6935 (N_6935,N_6785,N_6841);
and U6936 (N_6936,N_6792,N_6765);
xor U6937 (N_6937,N_6880,N_6835);
nand U6938 (N_6938,N_6801,N_6802);
and U6939 (N_6939,N_6846,N_6879);
and U6940 (N_6940,N_6779,N_6819);
nand U6941 (N_6941,N_6834,N_6762);
and U6942 (N_6942,N_6876,N_6763);
and U6943 (N_6943,N_6783,N_6806);
or U6944 (N_6944,N_6863,N_6761);
nand U6945 (N_6945,N_6760,N_6820);
and U6946 (N_6946,N_6849,N_6843);
xor U6947 (N_6947,N_6833,N_6824);
or U6948 (N_6948,N_6864,N_6812);
xnor U6949 (N_6949,N_6796,N_6855);
and U6950 (N_6950,N_6791,N_6780);
and U6951 (N_6951,N_6891,N_6836);
nor U6952 (N_6952,N_6868,N_6830);
or U6953 (N_6953,N_6822,N_6883);
or U6954 (N_6954,N_6754,N_6825);
and U6955 (N_6955,N_6804,N_6778);
nor U6956 (N_6956,N_6873,N_6777);
and U6957 (N_6957,N_6870,N_6759);
nor U6958 (N_6958,N_6794,N_6767);
and U6959 (N_6959,N_6793,N_6851);
xnor U6960 (N_6960,N_6782,N_6784);
xnor U6961 (N_6961,N_6769,N_6803);
nor U6962 (N_6962,N_6872,N_6807);
nand U6963 (N_6963,N_6881,N_6850);
and U6964 (N_6964,N_6772,N_6831);
nand U6965 (N_6965,N_6808,N_6888);
nor U6966 (N_6966,N_6781,N_6854);
and U6967 (N_6967,N_6884,N_6856);
nand U6968 (N_6968,N_6869,N_6821);
or U6969 (N_6969,N_6847,N_6810);
nand U6970 (N_6970,N_6853,N_6874);
xnor U6971 (N_6971,N_6752,N_6755);
nand U6972 (N_6972,N_6878,N_6790);
nand U6973 (N_6973,N_6889,N_6871);
or U6974 (N_6974,N_6832,N_6893);
and U6975 (N_6975,N_6811,N_6854);
nand U6976 (N_6976,N_6897,N_6820);
and U6977 (N_6977,N_6841,N_6812);
nand U6978 (N_6978,N_6839,N_6810);
nor U6979 (N_6979,N_6823,N_6805);
nor U6980 (N_6980,N_6755,N_6792);
and U6981 (N_6981,N_6890,N_6845);
and U6982 (N_6982,N_6859,N_6849);
or U6983 (N_6983,N_6763,N_6848);
xor U6984 (N_6984,N_6812,N_6843);
and U6985 (N_6985,N_6884,N_6814);
nor U6986 (N_6986,N_6797,N_6893);
nand U6987 (N_6987,N_6892,N_6779);
xnor U6988 (N_6988,N_6813,N_6860);
and U6989 (N_6989,N_6849,N_6890);
or U6990 (N_6990,N_6757,N_6859);
or U6991 (N_6991,N_6821,N_6794);
nand U6992 (N_6992,N_6798,N_6876);
nand U6993 (N_6993,N_6865,N_6843);
nand U6994 (N_6994,N_6856,N_6838);
or U6995 (N_6995,N_6801,N_6750);
xor U6996 (N_6996,N_6818,N_6875);
and U6997 (N_6997,N_6807,N_6810);
nor U6998 (N_6998,N_6847,N_6768);
xor U6999 (N_6999,N_6897,N_6871);
or U7000 (N_7000,N_6761,N_6764);
nand U7001 (N_7001,N_6758,N_6771);
nand U7002 (N_7002,N_6809,N_6849);
nand U7003 (N_7003,N_6764,N_6848);
or U7004 (N_7004,N_6846,N_6847);
nand U7005 (N_7005,N_6865,N_6893);
nand U7006 (N_7006,N_6814,N_6781);
xnor U7007 (N_7007,N_6824,N_6755);
nor U7008 (N_7008,N_6762,N_6892);
nand U7009 (N_7009,N_6849,N_6753);
xnor U7010 (N_7010,N_6809,N_6775);
nor U7011 (N_7011,N_6835,N_6885);
and U7012 (N_7012,N_6833,N_6792);
or U7013 (N_7013,N_6762,N_6871);
nand U7014 (N_7014,N_6789,N_6800);
xnor U7015 (N_7015,N_6775,N_6862);
and U7016 (N_7016,N_6824,N_6769);
xnor U7017 (N_7017,N_6750,N_6769);
xor U7018 (N_7018,N_6772,N_6882);
nand U7019 (N_7019,N_6809,N_6855);
nor U7020 (N_7020,N_6797,N_6784);
nand U7021 (N_7021,N_6755,N_6856);
and U7022 (N_7022,N_6805,N_6752);
and U7023 (N_7023,N_6785,N_6771);
or U7024 (N_7024,N_6854,N_6863);
nor U7025 (N_7025,N_6835,N_6876);
or U7026 (N_7026,N_6823,N_6757);
nor U7027 (N_7027,N_6812,N_6754);
nor U7028 (N_7028,N_6783,N_6779);
xor U7029 (N_7029,N_6771,N_6811);
or U7030 (N_7030,N_6807,N_6799);
and U7031 (N_7031,N_6762,N_6877);
and U7032 (N_7032,N_6824,N_6772);
or U7033 (N_7033,N_6891,N_6757);
or U7034 (N_7034,N_6873,N_6813);
xor U7035 (N_7035,N_6878,N_6899);
xor U7036 (N_7036,N_6768,N_6882);
nand U7037 (N_7037,N_6894,N_6897);
xnor U7038 (N_7038,N_6768,N_6789);
nand U7039 (N_7039,N_6762,N_6805);
and U7040 (N_7040,N_6816,N_6822);
nand U7041 (N_7041,N_6756,N_6775);
nor U7042 (N_7042,N_6807,N_6800);
nor U7043 (N_7043,N_6769,N_6873);
or U7044 (N_7044,N_6769,N_6892);
or U7045 (N_7045,N_6809,N_6840);
nor U7046 (N_7046,N_6838,N_6891);
nor U7047 (N_7047,N_6773,N_6819);
or U7048 (N_7048,N_6857,N_6754);
nand U7049 (N_7049,N_6899,N_6775);
or U7050 (N_7050,N_6938,N_6971);
and U7051 (N_7051,N_6983,N_6913);
or U7052 (N_7052,N_6951,N_6949);
nand U7053 (N_7053,N_6980,N_6984);
xor U7054 (N_7054,N_7021,N_6964);
or U7055 (N_7055,N_7023,N_6925);
xor U7056 (N_7056,N_7035,N_6995);
xnor U7057 (N_7057,N_6985,N_6915);
nand U7058 (N_7058,N_6909,N_7019);
and U7059 (N_7059,N_6968,N_6939);
nor U7060 (N_7060,N_7000,N_7040);
xnor U7061 (N_7061,N_6933,N_7034);
and U7062 (N_7062,N_7032,N_6910);
or U7063 (N_7063,N_6994,N_6959);
nor U7064 (N_7064,N_6936,N_6927);
and U7065 (N_7065,N_6976,N_6952);
nor U7066 (N_7066,N_7038,N_6967);
nor U7067 (N_7067,N_6911,N_6931);
or U7068 (N_7068,N_7001,N_6953);
and U7069 (N_7069,N_7005,N_7031);
nand U7070 (N_7070,N_6975,N_6978);
or U7071 (N_7071,N_7002,N_6986);
xnor U7072 (N_7072,N_6946,N_7016);
and U7073 (N_7073,N_6997,N_6907);
or U7074 (N_7074,N_6932,N_6900);
or U7075 (N_7075,N_6917,N_6906);
or U7076 (N_7076,N_7004,N_6996);
and U7077 (N_7077,N_6903,N_6973);
and U7078 (N_7078,N_6942,N_6916);
or U7079 (N_7079,N_6961,N_6935);
nand U7080 (N_7080,N_6914,N_6957);
or U7081 (N_7081,N_6923,N_7036);
and U7082 (N_7082,N_6991,N_6960);
nor U7083 (N_7083,N_6930,N_7029);
nor U7084 (N_7084,N_7044,N_6920);
xnor U7085 (N_7085,N_7008,N_6981);
nand U7086 (N_7086,N_6919,N_6993);
xnor U7087 (N_7087,N_7048,N_7028);
nor U7088 (N_7088,N_7009,N_6926);
nand U7089 (N_7089,N_7033,N_6965);
or U7090 (N_7090,N_6962,N_7043);
nand U7091 (N_7091,N_6992,N_7030);
xor U7092 (N_7092,N_7047,N_6929);
nand U7093 (N_7093,N_6934,N_6904);
or U7094 (N_7094,N_7027,N_7037);
xor U7095 (N_7095,N_7014,N_6990);
and U7096 (N_7096,N_6956,N_6974);
or U7097 (N_7097,N_6982,N_7026);
nor U7098 (N_7098,N_6977,N_6958);
nor U7099 (N_7099,N_7003,N_7042);
xnor U7100 (N_7100,N_7017,N_6905);
nor U7101 (N_7101,N_6969,N_6966);
or U7102 (N_7102,N_6979,N_7011);
nand U7103 (N_7103,N_6921,N_6972);
or U7104 (N_7104,N_6912,N_6999);
and U7105 (N_7105,N_6943,N_6944);
nand U7106 (N_7106,N_7025,N_6908);
nor U7107 (N_7107,N_7007,N_6928);
or U7108 (N_7108,N_6947,N_7018);
nand U7109 (N_7109,N_6901,N_6902);
nand U7110 (N_7110,N_6954,N_7015);
nand U7111 (N_7111,N_7013,N_6989);
xor U7112 (N_7112,N_6988,N_7006);
nor U7113 (N_7113,N_6998,N_6918);
or U7114 (N_7114,N_7045,N_7010);
or U7115 (N_7115,N_7039,N_6937);
nand U7116 (N_7116,N_7049,N_7020);
xnor U7117 (N_7117,N_6987,N_6950);
nor U7118 (N_7118,N_6948,N_6963);
nor U7119 (N_7119,N_7022,N_7024);
nor U7120 (N_7120,N_7046,N_6941);
and U7121 (N_7121,N_6940,N_6945);
and U7122 (N_7122,N_6922,N_6955);
nand U7123 (N_7123,N_6924,N_6970);
or U7124 (N_7124,N_7041,N_7012);
or U7125 (N_7125,N_6978,N_6993);
nor U7126 (N_7126,N_7008,N_6938);
nand U7127 (N_7127,N_7028,N_7036);
xor U7128 (N_7128,N_6965,N_7036);
nand U7129 (N_7129,N_7049,N_6958);
xor U7130 (N_7130,N_6946,N_7039);
nor U7131 (N_7131,N_7019,N_7025);
or U7132 (N_7132,N_6920,N_7021);
or U7133 (N_7133,N_7000,N_7009);
and U7134 (N_7134,N_6928,N_6995);
or U7135 (N_7135,N_7039,N_6929);
xor U7136 (N_7136,N_6966,N_7008);
nand U7137 (N_7137,N_6943,N_7003);
nor U7138 (N_7138,N_6994,N_7006);
nor U7139 (N_7139,N_6921,N_7024);
nand U7140 (N_7140,N_6996,N_6995);
and U7141 (N_7141,N_6923,N_6931);
xor U7142 (N_7142,N_6979,N_6921);
and U7143 (N_7143,N_6974,N_6933);
or U7144 (N_7144,N_6913,N_7012);
and U7145 (N_7145,N_7042,N_6958);
nand U7146 (N_7146,N_7043,N_6929);
nand U7147 (N_7147,N_7041,N_7016);
xnor U7148 (N_7148,N_6961,N_7024);
or U7149 (N_7149,N_7021,N_6917);
nand U7150 (N_7150,N_7022,N_7013);
nand U7151 (N_7151,N_7023,N_6984);
xor U7152 (N_7152,N_6996,N_7025);
nor U7153 (N_7153,N_6957,N_6959);
and U7154 (N_7154,N_7040,N_7024);
or U7155 (N_7155,N_7034,N_7026);
and U7156 (N_7156,N_7001,N_7006);
nand U7157 (N_7157,N_7039,N_6910);
nor U7158 (N_7158,N_7049,N_6984);
nor U7159 (N_7159,N_7029,N_7048);
and U7160 (N_7160,N_6924,N_7021);
or U7161 (N_7161,N_6934,N_6961);
or U7162 (N_7162,N_6952,N_6969);
nand U7163 (N_7163,N_7012,N_7023);
and U7164 (N_7164,N_7037,N_7041);
or U7165 (N_7165,N_6968,N_6983);
and U7166 (N_7166,N_6955,N_7022);
and U7167 (N_7167,N_7006,N_6921);
xnor U7168 (N_7168,N_6944,N_6978);
and U7169 (N_7169,N_7020,N_7033);
or U7170 (N_7170,N_6968,N_7040);
and U7171 (N_7171,N_6939,N_6921);
nand U7172 (N_7172,N_6946,N_6985);
nand U7173 (N_7173,N_6911,N_6946);
nand U7174 (N_7174,N_6936,N_6921);
or U7175 (N_7175,N_7018,N_6955);
and U7176 (N_7176,N_6970,N_7026);
nor U7177 (N_7177,N_7036,N_6942);
or U7178 (N_7178,N_7002,N_6918);
xor U7179 (N_7179,N_7014,N_6942);
xnor U7180 (N_7180,N_7001,N_6927);
or U7181 (N_7181,N_6992,N_6956);
or U7182 (N_7182,N_6900,N_6920);
or U7183 (N_7183,N_6932,N_6985);
and U7184 (N_7184,N_6984,N_6929);
nor U7185 (N_7185,N_6976,N_6902);
or U7186 (N_7186,N_7031,N_7047);
or U7187 (N_7187,N_7008,N_6969);
and U7188 (N_7188,N_6996,N_6975);
and U7189 (N_7189,N_6955,N_6958);
nor U7190 (N_7190,N_6995,N_6957);
and U7191 (N_7191,N_6922,N_7016);
xnor U7192 (N_7192,N_7002,N_6962);
nand U7193 (N_7193,N_7043,N_7034);
and U7194 (N_7194,N_6957,N_7015);
or U7195 (N_7195,N_6977,N_6991);
xor U7196 (N_7196,N_6987,N_7041);
nand U7197 (N_7197,N_6918,N_7036);
nand U7198 (N_7198,N_7048,N_6929);
nor U7199 (N_7199,N_7019,N_6958);
xnor U7200 (N_7200,N_7174,N_7084);
nor U7201 (N_7201,N_7135,N_7136);
nand U7202 (N_7202,N_7097,N_7173);
xor U7203 (N_7203,N_7079,N_7188);
or U7204 (N_7204,N_7118,N_7158);
or U7205 (N_7205,N_7182,N_7137);
nor U7206 (N_7206,N_7092,N_7057);
or U7207 (N_7207,N_7122,N_7155);
nor U7208 (N_7208,N_7167,N_7153);
xnor U7209 (N_7209,N_7056,N_7119);
xnor U7210 (N_7210,N_7109,N_7123);
nor U7211 (N_7211,N_7177,N_7141);
nand U7212 (N_7212,N_7114,N_7060);
and U7213 (N_7213,N_7140,N_7179);
xnor U7214 (N_7214,N_7164,N_7178);
nor U7215 (N_7215,N_7147,N_7061);
or U7216 (N_7216,N_7134,N_7159);
xor U7217 (N_7217,N_7098,N_7152);
nand U7218 (N_7218,N_7130,N_7161);
nand U7219 (N_7219,N_7183,N_7185);
or U7220 (N_7220,N_7193,N_7051);
xnor U7221 (N_7221,N_7090,N_7081);
or U7222 (N_7222,N_7063,N_7133);
or U7223 (N_7223,N_7148,N_7068);
nor U7224 (N_7224,N_7184,N_7072);
or U7225 (N_7225,N_7100,N_7074);
or U7226 (N_7226,N_7125,N_7059);
xnor U7227 (N_7227,N_7160,N_7050);
xor U7228 (N_7228,N_7149,N_7089);
nand U7229 (N_7229,N_7088,N_7181);
or U7230 (N_7230,N_7139,N_7094);
nor U7231 (N_7231,N_7082,N_7091);
or U7232 (N_7232,N_7099,N_7199);
nor U7233 (N_7233,N_7190,N_7126);
nor U7234 (N_7234,N_7106,N_7166);
nand U7235 (N_7235,N_7145,N_7078);
nor U7236 (N_7236,N_7162,N_7103);
or U7237 (N_7237,N_7154,N_7080);
nor U7238 (N_7238,N_7151,N_7107);
nand U7239 (N_7239,N_7127,N_7053);
and U7240 (N_7240,N_7062,N_7120);
nand U7241 (N_7241,N_7191,N_7058);
and U7242 (N_7242,N_7128,N_7085);
nor U7243 (N_7243,N_7175,N_7116);
nor U7244 (N_7244,N_7157,N_7064);
nor U7245 (N_7245,N_7195,N_7086);
and U7246 (N_7246,N_7170,N_7142);
nand U7247 (N_7247,N_7146,N_7192);
nor U7248 (N_7248,N_7197,N_7093);
xnor U7249 (N_7249,N_7129,N_7075);
nand U7250 (N_7250,N_7189,N_7108);
nor U7251 (N_7251,N_7156,N_7150);
nand U7252 (N_7252,N_7095,N_7132);
nand U7253 (N_7253,N_7101,N_7052);
nand U7254 (N_7254,N_7087,N_7110);
or U7255 (N_7255,N_7104,N_7169);
and U7256 (N_7256,N_7067,N_7143);
and U7257 (N_7257,N_7054,N_7172);
xor U7258 (N_7258,N_7124,N_7165);
and U7259 (N_7259,N_7071,N_7186);
nor U7260 (N_7260,N_7069,N_7102);
or U7261 (N_7261,N_7066,N_7198);
or U7262 (N_7262,N_7065,N_7073);
xor U7263 (N_7263,N_7163,N_7138);
and U7264 (N_7264,N_7112,N_7131);
or U7265 (N_7265,N_7117,N_7083);
nor U7266 (N_7266,N_7171,N_7121);
xnor U7267 (N_7267,N_7070,N_7196);
nand U7268 (N_7268,N_7076,N_7077);
nand U7269 (N_7269,N_7144,N_7180);
nor U7270 (N_7270,N_7105,N_7187);
and U7271 (N_7271,N_7055,N_7115);
xor U7272 (N_7272,N_7168,N_7111);
or U7273 (N_7273,N_7194,N_7176);
or U7274 (N_7274,N_7096,N_7113);
or U7275 (N_7275,N_7096,N_7162);
nand U7276 (N_7276,N_7112,N_7182);
nor U7277 (N_7277,N_7129,N_7083);
xnor U7278 (N_7278,N_7126,N_7145);
nand U7279 (N_7279,N_7141,N_7093);
nor U7280 (N_7280,N_7193,N_7129);
and U7281 (N_7281,N_7065,N_7066);
and U7282 (N_7282,N_7062,N_7052);
or U7283 (N_7283,N_7112,N_7117);
or U7284 (N_7284,N_7081,N_7050);
xnor U7285 (N_7285,N_7122,N_7176);
xnor U7286 (N_7286,N_7178,N_7078);
nand U7287 (N_7287,N_7142,N_7121);
nor U7288 (N_7288,N_7178,N_7158);
or U7289 (N_7289,N_7193,N_7149);
and U7290 (N_7290,N_7086,N_7154);
nor U7291 (N_7291,N_7063,N_7178);
and U7292 (N_7292,N_7050,N_7077);
nor U7293 (N_7293,N_7083,N_7170);
and U7294 (N_7294,N_7064,N_7137);
and U7295 (N_7295,N_7070,N_7097);
and U7296 (N_7296,N_7086,N_7104);
nand U7297 (N_7297,N_7157,N_7164);
xnor U7298 (N_7298,N_7162,N_7090);
and U7299 (N_7299,N_7091,N_7095);
or U7300 (N_7300,N_7116,N_7159);
xor U7301 (N_7301,N_7056,N_7156);
and U7302 (N_7302,N_7183,N_7169);
nor U7303 (N_7303,N_7154,N_7057);
nand U7304 (N_7304,N_7182,N_7138);
or U7305 (N_7305,N_7066,N_7196);
xnor U7306 (N_7306,N_7088,N_7094);
xor U7307 (N_7307,N_7132,N_7169);
nor U7308 (N_7308,N_7174,N_7109);
xnor U7309 (N_7309,N_7164,N_7085);
nand U7310 (N_7310,N_7176,N_7128);
nor U7311 (N_7311,N_7141,N_7084);
or U7312 (N_7312,N_7063,N_7183);
and U7313 (N_7313,N_7092,N_7194);
or U7314 (N_7314,N_7182,N_7145);
nand U7315 (N_7315,N_7154,N_7197);
or U7316 (N_7316,N_7167,N_7163);
and U7317 (N_7317,N_7174,N_7094);
xor U7318 (N_7318,N_7120,N_7167);
nand U7319 (N_7319,N_7199,N_7085);
and U7320 (N_7320,N_7051,N_7115);
nor U7321 (N_7321,N_7124,N_7062);
xor U7322 (N_7322,N_7178,N_7077);
or U7323 (N_7323,N_7196,N_7111);
nor U7324 (N_7324,N_7095,N_7121);
or U7325 (N_7325,N_7081,N_7086);
or U7326 (N_7326,N_7061,N_7066);
nor U7327 (N_7327,N_7159,N_7099);
xnor U7328 (N_7328,N_7053,N_7060);
xnor U7329 (N_7329,N_7160,N_7130);
xor U7330 (N_7330,N_7168,N_7192);
and U7331 (N_7331,N_7137,N_7196);
nor U7332 (N_7332,N_7164,N_7095);
and U7333 (N_7333,N_7104,N_7173);
or U7334 (N_7334,N_7050,N_7074);
or U7335 (N_7335,N_7100,N_7159);
nand U7336 (N_7336,N_7171,N_7125);
or U7337 (N_7337,N_7124,N_7095);
xor U7338 (N_7338,N_7155,N_7071);
nor U7339 (N_7339,N_7195,N_7185);
or U7340 (N_7340,N_7130,N_7171);
and U7341 (N_7341,N_7092,N_7164);
nand U7342 (N_7342,N_7074,N_7130);
and U7343 (N_7343,N_7082,N_7163);
xnor U7344 (N_7344,N_7073,N_7132);
nor U7345 (N_7345,N_7197,N_7112);
xor U7346 (N_7346,N_7174,N_7169);
or U7347 (N_7347,N_7198,N_7179);
xor U7348 (N_7348,N_7081,N_7197);
nor U7349 (N_7349,N_7099,N_7151);
nor U7350 (N_7350,N_7252,N_7327);
or U7351 (N_7351,N_7235,N_7322);
xor U7352 (N_7352,N_7310,N_7332);
and U7353 (N_7353,N_7244,N_7298);
and U7354 (N_7354,N_7204,N_7299);
nor U7355 (N_7355,N_7296,N_7214);
nor U7356 (N_7356,N_7262,N_7219);
or U7357 (N_7357,N_7254,N_7344);
nor U7358 (N_7358,N_7209,N_7256);
or U7359 (N_7359,N_7314,N_7258);
or U7360 (N_7360,N_7265,N_7257);
and U7361 (N_7361,N_7281,N_7249);
xor U7362 (N_7362,N_7291,N_7269);
xnor U7363 (N_7363,N_7305,N_7294);
and U7364 (N_7364,N_7241,N_7231);
and U7365 (N_7365,N_7284,N_7286);
nand U7366 (N_7366,N_7227,N_7316);
or U7367 (N_7367,N_7331,N_7321);
nor U7368 (N_7368,N_7230,N_7273);
nand U7369 (N_7369,N_7211,N_7279);
xor U7370 (N_7370,N_7313,N_7271);
and U7371 (N_7371,N_7290,N_7213);
nor U7372 (N_7372,N_7307,N_7232);
nand U7373 (N_7373,N_7222,N_7226);
or U7374 (N_7374,N_7240,N_7205);
and U7375 (N_7375,N_7301,N_7207);
nor U7376 (N_7376,N_7287,N_7263);
and U7377 (N_7377,N_7323,N_7308);
or U7378 (N_7378,N_7297,N_7234);
xnor U7379 (N_7379,N_7339,N_7202);
or U7380 (N_7380,N_7251,N_7300);
and U7381 (N_7381,N_7245,N_7319);
nor U7382 (N_7382,N_7318,N_7325);
and U7383 (N_7383,N_7340,N_7336);
nor U7384 (N_7384,N_7276,N_7341);
xnor U7385 (N_7385,N_7277,N_7218);
nor U7386 (N_7386,N_7280,N_7312);
or U7387 (N_7387,N_7225,N_7302);
nand U7388 (N_7388,N_7224,N_7238);
nor U7389 (N_7389,N_7348,N_7223);
nor U7390 (N_7390,N_7282,N_7229);
or U7391 (N_7391,N_7216,N_7255);
and U7392 (N_7392,N_7259,N_7288);
and U7393 (N_7393,N_7333,N_7320);
and U7394 (N_7394,N_7261,N_7309);
nand U7395 (N_7395,N_7346,N_7289);
or U7396 (N_7396,N_7347,N_7275);
and U7397 (N_7397,N_7342,N_7317);
nand U7398 (N_7398,N_7349,N_7250);
nand U7399 (N_7399,N_7233,N_7212);
and U7400 (N_7400,N_7266,N_7338);
and U7401 (N_7401,N_7330,N_7303);
nand U7402 (N_7402,N_7334,N_7345);
nand U7403 (N_7403,N_7278,N_7208);
nand U7404 (N_7404,N_7228,N_7237);
xor U7405 (N_7405,N_7328,N_7206);
nor U7406 (N_7406,N_7201,N_7203);
nand U7407 (N_7407,N_7293,N_7215);
nand U7408 (N_7408,N_7220,N_7200);
nand U7409 (N_7409,N_7264,N_7335);
nor U7410 (N_7410,N_7217,N_7274);
xor U7411 (N_7411,N_7304,N_7295);
nor U7412 (N_7412,N_7248,N_7292);
or U7413 (N_7413,N_7343,N_7270);
nand U7414 (N_7414,N_7324,N_7329);
xnor U7415 (N_7415,N_7315,N_7337);
or U7416 (N_7416,N_7260,N_7242);
nor U7417 (N_7417,N_7236,N_7285);
nor U7418 (N_7418,N_7247,N_7210);
xor U7419 (N_7419,N_7311,N_7243);
and U7420 (N_7420,N_7326,N_7221);
and U7421 (N_7421,N_7272,N_7253);
and U7422 (N_7422,N_7306,N_7267);
and U7423 (N_7423,N_7239,N_7246);
nand U7424 (N_7424,N_7283,N_7268);
nor U7425 (N_7425,N_7241,N_7270);
and U7426 (N_7426,N_7247,N_7244);
nor U7427 (N_7427,N_7230,N_7339);
xnor U7428 (N_7428,N_7303,N_7267);
and U7429 (N_7429,N_7284,N_7202);
xor U7430 (N_7430,N_7272,N_7330);
or U7431 (N_7431,N_7205,N_7254);
and U7432 (N_7432,N_7343,N_7289);
or U7433 (N_7433,N_7260,N_7312);
or U7434 (N_7434,N_7227,N_7344);
and U7435 (N_7435,N_7229,N_7233);
xnor U7436 (N_7436,N_7245,N_7327);
and U7437 (N_7437,N_7323,N_7332);
nand U7438 (N_7438,N_7300,N_7341);
nor U7439 (N_7439,N_7318,N_7252);
nand U7440 (N_7440,N_7343,N_7272);
nand U7441 (N_7441,N_7323,N_7241);
xnor U7442 (N_7442,N_7207,N_7204);
nand U7443 (N_7443,N_7237,N_7221);
nand U7444 (N_7444,N_7211,N_7201);
nand U7445 (N_7445,N_7306,N_7316);
and U7446 (N_7446,N_7246,N_7203);
nand U7447 (N_7447,N_7233,N_7210);
xnor U7448 (N_7448,N_7212,N_7294);
and U7449 (N_7449,N_7256,N_7219);
or U7450 (N_7450,N_7204,N_7210);
nand U7451 (N_7451,N_7253,N_7277);
and U7452 (N_7452,N_7287,N_7255);
nand U7453 (N_7453,N_7344,N_7339);
or U7454 (N_7454,N_7240,N_7317);
nor U7455 (N_7455,N_7335,N_7228);
and U7456 (N_7456,N_7255,N_7200);
or U7457 (N_7457,N_7303,N_7286);
and U7458 (N_7458,N_7308,N_7318);
or U7459 (N_7459,N_7264,N_7299);
nor U7460 (N_7460,N_7276,N_7271);
or U7461 (N_7461,N_7309,N_7241);
or U7462 (N_7462,N_7223,N_7237);
nor U7463 (N_7463,N_7345,N_7206);
xnor U7464 (N_7464,N_7340,N_7264);
nand U7465 (N_7465,N_7281,N_7245);
nor U7466 (N_7466,N_7261,N_7336);
and U7467 (N_7467,N_7248,N_7346);
nor U7468 (N_7468,N_7280,N_7265);
and U7469 (N_7469,N_7254,N_7340);
and U7470 (N_7470,N_7214,N_7331);
nor U7471 (N_7471,N_7276,N_7220);
nor U7472 (N_7472,N_7349,N_7297);
and U7473 (N_7473,N_7258,N_7268);
and U7474 (N_7474,N_7271,N_7344);
nand U7475 (N_7475,N_7242,N_7214);
and U7476 (N_7476,N_7236,N_7277);
or U7477 (N_7477,N_7276,N_7206);
or U7478 (N_7478,N_7224,N_7318);
or U7479 (N_7479,N_7295,N_7229);
nor U7480 (N_7480,N_7205,N_7325);
or U7481 (N_7481,N_7329,N_7261);
and U7482 (N_7482,N_7259,N_7251);
and U7483 (N_7483,N_7252,N_7322);
or U7484 (N_7484,N_7222,N_7225);
nor U7485 (N_7485,N_7230,N_7340);
nor U7486 (N_7486,N_7320,N_7268);
nand U7487 (N_7487,N_7262,N_7247);
xnor U7488 (N_7488,N_7310,N_7349);
xor U7489 (N_7489,N_7316,N_7347);
or U7490 (N_7490,N_7215,N_7255);
nand U7491 (N_7491,N_7282,N_7312);
xor U7492 (N_7492,N_7264,N_7305);
xnor U7493 (N_7493,N_7283,N_7308);
xor U7494 (N_7494,N_7224,N_7210);
nor U7495 (N_7495,N_7251,N_7262);
nor U7496 (N_7496,N_7281,N_7349);
xor U7497 (N_7497,N_7305,N_7332);
nand U7498 (N_7498,N_7297,N_7294);
xor U7499 (N_7499,N_7265,N_7222);
and U7500 (N_7500,N_7415,N_7475);
and U7501 (N_7501,N_7390,N_7468);
nor U7502 (N_7502,N_7466,N_7479);
and U7503 (N_7503,N_7464,N_7383);
nand U7504 (N_7504,N_7477,N_7350);
or U7505 (N_7505,N_7355,N_7451);
nand U7506 (N_7506,N_7362,N_7412);
and U7507 (N_7507,N_7419,N_7432);
or U7508 (N_7508,N_7483,N_7397);
nand U7509 (N_7509,N_7378,N_7457);
nand U7510 (N_7510,N_7495,N_7373);
xor U7511 (N_7511,N_7365,N_7394);
or U7512 (N_7512,N_7381,N_7488);
or U7513 (N_7513,N_7399,N_7380);
and U7514 (N_7514,N_7492,N_7471);
and U7515 (N_7515,N_7461,N_7361);
xor U7516 (N_7516,N_7452,N_7444);
nand U7517 (N_7517,N_7489,N_7474);
xnor U7518 (N_7518,N_7443,N_7476);
nand U7519 (N_7519,N_7429,N_7369);
nand U7520 (N_7520,N_7408,N_7382);
xnor U7521 (N_7521,N_7482,N_7422);
and U7522 (N_7522,N_7391,N_7487);
or U7523 (N_7523,N_7363,N_7438);
nand U7524 (N_7524,N_7354,N_7371);
nor U7525 (N_7525,N_7403,N_7370);
nand U7526 (N_7526,N_7486,N_7480);
or U7527 (N_7527,N_7435,N_7442);
nor U7528 (N_7528,N_7449,N_7459);
or U7529 (N_7529,N_7469,N_7379);
nor U7530 (N_7530,N_7454,N_7446);
nand U7531 (N_7531,N_7406,N_7426);
nor U7532 (N_7532,N_7404,N_7409);
nor U7533 (N_7533,N_7472,N_7490);
nor U7534 (N_7534,N_7400,N_7470);
or U7535 (N_7535,N_7401,N_7440);
or U7536 (N_7536,N_7389,N_7387);
or U7537 (N_7537,N_7456,N_7356);
or U7538 (N_7538,N_7427,N_7374);
xnor U7539 (N_7539,N_7467,N_7499);
and U7540 (N_7540,N_7364,N_7455);
and U7541 (N_7541,N_7441,N_7413);
nor U7542 (N_7542,N_7491,N_7386);
and U7543 (N_7543,N_7392,N_7463);
xor U7544 (N_7544,N_7393,N_7385);
nand U7545 (N_7545,N_7496,N_7367);
or U7546 (N_7546,N_7424,N_7377);
nor U7547 (N_7547,N_7410,N_7416);
or U7548 (N_7548,N_7458,N_7351);
nand U7549 (N_7549,N_7448,N_7436);
and U7550 (N_7550,N_7425,N_7497);
xnor U7551 (N_7551,N_7376,N_7494);
nor U7552 (N_7552,N_7433,N_7420);
nand U7553 (N_7553,N_7360,N_7450);
or U7554 (N_7554,N_7421,N_7366);
nor U7555 (N_7555,N_7430,N_7359);
nand U7556 (N_7556,N_7453,N_7437);
nor U7557 (N_7557,N_7352,N_7473);
nor U7558 (N_7558,N_7417,N_7407);
nand U7559 (N_7559,N_7445,N_7388);
and U7560 (N_7560,N_7398,N_7414);
and U7561 (N_7561,N_7358,N_7478);
nand U7562 (N_7562,N_7396,N_7353);
xor U7563 (N_7563,N_7384,N_7481);
nor U7564 (N_7564,N_7462,N_7428);
nand U7565 (N_7565,N_7485,N_7418);
or U7566 (N_7566,N_7372,N_7357);
nor U7567 (N_7567,N_7395,N_7439);
and U7568 (N_7568,N_7402,N_7423);
xnor U7569 (N_7569,N_7484,N_7434);
and U7570 (N_7570,N_7447,N_7405);
and U7571 (N_7571,N_7411,N_7431);
nor U7572 (N_7572,N_7498,N_7493);
xor U7573 (N_7573,N_7465,N_7460);
nor U7574 (N_7574,N_7375,N_7368);
and U7575 (N_7575,N_7375,N_7377);
xnor U7576 (N_7576,N_7487,N_7383);
and U7577 (N_7577,N_7388,N_7352);
xor U7578 (N_7578,N_7355,N_7391);
xnor U7579 (N_7579,N_7424,N_7459);
or U7580 (N_7580,N_7494,N_7364);
or U7581 (N_7581,N_7492,N_7396);
nand U7582 (N_7582,N_7486,N_7471);
nand U7583 (N_7583,N_7490,N_7365);
nand U7584 (N_7584,N_7407,N_7420);
or U7585 (N_7585,N_7420,N_7357);
or U7586 (N_7586,N_7461,N_7364);
xor U7587 (N_7587,N_7474,N_7393);
and U7588 (N_7588,N_7390,N_7382);
xnor U7589 (N_7589,N_7482,N_7364);
xor U7590 (N_7590,N_7477,N_7368);
xor U7591 (N_7591,N_7418,N_7478);
nand U7592 (N_7592,N_7471,N_7433);
nand U7593 (N_7593,N_7430,N_7474);
nor U7594 (N_7594,N_7369,N_7421);
or U7595 (N_7595,N_7365,N_7450);
nand U7596 (N_7596,N_7391,N_7362);
nand U7597 (N_7597,N_7364,N_7477);
or U7598 (N_7598,N_7364,N_7450);
or U7599 (N_7599,N_7371,N_7476);
and U7600 (N_7600,N_7410,N_7411);
nor U7601 (N_7601,N_7492,N_7359);
and U7602 (N_7602,N_7457,N_7381);
nand U7603 (N_7603,N_7454,N_7362);
and U7604 (N_7604,N_7382,N_7484);
and U7605 (N_7605,N_7405,N_7432);
nor U7606 (N_7606,N_7481,N_7439);
xor U7607 (N_7607,N_7377,N_7416);
nor U7608 (N_7608,N_7419,N_7490);
nand U7609 (N_7609,N_7460,N_7386);
xnor U7610 (N_7610,N_7397,N_7430);
nand U7611 (N_7611,N_7387,N_7437);
xor U7612 (N_7612,N_7447,N_7470);
or U7613 (N_7613,N_7395,N_7415);
nand U7614 (N_7614,N_7371,N_7418);
nand U7615 (N_7615,N_7446,N_7370);
nand U7616 (N_7616,N_7357,N_7356);
or U7617 (N_7617,N_7409,N_7455);
or U7618 (N_7618,N_7410,N_7390);
xor U7619 (N_7619,N_7422,N_7351);
or U7620 (N_7620,N_7449,N_7443);
or U7621 (N_7621,N_7365,N_7494);
nor U7622 (N_7622,N_7457,N_7352);
xor U7623 (N_7623,N_7383,N_7363);
xor U7624 (N_7624,N_7440,N_7459);
nand U7625 (N_7625,N_7378,N_7384);
xor U7626 (N_7626,N_7411,N_7361);
xor U7627 (N_7627,N_7474,N_7408);
nor U7628 (N_7628,N_7474,N_7365);
or U7629 (N_7629,N_7481,N_7350);
xor U7630 (N_7630,N_7390,N_7388);
xor U7631 (N_7631,N_7486,N_7419);
nor U7632 (N_7632,N_7486,N_7401);
nand U7633 (N_7633,N_7364,N_7457);
or U7634 (N_7634,N_7495,N_7365);
nand U7635 (N_7635,N_7360,N_7392);
nand U7636 (N_7636,N_7481,N_7462);
and U7637 (N_7637,N_7434,N_7460);
nor U7638 (N_7638,N_7494,N_7423);
nor U7639 (N_7639,N_7375,N_7370);
nor U7640 (N_7640,N_7452,N_7407);
and U7641 (N_7641,N_7478,N_7360);
nand U7642 (N_7642,N_7351,N_7480);
nor U7643 (N_7643,N_7496,N_7381);
nor U7644 (N_7644,N_7419,N_7395);
nand U7645 (N_7645,N_7485,N_7471);
xnor U7646 (N_7646,N_7423,N_7490);
or U7647 (N_7647,N_7468,N_7479);
nand U7648 (N_7648,N_7411,N_7481);
xor U7649 (N_7649,N_7422,N_7452);
or U7650 (N_7650,N_7503,N_7583);
nand U7651 (N_7651,N_7605,N_7531);
nand U7652 (N_7652,N_7540,N_7563);
or U7653 (N_7653,N_7569,N_7608);
nand U7654 (N_7654,N_7595,N_7534);
and U7655 (N_7655,N_7527,N_7588);
xnor U7656 (N_7656,N_7579,N_7623);
or U7657 (N_7657,N_7501,N_7602);
or U7658 (N_7658,N_7573,N_7541);
or U7659 (N_7659,N_7613,N_7636);
xor U7660 (N_7660,N_7559,N_7631);
or U7661 (N_7661,N_7598,N_7548);
nand U7662 (N_7662,N_7626,N_7571);
nand U7663 (N_7663,N_7622,N_7627);
xor U7664 (N_7664,N_7582,N_7547);
nand U7665 (N_7665,N_7610,N_7513);
and U7666 (N_7666,N_7643,N_7648);
nand U7667 (N_7667,N_7632,N_7630);
nand U7668 (N_7668,N_7570,N_7511);
nor U7669 (N_7669,N_7526,N_7586);
nor U7670 (N_7670,N_7624,N_7596);
nor U7671 (N_7671,N_7521,N_7529);
or U7672 (N_7672,N_7616,N_7600);
or U7673 (N_7673,N_7519,N_7647);
or U7674 (N_7674,N_7502,N_7543);
or U7675 (N_7675,N_7614,N_7590);
nor U7676 (N_7676,N_7620,N_7536);
nor U7677 (N_7677,N_7532,N_7589);
nand U7678 (N_7678,N_7615,N_7642);
nand U7679 (N_7679,N_7607,N_7506);
nor U7680 (N_7680,N_7567,N_7507);
or U7681 (N_7681,N_7585,N_7515);
nand U7682 (N_7682,N_7558,N_7524);
nand U7683 (N_7683,N_7522,N_7584);
nand U7684 (N_7684,N_7617,N_7562);
xor U7685 (N_7685,N_7634,N_7649);
and U7686 (N_7686,N_7603,N_7645);
nor U7687 (N_7687,N_7518,N_7560);
and U7688 (N_7688,N_7504,N_7564);
and U7689 (N_7689,N_7509,N_7594);
nor U7690 (N_7690,N_7606,N_7619);
xor U7691 (N_7691,N_7572,N_7565);
and U7692 (N_7692,N_7554,N_7539);
xnor U7693 (N_7693,N_7574,N_7508);
xor U7694 (N_7694,N_7530,N_7593);
and U7695 (N_7695,N_7581,N_7629);
or U7696 (N_7696,N_7546,N_7500);
and U7697 (N_7697,N_7555,N_7510);
xor U7698 (N_7698,N_7646,N_7621);
and U7699 (N_7699,N_7538,N_7523);
nand U7700 (N_7700,N_7633,N_7577);
xnor U7701 (N_7701,N_7575,N_7551);
xnor U7702 (N_7702,N_7552,N_7641);
nor U7703 (N_7703,N_7612,N_7604);
xor U7704 (N_7704,N_7640,N_7580);
nand U7705 (N_7705,N_7639,N_7635);
or U7706 (N_7706,N_7517,N_7514);
xnor U7707 (N_7707,N_7644,N_7637);
xnor U7708 (N_7708,N_7609,N_7533);
xor U7709 (N_7709,N_7587,N_7528);
or U7710 (N_7710,N_7525,N_7553);
or U7711 (N_7711,N_7578,N_7599);
or U7712 (N_7712,N_7542,N_7545);
xor U7713 (N_7713,N_7516,N_7520);
xnor U7714 (N_7714,N_7537,N_7544);
or U7715 (N_7715,N_7556,N_7557);
nand U7716 (N_7716,N_7591,N_7638);
xnor U7717 (N_7717,N_7566,N_7505);
nor U7718 (N_7718,N_7618,N_7549);
or U7719 (N_7719,N_7568,N_7597);
xnor U7720 (N_7720,N_7611,N_7535);
or U7721 (N_7721,N_7601,N_7512);
nor U7722 (N_7722,N_7628,N_7576);
or U7723 (N_7723,N_7592,N_7550);
or U7724 (N_7724,N_7561,N_7625);
xnor U7725 (N_7725,N_7527,N_7590);
nand U7726 (N_7726,N_7507,N_7607);
nand U7727 (N_7727,N_7597,N_7554);
or U7728 (N_7728,N_7636,N_7642);
nor U7729 (N_7729,N_7603,N_7622);
or U7730 (N_7730,N_7502,N_7542);
nand U7731 (N_7731,N_7534,N_7524);
and U7732 (N_7732,N_7508,N_7579);
nor U7733 (N_7733,N_7507,N_7531);
nand U7734 (N_7734,N_7503,N_7510);
xor U7735 (N_7735,N_7592,N_7566);
nand U7736 (N_7736,N_7628,N_7590);
nand U7737 (N_7737,N_7641,N_7583);
or U7738 (N_7738,N_7609,N_7630);
or U7739 (N_7739,N_7596,N_7511);
nor U7740 (N_7740,N_7600,N_7554);
and U7741 (N_7741,N_7592,N_7610);
nor U7742 (N_7742,N_7614,N_7552);
nand U7743 (N_7743,N_7514,N_7582);
nand U7744 (N_7744,N_7619,N_7594);
xor U7745 (N_7745,N_7500,N_7604);
nand U7746 (N_7746,N_7610,N_7593);
nor U7747 (N_7747,N_7583,N_7593);
xor U7748 (N_7748,N_7601,N_7629);
or U7749 (N_7749,N_7552,N_7603);
xor U7750 (N_7750,N_7606,N_7610);
nand U7751 (N_7751,N_7571,N_7606);
and U7752 (N_7752,N_7611,N_7583);
nand U7753 (N_7753,N_7528,N_7621);
nand U7754 (N_7754,N_7636,N_7532);
nor U7755 (N_7755,N_7610,N_7519);
and U7756 (N_7756,N_7551,N_7565);
nand U7757 (N_7757,N_7553,N_7579);
nor U7758 (N_7758,N_7599,N_7502);
or U7759 (N_7759,N_7507,N_7637);
nand U7760 (N_7760,N_7501,N_7500);
nand U7761 (N_7761,N_7546,N_7518);
nor U7762 (N_7762,N_7570,N_7587);
and U7763 (N_7763,N_7537,N_7628);
xor U7764 (N_7764,N_7611,N_7617);
and U7765 (N_7765,N_7543,N_7557);
nand U7766 (N_7766,N_7645,N_7629);
nor U7767 (N_7767,N_7538,N_7611);
nand U7768 (N_7768,N_7646,N_7594);
xnor U7769 (N_7769,N_7569,N_7560);
or U7770 (N_7770,N_7526,N_7536);
nor U7771 (N_7771,N_7544,N_7644);
xnor U7772 (N_7772,N_7633,N_7547);
xor U7773 (N_7773,N_7515,N_7580);
or U7774 (N_7774,N_7521,N_7579);
nand U7775 (N_7775,N_7633,N_7623);
and U7776 (N_7776,N_7624,N_7564);
and U7777 (N_7777,N_7553,N_7633);
nor U7778 (N_7778,N_7582,N_7585);
nor U7779 (N_7779,N_7509,N_7634);
xnor U7780 (N_7780,N_7583,N_7510);
xor U7781 (N_7781,N_7582,N_7596);
xor U7782 (N_7782,N_7622,N_7512);
nand U7783 (N_7783,N_7529,N_7540);
and U7784 (N_7784,N_7607,N_7583);
nor U7785 (N_7785,N_7574,N_7525);
xor U7786 (N_7786,N_7530,N_7592);
and U7787 (N_7787,N_7618,N_7577);
or U7788 (N_7788,N_7618,N_7524);
xnor U7789 (N_7789,N_7541,N_7574);
or U7790 (N_7790,N_7574,N_7623);
and U7791 (N_7791,N_7502,N_7608);
nand U7792 (N_7792,N_7615,N_7500);
nand U7793 (N_7793,N_7507,N_7603);
nor U7794 (N_7794,N_7616,N_7549);
xnor U7795 (N_7795,N_7577,N_7630);
nand U7796 (N_7796,N_7636,N_7544);
and U7797 (N_7797,N_7639,N_7536);
nand U7798 (N_7798,N_7578,N_7627);
nand U7799 (N_7799,N_7577,N_7524);
and U7800 (N_7800,N_7770,N_7786);
nor U7801 (N_7801,N_7772,N_7737);
nor U7802 (N_7802,N_7653,N_7747);
xnor U7803 (N_7803,N_7743,N_7736);
xnor U7804 (N_7804,N_7721,N_7700);
nor U7805 (N_7805,N_7680,N_7757);
nand U7806 (N_7806,N_7795,N_7776);
nor U7807 (N_7807,N_7669,N_7725);
or U7808 (N_7808,N_7759,N_7753);
and U7809 (N_7809,N_7738,N_7752);
and U7810 (N_7810,N_7662,N_7663);
nor U7811 (N_7811,N_7667,N_7788);
nand U7812 (N_7812,N_7657,N_7785);
nor U7813 (N_7813,N_7792,N_7678);
or U7814 (N_7814,N_7712,N_7664);
and U7815 (N_7815,N_7754,N_7748);
or U7816 (N_7816,N_7793,N_7665);
and U7817 (N_7817,N_7787,N_7727);
or U7818 (N_7818,N_7742,N_7693);
nand U7819 (N_7819,N_7778,N_7760);
nand U7820 (N_7820,N_7791,N_7782);
or U7821 (N_7821,N_7659,N_7698);
xor U7822 (N_7822,N_7689,N_7767);
or U7823 (N_7823,N_7658,N_7673);
xor U7824 (N_7824,N_7694,N_7774);
or U7825 (N_7825,N_7696,N_7728);
and U7826 (N_7826,N_7714,N_7756);
xnor U7827 (N_7827,N_7740,N_7686);
nor U7828 (N_7828,N_7764,N_7724);
or U7829 (N_7829,N_7726,N_7773);
nor U7830 (N_7830,N_7668,N_7682);
nor U7831 (N_7831,N_7794,N_7706);
nand U7832 (N_7832,N_7703,N_7710);
nor U7833 (N_7833,N_7719,N_7779);
or U7834 (N_7834,N_7715,N_7711);
and U7835 (N_7835,N_7758,N_7656);
or U7836 (N_7836,N_7708,N_7704);
or U7837 (N_7837,N_7730,N_7799);
and U7838 (N_7838,N_7707,N_7797);
and U7839 (N_7839,N_7745,N_7765);
nor U7840 (N_7840,N_7702,N_7784);
and U7841 (N_7841,N_7798,N_7697);
and U7842 (N_7842,N_7681,N_7762);
nor U7843 (N_7843,N_7683,N_7709);
nor U7844 (N_7844,N_7685,N_7763);
and U7845 (N_7845,N_7691,N_7671);
or U7846 (N_7846,N_7781,N_7679);
xnor U7847 (N_7847,N_7699,N_7768);
nand U7848 (N_7848,N_7729,N_7705);
nand U7849 (N_7849,N_7718,N_7790);
and U7850 (N_7850,N_7670,N_7723);
or U7851 (N_7851,N_7720,N_7750);
nand U7852 (N_7852,N_7695,N_7660);
nand U7853 (N_7853,N_7735,N_7684);
and U7854 (N_7854,N_7655,N_7677);
nor U7855 (N_7855,N_7746,N_7741);
or U7856 (N_7856,N_7651,N_7716);
nand U7857 (N_7857,N_7789,N_7796);
nor U7858 (N_7858,N_7701,N_7755);
or U7859 (N_7859,N_7713,N_7666);
or U7860 (N_7860,N_7688,N_7780);
nor U7861 (N_7861,N_7734,N_7687);
and U7862 (N_7862,N_7732,N_7777);
nor U7863 (N_7863,N_7717,N_7775);
nand U7864 (N_7864,N_7749,N_7771);
nand U7865 (N_7865,N_7769,N_7733);
nor U7866 (N_7866,N_7650,N_7739);
or U7867 (N_7867,N_7761,N_7652);
or U7868 (N_7868,N_7722,N_7751);
or U7869 (N_7869,N_7766,N_7692);
nand U7870 (N_7870,N_7654,N_7690);
and U7871 (N_7871,N_7672,N_7744);
nor U7872 (N_7872,N_7661,N_7731);
and U7873 (N_7873,N_7783,N_7676);
and U7874 (N_7874,N_7675,N_7674);
xnor U7875 (N_7875,N_7799,N_7724);
nor U7876 (N_7876,N_7718,N_7787);
nand U7877 (N_7877,N_7770,N_7684);
and U7878 (N_7878,N_7705,N_7717);
or U7879 (N_7879,N_7780,N_7657);
nor U7880 (N_7880,N_7769,N_7682);
nor U7881 (N_7881,N_7682,N_7775);
nand U7882 (N_7882,N_7688,N_7710);
or U7883 (N_7883,N_7673,N_7729);
nand U7884 (N_7884,N_7669,N_7723);
xnor U7885 (N_7885,N_7760,N_7694);
or U7886 (N_7886,N_7686,N_7752);
nand U7887 (N_7887,N_7780,N_7721);
nor U7888 (N_7888,N_7790,N_7709);
or U7889 (N_7889,N_7662,N_7664);
nor U7890 (N_7890,N_7747,N_7750);
nand U7891 (N_7891,N_7683,N_7704);
nand U7892 (N_7892,N_7755,N_7737);
nor U7893 (N_7893,N_7663,N_7691);
xnor U7894 (N_7894,N_7695,N_7721);
nor U7895 (N_7895,N_7680,N_7793);
nand U7896 (N_7896,N_7794,N_7656);
or U7897 (N_7897,N_7718,N_7710);
xnor U7898 (N_7898,N_7760,N_7650);
and U7899 (N_7899,N_7741,N_7728);
nor U7900 (N_7900,N_7773,N_7682);
and U7901 (N_7901,N_7651,N_7686);
and U7902 (N_7902,N_7756,N_7785);
and U7903 (N_7903,N_7654,N_7688);
nor U7904 (N_7904,N_7698,N_7755);
or U7905 (N_7905,N_7753,N_7711);
nand U7906 (N_7906,N_7770,N_7771);
nor U7907 (N_7907,N_7781,N_7759);
nor U7908 (N_7908,N_7782,N_7727);
and U7909 (N_7909,N_7705,N_7727);
and U7910 (N_7910,N_7795,N_7676);
nand U7911 (N_7911,N_7760,N_7739);
nor U7912 (N_7912,N_7760,N_7696);
nor U7913 (N_7913,N_7734,N_7779);
nand U7914 (N_7914,N_7727,N_7682);
xnor U7915 (N_7915,N_7687,N_7763);
nor U7916 (N_7916,N_7790,N_7758);
or U7917 (N_7917,N_7737,N_7757);
and U7918 (N_7918,N_7709,N_7785);
nand U7919 (N_7919,N_7724,N_7784);
or U7920 (N_7920,N_7656,N_7796);
nor U7921 (N_7921,N_7684,N_7707);
or U7922 (N_7922,N_7672,N_7794);
xnor U7923 (N_7923,N_7673,N_7706);
nor U7924 (N_7924,N_7750,N_7651);
xor U7925 (N_7925,N_7667,N_7733);
xor U7926 (N_7926,N_7765,N_7717);
nand U7927 (N_7927,N_7657,N_7670);
nor U7928 (N_7928,N_7754,N_7682);
nor U7929 (N_7929,N_7789,N_7711);
xnor U7930 (N_7930,N_7711,N_7723);
xnor U7931 (N_7931,N_7678,N_7764);
nor U7932 (N_7932,N_7690,N_7749);
nor U7933 (N_7933,N_7766,N_7674);
xor U7934 (N_7934,N_7790,N_7724);
xnor U7935 (N_7935,N_7726,N_7729);
xor U7936 (N_7936,N_7654,N_7793);
or U7937 (N_7937,N_7722,N_7763);
and U7938 (N_7938,N_7728,N_7737);
nor U7939 (N_7939,N_7708,N_7779);
xor U7940 (N_7940,N_7651,N_7742);
or U7941 (N_7941,N_7657,N_7759);
nor U7942 (N_7942,N_7650,N_7700);
nor U7943 (N_7943,N_7720,N_7744);
nor U7944 (N_7944,N_7751,N_7793);
and U7945 (N_7945,N_7791,N_7672);
nor U7946 (N_7946,N_7685,N_7673);
xor U7947 (N_7947,N_7667,N_7732);
nor U7948 (N_7948,N_7657,N_7754);
nand U7949 (N_7949,N_7776,N_7721);
and U7950 (N_7950,N_7805,N_7812);
nor U7951 (N_7951,N_7853,N_7926);
xor U7952 (N_7952,N_7806,N_7923);
nor U7953 (N_7953,N_7901,N_7931);
xor U7954 (N_7954,N_7819,N_7838);
nor U7955 (N_7955,N_7854,N_7811);
xor U7956 (N_7956,N_7884,N_7908);
xnor U7957 (N_7957,N_7914,N_7847);
or U7958 (N_7958,N_7810,N_7862);
xnor U7959 (N_7959,N_7915,N_7904);
or U7960 (N_7960,N_7876,N_7872);
nor U7961 (N_7961,N_7868,N_7946);
and U7962 (N_7962,N_7928,N_7800);
nand U7963 (N_7963,N_7940,N_7834);
nor U7964 (N_7964,N_7911,N_7947);
or U7965 (N_7965,N_7942,N_7830);
or U7966 (N_7966,N_7860,N_7945);
nand U7967 (N_7967,N_7867,N_7903);
nand U7968 (N_7968,N_7845,N_7827);
nor U7969 (N_7969,N_7822,N_7803);
nor U7970 (N_7970,N_7818,N_7918);
nand U7971 (N_7971,N_7930,N_7839);
or U7972 (N_7972,N_7837,N_7916);
or U7973 (N_7973,N_7869,N_7873);
or U7974 (N_7974,N_7937,N_7932);
nor U7975 (N_7975,N_7922,N_7870);
nor U7976 (N_7976,N_7897,N_7927);
or U7977 (N_7977,N_7949,N_7823);
nor U7978 (N_7978,N_7887,N_7809);
nor U7979 (N_7979,N_7841,N_7816);
or U7980 (N_7980,N_7885,N_7815);
nor U7981 (N_7981,N_7848,N_7859);
nand U7982 (N_7982,N_7829,N_7935);
and U7983 (N_7983,N_7943,N_7813);
xnor U7984 (N_7984,N_7910,N_7886);
or U7985 (N_7985,N_7907,N_7857);
xnor U7986 (N_7986,N_7936,N_7856);
or U7987 (N_7987,N_7880,N_7902);
nand U7988 (N_7988,N_7894,N_7891);
or U7989 (N_7989,N_7808,N_7882);
nand U7990 (N_7990,N_7896,N_7900);
xnor U7991 (N_7991,N_7804,N_7846);
or U7992 (N_7992,N_7840,N_7826);
nand U7993 (N_7993,N_7919,N_7835);
xor U7994 (N_7994,N_7821,N_7874);
xnor U7995 (N_7995,N_7842,N_7920);
xor U7996 (N_7996,N_7858,N_7801);
nor U7997 (N_7997,N_7906,N_7844);
nor U7998 (N_7998,N_7917,N_7939);
or U7999 (N_7999,N_7893,N_7913);
and U8000 (N_8000,N_7929,N_7881);
and U8001 (N_8001,N_7888,N_7851);
xor U8002 (N_8002,N_7820,N_7934);
and U8003 (N_8003,N_7875,N_7899);
xnor U8004 (N_8004,N_7852,N_7817);
or U8005 (N_8005,N_7824,N_7912);
and U8006 (N_8006,N_7924,N_7865);
xor U8007 (N_8007,N_7944,N_7850);
and U8008 (N_8008,N_7921,N_7828);
xnor U8009 (N_8009,N_7836,N_7807);
and U8010 (N_8010,N_7802,N_7938);
xnor U8011 (N_8011,N_7861,N_7833);
xor U8012 (N_8012,N_7879,N_7898);
or U8013 (N_8013,N_7871,N_7832);
or U8014 (N_8014,N_7905,N_7855);
xnor U8015 (N_8015,N_7814,N_7892);
or U8016 (N_8016,N_7948,N_7889);
xnor U8017 (N_8017,N_7866,N_7925);
nor U8018 (N_8018,N_7895,N_7831);
xnor U8019 (N_8019,N_7863,N_7933);
nor U8020 (N_8020,N_7890,N_7864);
xnor U8021 (N_8021,N_7843,N_7849);
and U8022 (N_8022,N_7878,N_7941);
and U8023 (N_8023,N_7825,N_7883);
nand U8024 (N_8024,N_7877,N_7909);
nor U8025 (N_8025,N_7826,N_7850);
or U8026 (N_8026,N_7896,N_7815);
or U8027 (N_8027,N_7891,N_7802);
xor U8028 (N_8028,N_7833,N_7913);
nor U8029 (N_8029,N_7855,N_7873);
and U8030 (N_8030,N_7813,N_7845);
nand U8031 (N_8031,N_7947,N_7844);
xnor U8032 (N_8032,N_7819,N_7879);
nor U8033 (N_8033,N_7829,N_7825);
nor U8034 (N_8034,N_7878,N_7817);
nor U8035 (N_8035,N_7877,N_7947);
and U8036 (N_8036,N_7935,N_7919);
and U8037 (N_8037,N_7868,N_7943);
xnor U8038 (N_8038,N_7904,N_7808);
or U8039 (N_8039,N_7812,N_7843);
nand U8040 (N_8040,N_7844,N_7853);
xnor U8041 (N_8041,N_7822,N_7877);
nand U8042 (N_8042,N_7867,N_7835);
xnor U8043 (N_8043,N_7817,N_7834);
xor U8044 (N_8044,N_7935,N_7937);
or U8045 (N_8045,N_7868,N_7835);
nand U8046 (N_8046,N_7946,N_7871);
nand U8047 (N_8047,N_7813,N_7818);
nor U8048 (N_8048,N_7869,N_7949);
nand U8049 (N_8049,N_7856,N_7840);
nor U8050 (N_8050,N_7899,N_7932);
nand U8051 (N_8051,N_7881,N_7902);
nor U8052 (N_8052,N_7817,N_7813);
or U8053 (N_8053,N_7885,N_7810);
nor U8054 (N_8054,N_7877,N_7855);
nand U8055 (N_8055,N_7903,N_7904);
nor U8056 (N_8056,N_7921,N_7859);
or U8057 (N_8057,N_7949,N_7891);
nand U8058 (N_8058,N_7861,N_7817);
or U8059 (N_8059,N_7909,N_7893);
nand U8060 (N_8060,N_7904,N_7843);
nand U8061 (N_8061,N_7873,N_7822);
nor U8062 (N_8062,N_7815,N_7804);
nor U8063 (N_8063,N_7903,N_7881);
nor U8064 (N_8064,N_7809,N_7929);
and U8065 (N_8065,N_7935,N_7887);
and U8066 (N_8066,N_7814,N_7807);
xnor U8067 (N_8067,N_7830,N_7844);
nand U8068 (N_8068,N_7823,N_7859);
nand U8069 (N_8069,N_7879,N_7930);
xor U8070 (N_8070,N_7863,N_7921);
and U8071 (N_8071,N_7822,N_7912);
nor U8072 (N_8072,N_7873,N_7868);
or U8073 (N_8073,N_7845,N_7926);
and U8074 (N_8074,N_7855,N_7888);
nor U8075 (N_8075,N_7862,N_7800);
and U8076 (N_8076,N_7899,N_7817);
xnor U8077 (N_8077,N_7889,N_7901);
or U8078 (N_8078,N_7827,N_7880);
nor U8079 (N_8079,N_7906,N_7849);
and U8080 (N_8080,N_7814,N_7908);
nor U8081 (N_8081,N_7936,N_7886);
xnor U8082 (N_8082,N_7819,N_7891);
nor U8083 (N_8083,N_7863,N_7856);
or U8084 (N_8084,N_7808,N_7830);
nand U8085 (N_8085,N_7894,N_7876);
xnor U8086 (N_8086,N_7807,N_7861);
and U8087 (N_8087,N_7925,N_7927);
nand U8088 (N_8088,N_7945,N_7866);
or U8089 (N_8089,N_7945,N_7830);
nor U8090 (N_8090,N_7935,N_7846);
nand U8091 (N_8091,N_7854,N_7932);
nand U8092 (N_8092,N_7821,N_7930);
nor U8093 (N_8093,N_7842,N_7837);
nand U8094 (N_8094,N_7947,N_7818);
and U8095 (N_8095,N_7825,N_7869);
nor U8096 (N_8096,N_7943,N_7927);
or U8097 (N_8097,N_7879,N_7834);
nor U8098 (N_8098,N_7852,N_7906);
and U8099 (N_8099,N_7884,N_7855);
nor U8100 (N_8100,N_8063,N_7976);
xnor U8101 (N_8101,N_7981,N_7994);
or U8102 (N_8102,N_7980,N_8064);
xor U8103 (N_8103,N_7950,N_8025);
and U8104 (N_8104,N_8026,N_8000);
xnor U8105 (N_8105,N_7986,N_8008);
nor U8106 (N_8106,N_7959,N_8076);
xnor U8107 (N_8107,N_8096,N_7993);
and U8108 (N_8108,N_7966,N_8074);
nand U8109 (N_8109,N_8016,N_8067);
nand U8110 (N_8110,N_8011,N_8001);
xor U8111 (N_8111,N_8081,N_7979);
nor U8112 (N_8112,N_7997,N_7961);
or U8113 (N_8113,N_7953,N_8093);
nor U8114 (N_8114,N_7958,N_8044);
and U8115 (N_8115,N_8070,N_8082);
xnor U8116 (N_8116,N_8037,N_8075);
nand U8117 (N_8117,N_8004,N_8003);
xor U8118 (N_8118,N_7974,N_7965);
xnor U8119 (N_8119,N_8041,N_8034);
or U8120 (N_8120,N_8073,N_7954);
nand U8121 (N_8121,N_7985,N_8043);
and U8122 (N_8122,N_8065,N_8014);
or U8123 (N_8123,N_8050,N_7964);
or U8124 (N_8124,N_8053,N_7951);
or U8125 (N_8125,N_8056,N_7978);
or U8126 (N_8126,N_8085,N_8068);
and U8127 (N_8127,N_8078,N_7960);
nand U8128 (N_8128,N_8009,N_8055);
and U8129 (N_8129,N_8042,N_7962);
nand U8130 (N_8130,N_7991,N_8086);
nor U8131 (N_8131,N_8022,N_8094);
nand U8132 (N_8132,N_8005,N_8089);
xnor U8133 (N_8133,N_8028,N_8069);
nor U8134 (N_8134,N_8030,N_7971);
nand U8135 (N_8135,N_8088,N_8020);
and U8136 (N_8136,N_8058,N_8092);
nor U8137 (N_8137,N_7984,N_7998);
and U8138 (N_8138,N_7957,N_8015);
nor U8139 (N_8139,N_7988,N_8035);
or U8140 (N_8140,N_8095,N_7992);
nand U8141 (N_8141,N_8060,N_7989);
xor U8142 (N_8142,N_8047,N_7990);
or U8143 (N_8143,N_7969,N_8019);
and U8144 (N_8144,N_8051,N_8099);
or U8145 (N_8145,N_8066,N_7982);
nor U8146 (N_8146,N_8072,N_7955);
or U8147 (N_8147,N_8087,N_8090);
nor U8148 (N_8148,N_7968,N_7987);
and U8149 (N_8149,N_8079,N_7970);
or U8150 (N_8150,N_8032,N_8038);
nor U8151 (N_8151,N_8007,N_8084);
and U8152 (N_8152,N_8052,N_8040);
nand U8153 (N_8153,N_8021,N_8023);
xnor U8154 (N_8154,N_8061,N_8033);
xor U8155 (N_8155,N_8098,N_8077);
xnor U8156 (N_8156,N_8036,N_8045);
xor U8157 (N_8157,N_8091,N_8062);
nor U8158 (N_8158,N_8049,N_7995);
and U8159 (N_8159,N_8057,N_7963);
xnor U8160 (N_8160,N_8071,N_7983);
xnor U8161 (N_8161,N_7977,N_8018);
nor U8162 (N_8162,N_8046,N_7996);
xnor U8163 (N_8163,N_8024,N_7975);
or U8164 (N_8164,N_8029,N_8027);
or U8165 (N_8165,N_8080,N_8097);
and U8166 (N_8166,N_7952,N_7972);
nand U8167 (N_8167,N_8039,N_8054);
nor U8168 (N_8168,N_8002,N_8031);
or U8169 (N_8169,N_7967,N_8048);
nand U8170 (N_8170,N_8017,N_7999);
or U8171 (N_8171,N_8059,N_8006);
or U8172 (N_8172,N_7956,N_8083);
and U8173 (N_8173,N_8010,N_8013);
or U8174 (N_8174,N_8012,N_7973);
nor U8175 (N_8175,N_8025,N_8076);
xnor U8176 (N_8176,N_7977,N_7956);
or U8177 (N_8177,N_8048,N_8014);
or U8178 (N_8178,N_8014,N_7970);
and U8179 (N_8179,N_8021,N_8038);
xor U8180 (N_8180,N_8025,N_8064);
nor U8181 (N_8181,N_8005,N_8038);
xnor U8182 (N_8182,N_8038,N_7952);
nor U8183 (N_8183,N_8011,N_8002);
or U8184 (N_8184,N_7962,N_8024);
or U8185 (N_8185,N_8034,N_8028);
or U8186 (N_8186,N_7976,N_8060);
nand U8187 (N_8187,N_7967,N_7982);
nor U8188 (N_8188,N_8066,N_7975);
or U8189 (N_8189,N_8090,N_8017);
nor U8190 (N_8190,N_7970,N_8077);
and U8191 (N_8191,N_8002,N_8089);
and U8192 (N_8192,N_7973,N_8011);
nand U8193 (N_8193,N_7981,N_8091);
xor U8194 (N_8194,N_7951,N_8026);
and U8195 (N_8195,N_8034,N_8008);
xor U8196 (N_8196,N_8068,N_8060);
nor U8197 (N_8197,N_8056,N_7971);
nor U8198 (N_8198,N_7955,N_8028);
or U8199 (N_8199,N_8016,N_8055);
nand U8200 (N_8200,N_8035,N_8033);
xnor U8201 (N_8201,N_8080,N_8069);
and U8202 (N_8202,N_7995,N_7958);
nor U8203 (N_8203,N_8039,N_7953);
and U8204 (N_8204,N_8039,N_8083);
nor U8205 (N_8205,N_8060,N_7982);
nor U8206 (N_8206,N_8047,N_8011);
nor U8207 (N_8207,N_7985,N_7992);
xor U8208 (N_8208,N_8080,N_8014);
nand U8209 (N_8209,N_7973,N_8086);
nor U8210 (N_8210,N_7975,N_8063);
or U8211 (N_8211,N_7970,N_7989);
nor U8212 (N_8212,N_7983,N_7956);
nand U8213 (N_8213,N_8026,N_7973);
xor U8214 (N_8214,N_8002,N_7967);
nor U8215 (N_8215,N_7954,N_8022);
nand U8216 (N_8216,N_8099,N_8010);
xor U8217 (N_8217,N_8028,N_8041);
nand U8218 (N_8218,N_8024,N_7955);
and U8219 (N_8219,N_8082,N_7966);
nor U8220 (N_8220,N_8087,N_7994);
xnor U8221 (N_8221,N_8056,N_7992);
or U8222 (N_8222,N_7963,N_8084);
nor U8223 (N_8223,N_8077,N_8044);
nor U8224 (N_8224,N_8041,N_8009);
nor U8225 (N_8225,N_8049,N_8047);
nand U8226 (N_8226,N_8070,N_8052);
nand U8227 (N_8227,N_8009,N_8006);
nor U8228 (N_8228,N_8021,N_7997);
and U8229 (N_8229,N_8062,N_8022);
and U8230 (N_8230,N_8029,N_8002);
xor U8231 (N_8231,N_8072,N_7970);
nand U8232 (N_8232,N_8003,N_8049);
or U8233 (N_8233,N_8049,N_8084);
nor U8234 (N_8234,N_7991,N_8033);
and U8235 (N_8235,N_7962,N_8076);
nor U8236 (N_8236,N_8003,N_8042);
or U8237 (N_8237,N_7983,N_8094);
xnor U8238 (N_8238,N_8017,N_7962);
or U8239 (N_8239,N_8086,N_8061);
nand U8240 (N_8240,N_8011,N_8086);
and U8241 (N_8241,N_7964,N_8099);
xnor U8242 (N_8242,N_8014,N_8040);
and U8243 (N_8243,N_7999,N_7954);
nand U8244 (N_8244,N_8027,N_8086);
xor U8245 (N_8245,N_8003,N_8063);
nand U8246 (N_8246,N_7982,N_8052);
nor U8247 (N_8247,N_8024,N_8089);
xor U8248 (N_8248,N_7962,N_7963);
nor U8249 (N_8249,N_8072,N_7991);
nor U8250 (N_8250,N_8131,N_8124);
nor U8251 (N_8251,N_8141,N_8166);
or U8252 (N_8252,N_8206,N_8103);
xor U8253 (N_8253,N_8165,N_8142);
nor U8254 (N_8254,N_8209,N_8248);
xor U8255 (N_8255,N_8168,N_8227);
or U8256 (N_8256,N_8200,N_8137);
or U8257 (N_8257,N_8205,N_8148);
xor U8258 (N_8258,N_8135,N_8202);
xnor U8259 (N_8259,N_8129,N_8163);
or U8260 (N_8260,N_8228,N_8222);
and U8261 (N_8261,N_8226,N_8212);
or U8262 (N_8262,N_8112,N_8244);
nor U8263 (N_8263,N_8119,N_8145);
nor U8264 (N_8264,N_8171,N_8100);
and U8265 (N_8265,N_8233,N_8246);
xnor U8266 (N_8266,N_8240,N_8109);
xnor U8267 (N_8267,N_8120,N_8185);
or U8268 (N_8268,N_8245,N_8132);
nor U8269 (N_8269,N_8224,N_8211);
or U8270 (N_8270,N_8217,N_8213);
xor U8271 (N_8271,N_8153,N_8161);
nand U8272 (N_8272,N_8218,N_8182);
nor U8273 (N_8273,N_8197,N_8180);
nand U8274 (N_8274,N_8221,N_8116);
xor U8275 (N_8275,N_8101,N_8104);
nor U8276 (N_8276,N_8249,N_8176);
and U8277 (N_8277,N_8239,N_8183);
nand U8278 (N_8278,N_8133,N_8220);
or U8279 (N_8279,N_8177,N_8178);
nand U8280 (N_8280,N_8242,N_8123);
xnor U8281 (N_8281,N_8122,N_8134);
nand U8282 (N_8282,N_8110,N_8146);
nand U8283 (N_8283,N_8238,N_8234);
nand U8284 (N_8284,N_8192,N_8196);
xor U8285 (N_8285,N_8230,N_8179);
or U8286 (N_8286,N_8241,N_8115);
or U8287 (N_8287,N_8154,N_8152);
xnor U8288 (N_8288,N_8199,N_8114);
xnor U8289 (N_8289,N_8243,N_8113);
xor U8290 (N_8290,N_8187,N_8223);
nand U8291 (N_8291,N_8121,N_8125);
and U8292 (N_8292,N_8175,N_8151);
nand U8293 (N_8293,N_8150,N_8147);
and U8294 (N_8294,N_8189,N_8174);
nor U8295 (N_8295,N_8106,N_8105);
xor U8296 (N_8296,N_8158,N_8172);
nor U8297 (N_8297,N_8195,N_8236);
xor U8298 (N_8298,N_8181,N_8235);
or U8299 (N_8299,N_8140,N_8102);
nand U8300 (N_8300,N_8117,N_8231);
nand U8301 (N_8301,N_8215,N_8169);
nand U8302 (N_8302,N_8156,N_8208);
xnor U8303 (N_8303,N_8193,N_8203);
and U8304 (N_8304,N_8162,N_8184);
or U8305 (N_8305,N_8108,N_8186);
or U8306 (N_8306,N_8216,N_8143);
xor U8307 (N_8307,N_8128,N_8130);
nor U8308 (N_8308,N_8107,N_8204);
and U8309 (N_8309,N_8225,N_8194);
and U8310 (N_8310,N_8111,N_8149);
nor U8311 (N_8311,N_8201,N_8219);
xnor U8312 (N_8312,N_8214,N_8191);
xnor U8313 (N_8313,N_8229,N_8118);
nor U8314 (N_8314,N_8173,N_8167);
and U8315 (N_8315,N_8237,N_8139);
nand U8316 (N_8316,N_8159,N_8232);
nor U8317 (N_8317,N_8144,N_8198);
or U8318 (N_8318,N_8188,N_8136);
nand U8319 (N_8319,N_8247,N_8138);
nor U8320 (N_8320,N_8207,N_8155);
or U8321 (N_8321,N_8170,N_8164);
nand U8322 (N_8322,N_8210,N_8190);
nor U8323 (N_8323,N_8126,N_8157);
nor U8324 (N_8324,N_8127,N_8160);
or U8325 (N_8325,N_8221,N_8174);
and U8326 (N_8326,N_8225,N_8226);
nor U8327 (N_8327,N_8183,N_8244);
nand U8328 (N_8328,N_8248,N_8199);
or U8329 (N_8329,N_8147,N_8189);
nand U8330 (N_8330,N_8243,N_8207);
xor U8331 (N_8331,N_8127,N_8179);
nor U8332 (N_8332,N_8147,N_8225);
or U8333 (N_8333,N_8112,N_8212);
xor U8334 (N_8334,N_8205,N_8101);
xor U8335 (N_8335,N_8113,N_8150);
and U8336 (N_8336,N_8198,N_8247);
nand U8337 (N_8337,N_8162,N_8183);
nand U8338 (N_8338,N_8105,N_8220);
nand U8339 (N_8339,N_8116,N_8194);
nor U8340 (N_8340,N_8152,N_8239);
xor U8341 (N_8341,N_8188,N_8181);
xor U8342 (N_8342,N_8210,N_8189);
or U8343 (N_8343,N_8109,N_8147);
or U8344 (N_8344,N_8140,N_8157);
nor U8345 (N_8345,N_8213,N_8122);
xnor U8346 (N_8346,N_8130,N_8132);
nor U8347 (N_8347,N_8214,N_8149);
or U8348 (N_8348,N_8101,N_8125);
nand U8349 (N_8349,N_8176,N_8237);
nor U8350 (N_8350,N_8154,N_8139);
nor U8351 (N_8351,N_8140,N_8136);
nor U8352 (N_8352,N_8180,N_8161);
or U8353 (N_8353,N_8248,N_8208);
or U8354 (N_8354,N_8153,N_8128);
and U8355 (N_8355,N_8219,N_8136);
nor U8356 (N_8356,N_8246,N_8185);
and U8357 (N_8357,N_8167,N_8184);
nand U8358 (N_8358,N_8208,N_8235);
and U8359 (N_8359,N_8143,N_8177);
and U8360 (N_8360,N_8113,N_8147);
nand U8361 (N_8361,N_8248,N_8225);
and U8362 (N_8362,N_8182,N_8107);
xor U8363 (N_8363,N_8210,N_8187);
xor U8364 (N_8364,N_8232,N_8218);
and U8365 (N_8365,N_8199,N_8112);
xnor U8366 (N_8366,N_8108,N_8112);
xor U8367 (N_8367,N_8217,N_8127);
and U8368 (N_8368,N_8113,N_8176);
and U8369 (N_8369,N_8185,N_8174);
and U8370 (N_8370,N_8223,N_8215);
and U8371 (N_8371,N_8242,N_8175);
nor U8372 (N_8372,N_8224,N_8207);
nand U8373 (N_8373,N_8222,N_8216);
xnor U8374 (N_8374,N_8183,N_8128);
or U8375 (N_8375,N_8175,N_8128);
nor U8376 (N_8376,N_8193,N_8180);
nand U8377 (N_8377,N_8205,N_8113);
nor U8378 (N_8378,N_8210,N_8131);
and U8379 (N_8379,N_8178,N_8155);
xnor U8380 (N_8380,N_8205,N_8192);
nand U8381 (N_8381,N_8170,N_8171);
xor U8382 (N_8382,N_8183,N_8112);
nand U8383 (N_8383,N_8107,N_8227);
nand U8384 (N_8384,N_8160,N_8247);
nor U8385 (N_8385,N_8117,N_8206);
nor U8386 (N_8386,N_8164,N_8240);
nor U8387 (N_8387,N_8126,N_8224);
nor U8388 (N_8388,N_8174,N_8202);
and U8389 (N_8389,N_8241,N_8239);
nor U8390 (N_8390,N_8240,N_8199);
or U8391 (N_8391,N_8143,N_8157);
and U8392 (N_8392,N_8161,N_8222);
and U8393 (N_8393,N_8165,N_8146);
and U8394 (N_8394,N_8195,N_8220);
and U8395 (N_8395,N_8113,N_8182);
nand U8396 (N_8396,N_8120,N_8149);
xnor U8397 (N_8397,N_8228,N_8158);
xnor U8398 (N_8398,N_8152,N_8210);
or U8399 (N_8399,N_8117,N_8208);
or U8400 (N_8400,N_8334,N_8328);
nor U8401 (N_8401,N_8266,N_8283);
nand U8402 (N_8402,N_8306,N_8363);
or U8403 (N_8403,N_8313,N_8377);
nor U8404 (N_8404,N_8388,N_8301);
and U8405 (N_8405,N_8329,N_8369);
and U8406 (N_8406,N_8302,N_8348);
xnor U8407 (N_8407,N_8275,N_8295);
and U8408 (N_8408,N_8258,N_8308);
xor U8409 (N_8409,N_8255,N_8290);
nand U8410 (N_8410,N_8385,N_8397);
or U8411 (N_8411,N_8286,N_8294);
and U8412 (N_8412,N_8299,N_8312);
nor U8413 (N_8413,N_8352,N_8394);
and U8414 (N_8414,N_8359,N_8370);
nor U8415 (N_8415,N_8292,N_8327);
nand U8416 (N_8416,N_8323,N_8260);
xnor U8417 (N_8417,N_8257,N_8321);
nand U8418 (N_8418,N_8261,N_8314);
xor U8419 (N_8419,N_8337,N_8395);
nand U8420 (N_8420,N_8361,N_8259);
nand U8421 (N_8421,N_8356,N_8364);
nand U8422 (N_8422,N_8303,N_8367);
nand U8423 (N_8423,N_8358,N_8333);
nand U8424 (N_8424,N_8262,N_8269);
or U8425 (N_8425,N_8322,N_8318);
or U8426 (N_8426,N_8298,N_8389);
and U8427 (N_8427,N_8251,N_8392);
and U8428 (N_8428,N_8391,N_8305);
or U8429 (N_8429,N_8274,N_8346);
or U8430 (N_8430,N_8355,N_8373);
and U8431 (N_8431,N_8325,N_8332);
nand U8432 (N_8432,N_8307,N_8343);
nand U8433 (N_8433,N_8287,N_8277);
and U8434 (N_8434,N_8324,N_8365);
nor U8435 (N_8435,N_8354,N_8317);
and U8436 (N_8436,N_8340,N_8282);
and U8437 (N_8437,N_8383,N_8335);
xor U8438 (N_8438,N_8375,N_8320);
nand U8439 (N_8439,N_8344,N_8368);
nor U8440 (N_8440,N_8326,N_8316);
nor U8441 (N_8441,N_8256,N_8252);
and U8442 (N_8442,N_8376,N_8366);
xnor U8443 (N_8443,N_8271,N_8304);
or U8444 (N_8444,N_8273,N_8382);
nor U8445 (N_8445,N_8300,N_8350);
xor U8446 (N_8446,N_8371,N_8264);
nand U8447 (N_8447,N_8393,N_8268);
and U8448 (N_8448,N_8372,N_8281);
nor U8449 (N_8449,N_8272,N_8341);
nor U8450 (N_8450,N_8278,N_8387);
or U8451 (N_8451,N_8331,N_8384);
nand U8452 (N_8452,N_8263,N_8254);
and U8453 (N_8453,N_8250,N_8360);
and U8454 (N_8454,N_8390,N_8379);
nor U8455 (N_8455,N_8357,N_8289);
or U8456 (N_8456,N_8284,N_8380);
nand U8457 (N_8457,N_8342,N_8293);
nand U8458 (N_8458,N_8310,N_8336);
or U8459 (N_8459,N_8338,N_8330);
nor U8460 (N_8460,N_8386,N_8351);
nor U8461 (N_8461,N_8378,N_8347);
nand U8462 (N_8462,N_8399,N_8276);
nor U8463 (N_8463,N_8253,N_8297);
nor U8464 (N_8464,N_8339,N_8309);
nand U8465 (N_8465,N_8291,N_8349);
nor U8466 (N_8466,N_8296,N_8280);
nor U8467 (N_8467,N_8288,N_8285);
or U8468 (N_8468,N_8345,N_8398);
and U8469 (N_8469,N_8315,N_8311);
or U8470 (N_8470,N_8279,N_8362);
nor U8471 (N_8471,N_8381,N_8353);
nand U8472 (N_8472,N_8265,N_8319);
nor U8473 (N_8473,N_8396,N_8270);
xnor U8474 (N_8474,N_8267,N_8374);
nand U8475 (N_8475,N_8258,N_8320);
xnor U8476 (N_8476,N_8253,N_8380);
xor U8477 (N_8477,N_8356,N_8304);
xor U8478 (N_8478,N_8389,N_8297);
nor U8479 (N_8479,N_8338,N_8297);
nand U8480 (N_8480,N_8317,N_8390);
and U8481 (N_8481,N_8251,N_8373);
xor U8482 (N_8482,N_8267,N_8275);
nand U8483 (N_8483,N_8285,N_8263);
and U8484 (N_8484,N_8347,N_8386);
nand U8485 (N_8485,N_8354,N_8278);
nor U8486 (N_8486,N_8254,N_8292);
nor U8487 (N_8487,N_8260,N_8328);
nor U8488 (N_8488,N_8302,N_8264);
nor U8489 (N_8489,N_8352,N_8260);
nand U8490 (N_8490,N_8361,N_8296);
xnor U8491 (N_8491,N_8335,N_8286);
and U8492 (N_8492,N_8364,N_8278);
xnor U8493 (N_8493,N_8299,N_8305);
nor U8494 (N_8494,N_8288,N_8320);
nor U8495 (N_8495,N_8258,N_8322);
nor U8496 (N_8496,N_8384,N_8267);
xor U8497 (N_8497,N_8375,N_8348);
or U8498 (N_8498,N_8302,N_8394);
nor U8499 (N_8499,N_8359,N_8323);
nor U8500 (N_8500,N_8305,N_8288);
or U8501 (N_8501,N_8361,N_8395);
nand U8502 (N_8502,N_8319,N_8271);
nand U8503 (N_8503,N_8318,N_8348);
nand U8504 (N_8504,N_8339,N_8314);
or U8505 (N_8505,N_8333,N_8365);
nand U8506 (N_8506,N_8316,N_8313);
nor U8507 (N_8507,N_8301,N_8376);
nor U8508 (N_8508,N_8268,N_8363);
nor U8509 (N_8509,N_8316,N_8309);
nand U8510 (N_8510,N_8357,N_8374);
or U8511 (N_8511,N_8290,N_8351);
nor U8512 (N_8512,N_8341,N_8311);
xnor U8513 (N_8513,N_8302,N_8374);
and U8514 (N_8514,N_8368,N_8329);
nand U8515 (N_8515,N_8251,N_8397);
and U8516 (N_8516,N_8396,N_8319);
nor U8517 (N_8517,N_8394,N_8310);
nor U8518 (N_8518,N_8396,N_8314);
xor U8519 (N_8519,N_8261,N_8365);
or U8520 (N_8520,N_8377,N_8367);
or U8521 (N_8521,N_8271,N_8380);
nor U8522 (N_8522,N_8314,N_8290);
xor U8523 (N_8523,N_8360,N_8345);
or U8524 (N_8524,N_8336,N_8304);
nor U8525 (N_8525,N_8386,N_8326);
nor U8526 (N_8526,N_8309,N_8283);
and U8527 (N_8527,N_8299,N_8393);
nor U8528 (N_8528,N_8380,N_8263);
or U8529 (N_8529,N_8397,N_8379);
xnor U8530 (N_8530,N_8340,N_8262);
or U8531 (N_8531,N_8316,N_8332);
or U8532 (N_8532,N_8321,N_8299);
nand U8533 (N_8533,N_8323,N_8351);
and U8534 (N_8534,N_8383,N_8350);
nor U8535 (N_8535,N_8374,N_8268);
nor U8536 (N_8536,N_8329,N_8287);
xor U8537 (N_8537,N_8266,N_8255);
or U8538 (N_8538,N_8376,N_8320);
or U8539 (N_8539,N_8364,N_8317);
or U8540 (N_8540,N_8385,N_8262);
xor U8541 (N_8541,N_8334,N_8320);
nor U8542 (N_8542,N_8377,N_8268);
nor U8543 (N_8543,N_8347,N_8304);
nand U8544 (N_8544,N_8387,N_8352);
nor U8545 (N_8545,N_8307,N_8256);
nand U8546 (N_8546,N_8352,N_8363);
xnor U8547 (N_8547,N_8328,N_8317);
or U8548 (N_8548,N_8341,N_8326);
and U8549 (N_8549,N_8250,N_8314);
nor U8550 (N_8550,N_8485,N_8440);
nand U8551 (N_8551,N_8437,N_8490);
xor U8552 (N_8552,N_8537,N_8518);
xor U8553 (N_8553,N_8482,N_8525);
nor U8554 (N_8554,N_8447,N_8543);
and U8555 (N_8555,N_8507,N_8468);
and U8556 (N_8556,N_8541,N_8546);
or U8557 (N_8557,N_8469,N_8523);
xnor U8558 (N_8558,N_8465,N_8516);
nor U8559 (N_8559,N_8467,N_8512);
xnor U8560 (N_8560,N_8427,N_8530);
and U8561 (N_8561,N_8446,N_8462);
xnor U8562 (N_8562,N_8488,N_8458);
or U8563 (N_8563,N_8422,N_8472);
xnor U8564 (N_8564,N_8545,N_8480);
and U8565 (N_8565,N_8453,N_8414);
xor U8566 (N_8566,N_8439,N_8419);
and U8567 (N_8567,N_8428,N_8544);
xnor U8568 (N_8568,N_8400,N_8466);
xor U8569 (N_8569,N_8442,N_8402);
or U8570 (N_8570,N_8505,N_8423);
nor U8571 (N_8571,N_8533,N_8548);
or U8572 (N_8572,N_8405,N_8521);
nor U8573 (N_8573,N_8509,N_8529);
and U8574 (N_8574,N_8535,N_8496);
and U8575 (N_8575,N_8476,N_8421);
and U8576 (N_8576,N_8460,N_8540);
or U8577 (N_8577,N_8409,N_8484);
nor U8578 (N_8578,N_8475,N_8435);
or U8579 (N_8579,N_8429,N_8418);
xnor U8580 (N_8580,N_8463,N_8497);
xor U8581 (N_8581,N_8517,N_8508);
and U8582 (N_8582,N_8445,N_8538);
xnor U8583 (N_8583,N_8431,N_8404);
nor U8584 (N_8584,N_8448,N_8515);
nor U8585 (N_8585,N_8450,N_8489);
xnor U8586 (N_8586,N_8464,N_8504);
nor U8587 (N_8587,N_8420,N_8425);
nor U8588 (N_8588,N_8491,N_8531);
nand U8589 (N_8589,N_8532,N_8434);
and U8590 (N_8590,N_8413,N_8454);
and U8591 (N_8591,N_8471,N_8470);
nor U8592 (N_8592,N_8506,N_8536);
and U8593 (N_8593,N_8456,N_8433);
nor U8594 (N_8594,N_8499,N_8455);
nand U8595 (N_8595,N_8524,N_8520);
xnor U8596 (N_8596,N_8438,N_8514);
and U8597 (N_8597,N_8451,N_8430);
nor U8598 (N_8598,N_8410,N_8459);
nor U8599 (N_8599,N_8452,N_8407);
nand U8600 (N_8600,N_8502,N_8478);
nand U8601 (N_8601,N_8401,N_8511);
xor U8602 (N_8602,N_8473,N_8415);
nand U8603 (N_8603,N_8444,N_8403);
and U8604 (N_8604,N_8494,N_8483);
or U8605 (N_8605,N_8487,N_8513);
nand U8606 (N_8606,N_8526,N_8492);
xor U8607 (N_8607,N_8486,N_8527);
nor U8608 (N_8608,N_8474,N_8539);
and U8609 (N_8609,N_8519,N_8426);
nand U8610 (N_8610,N_8416,N_8406);
and U8611 (N_8611,N_8411,N_8417);
nand U8612 (N_8612,N_8461,N_8441);
xor U8613 (N_8613,N_8436,N_8510);
and U8614 (N_8614,N_8424,N_8549);
or U8615 (N_8615,N_8432,N_8493);
nor U8616 (N_8616,N_8547,N_8500);
nand U8617 (N_8617,N_8449,N_8501);
and U8618 (N_8618,N_8495,N_8481);
and U8619 (N_8619,N_8503,N_8479);
nand U8620 (N_8620,N_8498,N_8412);
nor U8621 (N_8621,N_8542,N_8457);
nand U8622 (N_8622,N_8408,N_8477);
or U8623 (N_8623,N_8443,N_8528);
xor U8624 (N_8624,N_8534,N_8522);
nor U8625 (N_8625,N_8418,N_8509);
or U8626 (N_8626,N_8414,N_8454);
or U8627 (N_8627,N_8499,N_8504);
xnor U8628 (N_8628,N_8546,N_8545);
nand U8629 (N_8629,N_8512,N_8461);
and U8630 (N_8630,N_8466,N_8422);
and U8631 (N_8631,N_8484,N_8464);
and U8632 (N_8632,N_8477,N_8464);
nand U8633 (N_8633,N_8424,N_8418);
and U8634 (N_8634,N_8476,N_8403);
or U8635 (N_8635,N_8515,N_8423);
nand U8636 (N_8636,N_8491,N_8520);
nor U8637 (N_8637,N_8530,N_8513);
xnor U8638 (N_8638,N_8441,N_8400);
xor U8639 (N_8639,N_8525,N_8488);
or U8640 (N_8640,N_8469,N_8518);
xor U8641 (N_8641,N_8487,N_8449);
xnor U8642 (N_8642,N_8519,N_8438);
xnor U8643 (N_8643,N_8538,N_8457);
nand U8644 (N_8644,N_8526,N_8513);
and U8645 (N_8645,N_8429,N_8457);
or U8646 (N_8646,N_8441,N_8475);
nor U8647 (N_8647,N_8457,N_8459);
xnor U8648 (N_8648,N_8412,N_8467);
and U8649 (N_8649,N_8417,N_8540);
and U8650 (N_8650,N_8479,N_8435);
nor U8651 (N_8651,N_8431,N_8446);
xnor U8652 (N_8652,N_8536,N_8491);
nor U8653 (N_8653,N_8537,N_8498);
or U8654 (N_8654,N_8475,N_8485);
nor U8655 (N_8655,N_8456,N_8490);
nand U8656 (N_8656,N_8500,N_8417);
or U8657 (N_8657,N_8400,N_8517);
and U8658 (N_8658,N_8484,N_8431);
xnor U8659 (N_8659,N_8423,N_8548);
nor U8660 (N_8660,N_8466,N_8501);
or U8661 (N_8661,N_8422,N_8421);
or U8662 (N_8662,N_8541,N_8547);
or U8663 (N_8663,N_8506,N_8440);
and U8664 (N_8664,N_8467,N_8476);
or U8665 (N_8665,N_8452,N_8418);
nor U8666 (N_8666,N_8450,N_8527);
nor U8667 (N_8667,N_8491,N_8418);
or U8668 (N_8668,N_8543,N_8463);
nand U8669 (N_8669,N_8435,N_8541);
xnor U8670 (N_8670,N_8543,N_8540);
xor U8671 (N_8671,N_8404,N_8472);
nor U8672 (N_8672,N_8417,N_8412);
and U8673 (N_8673,N_8462,N_8476);
nand U8674 (N_8674,N_8522,N_8510);
and U8675 (N_8675,N_8473,N_8427);
and U8676 (N_8676,N_8485,N_8452);
or U8677 (N_8677,N_8410,N_8532);
nand U8678 (N_8678,N_8508,N_8472);
nand U8679 (N_8679,N_8490,N_8417);
nor U8680 (N_8680,N_8436,N_8524);
and U8681 (N_8681,N_8455,N_8547);
nand U8682 (N_8682,N_8518,N_8424);
xor U8683 (N_8683,N_8475,N_8424);
and U8684 (N_8684,N_8537,N_8496);
or U8685 (N_8685,N_8516,N_8526);
nand U8686 (N_8686,N_8449,N_8543);
xor U8687 (N_8687,N_8502,N_8531);
nor U8688 (N_8688,N_8495,N_8436);
and U8689 (N_8689,N_8408,N_8433);
nor U8690 (N_8690,N_8461,N_8478);
nor U8691 (N_8691,N_8499,N_8539);
nand U8692 (N_8692,N_8462,N_8436);
or U8693 (N_8693,N_8493,N_8458);
nand U8694 (N_8694,N_8476,N_8505);
nand U8695 (N_8695,N_8538,N_8408);
and U8696 (N_8696,N_8450,N_8532);
xnor U8697 (N_8697,N_8541,N_8417);
and U8698 (N_8698,N_8463,N_8481);
nand U8699 (N_8699,N_8503,N_8452);
nand U8700 (N_8700,N_8636,N_8596);
and U8701 (N_8701,N_8609,N_8593);
nor U8702 (N_8702,N_8604,N_8651);
xor U8703 (N_8703,N_8589,N_8662);
and U8704 (N_8704,N_8608,N_8692);
xnor U8705 (N_8705,N_8670,N_8697);
nor U8706 (N_8706,N_8659,N_8669);
nor U8707 (N_8707,N_8642,N_8590);
and U8708 (N_8708,N_8638,N_8574);
xnor U8709 (N_8709,N_8630,N_8623);
xnor U8710 (N_8710,N_8628,N_8591);
nand U8711 (N_8711,N_8677,N_8552);
and U8712 (N_8712,N_8621,N_8611);
nor U8713 (N_8713,N_8555,N_8640);
or U8714 (N_8714,N_8699,N_8579);
or U8715 (N_8715,N_8598,N_8647);
nand U8716 (N_8716,N_8633,N_8649);
nand U8717 (N_8717,N_8663,N_8625);
xnor U8718 (N_8718,N_8622,N_8678);
xnor U8719 (N_8719,N_8619,N_8569);
or U8720 (N_8720,N_8629,N_8553);
xor U8721 (N_8721,N_8680,N_8612);
and U8722 (N_8722,N_8603,N_8661);
and U8723 (N_8723,N_8685,N_8615);
xor U8724 (N_8724,N_8691,N_8646);
nor U8725 (N_8725,N_8644,N_8627);
nand U8726 (N_8726,N_8582,N_8580);
or U8727 (N_8727,N_8645,N_8551);
nor U8728 (N_8728,N_8639,N_8654);
and U8729 (N_8729,N_8602,N_8557);
nor U8730 (N_8730,N_8689,N_8564);
or U8731 (N_8731,N_8676,N_8687);
nand U8732 (N_8732,N_8634,N_8671);
and U8733 (N_8733,N_8556,N_8675);
nand U8734 (N_8734,N_8617,N_8667);
nand U8735 (N_8735,N_8588,N_8652);
nand U8736 (N_8736,N_8626,N_8658);
and U8737 (N_8737,N_8605,N_8656);
nand U8738 (N_8738,N_8694,N_8550);
nor U8739 (N_8739,N_8581,N_8610);
nand U8740 (N_8740,N_8683,N_8616);
or U8741 (N_8741,N_8575,N_8618);
and U8742 (N_8742,N_8565,N_8578);
or U8743 (N_8743,N_8601,N_8693);
and U8744 (N_8744,N_8686,N_8585);
nor U8745 (N_8745,N_8668,N_8635);
xor U8746 (N_8746,N_8592,N_8572);
xnor U8747 (N_8747,N_8554,N_8567);
xor U8748 (N_8748,N_8681,N_8587);
xor U8749 (N_8749,N_8624,N_8595);
nor U8750 (N_8750,N_8620,N_8606);
and U8751 (N_8751,N_8632,N_8586);
xor U8752 (N_8752,N_8566,N_8664);
and U8753 (N_8753,N_8560,N_8577);
nand U8754 (N_8754,N_8594,N_8614);
xnor U8755 (N_8755,N_8559,N_8679);
nor U8756 (N_8756,N_8666,N_8698);
xnor U8757 (N_8757,N_8672,N_8641);
nor U8758 (N_8758,N_8576,N_8688);
nor U8759 (N_8759,N_8695,N_8562);
xor U8760 (N_8760,N_8571,N_8584);
nand U8761 (N_8761,N_8690,N_8631);
nor U8762 (N_8762,N_8600,N_8657);
xor U8763 (N_8763,N_8573,N_8684);
or U8764 (N_8764,N_8673,N_8558);
or U8765 (N_8765,N_8563,N_8650);
xor U8766 (N_8766,N_8637,N_8568);
nand U8767 (N_8767,N_8599,N_8561);
xnor U8768 (N_8768,N_8655,N_8682);
nor U8769 (N_8769,N_8648,N_8660);
or U8770 (N_8770,N_8597,N_8570);
xor U8771 (N_8771,N_8607,N_8613);
xnor U8772 (N_8772,N_8583,N_8665);
or U8773 (N_8773,N_8653,N_8643);
or U8774 (N_8774,N_8674,N_8696);
xnor U8775 (N_8775,N_8670,N_8633);
nor U8776 (N_8776,N_8576,N_8584);
nor U8777 (N_8777,N_8567,N_8632);
or U8778 (N_8778,N_8645,N_8646);
xnor U8779 (N_8779,N_8606,N_8660);
and U8780 (N_8780,N_8657,N_8596);
nand U8781 (N_8781,N_8677,N_8624);
or U8782 (N_8782,N_8638,N_8635);
xnor U8783 (N_8783,N_8649,N_8607);
nand U8784 (N_8784,N_8677,N_8681);
nor U8785 (N_8785,N_8679,N_8641);
nand U8786 (N_8786,N_8663,N_8642);
xor U8787 (N_8787,N_8565,N_8653);
and U8788 (N_8788,N_8615,N_8658);
nor U8789 (N_8789,N_8695,N_8633);
xnor U8790 (N_8790,N_8570,N_8659);
or U8791 (N_8791,N_8663,N_8648);
and U8792 (N_8792,N_8612,N_8605);
nand U8793 (N_8793,N_8610,N_8623);
xnor U8794 (N_8794,N_8592,N_8624);
or U8795 (N_8795,N_8577,N_8592);
nand U8796 (N_8796,N_8666,N_8579);
nor U8797 (N_8797,N_8650,N_8687);
nor U8798 (N_8798,N_8615,N_8561);
xnor U8799 (N_8799,N_8558,N_8628);
and U8800 (N_8800,N_8660,N_8575);
xnor U8801 (N_8801,N_8630,N_8673);
and U8802 (N_8802,N_8641,N_8591);
nand U8803 (N_8803,N_8661,N_8599);
or U8804 (N_8804,N_8584,N_8563);
and U8805 (N_8805,N_8688,N_8575);
xor U8806 (N_8806,N_8659,N_8693);
nor U8807 (N_8807,N_8685,N_8646);
and U8808 (N_8808,N_8624,N_8604);
xnor U8809 (N_8809,N_8565,N_8559);
or U8810 (N_8810,N_8557,N_8681);
and U8811 (N_8811,N_8663,N_8620);
nand U8812 (N_8812,N_8615,N_8678);
nor U8813 (N_8813,N_8631,N_8633);
and U8814 (N_8814,N_8604,N_8633);
and U8815 (N_8815,N_8586,N_8565);
nand U8816 (N_8816,N_8642,N_8644);
and U8817 (N_8817,N_8583,N_8594);
nor U8818 (N_8818,N_8596,N_8643);
nand U8819 (N_8819,N_8666,N_8684);
and U8820 (N_8820,N_8636,N_8646);
nor U8821 (N_8821,N_8643,N_8597);
xor U8822 (N_8822,N_8693,N_8649);
and U8823 (N_8823,N_8619,N_8610);
and U8824 (N_8824,N_8585,N_8617);
and U8825 (N_8825,N_8623,N_8587);
nor U8826 (N_8826,N_8675,N_8584);
nor U8827 (N_8827,N_8637,N_8552);
nand U8828 (N_8828,N_8623,N_8650);
nor U8829 (N_8829,N_8551,N_8680);
nor U8830 (N_8830,N_8610,N_8616);
nand U8831 (N_8831,N_8611,N_8563);
xnor U8832 (N_8832,N_8689,N_8685);
nand U8833 (N_8833,N_8671,N_8581);
nor U8834 (N_8834,N_8559,N_8673);
nand U8835 (N_8835,N_8633,N_8667);
xnor U8836 (N_8836,N_8656,N_8631);
and U8837 (N_8837,N_8595,N_8568);
xor U8838 (N_8838,N_8558,N_8617);
xnor U8839 (N_8839,N_8583,N_8577);
nand U8840 (N_8840,N_8594,N_8679);
or U8841 (N_8841,N_8675,N_8696);
nor U8842 (N_8842,N_8550,N_8604);
and U8843 (N_8843,N_8598,N_8619);
nor U8844 (N_8844,N_8608,N_8660);
and U8845 (N_8845,N_8688,N_8571);
nor U8846 (N_8846,N_8615,N_8567);
or U8847 (N_8847,N_8620,N_8642);
or U8848 (N_8848,N_8677,N_8570);
nor U8849 (N_8849,N_8572,N_8660);
xor U8850 (N_8850,N_8761,N_8776);
or U8851 (N_8851,N_8766,N_8717);
nand U8852 (N_8852,N_8740,N_8812);
or U8853 (N_8853,N_8708,N_8784);
xnor U8854 (N_8854,N_8810,N_8836);
nand U8855 (N_8855,N_8790,N_8815);
nor U8856 (N_8856,N_8795,N_8765);
nor U8857 (N_8857,N_8732,N_8793);
or U8858 (N_8858,N_8734,N_8741);
or U8859 (N_8859,N_8835,N_8747);
or U8860 (N_8860,N_8788,N_8774);
and U8861 (N_8861,N_8822,N_8752);
and U8862 (N_8862,N_8735,N_8780);
nor U8863 (N_8863,N_8826,N_8799);
xnor U8864 (N_8864,N_8749,N_8701);
or U8865 (N_8865,N_8715,N_8827);
or U8866 (N_8866,N_8845,N_8779);
nor U8867 (N_8867,N_8820,N_8837);
and U8868 (N_8868,N_8825,N_8729);
or U8869 (N_8869,N_8757,N_8737);
xnor U8870 (N_8870,N_8731,N_8777);
and U8871 (N_8871,N_8726,N_8840);
xor U8872 (N_8872,N_8781,N_8802);
nand U8873 (N_8873,N_8814,N_8768);
nor U8874 (N_8874,N_8772,N_8706);
nor U8875 (N_8875,N_8755,N_8721);
and U8876 (N_8876,N_8759,N_8705);
xnor U8877 (N_8877,N_8733,N_8796);
or U8878 (N_8878,N_8787,N_8844);
xnor U8879 (N_8879,N_8838,N_8775);
nor U8880 (N_8880,N_8754,N_8829);
or U8881 (N_8881,N_8738,N_8739);
nand U8882 (N_8882,N_8762,N_8702);
xor U8883 (N_8883,N_8816,N_8778);
or U8884 (N_8884,N_8771,N_8834);
nand U8885 (N_8885,N_8723,N_8709);
and U8886 (N_8886,N_8830,N_8743);
nor U8887 (N_8887,N_8786,N_8800);
nand U8888 (N_8888,N_8707,N_8711);
or U8889 (N_8889,N_8828,N_8750);
xnor U8890 (N_8890,N_8832,N_8813);
nand U8891 (N_8891,N_8797,N_8849);
xnor U8892 (N_8892,N_8751,N_8817);
nor U8893 (N_8893,N_8744,N_8770);
xnor U8894 (N_8894,N_8718,N_8833);
nor U8895 (N_8895,N_8819,N_8841);
or U8896 (N_8896,N_8809,N_8798);
xor U8897 (N_8897,N_8806,N_8847);
or U8898 (N_8898,N_8725,N_8712);
xor U8899 (N_8899,N_8724,N_8794);
and U8900 (N_8900,N_8716,N_8818);
or U8901 (N_8901,N_8848,N_8736);
nand U8902 (N_8902,N_8842,N_8753);
or U8903 (N_8903,N_8821,N_8769);
or U8904 (N_8904,N_8791,N_8746);
or U8905 (N_8905,N_8710,N_8730);
xor U8906 (N_8906,N_8823,N_8801);
nand U8907 (N_8907,N_8764,N_8831);
and U8908 (N_8908,N_8824,N_8722);
or U8909 (N_8909,N_8727,N_8742);
xnor U8910 (N_8910,N_8804,N_8808);
xor U8911 (N_8911,N_8719,N_8846);
nor U8912 (N_8912,N_8714,N_8700);
nor U8913 (N_8913,N_8789,N_8843);
nand U8914 (N_8914,N_8720,N_8792);
xor U8915 (N_8915,N_8713,N_8811);
nand U8916 (N_8916,N_8756,N_8760);
and U8917 (N_8917,N_8728,N_8803);
xnor U8918 (N_8918,N_8805,N_8773);
nor U8919 (N_8919,N_8703,N_8704);
xor U8920 (N_8920,N_8767,N_8783);
nor U8921 (N_8921,N_8782,N_8763);
nor U8922 (N_8922,N_8748,N_8839);
nor U8923 (N_8923,N_8758,N_8785);
or U8924 (N_8924,N_8745,N_8807);
or U8925 (N_8925,N_8704,N_8824);
xor U8926 (N_8926,N_8810,N_8736);
or U8927 (N_8927,N_8766,N_8728);
xnor U8928 (N_8928,N_8752,N_8804);
xnor U8929 (N_8929,N_8762,N_8783);
nand U8930 (N_8930,N_8806,N_8782);
nand U8931 (N_8931,N_8835,N_8813);
xor U8932 (N_8932,N_8829,N_8809);
nor U8933 (N_8933,N_8726,N_8716);
or U8934 (N_8934,N_8707,N_8702);
and U8935 (N_8935,N_8759,N_8823);
nand U8936 (N_8936,N_8747,N_8818);
or U8937 (N_8937,N_8722,N_8845);
and U8938 (N_8938,N_8770,N_8849);
nor U8939 (N_8939,N_8788,N_8816);
xor U8940 (N_8940,N_8816,N_8807);
nor U8941 (N_8941,N_8818,N_8755);
nand U8942 (N_8942,N_8834,N_8726);
nand U8943 (N_8943,N_8703,N_8705);
or U8944 (N_8944,N_8711,N_8780);
xor U8945 (N_8945,N_8773,N_8836);
or U8946 (N_8946,N_8725,N_8817);
nand U8947 (N_8947,N_8733,N_8760);
nor U8948 (N_8948,N_8794,N_8833);
or U8949 (N_8949,N_8845,N_8777);
or U8950 (N_8950,N_8701,N_8753);
xor U8951 (N_8951,N_8838,N_8779);
xor U8952 (N_8952,N_8778,N_8790);
nand U8953 (N_8953,N_8792,N_8719);
xor U8954 (N_8954,N_8743,N_8783);
nand U8955 (N_8955,N_8705,N_8725);
xnor U8956 (N_8956,N_8730,N_8729);
nand U8957 (N_8957,N_8786,N_8759);
and U8958 (N_8958,N_8796,N_8848);
nor U8959 (N_8959,N_8742,N_8798);
nor U8960 (N_8960,N_8756,N_8746);
and U8961 (N_8961,N_8716,N_8807);
nor U8962 (N_8962,N_8833,N_8842);
nor U8963 (N_8963,N_8811,N_8717);
or U8964 (N_8964,N_8701,N_8761);
and U8965 (N_8965,N_8726,N_8813);
xnor U8966 (N_8966,N_8798,N_8709);
and U8967 (N_8967,N_8841,N_8796);
or U8968 (N_8968,N_8789,N_8838);
xor U8969 (N_8969,N_8714,N_8811);
and U8970 (N_8970,N_8846,N_8805);
or U8971 (N_8971,N_8725,N_8750);
xor U8972 (N_8972,N_8732,N_8846);
and U8973 (N_8973,N_8796,N_8792);
and U8974 (N_8974,N_8764,N_8778);
xor U8975 (N_8975,N_8751,N_8736);
and U8976 (N_8976,N_8745,N_8816);
and U8977 (N_8977,N_8790,N_8847);
nor U8978 (N_8978,N_8704,N_8723);
and U8979 (N_8979,N_8738,N_8771);
and U8980 (N_8980,N_8756,N_8741);
nor U8981 (N_8981,N_8718,N_8812);
or U8982 (N_8982,N_8790,N_8789);
nand U8983 (N_8983,N_8791,N_8834);
and U8984 (N_8984,N_8753,N_8782);
or U8985 (N_8985,N_8807,N_8813);
nand U8986 (N_8986,N_8774,N_8736);
and U8987 (N_8987,N_8742,N_8832);
nand U8988 (N_8988,N_8785,N_8729);
nor U8989 (N_8989,N_8724,N_8772);
or U8990 (N_8990,N_8703,N_8836);
nor U8991 (N_8991,N_8741,N_8768);
xor U8992 (N_8992,N_8726,N_8804);
xor U8993 (N_8993,N_8705,N_8832);
nand U8994 (N_8994,N_8746,N_8802);
or U8995 (N_8995,N_8711,N_8808);
or U8996 (N_8996,N_8812,N_8760);
nor U8997 (N_8997,N_8771,N_8749);
and U8998 (N_8998,N_8744,N_8709);
and U8999 (N_8999,N_8787,N_8841);
nand U9000 (N_9000,N_8922,N_8985);
xor U9001 (N_9001,N_8862,N_8861);
nand U9002 (N_9002,N_8872,N_8917);
or U9003 (N_9003,N_8994,N_8904);
or U9004 (N_9004,N_8868,N_8995);
nand U9005 (N_9005,N_8983,N_8859);
nand U9006 (N_9006,N_8938,N_8997);
or U9007 (N_9007,N_8908,N_8877);
or U9008 (N_9008,N_8918,N_8946);
and U9009 (N_9009,N_8858,N_8880);
nand U9010 (N_9010,N_8989,N_8889);
xnor U9011 (N_9011,N_8947,N_8970);
nor U9012 (N_9012,N_8950,N_8912);
xor U9013 (N_9013,N_8987,N_8936);
nor U9014 (N_9014,N_8900,N_8982);
or U9015 (N_9015,N_8948,N_8855);
nor U9016 (N_9016,N_8852,N_8945);
and U9017 (N_9017,N_8875,N_8935);
nand U9018 (N_9018,N_8897,N_8902);
and U9019 (N_9019,N_8911,N_8854);
and U9020 (N_9020,N_8886,N_8992);
nand U9021 (N_9021,N_8984,N_8933);
xnor U9022 (N_9022,N_8850,N_8878);
xnor U9023 (N_9023,N_8884,N_8873);
or U9024 (N_9024,N_8932,N_8891);
xnor U9025 (N_9025,N_8876,N_8980);
and U9026 (N_9026,N_8976,N_8999);
or U9027 (N_9027,N_8966,N_8954);
and U9028 (N_9028,N_8910,N_8962);
xnor U9029 (N_9029,N_8958,N_8863);
xnor U9030 (N_9030,N_8853,N_8923);
xor U9031 (N_9031,N_8971,N_8953);
xor U9032 (N_9032,N_8894,N_8981);
or U9033 (N_9033,N_8986,N_8998);
or U9034 (N_9034,N_8939,N_8871);
nand U9035 (N_9035,N_8996,N_8866);
xor U9036 (N_9036,N_8860,N_8856);
xnor U9037 (N_9037,N_8942,N_8934);
nor U9038 (N_9038,N_8892,N_8974);
xor U9039 (N_9039,N_8893,N_8914);
nand U9040 (N_9040,N_8916,N_8883);
and U9041 (N_9041,N_8979,N_8881);
nor U9042 (N_9042,N_8909,N_8952);
xor U9043 (N_9043,N_8929,N_8921);
nand U9044 (N_9044,N_8956,N_8943);
nand U9045 (N_9045,N_8951,N_8960);
nand U9046 (N_9046,N_8864,N_8920);
xnor U9047 (N_9047,N_8957,N_8993);
or U9048 (N_9048,N_8867,N_8977);
and U9049 (N_9049,N_8969,N_8890);
xnor U9050 (N_9050,N_8903,N_8851);
and U9051 (N_9051,N_8991,N_8944);
or U9052 (N_9052,N_8967,N_8887);
xnor U9053 (N_9053,N_8955,N_8899);
and U9054 (N_9054,N_8879,N_8973);
xnor U9055 (N_9055,N_8869,N_8972);
nor U9056 (N_9056,N_8888,N_8901);
and U9057 (N_9057,N_8941,N_8898);
xor U9058 (N_9058,N_8959,N_8865);
xnor U9059 (N_9059,N_8937,N_8913);
xnor U9060 (N_9060,N_8895,N_8907);
nand U9061 (N_9061,N_8990,N_8882);
nor U9062 (N_9062,N_8925,N_8963);
and U9063 (N_9063,N_8930,N_8857);
nor U9064 (N_9064,N_8874,N_8915);
or U9065 (N_9065,N_8924,N_8905);
or U9066 (N_9066,N_8870,N_8988);
xor U9067 (N_9067,N_8949,N_8919);
or U9068 (N_9068,N_8961,N_8965);
nand U9069 (N_9069,N_8928,N_8964);
nor U9070 (N_9070,N_8906,N_8927);
nand U9071 (N_9071,N_8968,N_8975);
or U9072 (N_9072,N_8931,N_8885);
or U9073 (N_9073,N_8978,N_8926);
nor U9074 (N_9074,N_8896,N_8940);
or U9075 (N_9075,N_8885,N_8952);
nand U9076 (N_9076,N_8922,N_8904);
and U9077 (N_9077,N_8943,N_8883);
or U9078 (N_9078,N_8959,N_8868);
or U9079 (N_9079,N_8857,N_8983);
nor U9080 (N_9080,N_8948,N_8991);
or U9081 (N_9081,N_8929,N_8930);
xnor U9082 (N_9082,N_8928,N_8911);
nand U9083 (N_9083,N_8910,N_8875);
nor U9084 (N_9084,N_8852,N_8991);
nand U9085 (N_9085,N_8977,N_8887);
and U9086 (N_9086,N_8937,N_8969);
nor U9087 (N_9087,N_8852,N_8985);
xnor U9088 (N_9088,N_8931,N_8991);
xnor U9089 (N_9089,N_8893,N_8912);
and U9090 (N_9090,N_8855,N_8854);
xor U9091 (N_9091,N_8885,N_8891);
xnor U9092 (N_9092,N_8974,N_8968);
nand U9093 (N_9093,N_8931,N_8879);
nand U9094 (N_9094,N_8967,N_8974);
and U9095 (N_9095,N_8888,N_8895);
nand U9096 (N_9096,N_8872,N_8866);
nand U9097 (N_9097,N_8880,N_8983);
nand U9098 (N_9098,N_8909,N_8996);
or U9099 (N_9099,N_8963,N_8897);
or U9100 (N_9100,N_8968,N_8873);
and U9101 (N_9101,N_8993,N_8898);
or U9102 (N_9102,N_8962,N_8896);
xor U9103 (N_9103,N_8872,N_8971);
or U9104 (N_9104,N_8897,N_8936);
or U9105 (N_9105,N_8908,N_8874);
or U9106 (N_9106,N_8936,N_8895);
xnor U9107 (N_9107,N_8999,N_8948);
nor U9108 (N_9108,N_8992,N_8986);
or U9109 (N_9109,N_8920,N_8924);
and U9110 (N_9110,N_8885,N_8942);
or U9111 (N_9111,N_8970,N_8896);
nor U9112 (N_9112,N_8986,N_8947);
and U9113 (N_9113,N_8850,N_8887);
nand U9114 (N_9114,N_8881,N_8919);
or U9115 (N_9115,N_8906,N_8865);
xnor U9116 (N_9116,N_8929,N_8901);
nand U9117 (N_9117,N_8862,N_8890);
nand U9118 (N_9118,N_8889,N_8995);
nand U9119 (N_9119,N_8938,N_8888);
xnor U9120 (N_9120,N_8993,N_8911);
nand U9121 (N_9121,N_8892,N_8958);
xnor U9122 (N_9122,N_8944,N_8989);
or U9123 (N_9123,N_8986,N_8991);
xor U9124 (N_9124,N_8942,N_8957);
nand U9125 (N_9125,N_8963,N_8874);
nor U9126 (N_9126,N_8927,N_8996);
xor U9127 (N_9127,N_8984,N_8919);
nand U9128 (N_9128,N_8896,N_8965);
xor U9129 (N_9129,N_8938,N_8924);
nand U9130 (N_9130,N_8979,N_8904);
xor U9131 (N_9131,N_8878,N_8876);
nand U9132 (N_9132,N_8892,N_8983);
or U9133 (N_9133,N_8957,N_8862);
or U9134 (N_9134,N_8916,N_8921);
nand U9135 (N_9135,N_8987,N_8970);
nand U9136 (N_9136,N_8932,N_8907);
xnor U9137 (N_9137,N_8895,N_8856);
and U9138 (N_9138,N_8850,N_8855);
and U9139 (N_9139,N_8908,N_8878);
or U9140 (N_9140,N_8967,N_8993);
and U9141 (N_9141,N_8998,N_8989);
or U9142 (N_9142,N_8937,N_8858);
xnor U9143 (N_9143,N_8878,N_8859);
xor U9144 (N_9144,N_8962,N_8854);
nor U9145 (N_9145,N_8910,N_8902);
and U9146 (N_9146,N_8949,N_8888);
and U9147 (N_9147,N_8938,N_8968);
nand U9148 (N_9148,N_8932,N_8924);
or U9149 (N_9149,N_8886,N_8896);
nand U9150 (N_9150,N_9044,N_9109);
xnor U9151 (N_9151,N_9056,N_9079);
nand U9152 (N_9152,N_9113,N_9147);
nand U9153 (N_9153,N_9080,N_9055);
or U9154 (N_9154,N_9035,N_9002);
nand U9155 (N_9155,N_9128,N_9018);
and U9156 (N_9156,N_9095,N_9136);
nor U9157 (N_9157,N_9012,N_9137);
or U9158 (N_9158,N_9001,N_9017);
and U9159 (N_9159,N_9023,N_9141);
and U9160 (N_9160,N_9059,N_9065);
and U9161 (N_9161,N_9029,N_9062);
or U9162 (N_9162,N_9097,N_9084);
xnor U9163 (N_9163,N_9130,N_9078);
or U9164 (N_9164,N_9054,N_9116);
xnor U9165 (N_9165,N_9005,N_9073);
nand U9166 (N_9166,N_9104,N_9072);
xnor U9167 (N_9167,N_9125,N_9094);
and U9168 (N_9168,N_9006,N_9142);
xor U9169 (N_9169,N_9036,N_9042);
xor U9170 (N_9170,N_9091,N_9088);
and U9171 (N_9171,N_9112,N_9131);
nand U9172 (N_9172,N_9010,N_9081);
nor U9173 (N_9173,N_9037,N_9134);
xor U9174 (N_9174,N_9077,N_9066);
nor U9175 (N_9175,N_9060,N_9020);
or U9176 (N_9176,N_9108,N_9047);
nor U9177 (N_9177,N_9046,N_9016);
xnor U9178 (N_9178,N_9118,N_9045);
nor U9179 (N_9179,N_9048,N_9129);
nor U9180 (N_9180,N_9148,N_9107);
nor U9181 (N_9181,N_9015,N_9025);
nor U9182 (N_9182,N_9024,N_9027);
nor U9183 (N_9183,N_9149,N_9132);
xor U9184 (N_9184,N_9135,N_9011);
and U9185 (N_9185,N_9049,N_9068);
and U9186 (N_9186,N_9071,N_9143);
and U9187 (N_9187,N_9028,N_9019);
and U9188 (N_9188,N_9013,N_9086);
and U9189 (N_9189,N_9039,N_9089);
or U9190 (N_9190,N_9050,N_9034);
or U9191 (N_9191,N_9145,N_9096);
and U9192 (N_9192,N_9061,N_9117);
or U9193 (N_9193,N_9082,N_9140);
and U9194 (N_9194,N_9022,N_9067);
nor U9195 (N_9195,N_9000,N_9119);
nand U9196 (N_9196,N_9026,N_9031);
nand U9197 (N_9197,N_9074,N_9093);
xnor U9198 (N_9198,N_9038,N_9040);
or U9199 (N_9199,N_9053,N_9102);
or U9200 (N_9200,N_9120,N_9070);
nor U9201 (N_9201,N_9090,N_9139);
nor U9202 (N_9202,N_9032,N_9114);
nand U9203 (N_9203,N_9052,N_9111);
xnor U9204 (N_9204,N_9057,N_9030);
or U9205 (N_9205,N_9127,N_9146);
and U9206 (N_9206,N_9144,N_9087);
xor U9207 (N_9207,N_9051,N_9115);
nand U9208 (N_9208,N_9098,N_9014);
nor U9209 (N_9209,N_9003,N_9138);
nand U9210 (N_9210,N_9041,N_9133);
nand U9211 (N_9211,N_9064,N_9069);
xor U9212 (N_9212,N_9083,N_9004);
xnor U9213 (N_9213,N_9092,N_9021);
and U9214 (N_9214,N_9110,N_9124);
or U9215 (N_9215,N_9075,N_9009);
xnor U9216 (N_9216,N_9103,N_9099);
nor U9217 (N_9217,N_9076,N_9063);
or U9218 (N_9218,N_9043,N_9106);
or U9219 (N_9219,N_9123,N_9007);
or U9220 (N_9220,N_9058,N_9121);
nor U9221 (N_9221,N_9008,N_9126);
or U9222 (N_9222,N_9105,N_9100);
xor U9223 (N_9223,N_9101,N_9033);
and U9224 (N_9224,N_9085,N_9122);
nand U9225 (N_9225,N_9051,N_9047);
nor U9226 (N_9226,N_9132,N_9061);
or U9227 (N_9227,N_9126,N_9055);
or U9228 (N_9228,N_9026,N_9126);
xnor U9229 (N_9229,N_9064,N_9039);
xnor U9230 (N_9230,N_9026,N_9134);
nand U9231 (N_9231,N_9033,N_9003);
nand U9232 (N_9232,N_9096,N_9050);
or U9233 (N_9233,N_9084,N_9035);
and U9234 (N_9234,N_9026,N_9037);
or U9235 (N_9235,N_9016,N_9012);
nand U9236 (N_9236,N_9049,N_9118);
nand U9237 (N_9237,N_9149,N_9006);
and U9238 (N_9238,N_9149,N_9005);
and U9239 (N_9239,N_9083,N_9120);
nor U9240 (N_9240,N_9003,N_9027);
xnor U9241 (N_9241,N_9084,N_9147);
nor U9242 (N_9242,N_9037,N_9118);
nand U9243 (N_9243,N_9078,N_9100);
and U9244 (N_9244,N_9118,N_9080);
xnor U9245 (N_9245,N_9098,N_9043);
and U9246 (N_9246,N_9055,N_9110);
xor U9247 (N_9247,N_9021,N_9124);
xor U9248 (N_9248,N_9136,N_9129);
and U9249 (N_9249,N_9066,N_9045);
xor U9250 (N_9250,N_9011,N_9146);
nand U9251 (N_9251,N_9113,N_9079);
nand U9252 (N_9252,N_9030,N_9110);
nand U9253 (N_9253,N_9046,N_9052);
xnor U9254 (N_9254,N_9071,N_9140);
or U9255 (N_9255,N_9138,N_9069);
xor U9256 (N_9256,N_9057,N_9006);
xnor U9257 (N_9257,N_9060,N_9108);
xnor U9258 (N_9258,N_9026,N_9146);
nor U9259 (N_9259,N_9053,N_9132);
or U9260 (N_9260,N_9032,N_9144);
nand U9261 (N_9261,N_9045,N_9094);
nand U9262 (N_9262,N_9143,N_9137);
xnor U9263 (N_9263,N_9030,N_9102);
or U9264 (N_9264,N_9088,N_9107);
or U9265 (N_9265,N_9079,N_9085);
nand U9266 (N_9266,N_9099,N_9136);
and U9267 (N_9267,N_9064,N_9141);
nand U9268 (N_9268,N_9016,N_9128);
nand U9269 (N_9269,N_9021,N_9107);
nand U9270 (N_9270,N_9032,N_9055);
nor U9271 (N_9271,N_9010,N_9126);
nand U9272 (N_9272,N_9131,N_9111);
and U9273 (N_9273,N_9098,N_9007);
nor U9274 (N_9274,N_9111,N_9080);
xor U9275 (N_9275,N_9111,N_9087);
or U9276 (N_9276,N_9045,N_9070);
xor U9277 (N_9277,N_9071,N_9056);
or U9278 (N_9278,N_9040,N_9016);
nor U9279 (N_9279,N_9149,N_9143);
and U9280 (N_9280,N_9029,N_9104);
and U9281 (N_9281,N_9113,N_9058);
nor U9282 (N_9282,N_9096,N_9124);
nor U9283 (N_9283,N_9117,N_9030);
or U9284 (N_9284,N_9049,N_9024);
xor U9285 (N_9285,N_9040,N_9130);
xnor U9286 (N_9286,N_9109,N_9089);
and U9287 (N_9287,N_9011,N_9046);
nor U9288 (N_9288,N_9032,N_9006);
nor U9289 (N_9289,N_9040,N_9053);
and U9290 (N_9290,N_9020,N_9023);
and U9291 (N_9291,N_9111,N_9021);
and U9292 (N_9292,N_9122,N_9137);
or U9293 (N_9293,N_9071,N_9130);
nand U9294 (N_9294,N_9012,N_9099);
and U9295 (N_9295,N_9019,N_9078);
nor U9296 (N_9296,N_9004,N_9003);
xor U9297 (N_9297,N_9148,N_9065);
and U9298 (N_9298,N_9098,N_9019);
nor U9299 (N_9299,N_9081,N_9129);
nand U9300 (N_9300,N_9266,N_9212);
and U9301 (N_9301,N_9278,N_9287);
and U9302 (N_9302,N_9158,N_9208);
or U9303 (N_9303,N_9210,N_9220);
nand U9304 (N_9304,N_9165,N_9290);
nor U9305 (N_9305,N_9298,N_9192);
nor U9306 (N_9306,N_9260,N_9226);
nor U9307 (N_9307,N_9207,N_9197);
nand U9308 (N_9308,N_9180,N_9292);
nand U9309 (N_9309,N_9252,N_9228);
xor U9310 (N_9310,N_9250,N_9150);
xnor U9311 (N_9311,N_9233,N_9224);
and U9312 (N_9312,N_9172,N_9241);
or U9313 (N_9313,N_9234,N_9257);
xnor U9314 (N_9314,N_9268,N_9238);
and U9315 (N_9315,N_9201,N_9263);
or U9316 (N_9316,N_9178,N_9277);
xnor U9317 (N_9317,N_9262,N_9198);
xor U9318 (N_9318,N_9256,N_9244);
nor U9319 (N_9319,N_9194,N_9171);
nor U9320 (N_9320,N_9232,N_9272);
nor U9321 (N_9321,N_9236,N_9254);
nor U9322 (N_9322,N_9281,N_9274);
xnor U9323 (N_9323,N_9296,N_9259);
or U9324 (N_9324,N_9229,N_9255);
nand U9325 (N_9325,N_9291,N_9209);
nand U9326 (N_9326,N_9285,N_9221);
xnor U9327 (N_9327,N_9168,N_9230);
nand U9328 (N_9328,N_9190,N_9294);
nand U9329 (N_9329,N_9216,N_9204);
nand U9330 (N_9330,N_9174,N_9243);
nor U9331 (N_9331,N_9185,N_9289);
nor U9332 (N_9332,N_9184,N_9156);
xor U9333 (N_9333,N_9218,N_9269);
xnor U9334 (N_9334,N_9205,N_9248);
xor U9335 (N_9335,N_9242,N_9187);
nor U9336 (N_9336,N_9223,N_9200);
and U9337 (N_9337,N_9155,N_9239);
and U9338 (N_9338,N_9211,N_9203);
nand U9339 (N_9339,N_9153,N_9275);
nand U9340 (N_9340,N_9227,N_9240);
nor U9341 (N_9341,N_9251,N_9151);
xor U9342 (N_9342,N_9293,N_9264);
nor U9343 (N_9343,N_9191,N_9267);
nor U9344 (N_9344,N_9297,N_9282);
and U9345 (N_9345,N_9199,N_9152);
or U9346 (N_9346,N_9213,N_9261);
xor U9347 (N_9347,N_9154,N_9169);
or U9348 (N_9348,N_9286,N_9271);
or U9349 (N_9349,N_9237,N_9225);
and U9350 (N_9350,N_9161,N_9247);
xor U9351 (N_9351,N_9245,N_9163);
xor U9352 (N_9352,N_9182,N_9258);
and U9353 (N_9353,N_9177,N_9276);
nor U9354 (N_9354,N_9188,N_9219);
nor U9355 (N_9355,N_9280,N_9173);
nor U9356 (N_9356,N_9235,N_9295);
nand U9357 (N_9357,N_9288,N_9279);
or U9358 (N_9358,N_9195,N_9157);
nand U9359 (N_9359,N_9206,N_9299);
and U9360 (N_9360,N_9246,N_9189);
xnor U9361 (N_9361,N_9181,N_9175);
nand U9362 (N_9362,N_9183,N_9202);
nor U9363 (N_9363,N_9284,N_9176);
and U9364 (N_9364,N_9270,N_9179);
xnor U9365 (N_9365,N_9166,N_9273);
xnor U9366 (N_9366,N_9265,N_9222);
nor U9367 (N_9367,N_9193,N_9217);
or U9368 (N_9368,N_9215,N_9159);
xor U9369 (N_9369,N_9164,N_9162);
nor U9370 (N_9370,N_9214,N_9231);
and U9371 (N_9371,N_9167,N_9196);
xor U9372 (N_9372,N_9283,N_9186);
nand U9373 (N_9373,N_9170,N_9249);
or U9374 (N_9374,N_9253,N_9160);
nand U9375 (N_9375,N_9216,N_9252);
xor U9376 (N_9376,N_9207,N_9241);
or U9377 (N_9377,N_9269,N_9174);
xnor U9378 (N_9378,N_9167,N_9245);
or U9379 (N_9379,N_9268,N_9221);
xor U9380 (N_9380,N_9240,N_9281);
nor U9381 (N_9381,N_9221,N_9287);
and U9382 (N_9382,N_9245,N_9298);
or U9383 (N_9383,N_9271,N_9251);
or U9384 (N_9384,N_9253,N_9298);
nand U9385 (N_9385,N_9255,N_9210);
nand U9386 (N_9386,N_9186,N_9213);
xor U9387 (N_9387,N_9179,N_9168);
nor U9388 (N_9388,N_9253,N_9235);
nor U9389 (N_9389,N_9216,N_9219);
or U9390 (N_9390,N_9206,N_9252);
and U9391 (N_9391,N_9169,N_9177);
nor U9392 (N_9392,N_9163,N_9197);
and U9393 (N_9393,N_9293,N_9250);
xnor U9394 (N_9394,N_9297,N_9267);
and U9395 (N_9395,N_9230,N_9196);
or U9396 (N_9396,N_9264,N_9284);
xnor U9397 (N_9397,N_9231,N_9293);
and U9398 (N_9398,N_9203,N_9281);
nand U9399 (N_9399,N_9233,N_9213);
and U9400 (N_9400,N_9236,N_9256);
nand U9401 (N_9401,N_9269,N_9230);
nand U9402 (N_9402,N_9265,N_9179);
and U9403 (N_9403,N_9155,N_9201);
nor U9404 (N_9404,N_9162,N_9255);
or U9405 (N_9405,N_9155,N_9215);
or U9406 (N_9406,N_9173,N_9190);
xnor U9407 (N_9407,N_9278,N_9284);
or U9408 (N_9408,N_9247,N_9178);
or U9409 (N_9409,N_9264,N_9196);
and U9410 (N_9410,N_9231,N_9219);
xnor U9411 (N_9411,N_9151,N_9171);
xnor U9412 (N_9412,N_9223,N_9239);
nor U9413 (N_9413,N_9194,N_9191);
and U9414 (N_9414,N_9288,N_9176);
or U9415 (N_9415,N_9213,N_9195);
xor U9416 (N_9416,N_9277,N_9162);
nor U9417 (N_9417,N_9245,N_9202);
xnor U9418 (N_9418,N_9198,N_9154);
xor U9419 (N_9419,N_9205,N_9228);
and U9420 (N_9420,N_9198,N_9240);
or U9421 (N_9421,N_9163,N_9292);
xnor U9422 (N_9422,N_9232,N_9163);
and U9423 (N_9423,N_9294,N_9218);
nand U9424 (N_9424,N_9215,N_9188);
or U9425 (N_9425,N_9210,N_9172);
or U9426 (N_9426,N_9291,N_9285);
nand U9427 (N_9427,N_9250,N_9162);
and U9428 (N_9428,N_9261,N_9289);
nor U9429 (N_9429,N_9192,N_9228);
and U9430 (N_9430,N_9207,N_9245);
or U9431 (N_9431,N_9171,N_9197);
nor U9432 (N_9432,N_9199,N_9190);
nor U9433 (N_9433,N_9220,N_9299);
and U9434 (N_9434,N_9205,N_9271);
or U9435 (N_9435,N_9242,N_9236);
xor U9436 (N_9436,N_9196,N_9227);
and U9437 (N_9437,N_9250,N_9166);
nor U9438 (N_9438,N_9221,N_9156);
nor U9439 (N_9439,N_9197,N_9224);
nand U9440 (N_9440,N_9238,N_9162);
nand U9441 (N_9441,N_9224,N_9296);
nand U9442 (N_9442,N_9205,N_9180);
and U9443 (N_9443,N_9171,N_9156);
and U9444 (N_9444,N_9155,N_9237);
or U9445 (N_9445,N_9167,N_9244);
nor U9446 (N_9446,N_9286,N_9176);
nor U9447 (N_9447,N_9186,N_9217);
nor U9448 (N_9448,N_9158,N_9294);
xor U9449 (N_9449,N_9255,N_9278);
nand U9450 (N_9450,N_9351,N_9334);
and U9451 (N_9451,N_9359,N_9442);
xnor U9452 (N_9452,N_9439,N_9394);
and U9453 (N_9453,N_9366,N_9324);
xnor U9454 (N_9454,N_9312,N_9314);
or U9455 (N_9455,N_9399,N_9411);
xor U9456 (N_9456,N_9392,N_9319);
and U9457 (N_9457,N_9325,N_9414);
nor U9458 (N_9458,N_9331,N_9418);
xor U9459 (N_9459,N_9428,N_9430);
nand U9460 (N_9460,N_9333,N_9356);
nand U9461 (N_9461,N_9378,N_9385);
and U9462 (N_9462,N_9321,N_9374);
xnor U9463 (N_9463,N_9413,N_9322);
and U9464 (N_9464,N_9326,N_9307);
nand U9465 (N_9465,N_9383,N_9422);
nor U9466 (N_9466,N_9357,N_9305);
xor U9467 (N_9467,N_9363,N_9339);
nand U9468 (N_9468,N_9316,N_9429);
and U9469 (N_9469,N_9420,N_9407);
nand U9470 (N_9470,N_9310,N_9338);
xnor U9471 (N_9471,N_9346,N_9330);
nand U9472 (N_9472,N_9332,N_9303);
nor U9473 (N_9473,N_9401,N_9379);
and U9474 (N_9474,N_9387,N_9400);
nand U9475 (N_9475,N_9423,N_9449);
nand U9476 (N_9476,N_9358,N_9441);
xor U9477 (N_9477,N_9365,N_9302);
and U9478 (N_9478,N_9361,N_9354);
nor U9479 (N_9479,N_9349,N_9405);
nand U9480 (N_9480,N_9445,N_9438);
nor U9481 (N_9481,N_9433,N_9409);
nand U9482 (N_9482,N_9342,N_9373);
xor U9483 (N_9483,N_9415,N_9308);
nor U9484 (N_9484,N_9404,N_9353);
nand U9485 (N_9485,N_9448,N_9437);
or U9486 (N_9486,N_9444,N_9436);
xnor U9487 (N_9487,N_9388,N_9391);
and U9488 (N_9488,N_9397,N_9364);
nand U9489 (N_9489,N_9435,N_9380);
or U9490 (N_9490,N_9355,N_9390);
xor U9491 (N_9491,N_9304,N_9381);
nand U9492 (N_9492,N_9384,N_9336);
and U9493 (N_9493,N_9343,N_9377);
xor U9494 (N_9494,N_9306,N_9419);
and U9495 (N_9495,N_9375,N_9421);
and U9496 (N_9496,N_9382,N_9398);
and U9497 (N_9497,N_9403,N_9371);
nand U9498 (N_9498,N_9408,N_9406);
and U9499 (N_9499,N_9372,N_9309);
xnor U9500 (N_9500,N_9412,N_9410);
and U9501 (N_9501,N_9376,N_9301);
and U9502 (N_9502,N_9317,N_9431);
xor U9503 (N_9503,N_9386,N_9352);
and U9504 (N_9504,N_9323,N_9337);
xnor U9505 (N_9505,N_9335,N_9344);
nand U9506 (N_9506,N_9395,N_9440);
and U9507 (N_9507,N_9427,N_9315);
and U9508 (N_9508,N_9370,N_9327);
nor U9509 (N_9509,N_9362,N_9426);
and U9510 (N_9510,N_9417,N_9368);
and U9511 (N_9511,N_9443,N_9416);
and U9512 (N_9512,N_9432,N_9329);
or U9513 (N_9513,N_9350,N_9328);
or U9514 (N_9514,N_9396,N_9424);
or U9515 (N_9515,N_9320,N_9360);
or U9516 (N_9516,N_9425,N_9402);
xnor U9517 (N_9517,N_9393,N_9300);
xnor U9518 (N_9518,N_9447,N_9446);
nor U9519 (N_9519,N_9369,N_9311);
nor U9520 (N_9520,N_9348,N_9340);
or U9521 (N_9521,N_9347,N_9345);
and U9522 (N_9522,N_9434,N_9389);
and U9523 (N_9523,N_9318,N_9313);
and U9524 (N_9524,N_9341,N_9367);
or U9525 (N_9525,N_9358,N_9304);
nand U9526 (N_9526,N_9435,N_9335);
and U9527 (N_9527,N_9322,N_9444);
xor U9528 (N_9528,N_9422,N_9440);
xor U9529 (N_9529,N_9315,N_9412);
and U9530 (N_9530,N_9400,N_9437);
xor U9531 (N_9531,N_9405,N_9352);
or U9532 (N_9532,N_9443,N_9424);
xnor U9533 (N_9533,N_9371,N_9393);
xor U9534 (N_9534,N_9408,N_9383);
nand U9535 (N_9535,N_9432,N_9426);
xor U9536 (N_9536,N_9440,N_9329);
xor U9537 (N_9537,N_9356,N_9413);
nand U9538 (N_9538,N_9436,N_9334);
xor U9539 (N_9539,N_9393,N_9430);
or U9540 (N_9540,N_9427,N_9389);
xor U9541 (N_9541,N_9322,N_9393);
nand U9542 (N_9542,N_9411,N_9332);
xnor U9543 (N_9543,N_9382,N_9323);
xnor U9544 (N_9544,N_9322,N_9398);
nand U9545 (N_9545,N_9417,N_9303);
or U9546 (N_9546,N_9405,N_9433);
and U9547 (N_9547,N_9412,N_9426);
nand U9548 (N_9548,N_9338,N_9428);
xor U9549 (N_9549,N_9376,N_9350);
nor U9550 (N_9550,N_9342,N_9361);
xnor U9551 (N_9551,N_9339,N_9316);
nand U9552 (N_9552,N_9363,N_9350);
or U9553 (N_9553,N_9358,N_9330);
or U9554 (N_9554,N_9413,N_9426);
nor U9555 (N_9555,N_9309,N_9378);
nand U9556 (N_9556,N_9320,N_9342);
and U9557 (N_9557,N_9426,N_9302);
and U9558 (N_9558,N_9448,N_9326);
and U9559 (N_9559,N_9311,N_9348);
or U9560 (N_9560,N_9436,N_9304);
xnor U9561 (N_9561,N_9448,N_9325);
and U9562 (N_9562,N_9400,N_9409);
nor U9563 (N_9563,N_9301,N_9339);
and U9564 (N_9564,N_9310,N_9370);
and U9565 (N_9565,N_9309,N_9355);
xnor U9566 (N_9566,N_9314,N_9334);
or U9567 (N_9567,N_9385,N_9424);
xnor U9568 (N_9568,N_9312,N_9303);
nand U9569 (N_9569,N_9347,N_9393);
xnor U9570 (N_9570,N_9398,N_9307);
xnor U9571 (N_9571,N_9386,N_9411);
xor U9572 (N_9572,N_9400,N_9324);
and U9573 (N_9573,N_9438,N_9324);
nor U9574 (N_9574,N_9358,N_9394);
nor U9575 (N_9575,N_9342,N_9441);
and U9576 (N_9576,N_9305,N_9378);
and U9577 (N_9577,N_9316,N_9328);
or U9578 (N_9578,N_9336,N_9395);
nand U9579 (N_9579,N_9340,N_9449);
nor U9580 (N_9580,N_9418,N_9389);
and U9581 (N_9581,N_9441,N_9303);
xnor U9582 (N_9582,N_9325,N_9394);
nand U9583 (N_9583,N_9341,N_9445);
nand U9584 (N_9584,N_9402,N_9422);
nand U9585 (N_9585,N_9424,N_9384);
nand U9586 (N_9586,N_9339,N_9406);
nor U9587 (N_9587,N_9355,N_9439);
nand U9588 (N_9588,N_9361,N_9302);
or U9589 (N_9589,N_9425,N_9342);
xor U9590 (N_9590,N_9350,N_9425);
nor U9591 (N_9591,N_9404,N_9441);
nand U9592 (N_9592,N_9356,N_9360);
and U9593 (N_9593,N_9433,N_9348);
nor U9594 (N_9594,N_9344,N_9305);
and U9595 (N_9595,N_9448,N_9430);
xnor U9596 (N_9596,N_9310,N_9375);
nand U9597 (N_9597,N_9314,N_9355);
and U9598 (N_9598,N_9413,N_9306);
nor U9599 (N_9599,N_9444,N_9438);
nand U9600 (N_9600,N_9553,N_9518);
nand U9601 (N_9601,N_9515,N_9569);
nor U9602 (N_9602,N_9597,N_9501);
or U9603 (N_9603,N_9591,N_9592);
or U9604 (N_9604,N_9588,N_9546);
nand U9605 (N_9605,N_9551,N_9598);
nor U9606 (N_9606,N_9530,N_9468);
and U9607 (N_9607,N_9487,N_9581);
xor U9608 (N_9608,N_9472,N_9480);
nand U9609 (N_9609,N_9579,N_9478);
or U9610 (N_9610,N_9524,N_9491);
or U9611 (N_9611,N_9574,N_9525);
nand U9612 (N_9612,N_9458,N_9531);
nor U9613 (N_9613,N_9453,N_9513);
xor U9614 (N_9614,N_9482,N_9502);
or U9615 (N_9615,N_9547,N_9465);
or U9616 (N_9616,N_9532,N_9589);
nor U9617 (N_9617,N_9537,N_9507);
nand U9618 (N_9618,N_9457,N_9576);
nand U9619 (N_9619,N_9549,N_9466);
nor U9620 (N_9620,N_9464,N_9511);
xnor U9621 (N_9621,N_9490,N_9586);
and U9622 (N_9622,N_9562,N_9554);
or U9623 (N_9623,N_9583,N_9528);
xor U9624 (N_9624,N_9560,N_9508);
or U9625 (N_9625,N_9477,N_9523);
xnor U9626 (N_9626,N_9534,N_9595);
nand U9627 (N_9627,N_9570,N_9460);
nor U9628 (N_9628,N_9493,N_9454);
nor U9629 (N_9629,N_9517,N_9563);
nor U9630 (N_9630,N_9526,N_9527);
xnor U9631 (N_9631,N_9566,N_9559);
nor U9632 (N_9632,N_9471,N_9599);
xor U9633 (N_9633,N_9498,N_9486);
nand U9634 (N_9634,N_9473,N_9529);
and U9635 (N_9635,N_9536,N_9485);
nor U9636 (N_9636,N_9461,N_9594);
or U9637 (N_9637,N_9535,N_9561);
nor U9638 (N_9638,N_9555,N_9504);
and U9639 (N_9639,N_9481,N_9470);
and U9640 (N_9640,N_9548,N_9462);
xor U9641 (N_9641,N_9512,N_9575);
nand U9642 (N_9642,N_9538,N_9567);
nor U9643 (N_9643,N_9520,N_9488);
and U9644 (N_9644,N_9541,N_9494);
and U9645 (N_9645,N_9545,N_9483);
or U9646 (N_9646,N_9571,N_9543);
and U9647 (N_9647,N_9557,N_9542);
nand U9648 (N_9648,N_9452,N_9533);
nand U9649 (N_9649,N_9578,N_9587);
and U9650 (N_9650,N_9564,N_9556);
nor U9651 (N_9651,N_9585,N_9572);
nand U9652 (N_9652,N_9580,N_9476);
nor U9653 (N_9653,N_9474,N_9495);
nand U9654 (N_9654,N_9484,N_9496);
xnor U9655 (N_9655,N_9459,N_9497);
or U9656 (N_9656,N_9582,N_9514);
xor U9657 (N_9657,N_9467,N_9522);
xnor U9658 (N_9658,N_9584,N_9565);
xor U9659 (N_9659,N_9503,N_9521);
nand U9660 (N_9660,N_9463,N_9596);
and U9661 (N_9661,N_9455,N_9475);
xnor U9662 (N_9662,N_9544,N_9492);
or U9663 (N_9663,N_9509,N_9505);
xor U9664 (N_9664,N_9516,N_9519);
nand U9665 (N_9665,N_9577,N_9540);
nor U9666 (N_9666,N_9450,N_9593);
or U9667 (N_9667,N_9539,N_9590);
xnor U9668 (N_9668,N_9499,N_9456);
and U9669 (N_9669,N_9451,N_9552);
nand U9670 (N_9670,N_9568,N_9500);
xor U9671 (N_9671,N_9510,N_9469);
or U9672 (N_9672,N_9506,N_9489);
xor U9673 (N_9673,N_9573,N_9550);
xnor U9674 (N_9674,N_9479,N_9558);
or U9675 (N_9675,N_9452,N_9527);
nor U9676 (N_9676,N_9507,N_9541);
nor U9677 (N_9677,N_9465,N_9561);
and U9678 (N_9678,N_9599,N_9486);
xnor U9679 (N_9679,N_9555,N_9565);
xor U9680 (N_9680,N_9550,N_9560);
and U9681 (N_9681,N_9579,N_9556);
xor U9682 (N_9682,N_9491,N_9501);
nor U9683 (N_9683,N_9584,N_9567);
and U9684 (N_9684,N_9491,N_9451);
nor U9685 (N_9685,N_9542,N_9585);
and U9686 (N_9686,N_9551,N_9532);
and U9687 (N_9687,N_9497,N_9466);
xor U9688 (N_9688,N_9484,N_9471);
nor U9689 (N_9689,N_9468,N_9495);
nand U9690 (N_9690,N_9560,N_9599);
xor U9691 (N_9691,N_9585,N_9489);
nor U9692 (N_9692,N_9497,N_9533);
or U9693 (N_9693,N_9482,N_9596);
nor U9694 (N_9694,N_9482,N_9497);
and U9695 (N_9695,N_9554,N_9486);
nand U9696 (N_9696,N_9534,N_9553);
nor U9697 (N_9697,N_9487,N_9517);
or U9698 (N_9698,N_9450,N_9555);
nor U9699 (N_9699,N_9581,N_9481);
and U9700 (N_9700,N_9462,N_9510);
or U9701 (N_9701,N_9494,N_9549);
and U9702 (N_9702,N_9571,N_9506);
and U9703 (N_9703,N_9559,N_9588);
nand U9704 (N_9704,N_9569,N_9592);
nor U9705 (N_9705,N_9563,N_9562);
and U9706 (N_9706,N_9480,N_9464);
xnor U9707 (N_9707,N_9468,N_9594);
nand U9708 (N_9708,N_9481,N_9527);
xnor U9709 (N_9709,N_9592,N_9593);
nand U9710 (N_9710,N_9471,N_9475);
nand U9711 (N_9711,N_9538,N_9547);
xor U9712 (N_9712,N_9531,N_9467);
or U9713 (N_9713,N_9587,N_9527);
xnor U9714 (N_9714,N_9495,N_9565);
nand U9715 (N_9715,N_9543,N_9511);
xnor U9716 (N_9716,N_9467,N_9507);
or U9717 (N_9717,N_9596,N_9590);
xnor U9718 (N_9718,N_9598,N_9586);
nand U9719 (N_9719,N_9490,N_9567);
or U9720 (N_9720,N_9514,N_9533);
or U9721 (N_9721,N_9556,N_9558);
nand U9722 (N_9722,N_9565,N_9545);
nor U9723 (N_9723,N_9513,N_9516);
or U9724 (N_9724,N_9495,N_9473);
nand U9725 (N_9725,N_9599,N_9480);
and U9726 (N_9726,N_9549,N_9554);
nand U9727 (N_9727,N_9553,N_9450);
or U9728 (N_9728,N_9492,N_9519);
nand U9729 (N_9729,N_9535,N_9504);
nor U9730 (N_9730,N_9578,N_9576);
nand U9731 (N_9731,N_9467,N_9597);
and U9732 (N_9732,N_9574,N_9532);
or U9733 (N_9733,N_9552,N_9567);
or U9734 (N_9734,N_9501,N_9529);
xor U9735 (N_9735,N_9514,N_9597);
or U9736 (N_9736,N_9595,N_9477);
nand U9737 (N_9737,N_9464,N_9596);
nand U9738 (N_9738,N_9523,N_9484);
nand U9739 (N_9739,N_9549,N_9553);
nand U9740 (N_9740,N_9560,N_9501);
nand U9741 (N_9741,N_9547,N_9501);
nor U9742 (N_9742,N_9499,N_9523);
or U9743 (N_9743,N_9458,N_9520);
or U9744 (N_9744,N_9497,N_9523);
xnor U9745 (N_9745,N_9592,N_9557);
nor U9746 (N_9746,N_9512,N_9543);
xnor U9747 (N_9747,N_9582,N_9581);
nand U9748 (N_9748,N_9577,N_9508);
nand U9749 (N_9749,N_9463,N_9556);
nand U9750 (N_9750,N_9696,N_9749);
or U9751 (N_9751,N_9672,N_9730);
nor U9752 (N_9752,N_9745,N_9654);
and U9753 (N_9753,N_9665,N_9733);
nor U9754 (N_9754,N_9617,N_9616);
or U9755 (N_9755,N_9693,N_9661);
xor U9756 (N_9756,N_9604,N_9622);
xnor U9757 (N_9757,N_9653,N_9615);
xor U9758 (N_9758,N_9744,N_9664);
xor U9759 (N_9759,N_9704,N_9640);
xor U9760 (N_9760,N_9658,N_9729);
nor U9761 (N_9761,N_9614,N_9705);
xor U9762 (N_9762,N_9700,N_9692);
and U9763 (N_9763,N_9608,N_9699);
xnor U9764 (N_9764,N_9725,N_9674);
and U9765 (N_9765,N_9748,N_9621);
and U9766 (N_9766,N_9659,N_9600);
or U9767 (N_9767,N_9710,N_9723);
nor U9768 (N_9768,N_9635,N_9642);
or U9769 (N_9769,N_9734,N_9645);
nand U9770 (N_9770,N_9668,N_9629);
nand U9771 (N_9771,N_9686,N_9690);
and U9772 (N_9772,N_9666,N_9646);
xnor U9773 (N_9773,N_9721,N_9648);
or U9774 (N_9774,N_9619,N_9660);
or U9775 (N_9775,N_9667,N_9663);
nand U9776 (N_9776,N_9746,N_9689);
and U9777 (N_9777,N_9605,N_9650);
xor U9778 (N_9778,N_9682,N_9633);
or U9779 (N_9779,N_9630,N_9688);
nand U9780 (N_9780,N_9687,N_9694);
xor U9781 (N_9781,N_9740,N_9736);
xnor U9782 (N_9782,N_9739,N_9742);
nand U9783 (N_9783,N_9601,N_9631);
xnor U9784 (N_9784,N_9612,N_9683);
and U9785 (N_9785,N_9677,N_9670);
and U9786 (N_9786,N_9662,N_9716);
or U9787 (N_9787,N_9711,N_9675);
nor U9788 (N_9788,N_9735,N_9620);
nand U9789 (N_9789,N_9647,N_9657);
nand U9790 (N_9790,N_9634,N_9718);
xor U9791 (N_9791,N_9698,N_9644);
and U9792 (N_9792,N_9691,N_9623);
nor U9793 (N_9793,N_9606,N_9603);
or U9794 (N_9794,N_9697,N_9656);
xor U9795 (N_9795,N_9643,N_9714);
nand U9796 (N_9796,N_9715,N_9637);
or U9797 (N_9797,N_9717,N_9652);
and U9798 (N_9798,N_9673,N_9671);
xor U9799 (N_9799,N_9679,N_9624);
and U9800 (N_9800,N_9726,N_9607);
or U9801 (N_9801,N_9611,N_9722);
xor U9802 (N_9802,N_9706,N_9641);
nor U9803 (N_9803,N_9669,N_9684);
and U9804 (N_9804,N_9731,N_9713);
nand U9805 (N_9805,N_9685,N_9695);
or U9806 (N_9806,N_9732,N_9618);
xnor U9807 (N_9807,N_9639,N_9613);
or U9808 (N_9808,N_9627,N_9702);
nor U9809 (N_9809,N_9626,N_9708);
xor U9810 (N_9810,N_9727,N_9707);
xor U9811 (N_9811,N_9747,N_9712);
xor U9812 (N_9812,N_9709,N_9741);
xor U9813 (N_9813,N_9738,N_9681);
nand U9814 (N_9814,N_9720,N_9737);
nand U9815 (N_9815,N_9636,N_9676);
and U9816 (N_9816,N_9602,N_9743);
xnor U9817 (N_9817,N_9680,N_9609);
xor U9818 (N_9818,N_9678,N_9651);
nor U9819 (N_9819,N_9724,N_9649);
nor U9820 (N_9820,N_9701,N_9610);
nor U9821 (N_9821,N_9632,N_9703);
or U9822 (N_9822,N_9655,N_9625);
or U9823 (N_9823,N_9728,N_9719);
and U9824 (N_9824,N_9628,N_9638);
xnor U9825 (N_9825,N_9743,N_9722);
xnor U9826 (N_9826,N_9738,N_9711);
xnor U9827 (N_9827,N_9691,N_9708);
xor U9828 (N_9828,N_9689,N_9629);
xnor U9829 (N_9829,N_9661,N_9614);
xor U9830 (N_9830,N_9694,N_9742);
nor U9831 (N_9831,N_9649,N_9629);
xnor U9832 (N_9832,N_9700,N_9735);
and U9833 (N_9833,N_9616,N_9672);
or U9834 (N_9834,N_9642,N_9736);
nor U9835 (N_9835,N_9636,N_9741);
or U9836 (N_9836,N_9662,N_9651);
xor U9837 (N_9837,N_9744,N_9725);
nand U9838 (N_9838,N_9666,N_9738);
nand U9839 (N_9839,N_9666,N_9680);
and U9840 (N_9840,N_9635,N_9647);
or U9841 (N_9841,N_9720,N_9749);
or U9842 (N_9842,N_9741,N_9645);
nand U9843 (N_9843,N_9741,N_9640);
nand U9844 (N_9844,N_9611,N_9616);
xor U9845 (N_9845,N_9695,N_9623);
nor U9846 (N_9846,N_9602,N_9746);
or U9847 (N_9847,N_9617,N_9693);
nor U9848 (N_9848,N_9661,N_9680);
nor U9849 (N_9849,N_9742,N_9717);
xnor U9850 (N_9850,N_9691,N_9711);
or U9851 (N_9851,N_9696,N_9699);
and U9852 (N_9852,N_9607,N_9622);
and U9853 (N_9853,N_9734,N_9650);
nand U9854 (N_9854,N_9601,N_9713);
xor U9855 (N_9855,N_9627,N_9615);
nand U9856 (N_9856,N_9747,N_9624);
xnor U9857 (N_9857,N_9680,N_9603);
or U9858 (N_9858,N_9662,N_9626);
nand U9859 (N_9859,N_9624,N_9746);
and U9860 (N_9860,N_9613,N_9712);
nand U9861 (N_9861,N_9674,N_9717);
or U9862 (N_9862,N_9649,N_9610);
and U9863 (N_9863,N_9742,N_9740);
or U9864 (N_9864,N_9643,N_9716);
xnor U9865 (N_9865,N_9713,N_9728);
nand U9866 (N_9866,N_9608,N_9709);
or U9867 (N_9867,N_9651,N_9669);
nor U9868 (N_9868,N_9688,N_9641);
or U9869 (N_9869,N_9667,N_9652);
and U9870 (N_9870,N_9695,N_9702);
or U9871 (N_9871,N_9746,N_9728);
nor U9872 (N_9872,N_9712,N_9629);
xnor U9873 (N_9873,N_9617,N_9661);
or U9874 (N_9874,N_9605,N_9643);
and U9875 (N_9875,N_9624,N_9608);
nand U9876 (N_9876,N_9694,N_9659);
nor U9877 (N_9877,N_9715,N_9630);
nand U9878 (N_9878,N_9697,N_9647);
nand U9879 (N_9879,N_9696,N_9626);
and U9880 (N_9880,N_9647,N_9607);
xnor U9881 (N_9881,N_9722,N_9746);
or U9882 (N_9882,N_9728,N_9674);
xor U9883 (N_9883,N_9622,N_9749);
and U9884 (N_9884,N_9676,N_9656);
xor U9885 (N_9885,N_9629,N_9672);
or U9886 (N_9886,N_9630,N_9720);
or U9887 (N_9887,N_9749,N_9632);
xor U9888 (N_9888,N_9660,N_9704);
or U9889 (N_9889,N_9661,N_9741);
xnor U9890 (N_9890,N_9685,N_9610);
nor U9891 (N_9891,N_9640,N_9721);
or U9892 (N_9892,N_9685,N_9633);
or U9893 (N_9893,N_9627,N_9622);
nor U9894 (N_9894,N_9664,N_9722);
nor U9895 (N_9895,N_9716,N_9637);
xor U9896 (N_9896,N_9608,N_9706);
nor U9897 (N_9897,N_9611,N_9731);
or U9898 (N_9898,N_9714,N_9651);
nand U9899 (N_9899,N_9735,N_9627);
xnor U9900 (N_9900,N_9806,N_9801);
xnor U9901 (N_9901,N_9858,N_9846);
xor U9902 (N_9902,N_9898,N_9784);
nor U9903 (N_9903,N_9787,N_9766);
nor U9904 (N_9904,N_9881,N_9830);
nor U9905 (N_9905,N_9757,N_9767);
nor U9906 (N_9906,N_9793,N_9847);
xor U9907 (N_9907,N_9843,N_9820);
or U9908 (N_9908,N_9837,N_9781);
xor U9909 (N_9909,N_9796,N_9777);
and U9910 (N_9910,N_9782,N_9877);
nand U9911 (N_9911,N_9758,N_9822);
or U9912 (N_9912,N_9826,N_9788);
and U9913 (N_9913,N_9870,N_9809);
nor U9914 (N_9914,N_9896,N_9869);
nand U9915 (N_9915,N_9827,N_9761);
and U9916 (N_9916,N_9802,N_9867);
xor U9917 (N_9917,N_9885,N_9791);
or U9918 (N_9918,N_9813,N_9875);
xnor U9919 (N_9919,N_9855,N_9840);
or U9920 (N_9920,N_9882,N_9798);
nor U9921 (N_9921,N_9818,N_9889);
xor U9922 (N_9922,N_9799,N_9763);
or U9923 (N_9923,N_9841,N_9772);
nand U9924 (N_9924,N_9829,N_9751);
nand U9925 (N_9925,N_9764,N_9880);
or U9926 (N_9926,N_9895,N_9849);
xnor U9927 (N_9927,N_9862,N_9760);
or U9928 (N_9928,N_9828,N_9823);
xor U9929 (N_9929,N_9807,N_9783);
nand U9930 (N_9930,N_9871,N_9812);
nor U9931 (N_9931,N_9824,N_9831);
and U9932 (N_9932,N_9868,N_9892);
nand U9933 (N_9933,N_9842,N_9886);
and U9934 (N_9934,N_9794,N_9817);
xnor U9935 (N_9935,N_9861,N_9891);
xnor U9936 (N_9936,N_9883,N_9753);
or U9937 (N_9937,N_9863,N_9878);
or U9938 (N_9938,N_9851,N_9765);
nand U9939 (N_9939,N_9779,N_9859);
xnor U9940 (N_9940,N_9852,N_9810);
nand U9941 (N_9941,N_9775,N_9872);
and U9942 (N_9942,N_9771,N_9795);
and U9943 (N_9943,N_9884,N_9808);
or U9944 (N_9944,N_9857,N_9821);
or U9945 (N_9945,N_9769,N_9825);
nor U9946 (N_9946,N_9819,N_9792);
nor U9947 (N_9947,N_9897,N_9816);
nor U9948 (N_9948,N_9836,N_9768);
or U9949 (N_9949,N_9856,N_9860);
or U9950 (N_9950,N_9773,N_9845);
nand U9951 (N_9951,N_9879,N_9814);
or U9952 (N_9952,N_9864,N_9839);
nor U9953 (N_9953,N_9844,N_9759);
and U9954 (N_9954,N_9899,N_9838);
xnor U9955 (N_9955,N_9774,N_9850);
nand U9956 (N_9956,N_9754,N_9876);
nor U9957 (N_9957,N_9800,N_9832);
or U9958 (N_9958,N_9797,N_9805);
xnor U9959 (N_9959,N_9785,N_9887);
nor U9960 (N_9960,N_9894,N_9789);
nand U9961 (N_9961,N_9835,N_9890);
nand U9962 (N_9962,N_9755,N_9762);
and U9963 (N_9963,N_9815,N_9770);
nand U9964 (N_9964,N_9811,N_9803);
nor U9965 (N_9965,N_9848,N_9804);
xnor U9966 (N_9966,N_9874,N_9786);
xnor U9967 (N_9967,N_9752,N_9756);
xnor U9968 (N_9968,N_9778,N_9888);
and U9969 (N_9969,N_9854,N_9790);
nand U9970 (N_9970,N_9865,N_9893);
nand U9971 (N_9971,N_9833,N_9776);
nand U9972 (N_9972,N_9873,N_9780);
xnor U9973 (N_9973,N_9866,N_9834);
nand U9974 (N_9974,N_9750,N_9853);
or U9975 (N_9975,N_9839,N_9788);
nor U9976 (N_9976,N_9768,N_9779);
xnor U9977 (N_9977,N_9822,N_9886);
and U9978 (N_9978,N_9770,N_9810);
xor U9979 (N_9979,N_9870,N_9795);
nand U9980 (N_9980,N_9769,N_9805);
xor U9981 (N_9981,N_9856,N_9812);
nor U9982 (N_9982,N_9872,N_9810);
nand U9983 (N_9983,N_9805,N_9775);
nor U9984 (N_9984,N_9892,N_9894);
nand U9985 (N_9985,N_9751,N_9890);
nor U9986 (N_9986,N_9801,N_9856);
nor U9987 (N_9987,N_9875,N_9854);
and U9988 (N_9988,N_9805,N_9819);
nor U9989 (N_9989,N_9825,N_9883);
or U9990 (N_9990,N_9782,N_9887);
nor U9991 (N_9991,N_9888,N_9802);
nand U9992 (N_9992,N_9763,N_9856);
nor U9993 (N_9993,N_9784,N_9890);
or U9994 (N_9994,N_9830,N_9768);
nor U9995 (N_9995,N_9821,N_9756);
or U9996 (N_9996,N_9800,N_9835);
nor U9997 (N_9997,N_9824,N_9776);
xor U9998 (N_9998,N_9806,N_9868);
and U9999 (N_9999,N_9831,N_9757);
and U10000 (N_10000,N_9897,N_9810);
nand U10001 (N_10001,N_9864,N_9849);
and U10002 (N_10002,N_9817,N_9770);
nand U10003 (N_10003,N_9757,N_9827);
or U10004 (N_10004,N_9789,N_9760);
nand U10005 (N_10005,N_9879,N_9778);
xor U10006 (N_10006,N_9762,N_9780);
nor U10007 (N_10007,N_9814,N_9768);
nor U10008 (N_10008,N_9822,N_9862);
nand U10009 (N_10009,N_9861,N_9886);
and U10010 (N_10010,N_9787,N_9859);
or U10011 (N_10011,N_9837,N_9783);
xnor U10012 (N_10012,N_9814,N_9897);
xor U10013 (N_10013,N_9838,N_9780);
or U10014 (N_10014,N_9896,N_9755);
or U10015 (N_10015,N_9766,N_9827);
nor U10016 (N_10016,N_9769,N_9792);
and U10017 (N_10017,N_9839,N_9754);
and U10018 (N_10018,N_9845,N_9880);
nor U10019 (N_10019,N_9795,N_9878);
xor U10020 (N_10020,N_9750,N_9759);
nor U10021 (N_10021,N_9855,N_9853);
nor U10022 (N_10022,N_9828,N_9784);
and U10023 (N_10023,N_9834,N_9751);
nor U10024 (N_10024,N_9799,N_9766);
nor U10025 (N_10025,N_9841,N_9759);
and U10026 (N_10026,N_9776,N_9755);
or U10027 (N_10027,N_9797,N_9793);
or U10028 (N_10028,N_9846,N_9871);
and U10029 (N_10029,N_9828,N_9850);
xnor U10030 (N_10030,N_9856,N_9754);
or U10031 (N_10031,N_9791,N_9861);
nand U10032 (N_10032,N_9822,N_9776);
xor U10033 (N_10033,N_9850,N_9860);
nor U10034 (N_10034,N_9882,N_9850);
nor U10035 (N_10035,N_9886,N_9817);
nand U10036 (N_10036,N_9877,N_9838);
xnor U10037 (N_10037,N_9784,N_9873);
or U10038 (N_10038,N_9776,N_9843);
nor U10039 (N_10039,N_9812,N_9823);
nand U10040 (N_10040,N_9804,N_9761);
xor U10041 (N_10041,N_9765,N_9773);
nor U10042 (N_10042,N_9828,N_9795);
nand U10043 (N_10043,N_9828,N_9768);
nor U10044 (N_10044,N_9881,N_9866);
xnor U10045 (N_10045,N_9894,N_9874);
xor U10046 (N_10046,N_9876,N_9775);
or U10047 (N_10047,N_9870,N_9789);
nand U10048 (N_10048,N_9890,N_9758);
xor U10049 (N_10049,N_9780,N_9759);
nand U10050 (N_10050,N_9970,N_10020);
or U10051 (N_10051,N_10032,N_9916);
and U10052 (N_10052,N_9963,N_9959);
nand U10053 (N_10053,N_9977,N_9960);
and U10054 (N_10054,N_9902,N_10046);
xnor U10055 (N_10055,N_9929,N_10017);
and U10056 (N_10056,N_10021,N_9941);
xnor U10057 (N_10057,N_9913,N_9952);
and U10058 (N_10058,N_10004,N_9914);
xor U10059 (N_10059,N_9904,N_9987);
nand U10060 (N_10060,N_10009,N_9989);
and U10061 (N_10061,N_9974,N_9908);
and U10062 (N_10062,N_10002,N_10019);
or U10063 (N_10063,N_9969,N_9936);
nor U10064 (N_10064,N_10012,N_9957);
or U10065 (N_10065,N_10005,N_10043);
nand U10066 (N_10066,N_9967,N_9910);
nor U10067 (N_10067,N_9998,N_9915);
and U10068 (N_10068,N_9947,N_9938);
xnor U10069 (N_10069,N_9940,N_10047);
and U10070 (N_10070,N_10015,N_10029);
nor U10071 (N_10071,N_9925,N_10036);
nor U10072 (N_10072,N_9922,N_10006);
xor U10073 (N_10073,N_9921,N_10010);
or U10074 (N_10074,N_10023,N_9979);
and U10075 (N_10075,N_9971,N_9991);
nor U10076 (N_10076,N_9999,N_9958);
nor U10077 (N_10077,N_10022,N_9996);
xor U10078 (N_10078,N_9988,N_10007);
or U10079 (N_10079,N_9945,N_9911);
xnor U10080 (N_10080,N_9990,N_9964);
or U10081 (N_10081,N_9955,N_9939);
nor U10082 (N_10082,N_9912,N_9965);
nor U10083 (N_10083,N_9924,N_9909);
nand U10084 (N_10084,N_9944,N_9994);
nand U10085 (N_10085,N_10044,N_10041);
xnor U10086 (N_10086,N_9950,N_10033);
and U10087 (N_10087,N_10014,N_10045);
nor U10088 (N_10088,N_10024,N_10040);
and U10089 (N_10089,N_9997,N_9962);
xor U10090 (N_10090,N_9961,N_10027);
or U10091 (N_10091,N_9973,N_9978);
nor U10092 (N_10092,N_9932,N_10011);
or U10093 (N_10093,N_9901,N_9943);
or U10094 (N_10094,N_9927,N_10037);
or U10095 (N_10095,N_9907,N_9953);
xnor U10096 (N_10096,N_10035,N_9917);
or U10097 (N_10097,N_9949,N_9946);
or U10098 (N_10098,N_10016,N_10042);
nor U10099 (N_10099,N_10038,N_10018);
and U10100 (N_10100,N_9956,N_10049);
and U10101 (N_10101,N_9934,N_9951);
nand U10102 (N_10102,N_9900,N_10026);
xnor U10103 (N_10103,N_9972,N_9976);
xor U10104 (N_10104,N_9933,N_9948);
or U10105 (N_10105,N_9935,N_10028);
nand U10106 (N_10106,N_10001,N_9918);
or U10107 (N_10107,N_9923,N_9942);
and U10108 (N_10108,N_10000,N_9986);
nand U10109 (N_10109,N_9931,N_9995);
nand U10110 (N_10110,N_10031,N_9993);
xor U10111 (N_10111,N_9928,N_9937);
and U10112 (N_10112,N_9968,N_9982);
and U10113 (N_10113,N_9980,N_9905);
or U10114 (N_10114,N_9926,N_9985);
nand U10115 (N_10115,N_9975,N_10008);
nor U10116 (N_10116,N_9966,N_10003);
nor U10117 (N_10117,N_9903,N_9992);
or U10118 (N_10118,N_9930,N_10034);
and U10119 (N_10119,N_9984,N_10013);
nor U10120 (N_10120,N_9906,N_10039);
nor U10121 (N_10121,N_9983,N_10025);
or U10122 (N_10122,N_10048,N_9920);
xnor U10123 (N_10123,N_9981,N_10030);
and U10124 (N_10124,N_9919,N_9954);
nand U10125 (N_10125,N_10028,N_9961);
and U10126 (N_10126,N_9952,N_10011);
or U10127 (N_10127,N_9905,N_10030);
xor U10128 (N_10128,N_9990,N_9989);
nand U10129 (N_10129,N_9909,N_9995);
and U10130 (N_10130,N_9977,N_9943);
nor U10131 (N_10131,N_9900,N_9993);
and U10132 (N_10132,N_9911,N_9984);
nor U10133 (N_10133,N_10023,N_9923);
or U10134 (N_10134,N_10042,N_9952);
or U10135 (N_10135,N_10026,N_9907);
nor U10136 (N_10136,N_9956,N_10011);
and U10137 (N_10137,N_9990,N_9994);
nor U10138 (N_10138,N_10016,N_9906);
nand U10139 (N_10139,N_9975,N_9956);
and U10140 (N_10140,N_10000,N_10007);
and U10141 (N_10141,N_9953,N_9955);
nor U10142 (N_10142,N_10035,N_9925);
or U10143 (N_10143,N_10036,N_9986);
xnor U10144 (N_10144,N_9954,N_9943);
nand U10145 (N_10145,N_10037,N_9909);
or U10146 (N_10146,N_9903,N_9972);
and U10147 (N_10147,N_9906,N_9975);
nand U10148 (N_10148,N_9994,N_10005);
and U10149 (N_10149,N_9903,N_9934);
nor U10150 (N_10150,N_9985,N_10024);
nand U10151 (N_10151,N_10028,N_10043);
and U10152 (N_10152,N_9906,N_9961);
nand U10153 (N_10153,N_10009,N_10030);
xor U10154 (N_10154,N_9934,N_10036);
xnor U10155 (N_10155,N_9975,N_10043);
and U10156 (N_10156,N_9916,N_9929);
nor U10157 (N_10157,N_9982,N_9901);
and U10158 (N_10158,N_9964,N_9985);
nor U10159 (N_10159,N_10003,N_10006);
and U10160 (N_10160,N_9959,N_10015);
or U10161 (N_10161,N_10036,N_9960);
or U10162 (N_10162,N_9906,N_9909);
nor U10163 (N_10163,N_9986,N_9962);
nor U10164 (N_10164,N_10012,N_10006);
or U10165 (N_10165,N_10000,N_9978);
nand U10166 (N_10166,N_9955,N_9994);
nand U10167 (N_10167,N_10039,N_9971);
xor U10168 (N_10168,N_10037,N_9956);
or U10169 (N_10169,N_10039,N_9952);
nor U10170 (N_10170,N_9914,N_10023);
and U10171 (N_10171,N_10049,N_9998);
xor U10172 (N_10172,N_9925,N_9934);
or U10173 (N_10173,N_9979,N_10032);
nor U10174 (N_10174,N_9989,N_10046);
xnor U10175 (N_10175,N_10019,N_9997);
and U10176 (N_10176,N_9909,N_9923);
nand U10177 (N_10177,N_10032,N_9935);
and U10178 (N_10178,N_10021,N_9924);
xor U10179 (N_10179,N_9926,N_10017);
nand U10180 (N_10180,N_10035,N_10021);
xor U10181 (N_10181,N_9911,N_9946);
or U10182 (N_10182,N_9915,N_10047);
and U10183 (N_10183,N_9976,N_10000);
nand U10184 (N_10184,N_9928,N_9988);
and U10185 (N_10185,N_10038,N_9919);
nand U10186 (N_10186,N_10045,N_10025);
or U10187 (N_10187,N_9914,N_9954);
xor U10188 (N_10188,N_10046,N_9964);
xnor U10189 (N_10189,N_9949,N_9928);
or U10190 (N_10190,N_9969,N_9981);
nand U10191 (N_10191,N_9923,N_9962);
nand U10192 (N_10192,N_9925,N_9940);
xnor U10193 (N_10193,N_10007,N_9948);
and U10194 (N_10194,N_10019,N_10042);
nand U10195 (N_10195,N_9916,N_9997);
nand U10196 (N_10196,N_9943,N_9937);
nand U10197 (N_10197,N_10045,N_10041);
xor U10198 (N_10198,N_9975,N_9938);
and U10199 (N_10199,N_9926,N_10015);
nor U10200 (N_10200,N_10083,N_10162);
nor U10201 (N_10201,N_10126,N_10120);
or U10202 (N_10202,N_10087,N_10165);
or U10203 (N_10203,N_10081,N_10157);
and U10204 (N_10204,N_10089,N_10176);
nand U10205 (N_10205,N_10128,N_10102);
nor U10206 (N_10206,N_10186,N_10160);
nor U10207 (N_10207,N_10183,N_10057);
and U10208 (N_10208,N_10151,N_10148);
nor U10209 (N_10209,N_10194,N_10184);
and U10210 (N_10210,N_10132,N_10153);
nor U10211 (N_10211,N_10065,N_10054);
and U10212 (N_10212,N_10067,N_10117);
or U10213 (N_10213,N_10091,N_10105);
nand U10214 (N_10214,N_10191,N_10199);
nand U10215 (N_10215,N_10115,N_10170);
nand U10216 (N_10216,N_10075,N_10125);
and U10217 (N_10217,N_10171,N_10192);
and U10218 (N_10218,N_10173,N_10142);
and U10219 (N_10219,N_10150,N_10093);
xor U10220 (N_10220,N_10156,N_10103);
or U10221 (N_10221,N_10124,N_10071);
or U10222 (N_10222,N_10082,N_10174);
or U10223 (N_10223,N_10092,N_10088);
xnor U10224 (N_10224,N_10069,N_10052);
xor U10225 (N_10225,N_10146,N_10189);
and U10226 (N_10226,N_10064,N_10050);
nor U10227 (N_10227,N_10159,N_10090);
or U10228 (N_10228,N_10169,N_10154);
nand U10229 (N_10229,N_10053,N_10166);
or U10230 (N_10230,N_10136,N_10110);
and U10231 (N_10231,N_10073,N_10133);
or U10232 (N_10232,N_10195,N_10063);
and U10233 (N_10233,N_10118,N_10143);
nand U10234 (N_10234,N_10163,N_10056);
nor U10235 (N_10235,N_10196,N_10178);
xnor U10236 (N_10236,N_10061,N_10188);
nor U10237 (N_10237,N_10101,N_10155);
xnor U10238 (N_10238,N_10167,N_10070);
xnor U10239 (N_10239,N_10137,N_10068);
nor U10240 (N_10240,N_10127,N_10152);
nor U10241 (N_10241,N_10121,N_10185);
nand U10242 (N_10242,N_10084,N_10107);
xor U10243 (N_10243,N_10190,N_10198);
nand U10244 (N_10244,N_10175,N_10096);
nand U10245 (N_10245,N_10079,N_10119);
nor U10246 (N_10246,N_10085,N_10179);
nand U10247 (N_10247,N_10177,N_10197);
and U10248 (N_10248,N_10078,N_10180);
and U10249 (N_10249,N_10097,N_10145);
nand U10250 (N_10250,N_10076,N_10111);
nor U10251 (N_10251,N_10066,N_10086);
nand U10252 (N_10252,N_10099,N_10080);
or U10253 (N_10253,N_10140,N_10077);
or U10254 (N_10254,N_10181,N_10109);
xnor U10255 (N_10255,N_10116,N_10164);
nand U10256 (N_10256,N_10141,N_10072);
nor U10257 (N_10257,N_10074,N_10131);
and U10258 (N_10258,N_10193,N_10055);
or U10259 (N_10259,N_10134,N_10135);
or U10260 (N_10260,N_10123,N_10138);
or U10261 (N_10261,N_10095,N_10100);
or U10262 (N_10262,N_10113,N_10168);
or U10263 (N_10263,N_10108,N_10187);
nand U10264 (N_10264,N_10112,N_10147);
xnor U10265 (N_10265,N_10130,N_10161);
xor U10266 (N_10266,N_10062,N_10058);
nand U10267 (N_10267,N_10060,N_10158);
or U10268 (N_10268,N_10106,N_10051);
or U10269 (N_10269,N_10098,N_10139);
nor U10270 (N_10270,N_10149,N_10144);
or U10271 (N_10271,N_10129,N_10059);
and U10272 (N_10272,N_10172,N_10114);
xnor U10273 (N_10273,N_10122,N_10094);
xor U10274 (N_10274,N_10182,N_10104);
nor U10275 (N_10275,N_10111,N_10118);
nor U10276 (N_10276,N_10129,N_10186);
nand U10277 (N_10277,N_10077,N_10142);
nand U10278 (N_10278,N_10077,N_10194);
and U10279 (N_10279,N_10138,N_10098);
or U10280 (N_10280,N_10194,N_10172);
xor U10281 (N_10281,N_10070,N_10191);
and U10282 (N_10282,N_10162,N_10109);
xor U10283 (N_10283,N_10085,N_10073);
or U10284 (N_10284,N_10136,N_10120);
nand U10285 (N_10285,N_10101,N_10123);
xor U10286 (N_10286,N_10190,N_10090);
or U10287 (N_10287,N_10055,N_10068);
and U10288 (N_10288,N_10072,N_10063);
xor U10289 (N_10289,N_10163,N_10103);
or U10290 (N_10290,N_10124,N_10108);
and U10291 (N_10291,N_10052,N_10176);
or U10292 (N_10292,N_10191,N_10163);
or U10293 (N_10293,N_10056,N_10122);
and U10294 (N_10294,N_10096,N_10155);
xnor U10295 (N_10295,N_10111,N_10153);
or U10296 (N_10296,N_10173,N_10169);
or U10297 (N_10297,N_10137,N_10130);
and U10298 (N_10298,N_10123,N_10142);
and U10299 (N_10299,N_10173,N_10102);
xnor U10300 (N_10300,N_10144,N_10061);
or U10301 (N_10301,N_10059,N_10153);
xnor U10302 (N_10302,N_10053,N_10082);
nor U10303 (N_10303,N_10140,N_10065);
and U10304 (N_10304,N_10147,N_10130);
nand U10305 (N_10305,N_10072,N_10180);
nor U10306 (N_10306,N_10121,N_10123);
and U10307 (N_10307,N_10157,N_10130);
nor U10308 (N_10308,N_10132,N_10121);
xor U10309 (N_10309,N_10169,N_10072);
and U10310 (N_10310,N_10162,N_10145);
nor U10311 (N_10311,N_10100,N_10156);
or U10312 (N_10312,N_10090,N_10107);
or U10313 (N_10313,N_10140,N_10073);
and U10314 (N_10314,N_10172,N_10076);
xor U10315 (N_10315,N_10176,N_10162);
nand U10316 (N_10316,N_10195,N_10072);
and U10317 (N_10317,N_10111,N_10117);
or U10318 (N_10318,N_10181,N_10074);
xnor U10319 (N_10319,N_10112,N_10085);
or U10320 (N_10320,N_10106,N_10093);
nor U10321 (N_10321,N_10133,N_10075);
nor U10322 (N_10322,N_10111,N_10120);
or U10323 (N_10323,N_10170,N_10108);
nor U10324 (N_10324,N_10089,N_10187);
xnor U10325 (N_10325,N_10155,N_10146);
nand U10326 (N_10326,N_10054,N_10102);
xor U10327 (N_10327,N_10073,N_10157);
nand U10328 (N_10328,N_10134,N_10059);
or U10329 (N_10329,N_10176,N_10164);
nand U10330 (N_10330,N_10159,N_10107);
xor U10331 (N_10331,N_10066,N_10070);
or U10332 (N_10332,N_10169,N_10141);
and U10333 (N_10333,N_10095,N_10138);
xor U10334 (N_10334,N_10080,N_10064);
nand U10335 (N_10335,N_10131,N_10127);
and U10336 (N_10336,N_10071,N_10190);
nor U10337 (N_10337,N_10152,N_10173);
and U10338 (N_10338,N_10141,N_10129);
and U10339 (N_10339,N_10153,N_10197);
xnor U10340 (N_10340,N_10072,N_10115);
xnor U10341 (N_10341,N_10069,N_10089);
nand U10342 (N_10342,N_10106,N_10098);
or U10343 (N_10343,N_10067,N_10082);
nand U10344 (N_10344,N_10116,N_10119);
xor U10345 (N_10345,N_10121,N_10199);
nor U10346 (N_10346,N_10145,N_10139);
and U10347 (N_10347,N_10050,N_10173);
nor U10348 (N_10348,N_10052,N_10061);
nor U10349 (N_10349,N_10066,N_10146);
and U10350 (N_10350,N_10281,N_10285);
or U10351 (N_10351,N_10279,N_10231);
and U10352 (N_10352,N_10277,N_10245);
and U10353 (N_10353,N_10236,N_10322);
and U10354 (N_10354,N_10297,N_10326);
nor U10355 (N_10355,N_10293,N_10205);
and U10356 (N_10356,N_10233,N_10278);
nand U10357 (N_10357,N_10266,N_10229);
xor U10358 (N_10358,N_10310,N_10335);
or U10359 (N_10359,N_10291,N_10287);
xnor U10360 (N_10360,N_10305,N_10276);
or U10361 (N_10361,N_10252,N_10224);
and U10362 (N_10362,N_10201,N_10210);
and U10363 (N_10363,N_10349,N_10294);
or U10364 (N_10364,N_10346,N_10304);
and U10365 (N_10365,N_10308,N_10216);
and U10366 (N_10366,N_10272,N_10317);
nand U10367 (N_10367,N_10264,N_10341);
or U10368 (N_10368,N_10220,N_10257);
or U10369 (N_10369,N_10267,N_10269);
nand U10370 (N_10370,N_10323,N_10347);
nand U10371 (N_10371,N_10280,N_10241);
and U10372 (N_10372,N_10208,N_10213);
and U10373 (N_10373,N_10343,N_10222);
nor U10374 (N_10374,N_10235,N_10329);
and U10375 (N_10375,N_10274,N_10301);
xnor U10376 (N_10376,N_10265,N_10250);
nor U10377 (N_10377,N_10258,N_10237);
xor U10378 (N_10378,N_10290,N_10249);
and U10379 (N_10379,N_10284,N_10247);
xor U10380 (N_10380,N_10340,N_10311);
nor U10381 (N_10381,N_10270,N_10243);
and U10382 (N_10382,N_10282,N_10336);
nor U10383 (N_10383,N_10215,N_10260);
nor U10384 (N_10384,N_10342,N_10292);
or U10385 (N_10385,N_10331,N_10300);
and U10386 (N_10386,N_10324,N_10228);
and U10387 (N_10387,N_10314,N_10295);
or U10388 (N_10388,N_10226,N_10338);
or U10389 (N_10389,N_10321,N_10303);
nor U10390 (N_10390,N_10313,N_10253);
or U10391 (N_10391,N_10289,N_10223);
or U10392 (N_10392,N_10254,N_10327);
and U10393 (N_10393,N_10296,N_10307);
and U10394 (N_10394,N_10319,N_10217);
xnor U10395 (N_10395,N_10242,N_10232);
xor U10396 (N_10396,N_10244,N_10309);
or U10397 (N_10397,N_10334,N_10200);
nand U10398 (N_10398,N_10339,N_10221);
xnor U10399 (N_10399,N_10344,N_10345);
nor U10400 (N_10400,N_10239,N_10203);
and U10401 (N_10401,N_10225,N_10206);
and U10402 (N_10402,N_10298,N_10227);
or U10403 (N_10403,N_10268,N_10332);
or U10404 (N_10404,N_10271,N_10204);
xor U10405 (N_10405,N_10312,N_10230);
and U10406 (N_10406,N_10259,N_10320);
and U10407 (N_10407,N_10234,N_10246);
or U10408 (N_10408,N_10251,N_10248);
nand U10409 (N_10409,N_10348,N_10219);
nand U10410 (N_10410,N_10275,N_10325);
xnor U10411 (N_10411,N_10330,N_10283);
or U10412 (N_10412,N_10207,N_10328);
and U10413 (N_10413,N_10337,N_10286);
nor U10414 (N_10414,N_10333,N_10299);
nor U10415 (N_10415,N_10261,N_10316);
or U10416 (N_10416,N_10262,N_10318);
nand U10417 (N_10417,N_10214,N_10256);
nor U10418 (N_10418,N_10202,N_10306);
nor U10419 (N_10419,N_10212,N_10288);
or U10420 (N_10420,N_10238,N_10302);
xnor U10421 (N_10421,N_10255,N_10218);
nand U10422 (N_10422,N_10209,N_10315);
nor U10423 (N_10423,N_10211,N_10273);
xnor U10424 (N_10424,N_10240,N_10263);
or U10425 (N_10425,N_10232,N_10315);
or U10426 (N_10426,N_10260,N_10208);
nor U10427 (N_10427,N_10284,N_10256);
nor U10428 (N_10428,N_10282,N_10345);
xor U10429 (N_10429,N_10219,N_10253);
nor U10430 (N_10430,N_10236,N_10207);
nand U10431 (N_10431,N_10275,N_10233);
and U10432 (N_10432,N_10253,N_10338);
nand U10433 (N_10433,N_10256,N_10236);
or U10434 (N_10434,N_10213,N_10207);
and U10435 (N_10435,N_10213,N_10247);
xnor U10436 (N_10436,N_10273,N_10336);
nor U10437 (N_10437,N_10298,N_10235);
nand U10438 (N_10438,N_10326,N_10271);
nand U10439 (N_10439,N_10341,N_10303);
nand U10440 (N_10440,N_10307,N_10208);
or U10441 (N_10441,N_10263,N_10227);
xor U10442 (N_10442,N_10325,N_10294);
xor U10443 (N_10443,N_10300,N_10323);
nand U10444 (N_10444,N_10246,N_10237);
nor U10445 (N_10445,N_10313,N_10307);
xor U10446 (N_10446,N_10329,N_10292);
xor U10447 (N_10447,N_10258,N_10318);
nor U10448 (N_10448,N_10324,N_10323);
and U10449 (N_10449,N_10244,N_10245);
xor U10450 (N_10450,N_10314,N_10222);
xnor U10451 (N_10451,N_10252,N_10232);
or U10452 (N_10452,N_10229,N_10270);
nand U10453 (N_10453,N_10306,N_10242);
nor U10454 (N_10454,N_10280,N_10212);
nor U10455 (N_10455,N_10290,N_10224);
xnor U10456 (N_10456,N_10289,N_10312);
or U10457 (N_10457,N_10297,N_10309);
and U10458 (N_10458,N_10232,N_10238);
or U10459 (N_10459,N_10303,N_10327);
and U10460 (N_10460,N_10222,N_10224);
or U10461 (N_10461,N_10287,N_10205);
nor U10462 (N_10462,N_10221,N_10335);
nand U10463 (N_10463,N_10203,N_10283);
nor U10464 (N_10464,N_10285,N_10221);
or U10465 (N_10465,N_10201,N_10286);
or U10466 (N_10466,N_10317,N_10207);
or U10467 (N_10467,N_10322,N_10319);
nand U10468 (N_10468,N_10253,N_10208);
or U10469 (N_10469,N_10276,N_10320);
xor U10470 (N_10470,N_10215,N_10302);
xor U10471 (N_10471,N_10205,N_10274);
nor U10472 (N_10472,N_10320,N_10341);
nor U10473 (N_10473,N_10248,N_10308);
xor U10474 (N_10474,N_10330,N_10326);
nor U10475 (N_10475,N_10266,N_10221);
and U10476 (N_10476,N_10214,N_10347);
and U10477 (N_10477,N_10241,N_10211);
or U10478 (N_10478,N_10236,N_10231);
xor U10479 (N_10479,N_10339,N_10238);
nor U10480 (N_10480,N_10348,N_10344);
or U10481 (N_10481,N_10211,N_10342);
or U10482 (N_10482,N_10216,N_10291);
xor U10483 (N_10483,N_10211,N_10331);
and U10484 (N_10484,N_10257,N_10346);
nand U10485 (N_10485,N_10321,N_10228);
nand U10486 (N_10486,N_10315,N_10234);
and U10487 (N_10487,N_10314,N_10235);
or U10488 (N_10488,N_10275,N_10221);
nand U10489 (N_10489,N_10270,N_10200);
nand U10490 (N_10490,N_10210,N_10331);
xnor U10491 (N_10491,N_10205,N_10279);
xnor U10492 (N_10492,N_10232,N_10300);
or U10493 (N_10493,N_10282,N_10293);
xor U10494 (N_10494,N_10277,N_10287);
xnor U10495 (N_10495,N_10215,N_10233);
xnor U10496 (N_10496,N_10291,N_10230);
and U10497 (N_10497,N_10203,N_10278);
nand U10498 (N_10498,N_10209,N_10220);
nand U10499 (N_10499,N_10212,N_10338);
nor U10500 (N_10500,N_10434,N_10411);
or U10501 (N_10501,N_10357,N_10391);
xnor U10502 (N_10502,N_10370,N_10351);
nor U10503 (N_10503,N_10367,N_10442);
and U10504 (N_10504,N_10495,N_10364);
or U10505 (N_10505,N_10404,N_10372);
nor U10506 (N_10506,N_10483,N_10441);
or U10507 (N_10507,N_10361,N_10466);
xor U10508 (N_10508,N_10406,N_10490);
and U10509 (N_10509,N_10385,N_10392);
xor U10510 (N_10510,N_10407,N_10443);
or U10511 (N_10511,N_10428,N_10379);
or U10512 (N_10512,N_10453,N_10422);
nand U10513 (N_10513,N_10394,N_10444);
and U10514 (N_10514,N_10420,N_10447);
nor U10515 (N_10515,N_10402,N_10429);
xor U10516 (N_10516,N_10462,N_10396);
and U10517 (N_10517,N_10376,N_10414);
nor U10518 (N_10518,N_10381,N_10378);
nand U10519 (N_10519,N_10365,N_10405);
nand U10520 (N_10520,N_10496,N_10455);
and U10521 (N_10521,N_10486,N_10494);
and U10522 (N_10522,N_10452,N_10468);
and U10523 (N_10523,N_10399,N_10358);
xor U10524 (N_10524,N_10437,N_10427);
xor U10525 (N_10525,N_10460,N_10475);
nand U10526 (N_10526,N_10492,N_10491);
nor U10527 (N_10527,N_10493,N_10499);
nor U10528 (N_10528,N_10386,N_10446);
nand U10529 (N_10529,N_10374,N_10380);
xor U10530 (N_10530,N_10470,N_10369);
xnor U10531 (N_10531,N_10418,N_10363);
and U10532 (N_10532,N_10362,N_10477);
nand U10533 (N_10533,N_10448,N_10485);
nor U10534 (N_10534,N_10498,N_10397);
and U10535 (N_10535,N_10383,N_10408);
nor U10536 (N_10536,N_10465,N_10375);
xnor U10537 (N_10537,N_10360,N_10433);
nand U10538 (N_10538,N_10478,N_10395);
xnor U10539 (N_10539,N_10413,N_10353);
nand U10540 (N_10540,N_10484,N_10419);
or U10541 (N_10541,N_10426,N_10449);
nor U10542 (N_10542,N_10359,N_10435);
or U10543 (N_10543,N_10461,N_10488);
nand U10544 (N_10544,N_10354,N_10480);
nand U10545 (N_10545,N_10430,N_10384);
xor U10546 (N_10546,N_10355,N_10436);
and U10547 (N_10547,N_10350,N_10412);
nor U10548 (N_10548,N_10464,N_10409);
and U10549 (N_10549,N_10403,N_10356);
or U10550 (N_10550,N_10388,N_10431);
and U10551 (N_10551,N_10421,N_10410);
xnor U10552 (N_10552,N_10458,N_10459);
or U10553 (N_10553,N_10469,N_10389);
xnor U10554 (N_10554,N_10425,N_10400);
or U10555 (N_10555,N_10451,N_10423);
or U10556 (N_10556,N_10371,N_10497);
or U10557 (N_10557,N_10454,N_10471);
xnor U10558 (N_10558,N_10424,N_10401);
or U10559 (N_10559,N_10398,N_10457);
xor U10560 (N_10560,N_10368,N_10467);
nand U10561 (N_10561,N_10445,N_10373);
nand U10562 (N_10562,N_10476,N_10472);
nand U10563 (N_10563,N_10417,N_10482);
or U10564 (N_10564,N_10387,N_10481);
nand U10565 (N_10565,N_10438,N_10352);
and U10566 (N_10566,N_10479,N_10473);
nand U10567 (N_10567,N_10474,N_10440);
xor U10568 (N_10568,N_10366,N_10489);
nand U10569 (N_10569,N_10416,N_10377);
xnor U10570 (N_10570,N_10450,N_10415);
nor U10571 (N_10571,N_10456,N_10487);
nor U10572 (N_10572,N_10382,N_10463);
nand U10573 (N_10573,N_10390,N_10439);
or U10574 (N_10574,N_10432,N_10393);
xnor U10575 (N_10575,N_10451,N_10442);
and U10576 (N_10576,N_10449,N_10495);
nand U10577 (N_10577,N_10461,N_10383);
or U10578 (N_10578,N_10422,N_10430);
and U10579 (N_10579,N_10473,N_10447);
nand U10580 (N_10580,N_10381,N_10481);
nand U10581 (N_10581,N_10494,N_10453);
and U10582 (N_10582,N_10431,N_10443);
nand U10583 (N_10583,N_10371,N_10438);
nand U10584 (N_10584,N_10388,N_10499);
nand U10585 (N_10585,N_10401,N_10406);
xnor U10586 (N_10586,N_10372,N_10495);
xnor U10587 (N_10587,N_10441,N_10479);
and U10588 (N_10588,N_10449,N_10380);
xor U10589 (N_10589,N_10459,N_10426);
nor U10590 (N_10590,N_10395,N_10367);
and U10591 (N_10591,N_10498,N_10474);
nand U10592 (N_10592,N_10475,N_10479);
or U10593 (N_10593,N_10476,N_10369);
and U10594 (N_10594,N_10386,N_10471);
and U10595 (N_10595,N_10460,N_10413);
and U10596 (N_10596,N_10487,N_10438);
or U10597 (N_10597,N_10487,N_10451);
nor U10598 (N_10598,N_10415,N_10400);
or U10599 (N_10599,N_10369,N_10359);
and U10600 (N_10600,N_10427,N_10438);
nor U10601 (N_10601,N_10399,N_10447);
nor U10602 (N_10602,N_10414,N_10366);
and U10603 (N_10603,N_10393,N_10437);
and U10604 (N_10604,N_10405,N_10480);
and U10605 (N_10605,N_10449,N_10466);
and U10606 (N_10606,N_10461,N_10429);
xor U10607 (N_10607,N_10393,N_10412);
nor U10608 (N_10608,N_10382,N_10478);
nor U10609 (N_10609,N_10395,N_10470);
and U10610 (N_10610,N_10485,N_10396);
xor U10611 (N_10611,N_10463,N_10398);
or U10612 (N_10612,N_10498,N_10378);
and U10613 (N_10613,N_10475,N_10411);
nor U10614 (N_10614,N_10410,N_10428);
xnor U10615 (N_10615,N_10461,N_10368);
nor U10616 (N_10616,N_10472,N_10381);
nand U10617 (N_10617,N_10498,N_10492);
nor U10618 (N_10618,N_10400,N_10402);
nand U10619 (N_10619,N_10451,N_10383);
nand U10620 (N_10620,N_10382,N_10491);
or U10621 (N_10621,N_10477,N_10404);
xor U10622 (N_10622,N_10426,N_10443);
or U10623 (N_10623,N_10394,N_10417);
xnor U10624 (N_10624,N_10390,N_10362);
xor U10625 (N_10625,N_10380,N_10376);
and U10626 (N_10626,N_10424,N_10436);
nand U10627 (N_10627,N_10381,N_10395);
nor U10628 (N_10628,N_10482,N_10416);
nor U10629 (N_10629,N_10351,N_10481);
nand U10630 (N_10630,N_10476,N_10480);
nor U10631 (N_10631,N_10427,N_10478);
and U10632 (N_10632,N_10392,N_10452);
or U10633 (N_10633,N_10370,N_10429);
or U10634 (N_10634,N_10382,N_10425);
nor U10635 (N_10635,N_10423,N_10368);
xor U10636 (N_10636,N_10396,N_10359);
or U10637 (N_10637,N_10477,N_10448);
nand U10638 (N_10638,N_10494,N_10436);
and U10639 (N_10639,N_10359,N_10410);
or U10640 (N_10640,N_10410,N_10449);
nand U10641 (N_10641,N_10386,N_10428);
nand U10642 (N_10642,N_10395,N_10375);
or U10643 (N_10643,N_10410,N_10375);
and U10644 (N_10644,N_10452,N_10354);
or U10645 (N_10645,N_10457,N_10456);
xor U10646 (N_10646,N_10469,N_10442);
nand U10647 (N_10647,N_10390,N_10357);
xnor U10648 (N_10648,N_10499,N_10432);
and U10649 (N_10649,N_10350,N_10390);
nor U10650 (N_10650,N_10543,N_10626);
and U10651 (N_10651,N_10557,N_10501);
nand U10652 (N_10652,N_10578,N_10587);
xnor U10653 (N_10653,N_10569,N_10536);
xor U10654 (N_10654,N_10566,N_10644);
nor U10655 (N_10655,N_10526,N_10599);
xnor U10656 (N_10656,N_10508,N_10581);
and U10657 (N_10657,N_10603,N_10545);
xor U10658 (N_10658,N_10503,N_10518);
nor U10659 (N_10659,N_10629,N_10597);
xor U10660 (N_10660,N_10605,N_10541);
or U10661 (N_10661,N_10622,N_10500);
nor U10662 (N_10662,N_10571,N_10562);
xnor U10663 (N_10663,N_10627,N_10521);
nor U10664 (N_10664,N_10604,N_10631);
xor U10665 (N_10665,N_10642,N_10628);
nand U10666 (N_10666,N_10645,N_10636);
nor U10667 (N_10667,N_10609,N_10606);
nand U10668 (N_10668,N_10511,N_10515);
and U10669 (N_10669,N_10593,N_10574);
nor U10670 (N_10670,N_10547,N_10550);
nor U10671 (N_10671,N_10583,N_10590);
and U10672 (N_10672,N_10618,N_10594);
nor U10673 (N_10673,N_10509,N_10592);
xor U10674 (N_10674,N_10567,N_10540);
or U10675 (N_10675,N_10615,N_10546);
nand U10676 (N_10676,N_10610,N_10510);
xor U10677 (N_10677,N_10556,N_10551);
or U10678 (N_10678,N_10529,N_10607);
nor U10679 (N_10679,N_10595,N_10548);
and U10680 (N_10680,N_10635,N_10520);
or U10681 (N_10681,N_10639,N_10588);
nor U10682 (N_10682,N_10553,N_10563);
nand U10683 (N_10683,N_10602,N_10523);
and U10684 (N_10684,N_10619,N_10608);
and U10685 (N_10685,N_10585,N_10542);
and U10686 (N_10686,N_10559,N_10561);
or U10687 (N_10687,N_10648,N_10589);
nor U10688 (N_10688,N_10646,N_10565);
nor U10689 (N_10689,N_10572,N_10616);
and U10690 (N_10690,N_10506,N_10524);
or U10691 (N_10691,N_10533,N_10534);
or U10692 (N_10692,N_10568,N_10621);
or U10693 (N_10693,N_10573,N_10560);
nand U10694 (N_10694,N_10591,N_10532);
or U10695 (N_10695,N_10527,N_10596);
or U10696 (N_10696,N_10582,N_10620);
or U10697 (N_10697,N_10598,N_10537);
or U10698 (N_10698,N_10552,N_10502);
or U10699 (N_10699,N_10632,N_10580);
xnor U10700 (N_10700,N_10641,N_10577);
or U10701 (N_10701,N_10517,N_10625);
and U10702 (N_10702,N_10575,N_10623);
or U10703 (N_10703,N_10640,N_10584);
and U10704 (N_10704,N_10507,N_10538);
xnor U10705 (N_10705,N_10612,N_10586);
or U10706 (N_10706,N_10516,N_10643);
or U10707 (N_10707,N_10549,N_10617);
and U10708 (N_10708,N_10570,N_10579);
nand U10709 (N_10709,N_10513,N_10558);
and U10710 (N_10710,N_10522,N_10504);
nand U10711 (N_10711,N_10638,N_10512);
and U10712 (N_10712,N_10633,N_10634);
xor U10713 (N_10713,N_10564,N_10601);
xor U10714 (N_10714,N_10576,N_10519);
xor U10715 (N_10715,N_10611,N_10637);
nand U10716 (N_10716,N_10613,N_10535);
and U10717 (N_10717,N_10647,N_10614);
and U10718 (N_10718,N_10528,N_10544);
nand U10719 (N_10719,N_10530,N_10539);
and U10720 (N_10720,N_10514,N_10600);
and U10721 (N_10721,N_10649,N_10554);
nor U10722 (N_10722,N_10505,N_10525);
nor U10723 (N_10723,N_10624,N_10531);
nor U10724 (N_10724,N_10555,N_10630);
or U10725 (N_10725,N_10581,N_10524);
or U10726 (N_10726,N_10601,N_10575);
or U10727 (N_10727,N_10548,N_10510);
xnor U10728 (N_10728,N_10555,N_10515);
xnor U10729 (N_10729,N_10537,N_10516);
or U10730 (N_10730,N_10538,N_10518);
xnor U10731 (N_10731,N_10578,N_10508);
nor U10732 (N_10732,N_10619,N_10529);
nor U10733 (N_10733,N_10607,N_10587);
and U10734 (N_10734,N_10543,N_10579);
xnor U10735 (N_10735,N_10631,N_10576);
or U10736 (N_10736,N_10592,N_10597);
nand U10737 (N_10737,N_10598,N_10579);
xnor U10738 (N_10738,N_10598,N_10517);
nor U10739 (N_10739,N_10562,N_10574);
or U10740 (N_10740,N_10595,N_10597);
and U10741 (N_10741,N_10525,N_10603);
or U10742 (N_10742,N_10529,N_10617);
xnor U10743 (N_10743,N_10584,N_10532);
nand U10744 (N_10744,N_10595,N_10645);
nand U10745 (N_10745,N_10606,N_10647);
or U10746 (N_10746,N_10550,N_10533);
xnor U10747 (N_10747,N_10644,N_10510);
nor U10748 (N_10748,N_10544,N_10543);
or U10749 (N_10749,N_10585,N_10560);
nand U10750 (N_10750,N_10518,N_10519);
xnor U10751 (N_10751,N_10563,N_10649);
nor U10752 (N_10752,N_10637,N_10593);
and U10753 (N_10753,N_10638,N_10557);
xnor U10754 (N_10754,N_10641,N_10516);
nor U10755 (N_10755,N_10568,N_10549);
or U10756 (N_10756,N_10601,N_10621);
or U10757 (N_10757,N_10545,N_10591);
xnor U10758 (N_10758,N_10554,N_10575);
or U10759 (N_10759,N_10528,N_10614);
or U10760 (N_10760,N_10606,N_10636);
nor U10761 (N_10761,N_10563,N_10634);
nor U10762 (N_10762,N_10515,N_10647);
nor U10763 (N_10763,N_10567,N_10518);
nand U10764 (N_10764,N_10593,N_10618);
nor U10765 (N_10765,N_10520,N_10529);
xor U10766 (N_10766,N_10548,N_10536);
or U10767 (N_10767,N_10599,N_10613);
nor U10768 (N_10768,N_10613,N_10646);
xnor U10769 (N_10769,N_10599,N_10631);
nor U10770 (N_10770,N_10524,N_10585);
nand U10771 (N_10771,N_10604,N_10505);
and U10772 (N_10772,N_10513,N_10593);
or U10773 (N_10773,N_10636,N_10598);
xnor U10774 (N_10774,N_10644,N_10538);
xnor U10775 (N_10775,N_10640,N_10592);
or U10776 (N_10776,N_10600,N_10527);
or U10777 (N_10777,N_10510,N_10503);
nand U10778 (N_10778,N_10633,N_10523);
xor U10779 (N_10779,N_10507,N_10620);
and U10780 (N_10780,N_10555,N_10536);
xor U10781 (N_10781,N_10520,N_10532);
or U10782 (N_10782,N_10614,N_10538);
xnor U10783 (N_10783,N_10539,N_10630);
xnor U10784 (N_10784,N_10554,N_10548);
xor U10785 (N_10785,N_10514,N_10648);
nand U10786 (N_10786,N_10587,N_10509);
nor U10787 (N_10787,N_10535,N_10511);
xor U10788 (N_10788,N_10620,N_10602);
nor U10789 (N_10789,N_10635,N_10536);
nor U10790 (N_10790,N_10537,N_10501);
xor U10791 (N_10791,N_10525,N_10608);
nor U10792 (N_10792,N_10569,N_10637);
nand U10793 (N_10793,N_10585,N_10625);
nor U10794 (N_10794,N_10533,N_10622);
nand U10795 (N_10795,N_10502,N_10539);
and U10796 (N_10796,N_10598,N_10608);
or U10797 (N_10797,N_10504,N_10538);
and U10798 (N_10798,N_10595,N_10636);
xor U10799 (N_10799,N_10600,N_10608);
and U10800 (N_10800,N_10683,N_10691);
nor U10801 (N_10801,N_10796,N_10787);
nor U10802 (N_10802,N_10740,N_10710);
xnor U10803 (N_10803,N_10789,N_10668);
and U10804 (N_10804,N_10723,N_10775);
nand U10805 (N_10805,N_10737,N_10674);
xor U10806 (N_10806,N_10713,N_10794);
or U10807 (N_10807,N_10770,N_10661);
and U10808 (N_10808,N_10690,N_10689);
nor U10809 (N_10809,N_10782,N_10667);
or U10810 (N_10810,N_10653,N_10658);
and U10811 (N_10811,N_10654,N_10672);
and U10812 (N_10812,N_10792,N_10772);
and U10813 (N_10813,N_10693,N_10697);
nand U10814 (N_10814,N_10733,N_10657);
xor U10815 (N_10815,N_10703,N_10748);
nand U10816 (N_10816,N_10705,N_10721);
and U10817 (N_10817,N_10764,N_10708);
xor U10818 (N_10818,N_10719,N_10694);
and U10819 (N_10819,N_10735,N_10725);
or U10820 (N_10820,N_10715,N_10744);
nor U10821 (N_10821,N_10687,N_10790);
or U10822 (N_10822,N_10798,N_10729);
nand U10823 (N_10823,N_10738,N_10701);
xor U10824 (N_10824,N_10743,N_10747);
and U10825 (N_10825,N_10681,N_10712);
nor U10826 (N_10826,N_10783,N_10679);
nor U10827 (N_10827,N_10659,N_10763);
nand U10828 (N_10828,N_10753,N_10651);
nand U10829 (N_10829,N_10793,N_10779);
xnor U10830 (N_10830,N_10695,N_10720);
or U10831 (N_10831,N_10739,N_10760);
or U10832 (N_10832,N_10696,N_10762);
nor U10833 (N_10833,N_10791,N_10652);
or U10834 (N_10834,N_10774,N_10754);
nor U10835 (N_10835,N_10670,N_10682);
xor U10836 (N_10836,N_10734,N_10785);
xor U10837 (N_10837,N_10685,N_10752);
nor U10838 (N_10838,N_10711,N_10765);
or U10839 (N_10839,N_10788,N_10664);
nand U10840 (N_10840,N_10655,N_10660);
nand U10841 (N_10841,N_10736,N_10780);
and U10842 (N_10842,N_10769,N_10688);
nand U10843 (N_10843,N_10666,N_10706);
and U10844 (N_10844,N_10799,N_10797);
nor U10845 (N_10845,N_10678,N_10692);
nand U10846 (N_10846,N_10795,N_10781);
xor U10847 (N_10847,N_10686,N_10704);
nor U10848 (N_10848,N_10741,N_10718);
xnor U10849 (N_10849,N_10650,N_10786);
xnor U10850 (N_10850,N_10745,N_10699);
and U10851 (N_10851,N_10671,N_10767);
or U10852 (N_10852,N_10777,N_10758);
and U10853 (N_10853,N_10698,N_10714);
or U10854 (N_10854,N_10669,N_10709);
xor U10855 (N_10855,N_10724,N_10676);
xnor U10856 (N_10856,N_10766,N_10761);
nor U10857 (N_10857,N_10759,N_10751);
nor U10858 (N_10858,N_10742,N_10684);
or U10859 (N_10859,N_10750,N_10707);
xnor U10860 (N_10860,N_10663,N_10756);
or U10861 (N_10861,N_10746,N_10656);
and U10862 (N_10862,N_10768,N_10757);
and U10863 (N_10863,N_10700,N_10731);
or U10864 (N_10864,N_10784,N_10730);
nand U10865 (N_10865,N_10680,N_10773);
xnor U10866 (N_10866,N_10702,N_10675);
nand U10867 (N_10867,N_10732,N_10673);
or U10868 (N_10868,N_10722,N_10778);
xor U10869 (N_10869,N_10728,N_10776);
xor U10870 (N_10870,N_10755,N_10749);
and U10871 (N_10871,N_10727,N_10717);
nand U10872 (N_10872,N_10716,N_10726);
nor U10873 (N_10873,N_10677,N_10771);
xnor U10874 (N_10874,N_10665,N_10662);
and U10875 (N_10875,N_10662,N_10687);
nor U10876 (N_10876,N_10694,N_10678);
xor U10877 (N_10877,N_10736,N_10700);
nand U10878 (N_10878,N_10734,N_10685);
nand U10879 (N_10879,N_10762,N_10761);
and U10880 (N_10880,N_10710,N_10798);
nand U10881 (N_10881,N_10751,N_10744);
or U10882 (N_10882,N_10765,N_10668);
nand U10883 (N_10883,N_10666,N_10716);
nand U10884 (N_10884,N_10724,N_10736);
or U10885 (N_10885,N_10737,N_10757);
and U10886 (N_10886,N_10730,N_10725);
nand U10887 (N_10887,N_10752,N_10794);
or U10888 (N_10888,N_10751,N_10673);
and U10889 (N_10889,N_10745,N_10797);
or U10890 (N_10890,N_10769,N_10719);
nor U10891 (N_10891,N_10716,N_10675);
nand U10892 (N_10892,N_10783,N_10711);
xnor U10893 (N_10893,N_10798,N_10683);
or U10894 (N_10894,N_10785,N_10687);
xor U10895 (N_10895,N_10745,N_10662);
or U10896 (N_10896,N_10725,N_10793);
xor U10897 (N_10897,N_10655,N_10712);
nor U10898 (N_10898,N_10701,N_10693);
and U10899 (N_10899,N_10676,N_10746);
xnor U10900 (N_10900,N_10709,N_10668);
or U10901 (N_10901,N_10664,N_10743);
xnor U10902 (N_10902,N_10745,N_10760);
xor U10903 (N_10903,N_10711,N_10696);
xor U10904 (N_10904,N_10666,N_10684);
and U10905 (N_10905,N_10791,N_10682);
xor U10906 (N_10906,N_10774,N_10791);
and U10907 (N_10907,N_10757,N_10730);
or U10908 (N_10908,N_10754,N_10676);
or U10909 (N_10909,N_10668,N_10744);
nor U10910 (N_10910,N_10736,N_10727);
or U10911 (N_10911,N_10694,N_10765);
nor U10912 (N_10912,N_10764,N_10722);
and U10913 (N_10913,N_10671,N_10676);
and U10914 (N_10914,N_10768,N_10774);
and U10915 (N_10915,N_10720,N_10662);
nand U10916 (N_10916,N_10684,N_10689);
nor U10917 (N_10917,N_10714,N_10770);
xor U10918 (N_10918,N_10731,N_10764);
nor U10919 (N_10919,N_10722,N_10744);
nand U10920 (N_10920,N_10701,N_10687);
and U10921 (N_10921,N_10759,N_10793);
nor U10922 (N_10922,N_10762,N_10766);
or U10923 (N_10923,N_10659,N_10751);
xor U10924 (N_10924,N_10700,N_10763);
nand U10925 (N_10925,N_10675,N_10705);
xnor U10926 (N_10926,N_10664,N_10751);
nor U10927 (N_10927,N_10691,N_10675);
or U10928 (N_10928,N_10793,N_10711);
or U10929 (N_10929,N_10784,N_10650);
nor U10930 (N_10930,N_10653,N_10734);
xor U10931 (N_10931,N_10669,N_10786);
xor U10932 (N_10932,N_10700,N_10683);
or U10933 (N_10933,N_10770,N_10679);
nor U10934 (N_10934,N_10757,N_10657);
or U10935 (N_10935,N_10669,N_10792);
and U10936 (N_10936,N_10696,N_10664);
and U10937 (N_10937,N_10693,N_10758);
nand U10938 (N_10938,N_10696,N_10757);
and U10939 (N_10939,N_10794,N_10694);
nor U10940 (N_10940,N_10745,N_10650);
or U10941 (N_10941,N_10710,N_10651);
or U10942 (N_10942,N_10669,N_10711);
nor U10943 (N_10943,N_10657,N_10673);
nand U10944 (N_10944,N_10768,N_10704);
nand U10945 (N_10945,N_10677,N_10687);
and U10946 (N_10946,N_10777,N_10722);
xor U10947 (N_10947,N_10705,N_10698);
nand U10948 (N_10948,N_10709,N_10718);
xor U10949 (N_10949,N_10708,N_10770);
or U10950 (N_10950,N_10922,N_10825);
and U10951 (N_10951,N_10898,N_10810);
or U10952 (N_10952,N_10946,N_10821);
and U10953 (N_10953,N_10832,N_10826);
and U10954 (N_10954,N_10873,N_10903);
and U10955 (N_10955,N_10929,N_10851);
and U10956 (N_10956,N_10853,N_10888);
and U10957 (N_10957,N_10828,N_10862);
xor U10958 (N_10958,N_10904,N_10908);
and U10959 (N_10959,N_10887,N_10830);
or U10960 (N_10960,N_10837,N_10924);
nor U10961 (N_10961,N_10893,N_10845);
and U10962 (N_10962,N_10822,N_10865);
nand U10963 (N_10963,N_10859,N_10852);
and U10964 (N_10964,N_10829,N_10905);
nor U10965 (N_10965,N_10838,N_10880);
xnor U10966 (N_10966,N_10886,N_10919);
nand U10967 (N_10967,N_10833,N_10803);
nand U10968 (N_10968,N_10942,N_10879);
nor U10969 (N_10969,N_10876,N_10813);
or U10970 (N_10970,N_10885,N_10835);
or U10971 (N_10971,N_10928,N_10940);
nor U10972 (N_10972,N_10863,N_10844);
xor U10973 (N_10973,N_10890,N_10819);
and U10974 (N_10974,N_10882,N_10814);
or U10975 (N_10975,N_10900,N_10897);
or U10976 (N_10976,N_10846,N_10930);
xnor U10977 (N_10977,N_10912,N_10932);
nand U10978 (N_10978,N_10843,N_10923);
nor U10979 (N_10979,N_10917,N_10947);
or U10980 (N_10980,N_10914,N_10834);
xnor U10981 (N_10981,N_10937,N_10872);
xor U10982 (N_10982,N_10861,N_10938);
nand U10983 (N_10983,N_10883,N_10849);
or U10984 (N_10984,N_10933,N_10817);
xnor U10985 (N_10985,N_10856,N_10892);
nor U10986 (N_10986,N_10836,N_10875);
nand U10987 (N_10987,N_10841,N_10948);
nor U10988 (N_10988,N_10827,N_10910);
nor U10989 (N_10989,N_10807,N_10801);
or U10990 (N_10990,N_10944,N_10823);
or U10991 (N_10991,N_10870,N_10868);
nor U10992 (N_10992,N_10889,N_10869);
nand U10993 (N_10993,N_10864,N_10939);
nor U10994 (N_10994,N_10895,N_10927);
or U10995 (N_10995,N_10935,N_10871);
nor U10996 (N_10996,N_10804,N_10949);
or U10997 (N_10997,N_10907,N_10911);
nand U10998 (N_10998,N_10891,N_10877);
and U10999 (N_10999,N_10824,N_10943);
nand U11000 (N_11000,N_10816,N_10857);
xor U11001 (N_11001,N_10925,N_10866);
and U11002 (N_11002,N_10936,N_10874);
and U11003 (N_11003,N_10818,N_10858);
xnor U11004 (N_11004,N_10831,N_10820);
nor U11005 (N_11005,N_10800,N_10941);
xnor U11006 (N_11006,N_10894,N_10899);
or U11007 (N_11007,N_10916,N_10918);
nand U11008 (N_11008,N_10896,N_10812);
nor U11009 (N_11009,N_10860,N_10926);
and U11010 (N_11010,N_10920,N_10901);
and U11011 (N_11011,N_10921,N_10884);
xnor U11012 (N_11012,N_10867,N_10839);
nor U11013 (N_11013,N_10915,N_10811);
nor U11014 (N_11014,N_10805,N_10881);
or U11015 (N_11015,N_10931,N_10878);
xnor U11016 (N_11016,N_10815,N_10802);
xor U11017 (N_11017,N_10847,N_10854);
nor U11018 (N_11018,N_10850,N_10909);
or U11019 (N_11019,N_10855,N_10906);
or U11020 (N_11020,N_10945,N_10842);
nand U11021 (N_11021,N_10809,N_10808);
and U11022 (N_11022,N_10806,N_10840);
nor U11023 (N_11023,N_10913,N_10902);
xnor U11024 (N_11024,N_10848,N_10934);
and U11025 (N_11025,N_10900,N_10903);
nand U11026 (N_11026,N_10905,N_10949);
nand U11027 (N_11027,N_10844,N_10842);
and U11028 (N_11028,N_10938,N_10875);
or U11029 (N_11029,N_10935,N_10818);
nand U11030 (N_11030,N_10864,N_10940);
nand U11031 (N_11031,N_10804,N_10839);
and U11032 (N_11032,N_10916,N_10861);
or U11033 (N_11033,N_10899,N_10922);
and U11034 (N_11034,N_10845,N_10851);
nor U11035 (N_11035,N_10920,N_10882);
and U11036 (N_11036,N_10924,N_10858);
or U11037 (N_11037,N_10810,N_10823);
xor U11038 (N_11038,N_10920,N_10815);
or U11039 (N_11039,N_10874,N_10811);
nor U11040 (N_11040,N_10920,N_10881);
and U11041 (N_11041,N_10889,N_10924);
nor U11042 (N_11042,N_10859,N_10842);
or U11043 (N_11043,N_10839,N_10926);
nor U11044 (N_11044,N_10830,N_10815);
nor U11045 (N_11045,N_10919,N_10860);
or U11046 (N_11046,N_10926,N_10897);
nor U11047 (N_11047,N_10867,N_10819);
nor U11048 (N_11048,N_10808,N_10901);
nor U11049 (N_11049,N_10852,N_10921);
xnor U11050 (N_11050,N_10800,N_10808);
nand U11051 (N_11051,N_10812,N_10876);
nor U11052 (N_11052,N_10841,N_10837);
or U11053 (N_11053,N_10803,N_10894);
and U11054 (N_11054,N_10930,N_10840);
and U11055 (N_11055,N_10900,N_10814);
or U11056 (N_11056,N_10846,N_10929);
nand U11057 (N_11057,N_10874,N_10911);
nor U11058 (N_11058,N_10814,N_10877);
nor U11059 (N_11059,N_10832,N_10901);
and U11060 (N_11060,N_10809,N_10933);
nor U11061 (N_11061,N_10899,N_10839);
and U11062 (N_11062,N_10834,N_10929);
or U11063 (N_11063,N_10826,N_10882);
and U11064 (N_11064,N_10864,N_10823);
xor U11065 (N_11065,N_10847,N_10848);
or U11066 (N_11066,N_10840,N_10849);
nand U11067 (N_11067,N_10870,N_10889);
nand U11068 (N_11068,N_10832,N_10854);
xor U11069 (N_11069,N_10883,N_10822);
nand U11070 (N_11070,N_10928,N_10896);
nand U11071 (N_11071,N_10801,N_10818);
xor U11072 (N_11072,N_10885,N_10870);
nand U11073 (N_11073,N_10835,N_10852);
or U11074 (N_11074,N_10816,N_10921);
and U11075 (N_11075,N_10880,N_10937);
xor U11076 (N_11076,N_10859,N_10836);
nor U11077 (N_11077,N_10860,N_10884);
nand U11078 (N_11078,N_10910,N_10896);
nor U11079 (N_11079,N_10942,N_10830);
and U11080 (N_11080,N_10820,N_10826);
or U11081 (N_11081,N_10810,N_10880);
or U11082 (N_11082,N_10895,N_10812);
xnor U11083 (N_11083,N_10896,N_10933);
nor U11084 (N_11084,N_10832,N_10899);
xnor U11085 (N_11085,N_10878,N_10874);
nor U11086 (N_11086,N_10848,N_10918);
and U11087 (N_11087,N_10871,N_10812);
nand U11088 (N_11088,N_10897,N_10929);
xnor U11089 (N_11089,N_10901,N_10829);
nor U11090 (N_11090,N_10810,N_10903);
or U11091 (N_11091,N_10902,N_10877);
xnor U11092 (N_11092,N_10842,N_10922);
and U11093 (N_11093,N_10938,N_10914);
xor U11094 (N_11094,N_10940,N_10887);
and U11095 (N_11095,N_10822,N_10913);
or U11096 (N_11096,N_10859,N_10862);
xnor U11097 (N_11097,N_10813,N_10910);
or U11098 (N_11098,N_10925,N_10813);
or U11099 (N_11099,N_10811,N_10899);
nor U11100 (N_11100,N_11033,N_11031);
nor U11101 (N_11101,N_11010,N_10993);
nand U11102 (N_11102,N_11027,N_10971);
xnor U11103 (N_11103,N_11063,N_11057);
xor U11104 (N_11104,N_10990,N_11069);
or U11105 (N_11105,N_10962,N_11060);
nor U11106 (N_11106,N_11076,N_11025);
or U11107 (N_11107,N_11012,N_10955);
and U11108 (N_11108,N_11032,N_10998);
nand U11109 (N_11109,N_10950,N_11045);
nand U11110 (N_11110,N_11077,N_11068);
and U11111 (N_11111,N_10997,N_10952);
and U11112 (N_11112,N_10961,N_10974);
xnor U11113 (N_11113,N_11070,N_10968);
nand U11114 (N_11114,N_11090,N_11002);
or U11115 (N_11115,N_10988,N_11038);
nor U11116 (N_11116,N_11061,N_11049);
nor U11117 (N_11117,N_10957,N_11001);
nor U11118 (N_11118,N_11091,N_11054);
xor U11119 (N_11119,N_11016,N_11080);
and U11120 (N_11120,N_11005,N_10969);
xnor U11121 (N_11121,N_11062,N_11098);
or U11122 (N_11122,N_11042,N_11047);
xor U11123 (N_11123,N_11084,N_10973);
and U11124 (N_11124,N_11055,N_10975);
nor U11125 (N_11125,N_11082,N_10991);
xnor U11126 (N_11126,N_10982,N_11022);
nor U11127 (N_11127,N_11011,N_10983);
nand U11128 (N_11128,N_11079,N_10995);
nand U11129 (N_11129,N_11009,N_11088);
nor U11130 (N_11130,N_11092,N_11089);
nand U11131 (N_11131,N_11058,N_11099);
or U11132 (N_11132,N_11097,N_11020);
xor U11133 (N_11133,N_11066,N_11052);
or U11134 (N_11134,N_11008,N_11059);
xor U11135 (N_11135,N_11028,N_11093);
xnor U11136 (N_11136,N_10989,N_11095);
nor U11137 (N_11137,N_10960,N_10977);
xor U11138 (N_11138,N_11051,N_10976);
and U11139 (N_11139,N_11043,N_11035);
nor U11140 (N_11140,N_10999,N_10984);
nand U11141 (N_11141,N_11056,N_11096);
nand U11142 (N_11142,N_11044,N_10951);
and U11143 (N_11143,N_11067,N_11021);
or U11144 (N_11144,N_11083,N_11078);
nor U11145 (N_11145,N_11071,N_10972);
nand U11146 (N_11146,N_10994,N_11050);
nor U11147 (N_11147,N_11017,N_11023);
and U11148 (N_11148,N_11026,N_11073);
nand U11149 (N_11149,N_10986,N_11074);
xnor U11150 (N_11150,N_10992,N_11030);
nor U11151 (N_11151,N_11034,N_10965);
xor U11152 (N_11152,N_11003,N_11029);
nor U11153 (N_11153,N_10978,N_10996);
nand U11154 (N_11154,N_10956,N_10963);
and U11155 (N_11155,N_11046,N_11007);
or U11156 (N_11156,N_10959,N_11065);
nand U11157 (N_11157,N_11041,N_11019);
xnor U11158 (N_11158,N_10979,N_10980);
nor U11159 (N_11159,N_11004,N_11036);
or U11160 (N_11160,N_11064,N_10953);
or U11161 (N_11161,N_10970,N_10967);
xnor U11162 (N_11162,N_11094,N_10981);
or U11163 (N_11163,N_11024,N_10958);
or U11164 (N_11164,N_11039,N_11006);
nand U11165 (N_11165,N_10964,N_11000);
nand U11166 (N_11166,N_11053,N_11040);
or U11167 (N_11167,N_10985,N_10954);
xor U11168 (N_11168,N_11075,N_10966);
nor U11169 (N_11169,N_11087,N_11072);
or U11170 (N_11170,N_11015,N_11081);
nor U11171 (N_11171,N_11086,N_11048);
or U11172 (N_11172,N_11014,N_11013);
nand U11173 (N_11173,N_11018,N_10987);
xor U11174 (N_11174,N_11037,N_11085);
and U11175 (N_11175,N_11025,N_11044);
or U11176 (N_11176,N_11062,N_11068);
nand U11177 (N_11177,N_10982,N_11036);
xnor U11178 (N_11178,N_11065,N_11012);
or U11179 (N_11179,N_10975,N_11070);
nor U11180 (N_11180,N_10958,N_10964);
nand U11181 (N_11181,N_11086,N_11062);
xnor U11182 (N_11182,N_11046,N_11069);
and U11183 (N_11183,N_10989,N_11091);
nand U11184 (N_11184,N_11073,N_11053);
nor U11185 (N_11185,N_11029,N_10970);
nor U11186 (N_11186,N_11053,N_10968);
xnor U11187 (N_11187,N_11021,N_11055);
nand U11188 (N_11188,N_10960,N_10962);
nor U11189 (N_11189,N_11015,N_11096);
and U11190 (N_11190,N_11016,N_11059);
xor U11191 (N_11191,N_11012,N_11079);
nand U11192 (N_11192,N_11011,N_11029);
nand U11193 (N_11193,N_10985,N_11026);
nor U11194 (N_11194,N_11065,N_11096);
nand U11195 (N_11195,N_11018,N_10992);
nand U11196 (N_11196,N_11061,N_10955);
and U11197 (N_11197,N_11038,N_10985);
and U11198 (N_11198,N_11097,N_11034);
or U11199 (N_11199,N_11034,N_10958);
nor U11200 (N_11200,N_10991,N_10980);
xor U11201 (N_11201,N_11041,N_11065);
nor U11202 (N_11202,N_10979,N_11055);
and U11203 (N_11203,N_11076,N_11066);
xnor U11204 (N_11204,N_10976,N_11035);
nand U11205 (N_11205,N_10957,N_11073);
or U11206 (N_11206,N_10990,N_11089);
nand U11207 (N_11207,N_10973,N_10952);
or U11208 (N_11208,N_10969,N_11020);
nand U11209 (N_11209,N_11026,N_11039);
or U11210 (N_11210,N_10995,N_11038);
and U11211 (N_11211,N_11095,N_10959);
xor U11212 (N_11212,N_11007,N_11011);
nor U11213 (N_11213,N_10985,N_10969);
xor U11214 (N_11214,N_10962,N_11000);
nand U11215 (N_11215,N_11089,N_11012);
or U11216 (N_11216,N_10977,N_11040);
xor U11217 (N_11217,N_10956,N_11042);
and U11218 (N_11218,N_10992,N_10956);
nand U11219 (N_11219,N_11075,N_10985);
and U11220 (N_11220,N_10964,N_11066);
xor U11221 (N_11221,N_10973,N_11030);
xnor U11222 (N_11222,N_11049,N_10997);
xnor U11223 (N_11223,N_11066,N_11069);
nand U11224 (N_11224,N_11037,N_11090);
nand U11225 (N_11225,N_11035,N_10977);
nor U11226 (N_11226,N_11084,N_10966);
nor U11227 (N_11227,N_11030,N_11048);
nand U11228 (N_11228,N_11011,N_10981);
xnor U11229 (N_11229,N_11020,N_11071);
nor U11230 (N_11230,N_10974,N_10959);
or U11231 (N_11231,N_11025,N_11043);
xnor U11232 (N_11232,N_10985,N_11093);
and U11233 (N_11233,N_11053,N_10973);
or U11234 (N_11234,N_10958,N_11026);
xnor U11235 (N_11235,N_11067,N_11079);
nor U11236 (N_11236,N_11065,N_10977);
or U11237 (N_11237,N_11044,N_11077);
or U11238 (N_11238,N_11006,N_11089);
nor U11239 (N_11239,N_11097,N_11023);
xnor U11240 (N_11240,N_11001,N_11055);
nor U11241 (N_11241,N_11085,N_11039);
xor U11242 (N_11242,N_10976,N_11020);
nor U11243 (N_11243,N_11008,N_11018);
xnor U11244 (N_11244,N_10954,N_11054);
or U11245 (N_11245,N_11025,N_11040);
nor U11246 (N_11246,N_11095,N_10991);
nor U11247 (N_11247,N_11088,N_10983);
and U11248 (N_11248,N_10973,N_10963);
xor U11249 (N_11249,N_11009,N_11098);
xor U11250 (N_11250,N_11248,N_11218);
and U11251 (N_11251,N_11220,N_11153);
nor U11252 (N_11252,N_11177,N_11173);
nand U11253 (N_11253,N_11137,N_11238);
xnor U11254 (N_11254,N_11168,N_11205);
xnor U11255 (N_11255,N_11163,N_11126);
nand U11256 (N_11256,N_11132,N_11164);
nor U11257 (N_11257,N_11228,N_11145);
or U11258 (N_11258,N_11107,N_11213);
nor U11259 (N_11259,N_11206,N_11135);
xor U11260 (N_11260,N_11225,N_11224);
and U11261 (N_11261,N_11113,N_11235);
nor U11262 (N_11262,N_11148,N_11130);
nand U11263 (N_11263,N_11109,N_11117);
nand U11264 (N_11264,N_11208,N_11201);
and U11265 (N_11265,N_11156,N_11110);
or U11266 (N_11266,N_11222,N_11158);
or U11267 (N_11267,N_11142,N_11127);
and U11268 (N_11268,N_11155,N_11202);
xor U11269 (N_11269,N_11101,N_11192);
and U11270 (N_11270,N_11169,N_11242);
nor U11271 (N_11271,N_11232,N_11147);
and U11272 (N_11272,N_11118,N_11176);
or U11273 (N_11273,N_11226,N_11245);
xor U11274 (N_11274,N_11239,N_11180);
and U11275 (N_11275,N_11187,N_11151);
xnor U11276 (N_11276,N_11140,N_11179);
xnor U11277 (N_11277,N_11236,N_11112);
or U11278 (N_11278,N_11215,N_11111);
or U11279 (N_11279,N_11181,N_11139);
and U11280 (N_11280,N_11141,N_11197);
xnor U11281 (N_11281,N_11170,N_11157);
nand U11282 (N_11282,N_11152,N_11167);
or U11283 (N_11283,N_11193,N_11178);
nand U11284 (N_11284,N_11183,N_11247);
or U11285 (N_11285,N_11243,N_11150);
xor U11286 (N_11286,N_11203,N_11221);
nor U11287 (N_11287,N_11191,N_11199);
nand U11288 (N_11288,N_11120,N_11161);
nor U11289 (N_11289,N_11108,N_11104);
nand U11290 (N_11290,N_11219,N_11119);
nor U11291 (N_11291,N_11229,N_11122);
nor U11292 (N_11292,N_11166,N_11184);
or U11293 (N_11293,N_11144,N_11223);
xnor U11294 (N_11294,N_11196,N_11241);
xor U11295 (N_11295,N_11214,N_11227);
nor U11296 (N_11296,N_11106,N_11190);
or U11297 (N_11297,N_11233,N_11100);
xor U11298 (N_11298,N_11103,N_11143);
nand U11299 (N_11299,N_11231,N_11165);
nor U11300 (N_11300,N_11114,N_11207);
xnor U11301 (N_11301,N_11131,N_11125);
xnor U11302 (N_11302,N_11171,N_11230);
xnor U11303 (N_11303,N_11105,N_11195);
xor U11304 (N_11304,N_11124,N_11186);
nor U11305 (N_11305,N_11188,N_11216);
and U11306 (N_11306,N_11134,N_11172);
or U11307 (N_11307,N_11149,N_11209);
xnor U11308 (N_11308,N_11182,N_11128);
nor U11309 (N_11309,N_11129,N_11159);
xor U11310 (N_11310,N_11162,N_11211);
or U11311 (N_11311,N_11138,N_11244);
nand U11312 (N_11312,N_11136,N_11212);
nor U11313 (N_11313,N_11246,N_11123);
and U11314 (N_11314,N_11185,N_11240);
or U11315 (N_11315,N_11175,N_11146);
nor U11316 (N_11316,N_11160,N_11115);
xor U11317 (N_11317,N_11249,N_11194);
nor U11318 (N_11318,N_11102,N_11200);
xor U11319 (N_11319,N_11198,N_11234);
nand U11320 (N_11320,N_11121,N_11116);
or U11321 (N_11321,N_11174,N_11133);
and U11322 (N_11322,N_11217,N_11237);
and U11323 (N_11323,N_11210,N_11189);
xor U11324 (N_11324,N_11204,N_11154);
or U11325 (N_11325,N_11177,N_11234);
or U11326 (N_11326,N_11122,N_11113);
or U11327 (N_11327,N_11193,N_11136);
xor U11328 (N_11328,N_11189,N_11125);
or U11329 (N_11329,N_11144,N_11150);
nand U11330 (N_11330,N_11126,N_11113);
or U11331 (N_11331,N_11125,N_11188);
and U11332 (N_11332,N_11225,N_11244);
or U11333 (N_11333,N_11234,N_11186);
xor U11334 (N_11334,N_11130,N_11189);
and U11335 (N_11335,N_11236,N_11180);
nand U11336 (N_11336,N_11190,N_11102);
and U11337 (N_11337,N_11126,N_11114);
nor U11338 (N_11338,N_11148,N_11182);
xnor U11339 (N_11339,N_11134,N_11200);
nor U11340 (N_11340,N_11128,N_11215);
and U11341 (N_11341,N_11196,N_11193);
or U11342 (N_11342,N_11205,N_11101);
nand U11343 (N_11343,N_11130,N_11125);
nand U11344 (N_11344,N_11241,N_11176);
or U11345 (N_11345,N_11242,N_11104);
nor U11346 (N_11346,N_11219,N_11187);
and U11347 (N_11347,N_11120,N_11226);
or U11348 (N_11348,N_11102,N_11165);
xnor U11349 (N_11349,N_11191,N_11139);
nor U11350 (N_11350,N_11203,N_11179);
nor U11351 (N_11351,N_11205,N_11139);
and U11352 (N_11352,N_11210,N_11197);
nor U11353 (N_11353,N_11120,N_11179);
nand U11354 (N_11354,N_11159,N_11157);
nor U11355 (N_11355,N_11235,N_11164);
and U11356 (N_11356,N_11194,N_11210);
and U11357 (N_11357,N_11104,N_11119);
and U11358 (N_11358,N_11223,N_11229);
and U11359 (N_11359,N_11182,N_11165);
xnor U11360 (N_11360,N_11124,N_11129);
nor U11361 (N_11361,N_11221,N_11241);
and U11362 (N_11362,N_11219,N_11207);
and U11363 (N_11363,N_11241,N_11117);
nand U11364 (N_11364,N_11109,N_11243);
or U11365 (N_11365,N_11143,N_11202);
xor U11366 (N_11366,N_11187,N_11227);
nand U11367 (N_11367,N_11205,N_11173);
nand U11368 (N_11368,N_11110,N_11121);
or U11369 (N_11369,N_11153,N_11183);
nor U11370 (N_11370,N_11183,N_11181);
nor U11371 (N_11371,N_11141,N_11102);
nor U11372 (N_11372,N_11225,N_11183);
xnor U11373 (N_11373,N_11183,N_11144);
nand U11374 (N_11374,N_11201,N_11222);
or U11375 (N_11375,N_11150,N_11229);
nor U11376 (N_11376,N_11110,N_11128);
and U11377 (N_11377,N_11173,N_11180);
and U11378 (N_11378,N_11134,N_11206);
nor U11379 (N_11379,N_11243,N_11193);
xnor U11380 (N_11380,N_11152,N_11212);
or U11381 (N_11381,N_11154,N_11225);
and U11382 (N_11382,N_11164,N_11118);
xnor U11383 (N_11383,N_11222,N_11155);
or U11384 (N_11384,N_11163,N_11145);
and U11385 (N_11385,N_11235,N_11221);
or U11386 (N_11386,N_11211,N_11203);
or U11387 (N_11387,N_11204,N_11125);
nand U11388 (N_11388,N_11117,N_11239);
nor U11389 (N_11389,N_11184,N_11140);
nor U11390 (N_11390,N_11156,N_11166);
xor U11391 (N_11391,N_11221,N_11120);
or U11392 (N_11392,N_11115,N_11131);
or U11393 (N_11393,N_11245,N_11117);
nand U11394 (N_11394,N_11148,N_11102);
and U11395 (N_11395,N_11166,N_11220);
xnor U11396 (N_11396,N_11153,N_11221);
nand U11397 (N_11397,N_11230,N_11172);
xnor U11398 (N_11398,N_11158,N_11227);
and U11399 (N_11399,N_11238,N_11180);
and U11400 (N_11400,N_11273,N_11304);
nand U11401 (N_11401,N_11330,N_11263);
or U11402 (N_11402,N_11329,N_11283);
or U11403 (N_11403,N_11396,N_11317);
nand U11404 (N_11404,N_11319,N_11335);
nor U11405 (N_11405,N_11305,N_11256);
nor U11406 (N_11406,N_11261,N_11265);
xor U11407 (N_11407,N_11302,N_11279);
nand U11408 (N_11408,N_11352,N_11311);
xnor U11409 (N_11409,N_11251,N_11376);
or U11410 (N_11410,N_11285,N_11362);
nor U11411 (N_11411,N_11374,N_11277);
nor U11412 (N_11412,N_11295,N_11303);
or U11413 (N_11413,N_11388,N_11339);
or U11414 (N_11414,N_11262,N_11250);
or U11415 (N_11415,N_11340,N_11328);
xor U11416 (N_11416,N_11350,N_11254);
nand U11417 (N_11417,N_11292,N_11392);
nor U11418 (N_11418,N_11391,N_11320);
and U11419 (N_11419,N_11366,N_11397);
nor U11420 (N_11420,N_11346,N_11269);
nand U11421 (N_11421,N_11382,N_11358);
nand U11422 (N_11422,N_11383,N_11378);
or U11423 (N_11423,N_11375,N_11289);
nand U11424 (N_11424,N_11298,N_11314);
nor U11425 (N_11425,N_11343,N_11370);
xnor U11426 (N_11426,N_11258,N_11372);
or U11427 (N_11427,N_11338,N_11360);
xor U11428 (N_11428,N_11337,N_11342);
or U11429 (N_11429,N_11348,N_11336);
nand U11430 (N_11430,N_11299,N_11290);
nand U11431 (N_11431,N_11308,N_11294);
xor U11432 (N_11432,N_11288,N_11260);
xor U11433 (N_11433,N_11291,N_11280);
nand U11434 (N_11434,N_11313,N_11377);
and U11435 (N_11435,N_11268,N_11356);
and U11436 (N_11436,N_11345,N_11384);
nor U11437 (N_11437,N_11363,N_11393);
nand U11438 (N_11438,N_11264,N_11274);
and U11439 (N_11439,N_11322,N_11257);
xnor U11440 (N_11440,N_11287,N_11318);
nor U11441 (N_11441,N_11259,N_11389);
nand U11442 (N_11442,N_11316,N_11398);
nand U11443 (N_11443,N_11325,N_11296);
nand U11444 (N_11444,N_11399,N_11275);
and U11445 (N_11445,N_11349,N_11300);
or U11446 (N_11446,N_11286,N_11379);
or U11447 (N_11447,N_11347,N_11334);
nand U11448 (N_11448,N_11315,N_11381);
nor U11449 (N_11449,N_11365,N_11359);
nor U11450 (N_11450,N_11371,N_11293);
and U11451 (N_11451,N_11327,N_11357);
nand U11452 (N_11452,N_11341,N_11331);
or U11453 (N_11453,N_11361,N_11321);
nor U11454 (N_11454,N_11373,N_11270);
nand U11455 (N_11455,N_11390,N_11369);
and U11456 (N_11456,N_11355,N_11306);
xor U11457 (N_11457,N_11276,N_11353);
or U11458 (N_11458,N_11307,N_11266);
and U11459 (N_11459,N_11351,N_11309);
nand U11460 (N_11460,N_11252,N_11368);
nand U11461 (N_11461,N_11395,N_11385);
nand U11462 (N_11462,N_11394,N_11282);
nor U11463 (N_11463,N_11364,N_11297);
nand U11464 (N_11464,N_11367,N_11387);
nand U11465 (N_11465,N_11332,N_11284);
nand U11466 (N_11466,N_11333,N_11267);
nor U11467 (N_11467,N_11326,N_11278);
or U11468 (N_11468,N_11312,N_11344);
and U11469 (N_11469,N_11380,N_11253);
nand U11470 (N_11470,N_11301,N_11271);
xor U11471 (N_11471,N_11272,N_11281);
or U11472 (N_11472,N_11354,N_11323);
nor U11473 (N_11473,N_11324,N_11386);
xnor U11474 (N_11474,N_11255,N_11310);
xnor U11475 (N_11475,N_11343,N_11372);
nor U11476 (N_11476,N_11397,N_11250);
and U11477 (N_11477,N_11288,N_11357);
and U11478 (N_11478,N_11269,N_11387);
nor U11479 (N_11479,N_11299,N_11355);
and U11480 (N_11480,N_11395,N_11392);
xor U11481 (N_11481,N_11320,N_11295);
nor U11482 (N_11482,N_11350,N_11359);
and U11483 (N_11483,N_11380,N_11265);
and U11484 (N_11484,N_11255,N_11361);
xnor U11485 (N_11485,N_11355,N_11396);
nand U11486 (N_11486,N_11388,N_11357);
nand U11487 (N_11487,N_11276,N_11309);
and U11488 (N_11488,N_11381,N_11268);
xor U11489 (N_11489,N_11368,N_11372);
or U11490 (N_11490,N_11397,N_11378);
and U11491 (N_11491,N_11306,N_11382);
nand U11492 (N_11492,N_11327,N_11252);
or U11493 (N_11493,N_11327,N_11255);
or U11494 (N_11494,N_11254,N_11340);
nor U11495 (N_11495,N_11349,N_11366);
nor U11496 (N_11496,N_11274,N_11282);
nand U11497 (N_11497,N_11398,N_11267);
xor U11498 (N_11498,N_11353,N_11376);
nand U11499 (N_11499,N_11303,N_11382);
and U11500 (N_11500,N_11370,N_11307);
and U11501 (N_11501,N_11310,N_11266);
nor U11502 (N_11502,N_11254,N_11278);
or U11503 (N_11503,N_11341,N_11366);
nor U11504 (N_11504,N_11255,N_11354);
xnor U11505 (N_11505,N_11294,N_11383);
nor U11506 (N_11506,N_11283,N_11279);
and U11507 (N_11507,N_11274,N_11263);
nor U11508 (N_11508,N_11369,N_11355);
nand U11509 (N_11509,N_11313,N_11399);
xor U11510 (N_11510,N_11260,N_11325);
or U11511 (N_11511,N_11323,N_11360);
nor U11512 (N_11512,N_11258,N_11353);
xor U11513 (N_11513,N_11252,N_11339);
xnor U11514 (N_11514,N_11279,N_11258);
nand U11515 (N_11515,N_11397,N_11396);
nand U11516 (N_11516,N_11265,N_11293);
nor U11517 (N_11517,N_11300,N_11395);
and U11518 (N_11518,N_11331,N_11251);
or U11519 (N_11519,N_11333,N_11332);
xnor U11520 (N_11520,N_11255,N_11279);
nor U11521 (N_11521,N_11356,N_11340);
or U11522 (N_11522,N_11319,N_11292);
nor U11523 (N_11523,N_11372,N_11398);
or U11524 (N_11524,N_11332,N_11327);
nor U11525 (N_11525,N_11282,N_11349);
nand U11526 (N_11526,N_11337,N_11262);
nor U11527 (N_11527,N_11358,N_11303);
or U11528 (N_11528,N_11299,N_11366);
xor U11529 (N_11529,N_11331,N_11304);
or U11530 (N_11530,N_11399,N_11277);
xor U11531 (N_11531,N_11264,N_11283);
and U11532 (N_11532,N_11388,N_11364);
or U11533 (N_11533,N_11285,N_11393);
xor U11534 (N_11534,N_11310,N_11384);
or U11535 (N_11535,N_11383,N_11318);
nand U11536 (N_11536,N_11354,N_11325);
and U11537 (N_11537,N_11377,N_11354);
nand U11538 (N_11538,N_11311,N_11398);
xor U11539 (N_11539,N_11366,N_11395);
nor U11540 (N_11540,N_11384,N_11299);
nor U11541 (N_11541,N_11261,N_11351);
and U11542 (N_11542,N_11379,N_11254);
nand U11543 (N_11543,N_11251,N_11337);
or U11544 (N_11544,N_11313,N_11296);
nor U11545 (N_11545,N_11351,N_11294);
and U11546 (N_11546,N_11274,N_11311);
and U11547 (N_11547,N_11261,N_11281);
or U11548 (N_11548,N_11328,N_11263);
or U11549 (N_11549,N_11329,N_11313);
nand U11550 (N_11550,N_11411,N_11528);
nand U11551 (N_11551,N_11533,N_11457);
xor U11552 (N_11552,N_11415,N_11531);
nand U11553 (N_11553,N_11444,N_11450);
nand U11554 (N_11554,N_11493,N_11540);
nor U11555 (N_11555,N_11471,N_11490);
and U11556 (N_11556,N_11539,N_11440);
xor U11557 (N_11557,N_11460,N_11433);
nand U11558 (N_11558,N_11402,N_11547);
nor U11559 (N_11559,N_11403,N_11532);
nor U11560 (N_11560,N_11529,N_11487);
xor U11561 (N_11561,N_11515,N_11431);
and U11562 (N_11562,N_11482,N_11510);
xor U11563 (N_11563,N_11521,N_11489);
xnor U11564 (N_11564,N_11545,N_11409);
xnor U11565 (N_11565,N_11452,N_11435);
nor U11566 (N_11566,N_11463,N_11478);
or U11567 (N_11567,N_11498,N_11430);
nor U11568 (N_11568,N_11494,N_11511);
nor U11569 (N_11569,N_11448,N_11474);
and U11570 (N_11570,N_11462,N_11400);
or U11571 (N_11571,N_11502,N_11479);
and U11572 (N_11572,N_11500,N_11537);
xor U11573 (N_11573,N_11473,N_11512);
and U11574 (N_11574,N_11486,N_11543);
or U11575 (N_11575,N_11416,N_11507);
nor U11576 (N_11576,N_11447,N_11456);
and U11577 (N_11577,N_11509,N_11432);
nand U11578 (N_11578,N_11475,N_11527);
nor U11579 (N_11579,N_11441,N_11434);
and U11580 (N_11580,N_11436,N_11445);
xnor U11581 (N_11581,N_11519,N_11520);
xnor U11582 (N_11582,N_11404,N_11438);
nor U11583 (N_11583,N_11548,N_11405);
nor U11584 (N_11584,N_11499,N_11477);
nand U11585 (N_11585,N_11483,N_11401);
or U11586 (N_11586,N_11413,N_11454);
nor U11587 (N_11587,N_11484,N_11427);
xnor U11588 (N_11588,N_11549,N_11455);
nor U11589 (N_11589,N_11418,N_11513);
nor U11590 (N_11590,N_11536,N_11458);
xnor U11591 (N_11591,N_11469,N_11408);
nor U11592 (N_11592,N_11446,N_11443);
nor U11593 (N_11593,N_11538,N_11535);
and U11594 (N_11594,N_11428,N_11544);
nand U11595 (N_11595,N_11504,N_11406);
xnor U11596 (N_11596,N_11468,N_11451);
nor U11597 (N_11597,N_11476,N_11503);
nand U11598 (N_11598,N_11424,N_11495);
xor U11599 (N_11599,N_11426,N_11467);
nand U11600 (N_11600,N_11453,N_11485);
or U11601 (N_11601,N_11541,N_11423);
or U11602 (N_11602,N_11466,N_11472);
nor U11603 (N_11603,N_11464,N_11488);
and U11604 (N_11604,N_11425,N_11481);
and U11605 (N_11605,N_11523,N_11492);
xor U11606 (N_11606,N_11439,N_11497);
nor U11607 (N_11607,N_11505,N_11437);
or U11608 (N_11608,N_11501,N_11442);
nor U11609 (N_11609,N_11525,N_11496);
nand U11610 (N_11610,N_11526,N_11421);
xor U11611 (N_11611,N_11480,N_11422);
nand U11612 (N_11612,N_11518,N_11420);
and U11613 (N_11613,N_11506,N_11417);
xor U11614 (N_11614,N_11470,N_11516);
nand U11615 (N_11615,N_11465,N_11429);
and U11616 (N_11616,N_11534,N_11449);
xor U11617 (N_11617,N_11508,N_11410);
or U11618 (N_11618,N_11514,N_11412);
xor U11619 (N_11619,N_11530,N_11542);
nand U11620 (N_11620,N_11459,N_11461);
xnor U11621 (N_11621,N_11546,N_11517);
nor U11622 (N_11622,N_11522,N_11491);
or U11623 (N_11623,N_11524,N_11419);
xnor U11624 (N_11624,N_11407,N_11414);
nor U11625 (N_11625,N_11547,N_11423);
xor U11626 (N_11626,N_11459,N_11413);
nand U11627 (N_11627,N_11487,N_11427);
xnor U11628 (N_11628,N_11490,N_11421);
nand U11629 (N_11629,N_11494,N_11424);
nor U11630 (N_11630,N_11410,N_11447);
or U11631 (N_11631,N_11476,N_11433);
or U11632 (N_11632,N_11477,N_11486);
or U11633 (N_11633,N_11448,N_11467);
nor U11634 (N_11634,N_11480,N_11473);
or U11635 (N_11635,N_11452,N_11467);
or U11636 (N_11636,N_11437,N_11429);
or U11637 (N_11637,N_11510,N_11531);
xor U11638 (N_11638,N_11411,N_11417);
and U11639 (N_11639,N_11411,N_11493);
and U11640 (N_11640,N_11438,N_11534);
nor U11641 (N_11641,N_11501,N_11463);
and U11642 (N_11642,N_11419,N_11455);
nor U11643 (N_11643,N_11489,N_11403);
nand U11644 (N_11644,N_11426,N_11481);
or U11645 (N_11645,N_11495,N_11474);
and U11646 (N_11646,N_11523,N_11464);
nand U11647 (N_11647,N_11418,N_11497);
or U11648 (N_11648,N_11424,N_11413);
and U11649 (N_11649,N_11530,N_11423);
and U11650 (N_11650,N_11418,N_11533);
or U11651 (N_11651,N_11489,N_11458);
or U11652 (N_11652,N_11524,N_11512);
nor U11653 (N_11653,N_11521,N_11537);
and U11654 (N_11654,N_11523,N_11540);
nor U11655 (N_11655,N_11491,N_11434);
and U11656 (N_11656,N_11405,N_11524);
nor U11657 (N_11657,N_11478,N_11542);
nand U11658 (N_11658,N_11480,N_11430);
xor U11659 (N_11659,N_11454,N_11462);
xor U11660 (N_11660,N_11438,N_11479);
xor U11661 (N_11661,N_11470,N_11540);
and U11662 (N_11662,N_11430,N_11487);
or U11663 (N_11663,N_11514,N_11473);
and U11664 (N_11664,N_11517,N_11507);
and U11665 (N_11665,N_11495,N_11472);
nand U11666 (N_11666,N_11440,N_11409);
and U11667 (N_11667,N_11450,N_11518);
or U11668 (N_11668,N_11494,N_11455);
and U11669 (N_11669,N_11424,N_11484);
and U11670 (N_11670,N_11495,N_11417);
nor U11671 (N_11671,N_11473,N_11409);
or U11672 (N_11672,N_11495,N_11483);
nand U11673 (N_11673,N_11501,N_11430);
or U11674 (N_11674,N_11472,N_11545);
xor U11675 (N_11675,N_11474,N_11457);
xnor U11676 (N_11676,N_11436,N_11522);
xnor U11677 (N_11677,N_11548,N_11442);
or U11678 (N_11678,N_11510,N_11409);
nor U11679 (N_11679,N_11435,N_11415);
or U11680 (N_11680,N_11492,N_11531);
and U11681 (N_11681,N_11523,N_11496);
xor U11682 (N_11682,N_11466,N_11528);
and U11683 (N_11683,N_11439,N_11483);
nand U11684 (N_11684,N_11532,N_11523);
or U11685 (N_11685,N_11449,N_11454);
or U11686 (N_11686,N_11472,N_11450);
nand U11687 (N_11687,N_11437,N_11538);
nand U11688 (N_11688,N_11493,N_11499);
or U11689 (N_11689,N_11491,N_11514);
nand U11690 (N_11690,N_11418,N_11485);
or U11691 (N_11691,N_11400,N_11425);
nand U11692 (N_11692,N_11526,N_11520);
xor U11693 (N_11693,N_11536,N_11530);
and U11694 (N_11694,N_11434,N_11548);
or U11695 (N_11695,N_11538,N_11435);
nor U11696 (N_11696,N_11436,N_11468);
and U11697 (N_11697,N_11421,N_11542);
nor U11698 (N_11698,N_11484,N_11440);
nand U11699 (N_11699,N_11458,N_11511);
xnor U11700 (N_11700,N_11604,N_11620);
and U11701 (N_11701,N_11621,N_11662);
nand U11702 (N_11702,N_11551,N_11605);
and U11703 (N_11703,N_11645,N_11582);
nor U11704 (N_11704,N_11660,N_11612);
and U11705 (N_11705,N_11656,N_11590);
or U11706 (N_11706,N_11583,N_11692);
nor U11707 (N_11707,N_11616,N_11591);
or U11708 (N_11708,N_11635,N_11668);
and U11709 (N_11709,N_11599,N_11569);
or U11710 (N_11710,N_11588,N_11560);
or U11711 (N_11711,N_11696,N_11699);
or U11712 (N_11712,N_11683,N_11570);
xor U11713 (N_11713,N_11553,N_11644);
xnor U11714 (N_11714,N_11657,N_11653);
and U11715 (N_11715,N_11650,N_11681);
or U11716 (N_11716,N_11623,N_11586);
or U11717 (N_11717,N_11685,N_11627);
nor U11718 (N_11718,N_11587,N_11663);
xnor U11719 (N_11719,N_11563,N_11558);
or U11720 (N_11720,N_11584,N_11694);
nor U11721 (N_11721,N_11684,N_11658);
xnor U11722 (N_11722,N_11652,N_11671);
nand U11723 (N_11723,N_11610,N_11594);
or U11724 (N_11724,N_11608,N_11638);
nor U11725 (N_11725,N_11646,N_11597);
nor U11726 (N_11726,N_11682,N_11667);
and U11727 (N_11727,N_11614,N_11698);
and U11728 (N_11728,N_11555,N_11626);
nor U11729 (N_11729,N_11672,N_11637);
and U11730 (N_11730,N_11617,N_11665);
xnor U11731 (N_11731,N_11554,N_11559);
nor U11732 (N_11732,N_11691,N_11648);
and U11733 (N_11733,N_11647,N_11565);
xor U11734 (N_11734,N_11581,N_11598);
xor U11735 (N_11735,N_11592,N_11589);
and U11736 (N_11736,N_11550,N_11639);
nand U11737 (N_11737,N_11628,N_11634);
or U11738 (N_11738,N_11571,N_11643);
nand U11739 (N_11739,N_11636,N_11689);
and U11740 (N_11740,N_11651,N_11673);
xnor U11741 (N_11741,N_11675,N_11687);
or U11742 (N_11742,N_11686,N_11697);
xnor U11743 (N_11743,N_11602,N_11625);
nor U11744 (N_11744,N_11601,N_11659);
nand U11745 (N_11745,N_11611,N_11572);
and U11746 (N_11746,N_11661,N_11688);
nor U11747 (N_11747,N_11593,N_11670);
nand U11748 (N_11748,N_11679,N_11640);
xnor U11749 (N_11749,N_11566,N_11561);
nand U11750 (N_11750,N_11632,N_11624);
nor U11751 (N_11751,N_11690,N_11630);
nand U11752 (N_11752,N_11654,N_11595);
nor U11753 (N_11753,N_11603,N_11655);
or U11754 (N_11754,N_11633,N_11578);
or U11755 (N_11755,N_11577,N_11556);
or U11756 (N_11756,N_11573,N_11600);
and U11757 (N_11757,N_11585,N_11609);
or U11758 (N_11758,N_11552,N_11677);
nor U11759 (N_11759,N_11580,N_11574);
or U11760 (N_11760,N_11606,N_11596);
and U11761 (N_11761,N_11674,N_11618);
and U11762 (N_11762,N_11693,N_11615);
and U11763 (N_11763,N_11619,N_11579);
nor U11764 (N_11764,N_11629,N_11641);
nor U11765 (N_11765,N_11564,N_11695);
nor U11766 (N_11766,N_11613,N_11669);
and U11767 (N_11767,N_11680,N_11622);
and U11768 (N_11768,N_11649,N_11576);
or U11769 (N_11769,N_11568,N_11631);
nand U11770 (N_11770,N_11678,N_11664);
nor U11771 (N_11771,N_11666,N_11562);
and U11772 (N_11772,N_11642,N_11607);
or U11773 (N_11773,N_11567,N_11557);
nand U11774 (N_11774,N_11676,N_11575);
nand U11775 (N_11775,N_11579,N_11592);
nand U11776 (N_11776,N_11679,N_11670);
nor U11777 (N_11777,N_11598,N_11592);
nand U11778 (N_11778,N_11594,N_11618);
nand U11779 (N_11779,N_11641,N_11694);
nand U11780 (N_11780,N_11574,N_11661);
xor U11781 (N_11781,N_11607,N_11632);
or U11782 (N_11782,N_11655,N_11573);
and U11783 (N_11783,N_11595,N_11559);
and U11784 (N_11784,N_11694,N_11681);
nor U11785 (N_11785,N_11597,N_11618);
nand U11786 (N_11786,N_11567,N_11651);
and U11787 (N_11787,N_11559,N_11630);
or U11788 (N_11788,N_11655,N_11560);
and U11789 (N_11789,N_11562,N_11617);
nand U11790 (N_11790,N_11620,N_11654);
xnor U11791 (N_11791,N_11639,N_11562);
or U11792 (N_11792,N_11565,N_11615);
or U11793 (N_11793,N_11575,N_11597);
xnor U11794 (N_11794,N_11634,N_11648);
xor U11795 (N_11795,N_11563,N_11667);
or U11796 (N_11796,N_11588,N_11686);
and U11797 (N_11797,N_11594,N_11617);
nand U11798 (N_11798,N_11553,N_11698);
nor U11799 (N_11799,N_11573,N_11565);
or U11800 (N_11800,N_11621,N_11553);
or U11801 (N_11801,N_11581,N_11606);
xnor U11802 (N_11802,N_11630,N_11580);
and U11803 (N_11803,N_11699,N_11638);
nor U11804 (N_11804,N_11581,N_11672);
nand U11805 (N_11805,N_11597,N_11599);
xnor U11806 (N_11806,N_11667,N_11678);
or U11807 (N_11807,N_11599,N_11636);
nand U11808 (N_11808,N_11684,N_11674);
nor U11809 (N_11809,N_11652,N_11639);
xnor U11810 (N_11810,N_11611,N_11567);
nand U11811 (N_11811,N_11605,N_11604);
xnor U11812 (N_11812,N_11618,N_11644);
nor U11813 (N_11813,N_11630,N_11562);
nor U11814 (N_11814,N_11633,N_11667);
nor U11815 (N_11815,N_11649,N_11640);
and U11816 (N_11816,N_11616,N_11655);
nor U11817 (N_11817,N_11629,N_11604);
or U11818 (N_11818,N_11624,N_11616);
xnor U11819 (N_11819,N_11576,N_11678);
xnor U11820 (N_11820,N_11670,N_11572);
xor U11821 (N_11821,N_11619,N_11661);
and U11822 (N_11822,N_11667,N_11623);
xor U11823 (N_11823,N_11669,N_11662);
xor U11824 (N_11824,N_11598,N_11557);
nor U11825 (N_11825,N_11558,N_11617);
nor U11826 (N_11826,N_11676,N_11571);
and U11827 (N_11827,N_11569,N_11554);
or U11828 (N_11828,N_11560,N_11589);
and U11829 (N_11829,N_11564,N_11560);
or U11830 (N_11830,N_11641,N_11602);
nor U11831 (N_11831,N_11569,N_11634);
xor U11832 (N_11832,N_11643,N_11576);
nand U11833 (N_11833,N_11628,N_11674);
nand U11834 (N_11834,N_11568,N_11620);
xor U11835 (N_11835,N_11652,N_11617);
and U11836 (N_11836,N_11669,N_11630);
nand U11837 (N_11837,N_11694,N_11657);
nor U11838 (N_11838,N_11667,N_11637);
and U11839 (N_11839,N_11609,N_11631);
nor U11840 (N_11840,N_11553,N_11647);
nor U11841 (N_11841,N_11573,N_11566);
nor U11842 (N_11842,N_11621,N_11679);
xor U11843 (N_11843,N_11580,N_11572);
xnor U11844 (N_11844,N_11683,N_11658);
nand U11845 (N_11845,N_11578,N_11677);
nor U11846 (N_11846,N_11580,N_11662);
or U11847 (N_11847,N_11588,N_11580);
nand U11848 (N_11848,N_11610,N_11650);
xnor U11849 (N_11849,N_11580,N_11589);
and U11850 (N_11850,N_11772,N_11797);
xor U11851 (N_11851,N_11704,N_11796);
xnor U11852 (N_11852,N_11701,N_11751);
nand U11853 (N_11853,N_11725,N_11821);
nand U11854 (N_11854,N_11744,N_11803);
or U11855 (N_11855,N_11716,N_11711);
and U11856 (N_11856,N_11741,N_11707);
xnor U11857 (N_11857,N_11732,N_11739);
or U11858 (N_11858,N_11777,N_11717);
xnor U11859 (N_11859,N_11748,N_11786);
xor U11860 (N_11860,N_11802,N_11763);
xor U11861 (N_11861,N_11767,N_11815);
nor U11862 (N_11862,N_11787,N_11849);
xor U11863 (N_11863,N_11708,N_11747);
and U11864 (N_11864,N_11773,N_11793);
nand U11865 (N_11865,N_11820,N_11718);
and U11866 (N_11866,N_11722,N_11745);
and U11867 (N_11867,N_11844,N_11781);
nor U11868 (N_11868,N_11771,N_11749);
and U11869 (N_11869,N_11761,N_11729);
nor U11870 (N_11870,N_11835,N_11733);
xnor U11871 (N_11871,N_11789,N_11715);
nand U11872 (N_11872,N_11834,N_11798);
nand U11873 (N_11873,N_11764,N_11782);
nor U11874 (N_11874,N_11770,N_11847);
nor U11875 (N_11875,N_11817,N_11780);
and U11876 (N_11876,N_11827,N_11814);
nand U11877 (N_11877,N_11736,N_11700);
or U11878 (N_11878,N_11728,N_11735);
and U11879 (N_11879,N_11848,N_11709);
xnor U11880 (N_11880,N_11843,N_11734);
nor U11881 (N_11881,N_11775,N_11792);
xnor U11882 (N_11882,N_11737,N_11810);
nor U11883 (N_11883,N_11833,N_11731);
and U11884 (N_11884,N_11774,N_11723);
nand U11885 (N_11885,N_11839,N_11762);
nand U11886 (N_11886,N_11742,N_11807);
nand U11887 (N_11887,N_11738,N_11829);
and U11888 (N_11888,N_11754,N_11826);
or U11889 (N_11889,N_11705,N_11808);
nand U11890 (N_11890,N_11765,N_11750);
or U11891 (N_11891,N_11769,N_11788);
nor U11892 (N_11892,N_11753,N_11719);
nand U11893 (N_11893,N_11778,N_11818);
xor U11894 (N_11894,N_11743,N_11783);
and U11895 (N_11895,N_11756,N_11760);
nor U11896 (N_11896,N_11813,N_11779);
nor U11897 (N_11897,N_11846,N_11811);
nand U11898 (N_11898,N_11816,N_11812);
or U11899 (N_11899,N_11819,N_11713);
nand U11900 (N_11900,N_11804,N_11785);
xor U11901 (N_11901,N_11831,N_11795);
nand U11902 (N_11902,N_11720,N_11836);
or U11903 (N_11903,N_11824,N_11805);
nor U11904 (N_11904,N_11766,N_11830);
and U11905 (N_11905,N_11740,N_11721);
nand U11906 (N_11906,N_11825,N_11710);
and U11907 (N_11907,N_11706,N_11790);
nor U11908 (N_11908,N_11759,N_11758);
nand U11909 (N_11909,N_11791,N_11832);
nand U11910 (N_11910,N_11806,N_11837);
or U11911 (N_11911,N_11822,N_11752);
xor U11912 (N_11912,N_11712,N_11838);
nor U11913 (N_11913,N_11730,N_11784);
xor U11914 (N_11914,N_11768,N_11801);
nor U11915 (N_11915,N_11757,N_11799);
or U11916 (N_11916,N_11841,N_11823);
and U11917 (N_11917,N_11714,N_11726);
nand U11918 (N_11918,N_11702,N_11724);
or U11919 (N_11919,N_11776,N_11755);
or U11920 (N_11920,N_11746,N_11842);
nand U11921 (N_11921,N_11703,N_11809);
and U11922 (N_11922,N_11840,N_11800);
and U11923 (N_11923,N_11828,N_11727);
nand U11924 (N_11924,N_11794,N_11845);
nor U11925 (N_11925,N_11838,N_11782);
or U11926 (N_11926,N_11700,N_11779);
nand U11927 (N_11927,N_11846,N_11844);
xnor U11928 (N_11928,N_11773,N_11827);
xor U11929 (N_11929,N_11769,N_11807);
nor U11930 (N_11930,N_11778,N_11720);
and U11931 (N_11931,N_11846,N_11751);
or U11932 (N_11932,N_11740,N_11815);
or U11933 (N_11933,N_11752,N_11737);
nor U11934 (N_11934,N_11827,N_11807);
and U11935 (N_11935,N_11771,N_11709);
nor U11936 (N_11936,N_11709,N_11802);
or U11937 (N_11937,N_11730,N_11807);
or U11938 (N_11938,N_11712,N_11739);
xor U11939 (N_11939,N_11780,N_11723);
nand U11940 (N_11940,N_11819,N_11700);
or U11941 (N_11941,N_11846,N_11708);
or U11942 (N_11942,N_11803,N_11805);
and U11943 (N_11943,N_11734,N_11744);
xor U11944 (N_11944,N_11728,N_11805);
nand U11945 (N_11945,N_11712,N_11703);
and U11946 (N_11946,N_11737,N_11803);
and U11947 (N_11947,N_11777,N_11835);
nor U11948 (N_11948,N_11705,N_11831);
nor U11949 (N_11949,N_11717,N_11745);
xor U11950 (N_11950,N_11841,N_11781);
and U11951 (N_11951,N_11810,N_11719);
nand U11952 (N_11952,N_11791,N_11847);
xnor U11953 (N_11953,N_11757,N_11731);
and U11954 (N_11954,N_11730,N_11843);
nand U11955 (N_11955,N_11721,N_11709);
nor U11956 (N_11956,N_11762,N_11740);
nand U11957 (N_11957,N_11823,N_11748);
xnor U11958 (N_11958,N_11736,N_11718);
or U11959 (N_11959,N_11785,N_11783);
nand U11960 (N_11960,N_11767,N_11819);
nor U11961 (N_11961,N_11730,N_11767);
or U11962 (N_11962,N_11827,N_11793);
nand U11963 (N_11963,N_11799,N_11820);
and U11964 (N_11964,N_11804,N_11777);
or U11965 (N_11965,N_11838,N_11800);
nand U11966 (N_11966,N_11714,N_11829);
nor U11967 (N_11967,N_11728,N_11741);
or U11968 (N_11968,N_11730,N_11782);
and U11969 (N_11969,N_11756,N_11815);
xnor U11970 (N_11970,N_11818,N_11706);
or U11971 (N_11971,N_11739,N_11733);
or U11972 (N_11972,N_11771,N_11791);
xnor U11973 (N_11973,N_11731,N_11700);
nor U11974 (N_11974,N_11823,N_11710);
nand U11975 (N_11975,N_11759,N_11750);
xor U11976 (N_11976,N_11772,N_11734);
nor U11977 (N_11977,N_11775,N_11727);
xnor U11978 (N_11978,N_11770,N_11804);
nor U11979 (N_11979,N_11700,N_11809);
nand U11980 (N_11980,N_11763,N_11716);
or U11981 (N_11981,N_11803,N_11843);
or U11982 (N_11982,N_11832,N_11714);
and U11983 (N_11983,N_11711,N_11714);
or U11984 (N_11984,N_11749,N_11831);
nor U11985 (N_11985,N_11762,N_11705);
xnor U11986 (N_11986,N_11847,N_11743);
xnor U11987 (N_11987,N_11790,N_11827);
and U11988 (N_11988,N_11836,N_11829);
or U11989 (N_11989,N_11740,N_11826);
and U11990 (N_11990,N_11773,N_11706);
xnor U11991 (N_11991,N_11790,N_11787);
nor U11992 (N_11992,N_11705,N_11718);
and U11993 (N_11993,N_11821,N_11700);
nor U11994 (N_11994,N_11843,N_11827);
nand U11995 (N_11995,N_11815,N_11842);
and U11996 (N_11996,N_11781,N_11824);
xor U11997 (N_11997,N_11745,N_11726);
and U11998 (N_11998,N_11746,N_11806);
xor U11999 (N_11999,N_11810,N_11817);
and U12000 (N_12000,N_11985,N_11995);
xnor U12001 (N_12001,N_11881,N_11896);
xor U12002 (N_12002,N_11931,N_11935);
and U12003 (N_12003,N_11867,N_11928);
nor U12004 (N_12004,N_11877,N_11869);
or U12005 (N_12005,N_11893,N_11960);
nor U12006 (N_12006,N_11970,N_11929);
xnor U12007 (N_12007,N_11904,N_11964);
nand U12008 (N_12008,N_11954,N_11938);
nand U12009 (N_12009,N_11974,N_11897);
nor U12010 (N_12010,N_11882,N_11856);
nand U12011 (N_12011,N_11857,N_11955);
xnor U12012 (N_12012,N_11949,N_11965);
nand U12013 (N_12013,N_11959,N_11899);
xor U12014 (N_12014,N_11913,N_11933);
xor U12015 (N_12015,N_11875,N_11989);
nor U12016 (N_12016,N_11906,N_11879);
nand U12017 (N_12017,N_11924,N_11852);
xor U12018 (N_12018,N_11874,N_11982);
nor U12019 (N_12019,N_11914,N_11975);
nand U12020 (N_12020,N_11891,N_11939);
or U12021 (N_12021,N_11862,N_11866);
or U12022 (N_12022,N_11890,N_11872);
nor U12023 (N_12023,N_11968,N_11999);
nor U12024 (N_12024,N_11909,N_11947);
nor U12025 (N_12025,N_11958,N_11926);
nand U12026 (N_12026,N_11903,N_11851);
and U12027 (N_12027,N_11859,N_11957);
or U12028 (N_12028,N_11973,N_11981);
and U12029 (N_12029,N_11969,N_11988);
nor U12030 (N_12030,N_11894,N_11898);
nor U12031 (N_12031,N_11919,N_11977);
or U12032 (N_12032,N_11936,N_11943);
or U12033 (N_12033,N_11971,N_11868);
nand U12034 (N_12034,N_11983,N_11907);
or U12035 (N_12035,N_11997,N_11941);
and U12036 (N_12036,N_11887,N_11912);
xnor U12037 (N_12037,N_11861,N_11902);
nand U12038 (N_12038,N_11863,N_11873);
nor U12039 (N_12039,N_11987,N_11986);
nand U12040 (N_12040,N_11915,N_11900);
nor U12041 (N_12041,N_11910,N_11880);
and U12042 (N_12042,N_11916,N_11923);
and U12043 (N_12043,N_11911,N_11963);
nor U12044 (N_12044,N_11991,N_11972);
or U12045 (N_12045,N_11883,N_11967);
xnor U12046 (N_12046,N_11918,N_11922);
nor U12047 (N_12047,N_11876,N_11853);
nor U12048 (N_12048,N_11889,N_11864);
nor U12049 (N_12049,N_11961,N_11962);
nand U12050 (N_12050,N_11920,N_11990);
and U12051 (N_12051,N_11927,N_11950);
nor U12052 (N_12052,N_11858,N_11952);
nand U12053 (N_12053,N_11871,N_11886);
nand U12054 (N_12054,N_11895,N_11984);
nor U12055 (N_12055,N_11946,N_11951);
xor U12056 (N_12056,N_11937,N_11966);
nor U12057 (N_12057,N_11901,N_11878);
nand U12058 (N_12058,N_11932,N_11884);
or U12059 (N_12059,N_11992,N_11940);
nand U12060 (N_12060,N_11855,N_11953);
nor U12061 (N_12061,N_11944,N_11925);
or U12062 (N_12062,N_11948,N_11917);
nor U12063 (N_12063,N_11942,N_11850);
or U12064 (N_12064,N_11976,N_11934);
and U12065 (N_12065,N_11993,N_11956);
and U12066 (N_12066,N_11870,N_11854);
nor U12067 (N_12067,N_11980,N_11945);
nand U12068 (N_12068,N_11888,N_11885);
or U12069 (N_12069,N_11865,N_11996);
xnor U12070 (N_12070,N_11994,N_11998);
or U12071 (N_12071,N_11930,N_11905);
xnor U12072 (N_12072,N_11860,N_11979);
nor U12073 (N_12073,N_11978,N_11892);
nor U12074 (N_12074,N_11908,N_11921);
nor U12075 (N_12075,N_11922,N_11967);
nand U12076 (N_12076,N_11908,N_11864);
xnor U12077 (N_12077,N_11871,N_11960);
and U12078 (N_12078,N_11892,N_11887);
and U12079 (N_12079,N_11887,N_11888);
xor U12080 (N_12080,N_11976,N_11886);
and U12081 (N_12081,N_11855,N_11973);
xor U12082 (N_12082,N_11899,N_11966);
and U12083 (N_12083,N_11893,N_11870);
xnor U12084 (N_12084,N_11886,N_11917);
and U12085 (N_12085,N_11940,N_11934);
xnor U12086 (N_12086,N_11999,N_11950);
nor U12087 (N_12087,N_11976,N_11867);
nand U12088 (N_12088,N_11864,N_11854);
xnor U12089 (N_12089,N_11883,N_11914);
nor U12090 (N_12090,N_11867,N_11878);
and U12091 (N_12091,N_11993,N_11943);
xnor U12092 (N_12092,N_11878,N_11916);
xnor U12093 (N_12093,N_11874,N_11963);
or U12094 (N_12094,N_11885,N_11948);
or U12095 (N_12095,N_11966,N_11913);
or U12096 (N_12096,N_11987,N_11888);
nand U12097 (N_12097,N_11893,N_11909);
or U12098 (N_12098,N_11924,N_11883);
nand U12099 (N_12099,N_11944,N_11963);
and U12100 (N_12100,N_11851,N_11880);
nor U12101 (N_12101,N_11953,N_11904);
or U12102 (N_12102,N_11890,N_11927);
xor U12103 (N_12103,N_11914,N_11913);
and U12104 (N_12104,N_11983,N_11950);
xor U12105 (N_12105,N_11916,N_11902);
nor U12106 (N_12106,N_11961,N_11940);
and U12107 (N_12107,N_11900,N_11906);
xor U12108 (N_12108,N_11938,N_11893);
and U12109 (N_12109,N_11882,N_11854);
or U12110 (N_12110,N_11990,N_11912);
and U12111 (N_12111,N_11871,N_11876);
or U12112 (N_12112,N_11961,N_11958);
nand U12113 (N_12113,N_11872,N_11960);
nor U12114 (N_12114,N_11911,N_11973);
nor U12115 (N_12115,N_11918,N_11894);
nor U12116 (N_12116,N_11964,N_11991);
nand U12117 (N_12117,N_11851,N_11895);
or U12118 (N_12118,N_11982,N_11890);
xnor U12119 (N_12119,N_11994,N_11902);
xor U12120 (N_12120,N_11855,N_11969);
and U12121 (N_12121,N_11994,N_11922);
or U12122 (N_12122,N_11979,N_11974);
nor U12123 (N_12123,N_11874,N_11969);
xnor U12124 (N_12124,N_11953,N_11948);
nand U12125 (N_12125,N_11884,N_11966);
xor U12126 (N_12126,N_11925,N_11937);
nor U12127 (N_12127,N_11892,N_11993);
and U12128 (N_12128,N_11873,N_11969);
and U12129 (N_12129,N_11919,N_11950);
nand U12130 (N_12130,N_11911,N_11927);
nor U12131 (N_12131,N_11871,N_11866);
xnor U12132 (N_12132,N_11983,N_11915);
nor U12133 (N_12133,N_11933,N_11859);
nor U12134 (N_12134,N_11963,N_11929);
and U12135 (N_12135,N_11959,N_11884);
nor U12136 (N_12136,N_11944,N_11914);
and U12137 (N_12137,N_11854,N_11990);
xnor U12138 (N_12138,N_11929,N_11924);
or U12139 (N_12139,N_11856,N_11986);
and U12140 (N_12140,N_11896,N_11884);
or U12141 (N_12141,N_11992,N_11959);
and U12142 (N_12142,N_11857,N_11971);
nand U12143 (N_12143,N_11998,N_11907);
or U12144 (N_12144,N_11938,N_11947);
xnor U12145 (N_12145,N_11932,N_11881);
xor U12146 (N_12146,N_11893,N_11987);
and U12147 (N_12147,N_11987,N_11896);
and U12148 (N_12148,N_11982,N_11905);
or U12149 (N_12149,N_11973,N_11986);
nor U12150 (N_12150,N_12055,N_12132);
or U12151 (N_12151,N_12095,N_12082);
nor U12152 (N_12152,N_12036,N_12124);
nor U12153 (N_12153,N_12049,N_12080);
nand U12154 (N_12154,N_12064,N_12134);
nand U12155 (N_12155,N_12056,N_12065);
nand U12156 (N_12156,N_12106,N_12071);
nand U12157 (N_12157,N_12020,N_12072);
or U12158 (N_12158,N_12041,N_12146);
nand U12159 (N_12159,N_12089,N_12112);
nand U12160 (N_12160,N_12116,N_12048);
xnor U12161 (N_12161,N_12046,N_12047);
or U12162 (N_12162,N_12001,N_12085);
and U12163 (N_12163,N_12037,N_12032);
xnor U12164 (N_12164,N_12127,N_12052);
or U12165 (N_12165,N_12019,N_12137);
xnor U12166 (N_12166,N_12148,N_12029);
or U12167 (N_12167,N_12038,N_12119);
and U12168 (N_12168,N_12123,N_12003);
xnor U12169 (N_12169,N_12070,N_12053);
nand U12170 (N_12170,N_12060,N_12040);
nand U12171 (N_12171,N_12002,N_12147);
or U12172 (N_12172,N_12097,N_12111);
nor U12173 (N_12173,N_12098,N_12075);
and U12174 (N_12174,N_12028,N_12135);
nand U12175 (N_12175,N_12121,N_12078);
and U12176 (N_12176,N_12144,N_12043);
nor U12177 (N_12177,N_12073,N_12039);
or U12178 (N_12178,N_12079,N_12058);
xnor U12179 (N_12179,N_12015,N_12008);
xor U12180 (N_12180,N_12105,N_12012);
or U12181 (N_12181,N_12133,N_12027);
and U12182 (N_12182,N_12094,N_12013);
xor U12183 (N_12183,N_12061,N_12100);
xnor U12184 (N_12184,N_12118,N_12138);
and U12185 (N_12185,N_12125,N_12142);
xnor U12186 (N_12186,N_12074,N_12059);
or U12187 (N_12187,N_12129,N_12145);
or U12188 (N_12188,N_12107,N_12077);
nor U12189 (N_12189,N_12057,N_12050);
or U12190 (N_12190,N_12051,N_12113);
nand U12191 (N_12191,N_12131,N_12143);
xor U12192 (N_12192,N_12031,N_12025);
xor U12193 (N_12193,N_12130,N_12018);
nand U12194 (N_12194,N_12076,N_12005);
xor U12195 (N_12195,N_12045,N_12091);
and U12196 (N_12196,N_12021,N_12108);
or U12197 (N_12197,N_12092,N_12007);
or U12198 (N_12198,N_12000,N_12115);
xor U12199 (N_12199,N_12069,N_12011);
nor U12200 (N_12200,N_12068,N_12054);
nor U12201 (N_12201,N_12104,N_12030);
nand U12202 (N_12202,N_12033,N_12023);
or U12203 (N_12203,N_12103,N_12016);
xor U12204 (N_12204,N_12084,N_12004);
and U12205 (N_12205,N_12009,N_12026);
and U12206 (N_12206,N_12122,N_12126);
or U12207 (N_12207,N_12088,N_12022);
xor U12208 (N_12208,N_12141,N_12063);
or U12209 (N_12209,N_12110,N_12117);
and U12210 (N_12210,N_12114,N_12042);
or U12211 (N_12211,N_12149,N_12017);
nand U12212 (N_12212,N_12128,N_12102);
or U12213 (N_12213,N_12010,N_12024);
nor U12214 (N_12214,N_12087,N_12006);
and U12215 (N_12215,N_12044,N_12067);
xnor U12216 (N_12216,N_12034,N_12035);
nand U12217 (N_12217,N_12083,N_12066);
and U12218 (N_12218,N_12096,N_12062);
or U12219 (N_12219,N_12093,N_12136);
xor U12220 (N_12220,N_12086,N_12081);
or U12221 (N_12221,N_12140,N_12014);
xor U12222 (N_12222,N_12139,N_12101);
or U12223 (N_12223,N_12099,N_12120);
nand U12224 (N_12224,N_12109,N_12090);
nor U12225 (N_12225,N_12081,N_12111);
or U12226 (N_12226,N_12056,N_12059);
or U12227 (N_12227,N_12127,N_12032);
nand U12228 (N_12228,N_12137,N_12059);
or U12229 (N_12229,N_12146,N_12005);
xor U12230 (N_12230,N_12036,N_12055);
or U12231 (N_12231,N_12139,N_12079);
and U12232 (N_12232,N_12076,N_12095);
nand U12233 (N_12233,N_12051,N_12071);
or U12234 (N_12234,N_12090,N_12091);
nor U12235 (N_12235,N_12007,N_12002);
nand U12236 (N_12236,N_12048,N_12101);
xnor U12237 (N_12237,N_12095,N_12121);
nand U12238 (N_12238,N_12066,N_12073);
nor U12239 (N_12239,N_12070,N_12062);
nor U12240 (N_12240,N_12060,N_12056);
nor U12241 (N_12241,N_12085,N_12038);
and U12242 (N_12242,N_12080,N_12084);
or U12243 (N_12243,N_12003,N_12031);
nor U12244 (N_12244,N_12095,N_12024);
xor U12245 (N_12245,N_12147,N_12101);
xnor U12246 (N_12246,N_12116,N_12032);
xnor U12247 (N_12247,N_12072,N_12139);
or U12248 (N_12248,N_12048,N_12107);
or U12249 (N_12249,N_12128,N_12031);
and U12250 (N_12250,N_12000,N_12102);
xor U12251 (N_12251,N_12107,N_12012);
xnor U12252 (N_12252,N_12041,N_12068);
or U12253 (N_12253,N_12140,N_12113);
and U12254 (N_12254,N_12043,N_12146);
or U12255 (N_12255,N_12014,N_12065);
nand U12256 (N_12256,N_12095,N_12088);
nor U12257 (N_12257,N_12113,N_12146);
xnor U12258 (N_12258,N_12134,N_12116);
xor U12259 (N_12259,N_12047,N_12109);
xnor U12260 (N_12260,N_12013,N_12095);
xor U12261 (N_12261,N_12102,N_12062);
nand U12262 (N_12262,N_12089,N_12027);
nor U12263 (N_12263,N_12146,N_12025);
nand U12264 (N_12264,N_12057,N_12004);
or U12265 (N_12265,N_12077,N_12119);
nor U12266 (N_12266,N_12042,N_12067);
nand U12267 (N_12267,N_12046,N_12141);
nand U12268 (N_12268,N_12036,N_12069);
nor U12269 (N_12269,N_12105,N_12076);
or U12270 (N_12270,N_12033,N_12074);
nor U12271 (N_12271,N_12078,N_12081);
and U12272 (N_12272,N_12048,N_12031);
or U12273 (N_12273,N_12051,N_12068);
nand U12274 (N_12274,N_12119,N_12095);
nor U12275 (N_12275,N_12038,N_12008);
or U12276 (N_12276,N_12092,N_12053);
or U12277 (N_12277,N_12035,N_12005);
xnor U12278 (N_12278,N_12143,N_12089);
xnor U12279 (N_12279,N_12040,N_12075);
nand U12280 (N_12280,N_12086,N_12025);
nor U12281 (N_12281,N_12058,N_12090);
or U12282 (N_12282,N_12093,N_12069);
nand U12283 (N_12283,N_12021,N_12128);
nand U12284 (N_12284,N_12077,N_12109);
nand U12285 (N_12285,N_12013,N_12063);
or U12286 (N_12286,N_12084,N_12083);
nor U12287 (N_12287,N_12149,N_12004);
nor U12288 (N_12288,N_12062,N_12089);
and U12289 (N_12289,N_12128,N_12114);
nor U12290 (N_12290,N_12042,N_12008);
xnor U12291 (N_12291,N_12053,N_12147);
nor U12292 (N_12292,N_12106,N_12115);
nand U12293 (N_12293,N_12040,N_12112);
nor U12294 (N_12294,N_12062,N_12050);
xnor U12295 (N_12295,N_12129,N_12021);
nand U12296 (N_12296,N_12129,N_12013);
xor U12297 (N_12297,N_12021,N_12035);
nand U12298 (N_12298,N_12066,N_12076);
and U12299 (N_12299,N_12073,N_12131);
xnor U12300 (N_12300,N_12265,N_12226);
xnor U12301 (N_12301,N_12222,N_12180);
nand U12302 (N_12302,N_12295,N_12275);
nor U12303 (N_12303,N_12190,N_12266);
and U12304 (N_12304,N_12267,N_12168);
nand U12305 (N_12305,N_12291,N_12274);
or U12306 (N_12306,N_12280,N_12200);
nand U12307 (N_12307,N_12262,N_12175);
nand U12308 (N_12308,N_12252,N_12227);
and U12309 (N_12309,N_12297,N_12202);
and U12310 (N_12310,N_12238,N_12240);
and U12311 (N_12311,N_12272,N_12235);
nand U12312 (N_12312,N_12229,N_12296);
nand U12313 (N_12313,N_12203,N_12178);
nor U12314 (N_12314,N_12268,N_12153);
nor U12315 (N_12315,N_12288,N_12255);
or U12316 (N_12316,N_12273,N_12259);
nand U12317 (N_12317,N_12218,N_12276);
nand U12318 (N_12318,N_12177,N_12174);
nand U12319 (N_12319,N_12264,N_12209);
nor U12320 (N_12320,N_12208,N_12204);
xor U12321 (N_12321,N_12206,N_12198);
xor U12322 (N_12322,N_12160,N_12271);
nand U12323 (N_12323,N_12246,N_12199);
nand U12324 (N_12324,N_12249,N_12294);
nand U12325 (N_12325,N_12161,N_12152);
xor U12326 (N_12326,N_12283,N_12247);
xor U12327 (N_12327,N_12231,N_12224);
xnor U12328 (N_12328,N_12256,N_12181);
or U12329 (N_12329,N_12213,N_12292);
nor U12330 (N_12330,N_12170,N_12237);
nor U12331 (N_12331,N_12263,N_12269);
nor U12332 (N_12332,N_12156,N_12155);
xor U12333 (N_12333,N_12277,N_12233);
xor U12334 (N_12334,N_12228,N_12234);
nand U12335 (N_12335,N_12220,N_12197);
nand U12336 (N_12336,N_12164,N_12248);
nor U12337 (N_12337,N_12253,N_12225);
nor U12338 (N_12338,N_12282,N_12230);
or U12339 (N_12339,N_12214,N_12261);
and U12340 (N_12340,N_12165,N_12278);
xnor U12341 (N_12341,N_12167,N_12151);
xnor U12342 (N_12342,N_12254,N_12219);
nand U12343 (N_12343,N_12281,N_12195);
nand U12344 (N_12344,N_12290,N_12162);
or U12345 (N_12345,N_12211,N_12182);
nor U12346 (N_12346,N_12166,N_12194);
nor U12347 (N_12347,N_12286,N_12205);
nor U12348 (N_12348,N_12169,N_12287);
or U12349 (N_12349,N_12221,N_12207);
nand U12350 (N_12350,N_12158,N_12212);
nand U12351 (N_12351,N_12239,N_12258);
nand U12352 (N_12352,N_12216,N_12210);
or U12353 (N_12353,N_12201,N_12186);
xor U12354 (N_12354,N_12298,N_12223);
nand U12355 (N_12355,N_12251,N_12257);
nand U12356 (N_12356,N_12236,N_12184);
and U12357 (N_12357,N_12215,N_12243);
and U12358 (N_12358,N_12157,N_12173);
nor U12359 (N_12359,N_12260,N_12293);
or U12360 (N_12360,N_12244,N_12241);
or U12361 (N_12361,N_12284,N_12171);
nand U12362 (N_12362,N_12154,N_12192);
and U12363 (N_12363,N_12189,N_12188);
or U12364 (N_12364,N_12242,N_12289);
nor U12365 (N_12365,N_12232,N_12191);
nand U12366 (N_12366,N_12159,N_12299);
or U12367 (N_12367,N_12179,N_12185);
nor U12368 (N_12368,N_12176,N_12193);
xor U12369 (N_12369,N_12285,N_12150);
xor U12370 (N_12370,N_12279,N_12172);
or U12371 (N_12371,N_12163,N_12183);
nor U12372 (N_12372,N_12250,N_12196);
xor U12373 (N_12373,N_12187,N_12270);
nor U12374 (N_12374,N_12217,N_12245);
nor U12375 (N_12375,N_12166,N_12272);
and U12376 (N_12376,N_12255,N_12253);
and U12377 (N_12377,N_12255,N_12250);
or U12378 (N_12378,N_12253,N_12174);
xor U12379 (N_12379,N_12297,N_12178);
nand U12380 (N_12380,N_12267,N_12266);
xnor U12381 (N_12381,N_12227,N_12158);
nand U12382 (N_12382,N_12246,N_12299);
nand U12383 (N_12383,N_12223,N_12250);
nand U12384 (N_12384,N_12278,N_12251);
nor U12385 (N_12385,N_12175,N_12151);
xor U12386 (N_12386,N_12181,N_12235);
nor U12387 (N_12387,N_12194,N_12206);
nand U12388 (N_12388,N_12259,N_12154);
xnor U12389 (N_12389,N_12241,N_12248);
nor U12390 (N_12390,N_12169,N_12246);
xnor U12391 (N_12391,N_12285,N_12272);
nor U12392 (N_12392,N_12175,N_12196);
xor U12393 (N_12393,N_12252,N_12157);
and U12394 (N_12394,N_12227,N_12211);
or U12395 (N_12395,N_12192,N_12153);
and U12396 (N_12396,N_12199,N_12280);
nand U12397 (N_12397,N_12211,N_12255);
xor U12398 (N_12398,N_12206,N_12268);
nor U12399 (N_12399,N_12169,N_12171);
and U12400 (N_12400,N_12260,N_12152);
and U12401 (N_12401,N_12234,N_12227);
and U12402 (N_12402,N_12208,N_12253);
and U12403 (N_12403,N_12210,N_12284);
xnor U12404 (N_12404,N_12281,N_12238);
nand U12405 (N_12405,N_12175,N_12236);
and U12406 (N_12406,N_12177,N_12280);
nor U12407 (N_12407,N_12208,N_12179);
nand U12408 (N_12408,N_12156,N_12216);
nand U12409 (N_12409,N_12190,N_12291);
nand U12410 (N_12410,N_12252,N_12171);
and U12411 (N_12411,N_12221,N_12195);
and U12412 (N_12412,N_12239,N_12169);
nand U12413 (N_12413,N_12246,N_12214);
xor U12414 (N_12414,N_12241,N_12212);
or U12415 (N_12415,N_12168,N_12158);
nand U12416 (N_12416,N_12213,N_12245);
nor U12417 (N_12417,N_12207,N_12272);
nand U12418 (N_12418,N_12188,N_12295);
or U12419 (N_12419,N_12223,N_12271);
or U12420 (N_12420,N_12270,N_12258);
and U12421 (N_12421,N_12241,N_12238);
nor U12422 (N_12422,N_12189,N_12161);
and U12423 (N_12423,N_12194,N_12280);
xor U12424 (N_12424,N_12239,N_12161);
xor U12425 (N_12425,N_12182,N_12206);
or U12426 (N_12426,N_12157,N_12281);
nor U12427 (N_12427,N_12173,N_12251);
nand U12428 (N_12428,N_12175,N_12156);
or U12429 (N_12429,N_12202,N_12288);
nand U12430 (N_12430,N_12193,N_12184);
nand U12431 (N_12431,N_12237,N_12261);
or U12432 (N_12432,N_12151,N_12161);
xnor U12433 (N_12433,N_12206,N_12228);
or U12434 (N_12434,N_12220,N_12219);
nand U12435 (N_12435,N_12261,N_12188);
nor U12436 (N_12436,N_12193,N_12183);
or U12437 (N_12437,N_12201,N_12262);
and U12438 (N_12438,N_12289,N_12191);
nor U12439 (N_12439,N_12274,N_12222);
xor U12440 (N_12440,N_12229,N_12167);
nand U12441 (N_12441,N_12152,N_12186);
and U12442 (N_12442,N_12267,N_12196);
nand U12443 (N_12443,N_12264,N_12193);
or U12444 (N_12444,N_12274,N_12246);
and U12445 (N_12445,N_12170,N_12222);
or U12446 (N_12446,N_12258,N_12273);
nand U12447 (N_12447,N_12204,N_12247);
or U12448 (N_12448,N_12165,N_12184);
nor U12449 (N_12449,N_12176,N_12159);
xor U12450 (N_12450,N_12335,N_12393);
nor U12451 (N_12451,N_12375,N_12309);
nand U12452 (N_12452,N_12370,N_12443);
xor U12453 (N_12453,N_12429,N_12385);
and U12454 (N_12454,N_12420,N_12378);
and U12455 (N_12455,N_12361,N_12308);
or U12456 (N_12456,N_12306,N_12368);
nand U12457 (N_12457,N_12386,N_12310);
and U12458 (N_12458,N_12424,N_12421);
nor U12459 (N_12459,N_12374,N_12397);
or U12460 (N_12460,N_12373,N_12305);
and U12461 (N_12461,N_12339,N_12382);
or U12462 (N_12462,N_12355,N_12433);
and U12463 (N_12463,N_12332,N_12316);
nor U12464 (N_12464,N_12442,N_12388);
or U12465 (N_12465,N_12360,N_12413);
nor U12466 (N_12466,N_12337,N_12342);
nor U12467 (N_12467,N_12311,N_12427);
and U12468 (N_12468,N_12313,N_12323);
nor U12469 (N_12469,N_12405,N_12351);
nand U12470 (N_12470,N_12380,N_12389);
xnor U12471 (N_12471,N_12399,N_12329);
nor U12472 (N_12472,N_12330,N_12438);
xor U12473 (N_12473,N_12366,N_12381);
and U12474 (N_12474,N_12327,N_12445);
or U12475 (N_12475,N_12341,N_12395);
and U12476 (N_12476,N_12348,N_12364);
and U12477 (N_12477,N_12449,N_12369);
nor U12478 (N_12478,N_12447,N_12377);
and U12479 (N_12479,N_12358,N_12396);
or U12480 (N_12480,N_12432,N_12359);
and U12481 (N_12481,N_12372,N_12376);
nand U12482 (N_12482,N_12350,N_12347);
or U12483 (N_12483,N_12357,N_12415);
nand U12484 (N_12484,N_12383,N_12328);
nand U12485 (N_12485,N_12314,N_12390);
xnor U12486 (N_12486,N_12419,N_12336);
nand U12487 (N_12487,N_12440,N_12412);
and U12488 (N_12488,N_12317,N_12325);
nand U12489 (N_12489,N_12354,N_12319);
or U12490 (N_12490,N_12448,N_12322);
nand U12491 (N_12491,N_12352,N_12431);
and U12492 (N_12492,N_12425,N_12418);
xor U12493 (N_12493,N_12371,N_12320);
or U12494 (N_12494,N_12401,N_12437);
and U12495 (N_12495,N_12379,N_12312);
or U12496 (N_12496,N_12334,N_12414);
and U12497 (N_12497,N_12315,N_12353);
nand U12498 (N_12498,N_12402,N_12356);
or U12499 (N_12499,N_12436,N_12344);
or U12500 (N_12500,N_12406,N_12423);
nor U12501 (N_12501,N_12343,N_12307);
nor U12502 (N_12502,N_12417,N_12410);
xnor U12503 (N_12503,N_12422,N_12300);
and U12504 (N_12504,N_12349,N_12400);
or U12505 (N_12505,N_12426,N_12384);
nor U12506 (N_12506,N_12408,N_12331);
nand U12507 (N_12507,N_12303,N_12416);
and U12508 (N_12508,N_12338,N_12394);
or U12509 (N_12509,N_12318,N_12346);
xnor U12510 (N_12510,N_12387,N_12345);
nor U12511 (N_12511,N_12302,N_12333);
nor U12512 (N_12512,N_12392,N_12403);
nor U12513 (N_12513,N_12446,N_12321);
or U12514 (N_12514,N_12391,N_12362);
nor U12515 (N_12515,N_12435,N_12407);
or U12516 (N_12516,N_12324,N_12444);
xor U12517 (N_12517,N_12430,N_12304);
nand U12518 (N_12518,N_12365,N_12441);
xor U12519 (N_12519,N_12411,N_12340);
nor U12520 (N_12520,N_12367,N_12434);
nand U12521 (N_12521,N_12363,N_12398);
nor U12522 (N_12522,N_12404,N_12326);
nor U12523 (N_12523,N_12409,N_12428);
or U12524 (N_12524,N_12301,N_12439);
nor U12525 (N_12525,N_12385,N_12370);
and U12526 (N_12526,N_12348,N_12361);
and U12527 (N_12527,N_12330,N_12423);
xor U12528 (N_12528,N_12425,N_12397);
nor U12529 (N_12529,N_12382,N_12369);
nor U12530 (N_12530,N_12434,N_12410);
nor U12531 (N_12531,N_12329,N_12372);
and U12532 (N_12532,N_12408,N_12355);
or U12533 (N_12533,N_12440,N_12336);
xor U12534 (N_12534,N_12309,N_12346);
or U12535 (N_12535,N_12392,N_12411);
xnor U12536 (N_12536,N_12415,N_12327);
or U12537 (N_12537,N_12390,N_12337);
nand U12538 (N_12538,N_12417,N_12345);
and U12539 (N_12539,N_12326,N_12380);
nand U12540 (N_12540,N_12389,N_12376);
and U12541 (N_12541,N_12413,N_12387);
nor U12542 (N_12542,N_12367,N_12436);
xnor U12543 (N_12543,N_12428,N_12309);
or U12544 (N_12544,N_12376,N_12362);
xnor U12545 (N_12545,N_12415,N_12429);
nand U12546 (N_12546,N_12321,N_12316);
nand U12547 (N_12547,N_12417,N_12402);
nand U12548 (N_12548,N_12347,N_12300);
and U12549 (N_12549,N_12382,N_12420);
nor U12550 (N_12550,N_12442,N_12403);
or U12551 (N_12551,N_12376,N_12430);
or U12552 (N_12552,N_12367,N_12392);
nand U12553 (N_12553,N_12442,N_12304);
xnor U12554 (N_12554,N_12429,N_12352);
nor U12555 (N_12555,N_12418,N_12316);
or U12556 (N_12556,N_12361,N_12408);
and U12557 (N_12557,N_12392,N_12326);
or U12558 (N_12558,N_12363,N_12449);
nand U12559 (N_12559,N_12346,N_12306);
nor U12560 (N_12560,N_12370,N_12346);
nor U12561 (N_12561,N_12388,N_12379);
xnor U12562 (N_12562,N_12316,N_12358);
nand U12563 (N_12563,N_12393,N_12444);
or U12564 (N_12564,N_12414,N_12358);
xnor U12565 (N_12565,N_12330,N_12364);
nor U12566 (N_12566,N_12331,N_12403);
nor U12567 (N_12567,N_12426,N_12388);
nor U12568 (N_12568,N_12344,N_12398);
nor U12569 (N_12569,N_12390,N_12341);
nor U12570 (N_12570,N_12332,N_12421);
or U12571 (N_12571,N_12343,N_12435);
nor U12572 (N_12572,N_12412,N_12435);
nor U12573 (N_12573,N_12440,N_12399);
xor U12574 (N_12574,N_12398,N_12374);
xor U12575 (N_12575,N_12394,N_12423);
and U12576 (N_12576,N_12329,N_12302);
and U12577 (N_12577,N_12389,N_12409);
nor U12578 (N_12578,N_12436,N_12323);
or U12579 (N_12579,N_12370,N_12369);
or U12580 (N_12580,N_12315,N_12303);
and U12581 (N_12581,N_12364,N_12410);
xor U12582 (N_12582,N_12315,N_12431);
and U12583 (N_12583,N_12344,N_12438);
or U12584 (N_12584,N_12354,N_12360);
nand U12585 (N_12585,N_12359,N_12329);
nand U12586 (N_12586,N_12380,N_12364);
nand U12587 (N_12587,N_12355,N_12363);
nor U12588 (N_12588,N_12343,N_12424);
and U12589 (N_12589,N_12308,N_12397);
nand U12590 (N_12590,N_12317,N_12326);
nand U12591 (N_12591,N_12338,N_12420);
nor U12592 (N_12592,N_12429,N_12316);
or U12593 (N_12593,N_12361,N_12321);
or U12594 (N_12594,N_12343,N_12351);
or U12595 (N_12595,N_12380,N_12310);
and U12596 (N_12596,N_12313,N_12314);
nor U12597 (N_12597,N_12306,N_12338);
nand U12598 (N_12598,N_12412,N_12325);
and U12599 (N_12599,N_12423,N_12410);
nor U12600 (N_12600,N_12592,N_12507);
xor U12601 (N_12601,N_12500,N_12556);
nor U12602 (N_12602,N_12583,N_12536);
nand U12603 (N_12603,N_12575,N_12516);
or U12604 (N_12604,N_12502,N_12529);
xor U12605 (N_12605,N_12549,N_12538);
or U12606 (N_12606,N_12451,N_12484);
and U12607 (N_12607,N_12537,N_12471);
and U12608 (N_12608,N_12485,N_12581);
or U12609 (N_12609,N_12579,N_12459);
and U12610 (N_12610,N_12474,N_12452);
nand U12611 (N_12611,N_12584,N_12553);
nor U12612 (N_12612,N_12510,N_12535);
or U12613 (N_12613,N_12570,N_12532);
xor U12614 (N_12614,N_12503,N_12522);
and U12615 (N_12615,N_12525,N_12505);
or U12616 (N_12616,N_12506,N_12467);
nand U12617 (N_12617,N_12460,N_12524);
and U12618 (N_12618,N_12573,N_12561);
nand U12619 (N_12619,N_12567,N_12552);
nor U12620 (N_12620,N_12545,N_12453);
and U12621 (N_12621,N_12568,N_12468);
or U12622 (N_12622,N_12476,N_12574);
nor U12623 (N_12623,N_12499,N_12475);
and U12624 (N_12624,N_12595,N_12513);
or U12625 (N_12625,N_12494,N_12498);
nor U12626 (N_12626,N_12530,N_12548);
nand U12627 (N_12627,N_12539,N_12576);
nor U12628 (N_12628,N_12477,N_12456);
or U12629 (N_12629,N_12547,N_12521);
and U12630 (N_12630,N_12489,N_12585);
or U12631 (N_12631,N_12534,N_12497);
and U12632 (N_12632,N_12572,N_12555);
nor U12633 (N_12633,N_12515,N_12491);
xor U12634 (N_12634,N_12481,N_12540);
nor U12635 (N_12635,N_12565,N_12546);
xnor U12636 (N_12636,N_12486,N_12562);
or U12637 (N_12637,N_12564,N_12560);
or U12638 (N_12638,N_12558,N_12512);
and U12639 (N_12639,N_12465,N_12598);
xnor U12640 (N_12640,N_12461,N_12533);
and U12641 (N_12641,N_12483,N_12504);
and U12642 (N_12642,N_12508,N_12587);
nand U12643 (N_12643,N_12492,N_12457);
nand U12644 (N_12644,N_12590,N_12569);
nor U12645 (N_12645,N_12593,N_12520);
xnor U12646 (N_12646,N_12469,N_12531);
and U12647 (N_12647,N_12566,N_12588);
nor U12648 (N_12648,N_12473,N_12526);
and U12649 (N_12649,N_12478,N_12518);
xnor U12650 (N_12650,N_12523,N_12458);
or U12651 (N_12651,N_12488,N_12589);
nor U12652 (N_12652,N_12550,N_12554);
nand U12653 (N_12653,N_12514,N_12487);
and U12654 (N_12654,N_12509,N_12596);
nor U12655 (N_12655,N_12557,N_12578);
nand U12656 (N_12656,N_12594,N_12597);
or U12657 (N_12657,N_12582,N_12559);
xor U12658 (N_12658,N_12563,N_12551);
nor U12659 (N_12659,N_12580,N_12501);
nor U12660 (N_12660,N_12599,N_12544);
or U12661 (N_12661,N_12542,N_12454);
or U12662 (N_12662,N_12463,N_12482);
and U12663 (N_12663,N_12450,N_12517);
nand U12664 (N_12664,N_12470,N_12586);
xnor U12665 (N_12665,N_12591,N_12462);
and U12666 (N_12666,N_12496,N_12466);
or U12667 (N_12667,N_12480,N_12464);
nor U12668 (N_12668,N_12472,N_12571);
nand U12669 (N_12669,N_12519,N_12527);
xnor U12670 (N_12670,N_12541,N_12511);
or U12671 (N_12671,N_12543,N_12455);
or U12672 (N_12672,N_12528,N_12479);
nand U12673 (N_12673,N_12495,N_12493);
nor U12674 (N_12674,N_12577,N_12490);
or U12675 (N_12675,N_12597,N_12484);
or U12676 (N_12676,N_12599,N_12591);
or U12677 (N_12677,N_12478,N_12519);
nor U12678 (N_12678,N_12583,N_12530);
nor U12679 (N_12679,N_12459,N_12496);
nor U12680 (N_12680,N_12563,N_12457);
xor U12681 (N_12681,N_12508,N_12548);
nand U12682 (N_12682,N_12479,N_12567);
xnor U12683 (N_12683,N_12586,N_12504);
or U12684 (N_12684,N_12559,N_12469);
xnor U12685 (N_12685,N_12512,N_12555);
or U12686 (N_12686,N_12460,N_12530);
nor U12687 (N_12687,N_12593,N_12472);
nand U12688 (N_12688,N_12486,N_12579);
xor U12689 (N_12689,N_12583,N_12508);
nor U12690 (N_12690,N_12511,N_12554);
or U12691 (N_12691,N_12587,N_12496);
or U12692 (N_12692,N_12501,N_12483);
and U12693 (N_12693,N_12499,N_12452);
nor U12694 (N_12694,N_12547,N_12524);
and U12695 (N_12695,N_12553,N_12550);
and U12696 (N_12696,N_12496,N_12586);
nand U12697 (N_12697,N_12526,N_12596);
nand U12698 (N_12698,N_12545,N_12500);
and U12699 (N_12699,N_12489,N_12460);
nor U12700 (N_12700,N_12462,N_12519);
nand U12701 (N_12701,N_12554,N_12549);
nor U12702 (N_12702,N_12544,N_12569);
nand U12703 (N_12703,N_12548,N_12526);
and U12704 (N_12704,N_12592,N_12567);
and U12705 (N_12705,N_12461,N_12498);
xor U12706 (N_12706,N_12496,N_12560);
nand U12707 (N_12707,N_12534,N_12599);
nand U12708 (N_12708,N_12465,N_12517);
nand U12709 (N_12709,N_12587,N_12457);
or U12710 (N_12710,N_12526,N_12481);
and U12711 (N_12711,N_12513,N_12540);
or U12712 (N_12712,N_12480,N_12484);
nor U12713 (N_12713,N_12554,N_12517);
nand U12714 (N_12714,N_12458,N_12472);
xor U12715 (N_12715,N_12472,N_12578);
xnor U12716 (N_12716,N_12488,N_12452);
nor U12717 (N_12717,N_12459,N_12479);
nand U12718 (N_12718,N_12463,N_12487);
nand U12719 (N_12719,N_12545,N_12521);
nand U12720 (N_12720,N_12538,N_12514);
and U12721 (N_12721,N_12588,N_12505);
or U12722 (N_12722,N_12528,N_12530);
nand U12723 (N_12723,N_12497,N_12556);
and U12724 (N_12724,N_12509,N_12585);
and U12725 (N_12725,N_12547,N_12479);
or U12726 (N_12726,N_12481,N_12592);
xnor U12727 (N_12727,N_12554,N_12594);
and U12728 (N_12728,N_12589,N_12468);
nand U12729 (N_12729,N_12599,N_12562);
nor U12730 (N_12730,N_12475,N_12595);
nand U12731 (N_12731,N_12528,N_12476);
or U12732 (N_12732,N_12469,N_12485);
or U12733 (N_12733,N_12496,N_12551);
nand U12734 (N_12734,N_12497,N_12558);
or U12735 (N_12735,N_12596,N_12575);
or U12736 (N_12736,N_12595,N_12541);
nand U12737 (N_12737,N_12531,N_12470);
or U12738 (N_12738,N_12562,N_12520);
nor U12739 (N_12739,N_12540,N_12583);
nor U12740 (N_12740,N_12506,N_12505);
or U12741 (N_12741,N_12563,N_12599);
nand U12742 (N_12742,N_12458,N_12505);
and U12743 (N_12743,N_12575,N_12496);
or U12744 (N_12744,N_12473,N_12517);
nand U12745 (N_12745,N_12570,N_12507);
xnor U12746 (N_12746,N_12493,N_12489);
nor U12747 (N_12747,N_12571,N_12524);
xnor U12748 (N_12748,N_12580,N_12494);
and U12749 (N_12749,N_12534,N_12516);
and U12750 (N_12750,N_12644,N_12636);
nor U12751 (N_12751,N_12683,N_12695);
nand U12752 (N_12752,N_12697,N_12702);
or U12753 (N_12753,N_12660,N_12623);
nor U12754 (N_12754,N_12731,N_12632);
or U12755 (N_12755,N_12615,N_12609);
nand U12756 (N_12756,N_12628,N_12655);
nand U12757 (N_12757,N_12704,N_12661);
nand U12758 (N_12758,N_12601,N_12613);
nor U12759 (N_12759,N_12737,N_12610);
and U12760 (N_12760,N_12739,N_12639);
nand U12761 (N_12761,N_12707,N_12672);
nand U12762 (N_12762,N_12671,N_12719);
xnor U12763 (N_12763,N_12663,N_12606);
or U12764 (N_12764,N_12641,N_12692);
or U12765 (N_12765,N_12670,N_12614);
and U12766 (N_12766,N_12747,N_12648);
and U12767 (N_12767,N_12738,N_12673);
nand U12768 (N_12768,N_12645,N_12680);
and U12769 (N_12769,N_12675,N_12710);
or U12770 (N_12770,N_12646,N_12604);
xnor U12771 (N_12771,N_12682,N_12735);
or U12772 (N_12772,N_12669,N_12619);
and U12773 (N_12773,N_12718,N_12721);
nor U12774 (N_12774,N_12643,N_12629);
and U12775 (N_12775,N_12631,N_12626);
or U12776 (N_12776,N_12600,N_12608);
nor U12777 (N_12777,N_12685,N_12625);
and U12778 (N_12778,N_12730,N_12642);
nand U12779 (N_12779,N_12627,N_12679);
nor U12780 (N_12780,N_12741,N_12651);
and U12781 (N_12781,N_12630,N_12717);
nor U12782 (N_12782,N_12701,N_12633);
nor U12783 (N_12783,N_12622,N_12720);
and U12784 (N_12784,N_12603,N_12728);
xor U12785 (N_12785,N_12624,N_12658);
xor U12786 (N_12786,N_12722,N_12681);
or U12787 (N_12787,N_12726,N_12602);
and U12788 (N_12788,N_12611,N_12668);
and U12789 (N_12789,N_12686,N_12640);
nor U12790 (N_12790,N_12654,N_12659);
or U12791 (N_12791,N_12666,N_12724);
and U12792 (N_12792,N_12713,N_12618);
and U12793 (N_12793,N_12716,N_12647);
xnor U12794 (N_12794,N_12727,N_12733);
nand U12795 (N_12795,N_12706,N_12712);
and U12796 (N_12796,N_12746,N_12688);
nand U12797 (N_12797,N_12667,N_12684);
or U12798 (N_12798,N_12725,N_12708);
or U12799 (N_12799,N_12674,N_12634);
or U12800 (N_12800,N_12677,N_12734);
xor U12801 (N_12801,N_12621,N_12664);
and U12802 (N_12802,N_12678,N_12729);
and U12803 (N_12803,N_12637,N_12711);
xor U12804 (N_12804,N_12662,N_12693);
or U12805 (N_12805,N_12605,N_12748);
nand U12806 (N_12806,N_12714,N_12744);
nand U12807 (N_12807,N_12732,N_12635);
nand U12808 (N_12808,N_12616,N_12749);
xnor U12809 (N_12809,N_12612,N_12687);
nor U12810 (N_12810,N_12607,N_12740);
xnor U12811 (N_12811,N_12689,N_12705);
nand U12812 (N_12812,N_12715,N_12653);
nand U12813 (N_12813,N_12620,N_12652);
and U12814 (N_12814,N_12723,N_12649);
and U12815 (N_12815,N_12617,N_12694);
nor U12816 (N_12816,N_12656,N_12676);
nor U12817 (N_12817,N_12696,N_12691);
and U12818 (N_12818,N_12743,N_12699);
xnor U12819 (N_12819,N_12650,N_12700);
nand U12820 (N_12820,N_12698,N_12742);
xor U12821 (N_12821,N_12657,N_12736);
xnor U12822 (N_12822,N_12745,N_12665);
and U12823 (N_12823,N_12638,N_12709);
and U12824 (N_12824,N_12690,N_12703);
nand U12825 (N_12825,N_12632,N_12604);
xnor U12826 (N_12826,N_12679,N_12738);
xnor U12827 (N_12827,N_12726,N_12680);
xnor U12828 (N_12828,N_12733,N_12615);
nand U12829 (N_12829,N_12625,N_12603);
nand U12830 (N_12830,N_12650,N_12658);
nor U12831 (N_12831,N_12611,N_12696);
or U12832 (N_12832,N_12735,N_12687);
nand U12833 (N_12833,N_12711,N_12610);
nor U12834 (N_12834,N_12708,N_12731);
nand U12835 (N_12835,N_12642,N_12700);
nor U12836 (N_12836,N_12743,N_12721);
nor U12837 (N_12837,N_12609,N_12749);
nor U12838 (N_12838,N_12678,N_12695);
nand U12839 (N_12839,N_12740,N_12624);
nor U12840 (N_12840,N_12619,N_12613);
nor U12841 (N_12841,N_12726,N_12613);
and U12842 (N_12842,N_12662,N_12738);
nand U12843 (N_12843,N_12600,N_12735);
nand U12844 (N_12844,N_12662,N_12616);
or U12845 (N_12845,N_12685,N_12659);
or U12846 (N_12846,N_12701,N_12679);
xnor U12847 (N_12847,N_12618,N_12634);
or U12848 (N_12848,N_12713,N_12601);
nor U12849 (N_12849,N_12684,N_12663);
nand U12850 (N_12850,N_12655,N_12733);
xnor U12851 (N_12851,N_12698,N_12720);
or U12852 (N_12852,N_12650,N_12731);
or U12853 (N_12853,N_12745,N_12698);
nor U12854 (N_12854,N_12655,N_12729);
and U12855 (N_12855,N_12711,N_12723);
and U12856 (N_12856,N_12663,N_12672);
nor U12857 (N_12857,N_12607,N_12647);
or U12858 (N_12858,N_12632,N_12644);
or U12859 (N_12859,N_12666,N_12693);
and U12860 (N_12860,N_12709,N_12653);
and U12861 (N_12861,N_12600,N_12665);
or U12862 (N_12862,N_12640,N_12715);
or U12863 (N_12863,N_12747,N_12632);
nand U12864 (N_12864,N_12749,N_12690);
nand U12865 (N_12865,N_12674,N_12673);
and U12866 (N_12866,N_12722,N_12742);
or U12867 (N_12867,N_12717,N_12677);
and U12868 (N_12868,N_12696,N_12649);
nand U12869 (N_12869,N_12664,N_12634);
or U12870 (N_12870,N_12682,N_12730);
or U12871 (N_12871,N_12639,N_12624);
nand U12872 (N_12872,N_12656,N_12726);
nor U12873 (N_12873,N_12611,N_12622);
and U12874 (N_12874,N_12667,N_12717);
or U12875 (N_12875,N_12706,N_12725);
or U12876 (N_12876,N_12635,N_12604);
and U12877 (N_12877,N_12746,N_12739);
or U12878 (N_12878,N_12691,N_12604);
nand U12879 (N_12879,N_12623,N_12695);
xor U12880 (N_12880,N_12649,N_12607);
or U12881 (N_12881,N_12643,N_12608);
and U12882 (N_12882,N_12649,N_12747);
or U12883 (N_12883,N_12708,N_12674);
xor U12884 (N_12884,N_12608,N_12675);
xor U12885 (N_12885,N_12710,N_12637);
nor U12886 (N_12886,N_12632,N_12739);
xnor U12887 (N_12887,N_12717,N_12748);
nand U12888 (N_12888,N_12648,N_12604);
nand U12889 (N_12889,N_12619,N_12658);
or U12890 (N_12890,N_12705,N_12713);
and U12891 (N_12891,N_12681,N_12684);
nor U12892 (N_12892,N_12736,N_12676);
nor U12893 (N_12893,N_12738,N_12731);
xnor U12894 (N_12894,N_12655,N_12621);
nor U12895 (N_12895,N_12665,N_12700);
nor U12896 (N_12896,N_12725,N_12731);
or U12897 (N_12897,N_12624,N_12640);
nand U12898 (N_12898,N_12608,N_12624);
nand U12899 (N_12899,N_12625,N_12682);
and U12900 (N_12900,N_12827,N_12802);
nor U12901 (N_12901,N_12885,N_12891);
xnor U12902 (N_12902,N_12822,N_12840);
nor U12903 (N_12903,N_12772,N_12831);
nor U12904 (N_12904,N_12829,N_12899);
nor U12905 (N_12905,N_12842,N_12780);
xor U12906 (N_12906,N_12760,N_12809);
and U12907 (N_12907,N_12757,N_12771);
nand U12908 (N_12908,N_12798,N_12858);
xnor U12909 (N_12909,N_12884,N_12810);
or U12910 (N_12910,N_12869,N_12853);
nor U12911 (N_12911,N_12875,N_12787);
or U12912 (N_12912,N_12817,N_12855);
or U12913 (N_12913,N_12860,N_12774);
xnor U12914 (N_12914,N_12775,N_12892);
nor U12915 (N_12915,N_12818,N_12838);
and U12916 (N_12916,N_12754,N_12887);
nor U12917 (N_12917,N_12868,N_12784);
nor U12918 (N_12918,N_12761,N_12764);
or U12919 (N_12919,N_12866,N_12752);
nor U12920 (N_12920,N_12795,N_12786);
nand U12921 (N_12921,N_12876,N_12864);
nand U12922 (N_12922,N_12773,N_12896);
nand U12923 (N_12923,N_12828,N_12859);
nand U12924 (N_12924,N_12769,N_12851);
and U12925 (N_12925,N_12800,N_12750);
xor U12926 (N_12926,N_12766,N_12770);
and U12927 (N_12927,N_12898,N_12843);
and U12928 (N_12928,N_12832,N_12789);
nand U12929 (N_12929,N_12834,N_12889);
xnor U12930 (N_12930,N_12872,N_12796);
nor U12931 (N_12931,N_12816,N_12762);
and U12932 (N_12932,N_12805,N_12812);
xnor U12933 (N_12933,N_12835,N_12852);
nand U12934 (N_12934,N_12777,N_12841);
and U12935 (N_12935,N_12857,N_12801);
xnor U12936 (N_12936,N_12897,N_12871);
nand U12937 (N_12937,N_12895,N_12877);
and U12938 (N_12938,N_12790,N_12826);
and U12939 (N_12939,N_12825,N_12846);
xor U12940 (N_12940,N_12821,N_12836);
or U12941 (N_12941,N_12856,N_12833);
and U12942 (N_12942,N_12782,N_12758);
nor U12943 (N_12943,N_12854,N_12890);
and U12944 (N_12944,N_12778,N_12813);
nand U12945 (N_12945,N_12865,N_12797);
nor U12946 (N_12946,N_12863,N_12848);
and U12947 (N_12947,N_12824,N_12755);
nand U12948 (N_12948,N_12845,N_12888);
or U12949 (N_12949,N_12880,N_12847);
and U12950 (N_12950,N_12783,N_12791);
nor U12951 (N_12951,N_12879,N_12788);
nor U12952 (N_12952,N_12849,N_12781);
nand U12953 (N_12953,N_12839,N_12820);
and U12954 (N_12954,N_12823,N_12804);
xnor U12955 (N_12955,N_12893,N_12808);
nor U12956 (N_12956,N_12807,N_12886);
nor U12957 (N_12957,N_12785,N_12763);
or U12958 (N_12958,N_12873,N_12882);
nand U12959 (N_12959,N_12799,N_12811);
nor U12960 (N_12960,N_12830,N_12881);
nor U12961 (N_12961,N_12874,N_12894);
and U12962 (N_12962,N_12759,N_12861);
and U12963 (N_12963,N_12768,N_12803);
xor U12964 (N_12964,N_12751,N_12779);
nand U12965 (N_12965,N_12870,N_12776);
and U12966 (N_12966,N_12814,N_12806);
nor U12967 (N_12967,N_12819,N_12815);
nand U12968 (N_12968,N_12767,N_12837);
and U12969 (N_12969,N_12850,N_12883);
and U12970 (N_12970,N_12793,N_12756);
nand U12971 (N_12971,N_12844,N_12878);
nand U12972 (N_12972,N_12753,N_12867);
and U12973 (N_12973,N_12792,N_12862);
xnor U12974 (N_12974,N_12765,N_12794);
and U12975 (N_12975,N_12887,N_12782);
nand U12976 (N_12976,N_12759,N_12883);
xnor U12977 (N_12977,N_12798,N_12765);
or U12978 (N_12978,N_12773,N_12758);
or U12979 (N_12979,N_12772,N_12862);
xnor U12980 (N_12980,N_12786,N_12776);
xnor U12981 (N_12981,N_12768,N_12756);
or U12982 (N_12982,N_12861,N_12798);
and U12983 (N_12983,N_12826,N_12873);
xnor U12984 (N_12984,N_12894,N_12765);
nand U12985 (N_12985,N_12826,N_12791);
and U12986 (N_12986,N_12845,N_12848);
or U12987 (N_12987,N_12876,N_12762);
nor U12988 (N_12988,N_12751,N_12859);
and U12989 (N_12989,N_12769,N_12875);
xor U12990 (N_12990,N_12859,N_12750);
and U12991 (N_12991,N_12809,N_12771);
xnor U12992 (N_12992,N_12754,N_12834);
and U12993 (N_12993,N_12778,N_12816);
nand U12994 (N_12994,N_12839,N_12770);
nor U12995 (N_12995,N_12871,N_12760);
xor U12996 (N_12996,N_12830,N_12810);
or U12997 (N_12997,N_12846,N_12855);
nand U12998 (N_12998,N_12808,N_12810);
or U12999 (N_12999,N_12872,N_12765);
nor U13000 (N_13000,N_12878,N_12866);
nor U13001 (N_13001,N_12854,N_12810);
nand U13002 (N_13002,N_12867,N_12806);
or U13003 (N_13003,N_12789,N_12899);
nand U13004 (N_13004,N_12869,N_12787);
nand U13005 (N_13005,N_12839,N_12871);
nor U13006 (N_13006,N_12894,N_12766);
xnor U13007 (N_13007,N_12867,N_12811);
nand U13008 (N_13008,N_12881,N_12822);
nor U13009 (N_13009,N_12888,N_12765);
or U13010 (N_13010,N_12766,N_12872);
xor U13011 (N_13011,N_12807,N_12834);
xor U13012 (N_13012,N_12773,N_12813);
nand U13013 (N_13013,N_12802,N_12890);
or U13014 (N_13014,N_12773,N_12807);
or U13015 (N_13015,N_12897,N_12788);
and U13016 (N_13016,N_12870,N_12789);
and U13017 (N_13017,N_12775,N_12885);
and U13018 (N_13018,N_12898,N_12765);
nand U13019 (N_13019,N_12843,N_12844);
nand U13020 (N_13020,N_12893,N_12776);
and U13021 (N_13021,N_12790,N_12831);
and U13022 (N_13022,N_12753,N_12874);
or U13023 (N_13023,N_12787,N_12831);
xor U13024 (N_13024,N_12888,N_12822);
nor U13025 (N_13025,N_12822,N_12838);
and U13026 (N_13026,N_12867,N_12808);
nand U13027 (N_13027,N_12853,N_12840);
or U13028 (N_13028,N_12828,N_12885);
or U13029 (N_13029,N_12821,N_12772);
nor U13030 (N_13030,N_12791,N_12891);
or U13031 (N_13031,N_12751,N_12880);
and U13032 (N_13032,N_12761,N_12867);
nor U13033 (N_13033,N_12857,N_12899);
or U13034 (N_13034,N_12765,N_12776);
nor U13035 (N_13035,N_12797,N_12817);
xor U13036 (N_13036,N_12751,N_12803);
xnor U13037 (N_13037,N_12899,N_12878);
nor U13038 (N_13038,N_12795,N_12870);
and U13039 (N_13039,N_12832,N_12884);
and U13040 (N_13040,N_12853,N_12830);
and U13041 (N_13041,N_12752,N_12880);
xnor U13042 (N_13042,N_12898,N_12883);
xnor U13043 (N_13043,N_12776,N_12857);
nor U13044 (N_13044,N_12820,N_12812);
or U13045 (N_13045,N_12797,N_12896);
or U13046 (N_13046,N_12792,N_12787);
nor U13047 (N_13047,N_12880,N_12813);
nand U13048 (N_13048,N_12872,N_12841);
or U13049 (N_13049,N_12844,N_12792);
and U13050 (N_13050,N_12911,N_12917);
xor U13051 (N_13051,N_13009,N_12940);
nand U13052 (N_13052,N_12904,N_13023);
nor U13053 (N_13053,N_13031,N_12998);
nor U13054 (N_13054,N_13007,N_12966);
and U13055 (N_13055,N_12991,N_13046);
nor U13056 (N_13056,N_12928,N_13044);
nand U13057 (N_13057,N_12914,N_12900);
nor U13058 (N_13058,N_13018,N_13030);
or U13059 (N_13059,N_13004,N_12977);
nand U13060 (N_13060,N_13002,N_13033);
xnor U13061 (N_13061,N_12994,N_12988);
nand U13062 (N_13062,N_12950,N_12957);
and U13063 (N_13063,N_12922,N_12937);
and U13064 (N_13064,N_12927,N_12954);
and U13065 (N_13065,N_12908,N_12961);
or U13066 (N_13066,N_12912,N_12931);
nor U13067 (N_13067,N_13008,N_12983);
nor U13068 (N_13068,N_12948,N_13039);
and U13069 (N_13069,N_12973,N_12984);
and U13070 (N_13070,N_12985,N_13019);
nand U13071 (N_13071,N_12997,N_12943);
nor U13072 (N_13072,N_12933,N_12924);
nand U13073 (N_13073,N_12942,N_13032);
and U13074 (N_13074,N_13035,N_12969);
nand U13075 (N_13075,N_13016,N_12982);
nand U13076 (N_13076,N_12959,N_13034);
nand U13077 (N_13077,N_13020,N_13041);
nand U13078 (N_13078,N_12923,N_12995);
nor U13079 (N_13079,N_12967,N_12999);
or U13080 (N_13080,N_12956,N_12939);
nor U13081 (N_13081,N_13024,N_12918);
nand U13082 (N_13082,N_12996,N_13011);
or U13083 (N_13083,N_12972,N_13036);
nand U13084 (N_13084,N_12906,N_13010);
xor U13085 (N_13085,N_13003,N_12941);
or U13086 (N_13086,N_12910,N_12990);
nor U13087 (N_13087,N_12935,N_12947);
or U13088 (N_13088,N_13028,N_13040);
or U13089 (N_13089,N_12993,N_12953);
or U13090 (N_13090,N_12902,N_12974);
or U13091 (N_13091,N_12913,N_13025);
or U13092 (N_13092,N_13015,N_12925);
xnor U13093 (N_13093,N_13049,N_12989);
and U13094 (N_13094,N_12926,N_13017);
or U13095 (N_13095,N_12965,N_13013);
or U13096 (N_13096,N_12968,N_12981);
xor U13097 (N_13097,N_12936,N_13006);
nand U13098 (N_13098,N_13014,N_13027);
or U13099 (N_13099,N_12901,N_13038);
nand U13100 (N_13100,N_12958,N_13012);
and U13101 (N_13101,N_13001,N_13022);
and U13102 (N_13102,N_12945,N_12915);
xnor U13103 (N_13103,N_12938,N_13000);
nand U13104 (N_13104,N_13045,N_12978);
xor U13105 (N_13105,N_12949,N_13037);
xor U13106 (N_13106,N_12960,N_12907);
xor U13107 (N_13107,N_12929,N_12987);
or U13108 (N_13108,N_12951,N_13029);
xor U13109 (N_13109,N_13026,N_12920);
nor U13110 (N_13110,N_12962,N_12976);
nand U13111 (N_13111,N_12916,N_12975);
nor U13112 (N_13112,N_12971,N_12946);
and U13113 (N_13113,N_13043,N_12919);
nand U13114 (N_13114,N_12903,N_12964);
xor U13115 (N_13115,N_12921,N_12905);
or U13116 (N_13116,N_12952,N_12979);
and U13117 (N_13117,N_12934,N_13021);
nand U13118 (N_13118,N_12992,N_13005);
and U13119 (N_13119,N_12980,N_12970);
xor U13120 (N_13120,N_13042,N_12932);
or U13121 (N_13121,N_12909,N_12930);
nand U13122 (N_13122,N_12955,N_12963);
nand U13123 (N_13123,N_12986,N_12944);
nor U13124 (N_13124,N_13048,N_13047);
nor U13125 (N_13125,N_12979,N_12977);
xnor U13126 (N_13126,N_13018,N_12987);
and U13127 (N_13127,N_13048,N_12974);
nand U13128 (N_13128,N_12938,N_13041);
xor U13129 (N_13129,N_13023,N_12959);
nor U13130 (N_13130,N_13044,N_13034);
nand U13131 (N_13131,N_12988,N_13021);
xnor U13132 (N_13132,N_12966,N_13026);
xor U13133 (N_13133,N_13030,N_13009);
nand U13134 (N_13134,N_12986,N_13034);
nor U13135 (N_13135,N_13043,N_12974);
nand U13136 (N_13136,N_13048,N_12937);
xnor U13137 (N_13137,N_13005,N_12918);
and U13138 (N_13138,N_13019,N_12947);
nand U13139 (N_13139,N_12957,N_13036);
nor U13140 (N_13140,N_12996,N_12968);
and U13141 (N_13141,N_12973,N_13003);
nand U13142 (N_13142,N_13014,N_13045);
nor U13143 (N_13143,N_12922,N_13011);
nor U13144 (N_13144,N_12935,N_12908);
and U13145 (N_13145,N_13015,N_12958);
and U13146 (N_13146,N_12928,N_12929);
xnor U13147 (N_13147,N_13012,N_12935);
xnor U13148 (N_13148,N_13011,N_12920);
nand U13149 (N_13149,N_12978,N_13006);
xnor U13150 (N_13150,N_12960,N_12933);
nor U13151 (N_13151,N_12917,N_12945);
xnor U13152 (N_13152,N_13005,N_12964);
nor U13153 (N_13153,N_12975,N_13045);
nor U13154 (N_13154,N_12946,N_12999);
or U13155 (N_13155,N_12970,N_12929);
nor U13156 (N_13156,N_12968,N_13006);
and U13157 (N_13157,N_12911,N_12902);
xor U13158 (N_13158,N_13039,N_12928);
xnor U13159 (N_13159,N_12945,N_13047);
and U13160 (N_13160,N_12995,N_13012);
xnor U13161 (N_13161,N_13025,N_13037);
nand U13162 (N_13162,N_13016,N_12934);
nor U13163 (N_13163,N_12901,N_13017);
nand U13164 (N_13164,N_13043,N_13039);
and U13165 (N_13165,N_12961,N_12959);
xor U13166 (N_13166,N_12954,N_13010);
nor U13167 (N_13167,N_13021,N_12921);
nand U13168 (N_13168,N_12990,N_12930);
or U13169 (N_13169,N_12912,N_13031);
and U13170 (N_13170,N_13001,N_12917);
nand U13171 (N_13171,N_12956,N_13018);
nor U13172 (N_13172,N_13004,N_12972);
and U13173 (N_13173,N_13020,N_13028);
nor U13174 (N_13174,N_12929,N_12908);
or U13175 (N_13175,N_12935,N_12927);
or U13176 (N_13176,N_13002,N_13038);
nand U13177 (N_13177,N_13007,N_12989);
or U13178 (N_13178,N_13014,N_12944);
xnor U13179 (N_13179,N_13043,N_12942);
xor U13180 (N_13180,N_13030,N_12907);
xor U13181 (N_13181,N_13044,N_13015);
or U13182 (N_13182,N_12969,N_13036);
or U13183 (N_13183,N_12927,N_12974);
nor U13184 (N_13184,N_12975,N_12932);
xnor U13185 (N_13185,N_12951,N_12924);
and U13186 (N_13186,N_13031,N_12999);
nand U13187 (N_13187,N_12900,N_13044);
and U13188 (N_13188,N_12950,N_13000);
nor U13189 (N_13189,N_13007,N_12911);
xnor U13190 (N_13190,N_12937,N_12998);
and U13191 (N_13191,N_13031,N_12938);
xnor U13192 (N_13192,N_12993,N_12986);
nor U13193 (N_13193,N_12901,N_13045);
xnor U13194 (N_13194,N_13007,N_13006);
and U13195 (N_13195,N_13020,N_12988);
or U13196 (N_13196,N_13020,N_12991);
nand U13197 (N_13197,N_13023,N_13022);
and U13198 (N_13198,N_12947,N_12929);
nand U13199 (N_13199,N_12983,N_12939);
nand U13200 (N_13200,N_13119,N_13155);
or U13201 (N_13201,N_13182,N_13104);
nand U13202 (N_13202,N_13197,N_13164);
and U13203 (N_13203,N_13179,N_13100);
nand U13204 (N_13204,N_13144,N_13125);
nor U13205 (N_13205,N_13159,N_13143);
xnor U13206 (N_13206,N_13083,N_13065);
xor U13207 (N_13207,N_13085,N_13156);
or U13208 (N_13208,N_13102,N_13122);
nand U13209 (N_13209,N_13079,N_13055);
or U13210 (N_13210,N_13152,N_13103);
xnor U13211 (N_13211,N_13114,N_13071);
xor U13212 (N_13212,N_13165,N_13059);
and U13213 (N_13213,N_13166,N_13093);
nor U13214 (N_13214,N_13172,N_13196);
or U13215 (N_13215,N_13089,N_13177);
or U13216 (N_13216,N_13141,N_13163);
or U13217 (N_13217,N_13145,N_13066);
and U13218 (N_13218,N_13183,N_13082);
nand U13219 (N_13219,N_13139,N_13174);
nand U13220 (N_13220,N_13176,N_13084);
or U13221 (N_13221,N_13120,N_13094);
and U13222 (N_13222,N_13076,N_13069);
xor U13223 (N_13223,N_13160,N_13106);
xnor U13224 (N_13224,N_13115,N_13109);
and U13225 (N_13225,N_13050,N_13108);
nand U13226 (N_13226,N_13064,N_13067);
nand U13227 (N_13227,N_13126,N_13062);
xor U13228 (N_13228,N_13189,N_13137);
or U13229 (N_13229,N_13147,N_13099);
and U13230 (N_13230,N_13053,N_13056);
nand U13231 (N_13231,N_13192,N_13113);
nor U13232 (N_13232,N_13191,N_13068);
and U13233 (N_13233,N_13138,N_13148);
nand U13234 (N_13234,N_13157,N_13158);
xnor U13235 (N_13235,N_13097,N_13180);
xnor U13236 (N_13236,N_13060,N_13121);
nand U13237 (N_13237,N_13074,N_13150);
nor U13238 (N_13238,N_13190,N_13167);
and U13239 (N_13239,N_13111,N_13134);
xor U13240 (N_13240,N_13175,N_13151);
or U13241 (N_13241,N_13095,N_13135);
nor U13242 (N_13242,N_13184,N_13128);
xor U13243 (N_13243,N_13173,N_13075);
nor U13244 (N_13244,N_13107,N_13105);
or U13245 (N_13245,N_13153,N_13149);
or U13246 (N_13246,N_13091,N_13098);
nor U13247 (N_13247,N_13178,N_13187);
xnor U13248 (N_13248,N_13199,N_13136);
xor U13249 (N_13249,N_13129,N_13168);
nor U13250 (N_13250,N_13127,N_13181);
and U13251 (N_13251,N_13193,N_13169);
nand U13252 (N_13252,N_13054,N_13118);
nor U13253 (N_13253,N_13133,N_13101);
nor U13254 (N_13254,N_13078,N_13194);
nand U13255 (N_13255,N_13112,N_13146);
nand U13256 (N_13256,N_13057,N_13086);
and U13257 (N_13257,N_13092,N_13051);
nand U13258 (N_13258,N_13142,N_13188);
nor U13259 (N_13259,N_13070,N_13132);
nor U13260 (N_13260,N_13154,N_13140);
or U13261 (N_13261,N_13052,N_13170);
nand U13262 (N_13262,N_13186,N_13185);
nor U13263 (N_13263,N_13198,N_13162);
or U13264 (N_13264,N_13123,N_13063);
xnor U13265 (N_13265,N_13124,N_13058);
or U13266 (N_13266,N_13130,N_13061);
nand U13267 (N_13267,N_13195,N_13117);
or U13268 (N_13268,N_13090,N_13072);
xnor U13269 (N_13269,N_13077,N_13161);
and U13270 (N_13270,N_13116,N_13073);
and U13271 (N_13271,N_13088,N_13096);
nand U13272 (N_13272,N_13080,N_13131);
nand U13273 (N_13273,N_13110,N_13171);
and U13274 (N_13274,N_13081,N_13087);
and U13275 (N_13275,N_13195,N_13129);
nand U13276 (N_13276,N_13078,N_13074);
or U13277 (N_13277,N_13061,N_13142);
or U13278 (N_13278,N_13161,N_13171);
and U13279 (N_13279,N_13120,N_13093);
or U13280 (N_13280,N_13127,N_13128);
and U13281 (N_13281,N_13116,N_13092);
or U13282 (N_13282,N_13184,N_13129);
nor U13283 (N_13283,N_13156,N_13179);
xnor U13284 (N_13284,N_13109,N_13128);
nor U13285 (N_13285,N_13063,N_13080);
nor U13286 (N_13286,N_13056,N_13149);
or U13287 (N_13287,N_13090,N_13160);
nand U13288 (N_13288,N_13070,N_13100);
xnor U13289 (N_13289,N_13065,N_13078);
and U13290 (N_13290,N_13072,N_13115);
nor U13291 (N_13291,N_13156,N_13181);
nand U13292 (N_13292,N_13088,N_13111);
nor U13293 (N_13293,N_13170,N_13078);
and U13294 (N_13294,N_13189,N_13065);
xnor U13295 (N_13295,N_13074,N_13090);
nor U13296 (N_13296,N_13110,N_13128);
and U13297 (N_13297,N_13197,N_13050);
and U13298 (N_13298,N_13127,N_13053);
xor U13299 (N_13299,N_13075,N_13140);
nor U13300 (N_13300,N_13162,N_13052);
xnor U13301 (N_13301,N_13161,N_13115);
nor U13302 (N_13302,N_13117,N_13127);
nor U13303 (N_13303,N_13094,N_13089);
nand U13304 (N_13304,N_13140,N_13119);
or U13305 (N_13305,N_13095,N_13155);
or U13306 (N_13306,N_13188,N_13194);
nand U13307 (N_13307,N_13180,N_13116);
and U13308 (N_13308,N_13081,N_13178);
and U13309 (N_13309,N_13057,N_13050);
nand U13310 (N_13310,N_13106,N_13190);
and U13311 (N_13311,N_13142,N_13186);
xor U13312 (N_13312,N_13124,N_13194);
nand U13313 (N_13313,N_13064,N_13196);
and U13314 (N_13314,N_13162,N_13108);
nand U13315 (N_13315,N_13130,N_13195);
or U13316 (N_13316,N_13090,N_13123);
nor U13317 (N_13317,N_13089,N_13134);
or U13318 (N_13318,N_13061,N_13196);
xnor U13319 (N_13319,N_13170,N_13154);
or U13320 (N_13320,N_13126,N_13083);
or U13321 (N_13321,N_13143,N_13130);
and U13322 (N_13322,N_13126,N_13169);
nand U13323 (N_13323,N_13090,N_13082);
or U13324 (N_13324,N_13053,N_13112);
or U13325 (N_13325,N_13083,N_13087);
or U13326 (N_13326,N_13196,N_13128);
and U13327 (N_13327,N_13196,N_13050);
nand U13328 (N_13328,N_13133,N_13054);
and U13329 (N_13329,N_13179,N_13125);
or U13330 (N_13330,N_13080,N_13096);
and U13331 (N_13331,N_13120,N_13175);
xnor U13332 (N_13332,N_13078,N_13063);
nand U13333 (N_13333,N_13060,N_13066);
nor U13334 (N_13334,N_13093,N_13073);
nand U13335 (N_13335,N_13137,N_13156);
or U13336 (N_13336,N_13095,N_13171);
nor U13337 (N_13337,N_13061,N_13143);
nand U13338 (N_13338,N_13095,N_13190);
xnor U13339 (N_13339,N_13164,N_13194);
nand U13340 (N_13340,N_13063,N_13116);
or U13341 (N_13341,N_13109,N_13162);
or U13342 (N_13342,N_13119,N_13197);
nand U13343 (N_13343,N_13199,N_13162);
or U13344 (N_13344,N_13073,N_13069);
xor U13345 (N_13345,N_13080,N_13182);
nor U13346 (N_13346,N_13060,N_13168);
and U13347 (N_13347,N_13196,N_13156);
or U13348 (N_13348,N_13080,N_13174);
nor U13349 (N_13349,N_13076,N_13145);
nor U13350 (N_13350,N_13236,N_13276);
xnor U13351 (N_13351,N_13219,N_13221);
xnor U13352 (N_13352,N_13242,N_13312);
or U13353 (N_13353,N_13227,N_13345);
and U13354 (N_13354,N_13208,N_13207);
xor U13355 (N_13355,N_13230,N_13344);
nand U13356 (N_13356,N_13343,N_13209);
nand U13357 (N_13357,N_13288,N_13328);
xor U13358 (N_13358,N_13311,N_13298);
or U13359 (N_13359,N_13239,N_13278);
or U13360 (N_13360,N_13223,N_13292);
xnor U13361 (N_13361,N_13338,N_13244);
nand U13362 (N_13362,N_13327,N_13290);
nor U13363 (N_13363,N_13340,N_13225);
xor U13364 (N_13364,N_13264,N_13333);
xnor U13365 (N_13365,N_13205,N_13271);
and U13366 (N_13366,N_13331,N_13339);
nor U13367 (N_13367,N_13326,N_13201);
xnor U13368 (N_13368,N_13342,N_13218);
nor U13369 (N_13369,N_13269,N_13337);
nand U13370 (N_13370,N_13228,N_13211);
and U13371 (N_13371,N_13246,N_13284);
nor U13372 (N_13372,N_13296,N_13294);
nand U13373 (N_13373,N_13232,N_13286);
nand U13374 (N_13374,N_13258,N_13229);
nand U13375 (N_13375,N_13255,N_13277);
and U13376 (N_13376,N_13249,N_13226);
or U13377 (N_13377,N_13301,N_13237);
nor U13378 (N_13378,N_13293,N_13304);
and U13379 (N_13379,N_13248,N_13259);
xnor U13380 (N_13380,N_13322,N_13287);
nand U13381 (N_13381,N_13336,N_13233);
and U13382 (N_13382,N_13212,N_13210);
and U13383 (N_13383,N_13213,N_13349);
nor U13384 (N_13384,N_13325,N_13260);
or U13385 (N_13385,N_13216,N_13235);
and U13386 (N_13386,N_13268,N_13203);
and U13387 (N_13387,N_13320,N_13265);
and U13388 (N_13388,N_13285,N_13251);
nand U13389 (N_13389,N_13314,N_13305);
nor U13390 (N_13390,N_13217,N_13306);
nor U13391 (N_13391,N_13250,N_13319);
xnor U13392 (N_13392,N_13302,N_13220);
xnor U13393 (N_13393,N_13289,N_13222);
nor U13394 (N_13394,N_13261,N_13300);
xor U13395 (N_13395,N_13309,N_13241);
nand U13396 (N_13396,N_13341,N_13332);
xnor U13397 (N_13397,N_13346,N_13283);
nand U13398 (N_13398,N_13275,N_13282);
nor U13399 (N_13399,N_13281,N_13224);
nand U13400 (N_13400,N_13279,N_13295);
nand U13401 (N_13401,N_13215,N_13323);
or U13402 (N_13402,N_13231,N_13253);
and U13403 (N_13403,N_13262,N_13247);
or U13404 (N_13404,N_13252,N_13214);
and U13405 (N_13405,N_13243,N_13335);
or U13406 (N_13406,N_13348,N_13202);
nand U13407 (N_13407,N_13204,N_13313);
or U13408 (N_13408,N_13240,N_13330);
or U13409 (N_13409,N_13317,N_13273);
xnor U13410 (N_13410,N_13324,N_13238);
nor U13411 (N_13411,N_13267,N_13234);
nor U13412 (N_13412,N_13206,N_13299);
or U13413 (N_13413,N_13257,N_13291);
xor U13414 (N_13414,N_13297,N_13274);
xnor U13415 (N_13415,N_13318,N_13347);
and U13416 (N_13416,N_13200,N_13254);
or U13417 (N_13417,N_13303,N_13321);
nor U13418 (N_13418,N_13307,N_13245);
or U13419 (N_13419,N_13270,N_13272);
xnor U13420 (N_13420,N_13334,N_13263);
nand U13421 (N_13421,N_13308,N_13256);
or U13422 (N_13422,N_13316,N_13310);
or U13423 (N_13423,N_13329,N_13280);
and U13424 (N_13424,N_13266,N_13315);
and U13425 (N_13425,N_13320,N_13250);
or U13426 (N_13426,N_13344,N_13342);
nand U13427 (N_13427,N_13251,N_13269);
and U13428 (N_13428,N_13203,N_13218);
and U13429 (N_13429,N_13304,N_13331);
xor U13430 (N_13430,N_13224,N_13339);
nor U13431 (N_13431,N_13248,N_13255);
xnor U13432 (N_13432,N_13270,N_13203);
or U13433 (N_13433,N_13292,N_13216);
and U13434 (N_13434,N_13239,N_13267);
or U13435 (N_13435,N_13202,N_13235);
xor U13436 (N_13436,N_13344,N_13313);
nor U13437 (N_13437,N_13283,N_13281);
xnor U13438 (N_13438,N_13273,N_13278);
xnor U13439 (N_13439,N_13282,N_13203);
nor U13440 (N_13440,N_13231,N_13207);
or U13441 (N_13441,N_13267,N_13252);
and U13442 (N_13442,N_13343,N_13243);
nand U13443 (N_13443,N_13262,N_13269);
nand U13444 (N_13444,N_13219,N_13336);
xor U13445 (N_13445,N_13285,N_13275);
nand U13446 (N_13446,N_13219,N_13321);
nor U13447 (N_13447,N_13296,N_13235);
and U13448 (N_13448,N_13223,N_13210);
and U13449 (N_13449,N_13330,N_13262);
or U13450 (N_13450,N_13321,N_13324);
nand U13451 (N_13451,N_13329,N_13201);
nor U13452 (N_13452,N_13221,N_13271);
nor U13453 (N_13453,N_13253,N_13294);
or U13454 (N_13454,N_13326,N_13247);
and U13455 (N_13455,N_13219,N_13247);
xnor U13456 (N_13456,N_13328,N_13347);
nor U13457 (N_13457,N_13258,N_13338);
and U13458 (N_13458,N_13201,N_13248);
nand U13459 (N_13459,N_13349,N_13277);
nor U13460 (N_13460,N_13208,N_13320);
nand U13461 (N_13461,N_13267,N_13329);
and U13462 (N_13462,N_13258,N_13247);
xor U13463 (N_13463,N_13264,N_13298);
nor U13464 (N_13464,N_13248,N_13342);
and U13465 (N_13465,N_13269,N_13339);
or U13466 (N_13466,N_13223,N_13332);
or U13467 (N_13467,N_13221,N_13304);
and U13468 (N_13468,N_13330,N_13322);
nor U13469 (N_13469,N_13322,N_13239);
or U13470 (N_13470,N_13240,N_13333);
or U13471 (N_13471,N_13316,N_13341);
xor U13472 (N_13472,N_13201,N_13233);
nor U13473 (N_13473,N_13281,N_13341);
and U13474 (N_13474,N_13344,N_13238);
or U13475 (N_13475,N_13329,N_13294);
nand U13476 (N_13476,N_13257,N_13274);
and U13477 (N_13477,N_13216,N_13263);
nor U13478 (N_13478,N_13203,N_13272);
nor U13479 (N_13479,N_13239,N_13311);
nor U13480 (N_13480,N_13231,N_13255);
nand U13481 (N_13481,N_13211,N_13305);
nor U13482 (N_13482,N_13306,N_13340);
nor U13483 (N_13483,N_13225,N_13268);
xnor U13484 (N_13484,N_13310,N_13216);
xnor U13485 (N_13485,N_13207,N_13219);
nand U13486 (N_13486,N_13336,N_13314);
xor U13487 (N_13487,N_13293,N_13344);
or U13488 (N_13488,N_13331,N_13209);
xnor U13489 (N_13489,N_13294,N_13304);
nand U13490 (N_13490,N_13283,N_13238);
and U13491 (N_13491,N_13313,N_13226);
or U13492 (N_13492,N_13235,N_13308);
and U13493 (N_13493,N_13318,N_13320);
xnor U13494 (N_13494,N_13238,N_13293);
nor U13495 (N_13495,N_13200,N_13220);
and U13496 (N_13496,N_13344,N_13272);
xor U13497 (N_13497,N_13295,N_13269);
and U13498 (N_13498,N_13301,N_13324);
xnor U13499 (N_13499,N_13235,N_13272);
nor U13500 (N_13500,N_13415,N_13484);
or U13501 (N_13501,N_13352,N_13401);
or U13502 (N_13502,N_13398,N_13385);
nor U13503 (N_13503,N_13481,N_13428);
xnor U13504 (N_13504,N_13394,N_13351);
xor U13505 (N_13505,N_13480,N_13453);
xor U13506 (N_13506,N_13413,N_13466);
xor U13507 (N_13507,N_13362,N_13488);
and U13508 (N_13508,N_13442,N_13491);
or U13509 (N_13509,N_13465,N_13354);
or U13510 (N_13510,N_13443,N_13367);
nand U13511 (N_13511,N_13411,N_13475);
nand U13512 (N_13512,N_13364,N_13440);
xnor U13513 (N_13513,N_13422,N_13380);
or U13514 (N_13514,N_13355,N_13395);
and U13515 (N_13515,N_13496,N_13468);
nand U13516 (N_13516,N_13390,N_13433);
xnor U13517 (N_13517,N_13471,N_13366);
or U13518 (N_13518,N_13473,N_13486);
and U13519 (N_13519,N_13462,N_13497);
nor U13520 (N_13520,N_13448,N_13437);
nor U13521 (N_13521,N_13379,N_13425);
or U13522 (N_13522,N_13392,N_13464);
xnor U13523 (N_13523,N_13400,N_13461);
nor U13524 (N_13524,N_13386,N_13454);
and U13525 (N_13525,N_13419,N_13412);
nand U13526 (N_13526,N_13350,N_13388);
xnor U13527 (N_13527,N_13463,N_13397);
and U13528 (N_13528,N_13431,N_13424);
xor U13529 (N_13529,N_13459,N_13441);
or U13530 (N_13530,N_13490,N_13410);
xor U13531 (N_13531,N_13384,N_13447);
nand U13532 (N_13532,N_13375,N_13353);
or U13533 (N_13533,N_13477,N_13391);
nand U13534 (N_13534,N_13479,N_13495);
nand U13535 (N_13535,N_13474,N_13470);
nor U13536 (N_13536,N_13493,N_13365);
nand U13537 (N_13537,N_13378,N_13377);
nand U13538 (N_13538,N_13370,N_13357);
or U13539 (N_13539,N_13478,N_13404);
nand U13540 (N_13540,N_13387,N_13467);
nor U13541 (N_13541,N_13405,N_13450);
xor U13542 (N_13542,N_13492,N_13445);
nand U13543 (N_13543,N_13482,N_13356);
or U13544 (N_13544,N_13374,N_13476);
nand U13545 (N_13545,N_13358,N_13403);
nor U13546 (N_13546,N_13455,N_13487);
xnor U13547 (N_13547,N_13427,N_13438);
or U13548 (N_13548,N_13485,N_13363);
or U13549 (N_13549,N_13420,N_13359);
or U13550 (N_13550,N_13499,N_13489);
nor U13551 (N_13551,N_13389,N_13434);
or U13552 (N_13552,N_13429,N_13360);
or U13553 (N_13553,N_13452,N_13451);
xnor U13554 (N_13554,N_13406,N_13369);
or U13555 (N_13555,N_13396,N_13458);
and U13556 (N_13556,N_13483,N_13423);
or U13557 (N_13557,N_13399,N_13457);
xnor U13558 (N_13558,N_13498,N_13494);
and U13559 (N_13559,N_13376,N_13430);
nor U13560 (N_13560,N_13373,N_13381);
or U13561 (N_13561,N_13460,N_13417);
nand U13562 (N_13562,N_13449,N_13409);
and U13563 (N_13563,N_13426,N_13416);
and U13564 (N_13564,N_13469,N_13407);
xnor U13565 (N_13565,N_13439,N_13432);
xnor U13566 (N_13566,N_13383,N_13436);
nand U13567 (N_13567,N_13456,N_13361);
xor U13568 (N_13568,N_13368,N_13444);
and U13569 (N_13569,N_13414,N_13472);
nor U13570 (N_13570,N_13393,N_13408);
xor U13571 (N_13571,N_13382,N_13435);
or U13572 (N_13572,N_13371,N_13418);
or U13573 (N_13573,N_13421,N_13446);
or U13574 (N_13574,N_13372,N_13402);
and U13575 (N_13575,N_13442,N_13413);
nand U13576 (N_13576,N_13379,N_13494);
nand U13577 (N_13577,N_13438,N_13379);
and U13578 (N_13578,N_13472,N_13399);
and U13579 (N_13579,N_13412,N_13497);
nand U13580 (N_13580,N_13443,N_13406);
or U13581 (N_13581,N_13396,N_13493);
xnor U13582 (N_13582,N_13433,N_13441);
xor U13583 (N_13583,N_13353,N_13405);
nor U13584 (N_13584,N_13409,N_13420);
and U13585 (N_13585,N_13355,N_13358);
or U13586 (N_13586,N_13465,N_13428);
xnor U13587 (N_13587,N_13499,N_13451);
nand U13588 (N_13588,N_13494,N_13466);
and U13589 (N_13589,N_13359,N_13366);
xor U13590 (N_13590,N_13355,N_13440);
or U13591 (N_13591,N_13436,N_13449);
and U13592 (N_13592,N_13461,N_13447);
xor U13593 (N_13593,N_13393,N_13392);
xnor U13594 (N_13594,N_13495,N_13446);
nand U13595 (N_13595,N_13402,N_13352);
nor U13596 (N_13596,N_13401,N_13415);
nand U13597 (N_13597,N_13432,N_13351);
or U13598 (N_13598,N_13361,N_13350);
and U13599 (N_13599,N_13367,N_13495);
xor U13600 (N_13600,N_13457,N_13382);
nand U13601 (N_13601,N_13374,N_13362);
or U13602 (N_13602,N_13381,N_13379);
and U13603 (N_13603,N_13441,N_13458);
nand U13604 (N_13604,N_13364,N_13498);
and U13605 (N_13605,N_13383,N_13455);
or U13606 (N_13606,N_13469,N_13408);
and U13607 (N_13607,N_13468,N_13480);
nand U13608 (N_13608,N_13498,N_13367);
nand U13609 (N_13609,N_13459,N_13364);
and U13610 (N_13610,N_13494,N_13419);
nor U13611 (N_13611,N_13356,N_13490);
and U13612 (N_13612,N_13404,N_13482);
nand U13613 (N_13613,N_13387,N_13405);
xnor U13614 (N_13614,N_13468,N_13362);
xor U13615 (N_13615,N_13462,N_13461);
xor U13616 (N_13616,N_13367,N_13442);
and U13617 (N_13617,N_13393,N_13485);
or U13618 (N_13618,N_13361,N_13415);
or U13619 (N_13619,N_13466,N_13432);
and U13620 (N_13620,N_13464,N_13352);
and U13621 (N_13621,N_13383,N_13386);
nor U13622 (N_13622,N_13364,N_13411);
nor U13623 (N_13623,N_13431,N_13487);
xor U13624 (N_13624,N_13403,N_13460);
xnor U13625 (N_13625,N_13356,N_13496);
and U13626 (N_13626,N_13428,N_13377);
nand U13627 (N_13627,N_13394,N_13395);
or U13628 (N_13628,N_13473,N_13351);
or U13629 (N_13629,N_13450,N_13409);
nand U13630 (N_13630,N_13418,N_13411);
or U13631 (N_13631,N_13487,N_13436);
or U13632 (N_13632,N_13421,N_13387);
and U13633 (N_13633,N_13393,N_13468);
or U13634 (N_13634,N_13382,N_13473);
nand U13635 (N_13635,N_13395,N_13393);
xnor U13636 (N_13636,N_13377,N_13394);
nand U13637 (N_13637,N_13497,N_13360);
nand U13638 (N_13638,N_13472,N_13371);
and U13639 (N_13639,N_13377,N_13361);
or U13640 (N_13640,N_13477,N_13433);
and U13641 (N_13641,N_13352,N_13411);
and U13642 (N_13642,N_13493,N_13377);
or U13643 (N_13643,N_13490,N_13444);
nand U13644 (N_13644,N_13430,N_13384);
nor U13645 (N_13645,N_13372,N_13350);
nor U13646 (N_13646,N_13377,N_13436);
xnor U13647 (N_13647,N_13490,N_13441);
xnor U13648 (N_13648,N_13478,N_13496);
xor U13649 (N_13649,N_13351,N_13497);
nand U13650 (N_13650,N_13561,N_13538);
nor U13651 (N_13651,N_13531,N_13532);
and U13652 (N_13652,N_13593,N_13648);
nand U13653 (N_13653,N_13615,N_13548);
nor U13654 (N_13654,N_13586,N_13631);
xnor U13655 (N_13655,N_13595,N_13540);
or U13656 (N_13656,N_13638,N_13523);
or U13657 (N_13657,N_13501,N_13625);
nand U13658 (N_13658,N_13572,N_13633);
xnor U13659 (N_13659,N_13524,N_13643);
or U13660 (N_13660,N_13577,N_13554);
and U13661 (N_13661,N_13601,N_13629);
or U13662 (N_13662,N_13507,N_13530);
or U13663 (N_13663,N_13567,N_13649);
and U13664 (N_13664,N_13611,N_13632);
nand U13665 (N_13665,N_13591,N_13520);
and U13666 (N_13666,N_13587,N_13571);
or U13667 (N_13667,N_13590,N_13529);
or U13668 (N_13668,N_13550,N_13525);
nand U13669 (N_13669,N_13579,N_13605);
nor U13670 (N_13670,N_13535,N_13636);
nor U13671 (N_13671,N_13627,N_13618);
nand U13672 (N_13672,N_13619,N_13594);
or U13673 (N_13673,N_13521,N_13607);
nor U13674 (N_13674,N_13613,N_13564);
and U13675 (N_13675,N_13565,N_13589);
or U13676 (N_13676,N_13500,N_13526);
xnor U13677 (N_13677,N_13515,N_13573);
xnor U13678 (N_13678,N_13624,N_13517);
nand U13679 (N_13679,N_13646,N_13614);
or U13680 (N_13680,N_13562,N_13582);
nor U13681 (N_13681,N_13533,N_13616);
xor U13682 (N_13682,N_13552,N_13558);
nor U13683 (N_13683,N_13518,N_13612);
nor U13684 (N_13684,N_13522,N_13592);
xnor U13685 (N_13685,N_13574,N_13546);
and U13686 (N_13686,N_13505,N_13570);
or U13687 (N_13687,N_13557,N_13583);
nor U13688 (N_13688,N_13639,N_13637);
xor U13689 (N_13689,N_13560,N_13568);
xnor U13690 (N_13690,N_13634,N_13588);
xor U13691 (N_13691,N_13514,N_13512);
xnor U13692 (N_13692,N_13620,N_13534);
or U13693 (N_13693,N_13596,N_13536);
or U13694 (N_13694,N_13584,N_13599);
xnor U13695 (N_13695,N_13537,N_13603);
nor U13696 (N_13696,N_13539,N_13553);
nor U13697 (N_13697,N_13610,N_13623);
nor U13698 (N_13698,N_13510,N_13608);
xnor U13699 (N_13699,N_13641,N_13544);
nand U13700 (N_13700,N_13511,N_13602);
or U13701 (N_13701,N_13597,N_13549);
or U13702 (N_13702,N_13555,N_13516);
or U13703 (N_13703,N_13503,N_13622);
and U13704 (N_13704,N_13585,N_13630);
or U13705 (N_13705,N_13545,N_13547);
and U13706 (N_13706,N_13628,N_13566);
nor U13707 (N_13707,N_13645,N_13600);
xor U13708 (N_13708,N_13642,N_13569);
xnor U13709 (N_13709,N_13563,N_13519);
and U13710 (N_13710,N_13508,N_13644);
and U13711 (N_13711,N_13598,N_13647);
nor U13712 (N_13712,N_13621,N_13559);
and U13713 (N_13713,N_13606,N_13556);
or U13714 (N_13714,N_13541,N_13626);
xor U13715 (N_13715,N_13513,N_13617);
nand U13716 (N_13716,N_13502,N_13543);
or U13717 (N_13717,N_13581,N_13575);
or U13718 (N_13718,N_13551,N_13527);
xnor U13719 (N_13719,N_13528,N_13542);
or U13720 (N_13720,N_13509,N_13578);
nand U13721 (N_13721,N_13576,N_13506);
and U13722 (N_13722,N_13635,N_13580);
nor U13723 (N_13723,N_13609,N_13640);
xnor U13724 (N_13724,N_13504,N_13604);
or U13725 (N_13725,N_13548,N_13515);
and U13726 (N_13726,N_13537,N_13583);
or U13727 (N_13727,N_13508,N_13615);
nor U13728 (N_13728,N_13502,N_13603);
and U13729 (N_13729,N_13619,N_13649);
xor U13730 (N_13730,N_13583,N_13612);
nand U13731 (N_13731,N_13563,N_13590);
xor U13732 (N_13732,N_13606,N_13524);
nor U13733 (N_13733,N_13633,N_13649);
and U13734 (N_13734,N_13527,N_13605);
nor U13735 (N_13735,N_13511,N_13584);
or U13736 (N_13736,N_13594,N_13616);
nand U13737 (N_13737,N_13630,N_13511);
xnor U13738 (N_13738,N_13572,N_13545);
xnor U13739 (N_13739,N_13649,N_13577);
and U13740 (N_13740,N_13554,N_13559);
xor U13741 (N_13741,N_13553,N_13568);
nand U13742 (N_13742,N_13605,N_13504);
and U13743 (N_13743,N_13645,N_13637);
nor U13744 (N_13744,N_13580,N_13532);
or U13745 (N_13745,N_13552,N_13602);
or U13746 (N_13746,N_13520,N_13620);
and U13747 (N_13747,N_13640,N_13531);
xor U13748 (N_13748,N_13583,N_13647);
xor U13749 (N_13749,N_13588,N_13645);
and U13750 (N_13750,N_13557,N_13555);
and U13751 (N_13751,N_13567,N_13542);
nand U13752 (N_13752,N_13523,N_13586);
or U13753 (N_13753,N_13649,N_13584);
xor U13754 (N_13754,N_13514,N_13620);
nand U13755 (N_13755,N_13559,N_13618);
or U13756 (N_13756,N_13585,N_13584);
xnor U13757 (N_13757,N_13580,N_13506);
nand U13758 (N_13758,N_13602,N_13612);
nand U13759 (N_13759,N_13576,N_13641);
xor U13760 (N_13760,N_13536,N_13567);
nor U13761 (N_13761,N_13608,N_13647);
and U13762 (N_13762,N_13502,N_13637);
nand U13763 (N_13763,N_13597,N_13506);
nand U13764 (N_13764,N_13627,N_13642);
nand U13765 (N_13765,N_13571,N_13535);
nor U13766 (N_13766,N_13551,N_13537);
and U13767 (N_13767,N_13566,N_13600);
nand U13768 (N_13768,N_13606,N_13566);
or U13769 (N_13769,N_13635,N_13551);
and U13770 (N_13770,N_13594,N_13562);
nor U13771 (N_13771,N_13537,N_13576);
xor U13772 (N_13772,N_13613,N_13639);
and U13773 (N_13773,N_13510,N_13648);
nor U13774 (N_13774,N_13570,N_13611);
xor U13775 (N_13775,N_13554,N_13562);
nand U13776 (N_13776,N_13518,N_13579);
nand U13777 (N_13777,N_13559,N_13576);
nand U13778 (N_13778,N_13600,N_13580);
xnor U13779 (N_13779,N_13532,N_13502);
or U13780 (N_13780,N_13573,N_13595);
nand U13781 (N_13781,N_13576,N_13525);
xnor U13782 (N_13782,N_13529,N_13520);
xnor U13783 (N_13783,N_13571,N_13637);
or U13784 (N_13784,N_13587,N_13598);
nor U13785 (N_13785,N_13563,N_13537);
nor U13786 (N_13786,N_13642,N_13583);
xnor U13787 (N_13787,N_13612,N_13566);
nand U13788 (N_13788,N_13597,N_13569);
nand U13789 (N_13789,N_13606,N_13581);
nor U13790 (N_13790,N_13536,N_13513);
or U13791 (N_13791,N_13563,N_13565);
xor U13792 (N_13792,N_13591,N_13582);
or U13793 (N_13793,N_13638,N_13633);
or U13794 (N_13794,N_13587,N_13605);
nor U13795 (N_13795,N_13590,N_13593);
and U13796 (N_13796,N_13558,N_13522);
xnor U13797 (N_13797,N_13577,N_13540);
nor U13798 (N_13798,N_13623,N_13528);
xor U13799 (N_13799,N_13611,N_13630);
nand U13800 (N_13800,N_13726,N_13751);
nor U13801 (N_13801,N_13694,N_13686);
nand U13802 (N_13802,N_13719,N_13699);
nand U13803 (N_13803,N_13653,N_13754);
and U13804 (N_13804,N_13696,N_13765);
nor U13805 (N_13805,N_13766,N_13725);
xnor U13806 (N_13806,N_13675,N_13717);
nor U13807 (N_13807,N_13680,N_13741);
or U13808 (N_13808,N_13780,N_13791);
nand U13809 (N_13809,N_13703,N_13760);
nand U13810 (N_13810,N_13779,N_13666);
or U13811 (N_13811,N_13659,N_13728);
nor U13812 (N_13812,N_13656,N_13799);
nand U13813 (N_13813,N_13687,N_13664);
nand U13814 (N_13814,N_13693,N_13718);
nor U13815 (N_13815,N_13714,N_13738);
or U13816 (N_13816,N_13742,N_13715);
and U13817 (N_13817,N_13695,N_13785);
and U13818 (N_13818,N_13744,N_13690);
nor U13819 (N_13819,N_13735,N_13775);
xor U13820 (N_13820,N_13784,N_13792);
or U13821 (N_13821,N_13776,N_13730);
and U13822 (N_13822,N_13692,N_13685);
nor U13823 (N_13823,N_13722,N_13698);
nand U13824 (N_13824,N_13749,N_13764);
xor U13825 (N_13825,N_13716,N_13758);
nor U13826 (N_13826,N_13660,N_13790);
nor U13827 (N_13827,N_13743,N_13682);
xor U13828 (N_13828,N_13746,N_13684);
or U13829 (N_13829,N_13688,N_13713);
nor U13830 (N_13830,N_13721,N_13729);
xnor U13831 (N_13831,N_13769,N_13651);
or U13832 (N_13832,N_13762,N_13733);
and U13833 (N_13833,N_13672,N_13755);
xnor U13834 (N_13834,N_13676,N_13706);
or U13835 (N_13835,N_13771,N_13761);
xor U13836 (N_13836,N_13671,N_13670);
nand U13837 (N_13837,N_13669,N_13747);
nor U13838 (N_13838,N_13789,N_13770);
nand U13839 (N_13839,N_13674,N_13774);
or U13840 (N_13840,N_13677,N_13654);
nor U13841 (N_13841,N_13783,N_13748);
and U13842 (N_13842,N_13663,N_13657);
and U13843 (N_13843,N_13781,N_13734);
nand U13844 (N_13844,N_13745,N_13701);
xor U13845 (N_13845,N_13711,N_13795);
xnor U13846 (N_13846,N_13681,N_13652);
nand U13847 (N_13847,N_13665,N_13705);
and U13848 (N_13848,N_13732,N_13650);
xnor U13849 (N_13849,N_13667,N_13697);
and U13850 (N_13850,N_13661,N_13668);
nor U13851 (N_13851,N_13756,N_13704);
nand U13852 (N_13852,N_13757,N_13720);
xor U13853 (N_13853,N_13700,N_13736);
nand U13854 (N_13854,N_13727,N_13691);
nand U13855 (N_13855,N_13753,N_13739);
xor U13856 (N_13856,N_13724,N_13673);
xnor U13857 (N_13857,N_13778,N_13773);
xnor U13858 (N_13858,N_13709,N_13731);
or U13859 (N_13859,N_13678,N_13750);
xor U13860 (N_13860,N_13707,N_13798);
nor U13861 (N_13861,N_13662,N_13679);
nand U13862 (N_13862,N_13658,N_13772);
or U13863 (N_13863,N_13683,N_13655);
nand U13864 (N_13864,N_13723,N_13752);
nand U13865 (N_13865,N_13777,N_13710);
nor U13866 (N_13866,N_13786,N_13794);
or U13867 (N_13867,N_13788,N_13767);
and U13868 (N_13868,N_13796,N_13708);
and U13869 (N_13869,N_13763,N_13759);
or U13870 (N_13870,N_13737,N_13768);
or U13871 (N_13871,N_13797,N_13793);
or U13872 (N_13872,N_13712,N_13782);
xnor U13873 (N_13873,N_13787,N_13689);
xnor U13874 (N_13874,N_13702,N_13740);
and U13875 (N_13875,N_13791,N_13734);
nand U13876 (N_13876,N_13782,N_13732);
nand U13877 (N_13877,N_13781,N_13671);
xnor U13878 (N_13878,N_13780,N_13784);
xnor U13879 (N_13879,N_13682,N_13731);
xnor U13880 (N_13880,N_13681,N_13685);
or U13881 (N_13881,N_13777,N_13784);
xor U13882 (N_13882,N_13679,N_13691);
and U13883 (N_13883,N_13652,N_13695);
or U13884 (N_13884,N_13689,N_13711);
nor U13885 (N_13885,N_13727,N_13702);
nand U13886 (N_13886,N_13724,N_13721);
and U13887 (N_13887,N_13656,N_13741);
or U13888 (N_13888,N_13728,N_13763);
and U13889 (N_13889,N_13765,N_13747);
nand U13890 (N_13890,N_13692,N_13760);
or U13891 (N_13891,N_13732,N_13799);
and U13892 (N_13892,N_13770,N_13793);
or U13893 (N_13893,N_13666,N_13692);
or U13894 (N_13894,N_13676,N_13702);
xor U13895 (N_13895,N_13789,N_13787);
or U13896 (N_13896,N_13742,N_13670);
xnor U13897 (N_13897,N_13752,N_13796);
or U13898 (N_13898,N_13779,N_13707);
nand U13899 (N_13899,N_13699,N_13667);
and U13900 (N_13900,N_13787,N_13747);
or U13901 (N_13901,N_13686,N_13756);
and U13902 (N_13902,N_13661,N_13766);
xor U13903 (N_13903,N_13711,N_13780);
nor U13904 (N_13904,N_13770,N_13767);
nor U13905 (N_13905,N_13698,N_13706);
or U13906 (N_13906,N_13772,N_13795);
nand U13907 (N_13907,N_13695,N_13742);
nand U13908 (N_13908,N_13661,N_13787);
nor U13909 (N_13909,N_13673,N_13674);
nand U13910 (N_13910,N_13757,N_13666);
nand U13911 (N_13911,N_13662,N_13678);
nand U13912 (N_13912,N_13735,N_13682);
nand U13913 (N_13913,N_13717,N_13714);
and U13914 (N_13914,N_13724,N_13712);
or U13915 (N_13915,N_13732,N_13733);
nor U13916 (N_13916,N_13654,N_13754);
nor U13917 (N_13917,N_13784,N_13710);
xor U13918 (N_13918,N_13785,N_13739);
nor U13919 (N_13919,N_13730,N_13734);
or U13920 (N_13920,N_13762,N_13667);
or U13921 (N_13921,N_13666,N_13701);
nor U13922 (N_13922,N_13787,N_13666);
xor U13923 (N_13923,N_13755,N_13771);
nor U13924 (N_13924,N_13725,N_13742);
nor U13925 (N_13925,N_13746,N_13796);
and U13926 (N_13926,N_13655,N_13793);
and U13927 (N_13927,N_13762,N_13750);
xor U13928 (N_13928,N_13749,N_13727);
nor U13929 (N_13929,N_13769,N_13691);
nand U13930 (N_13930,N_13694,N_13791);
nor U13931 (N_13931,N_13717,N_13689);
xor U13932 (N_13932,N_13658,N_13784);
or U13933 (N_13933,N_13789,N_13661);
and U13934 (N_13934,N_13755,N_13714);
nor U13935 (N_13935,N_13746,N_13686);
xnor U13936 (N_13936,N_13751,N_13793);
and U13937 (N_13937,N_13782,N_13666);
or U13938 (N_13938,N_13706,N_13717);
nor U13939 (N_13939,N_13767,N_13650);
nor U13940 (N_13940,N_13693,N_13651);
or U13941 (N_13941,N_13676,N_13650);
nand U13942 (N_13942,N_13773,N_13722);
and U13943 (N_13943,N_13658,N_13709);
and U13944 (N_13944,N_13681,N_13739);
nor U13945 (N_13945,N_13699,N_13734);
xnor U13946 (N_13946,N_13730,N_13668);
nand U13947 (N_13947,N_13783,N_13732);
nand U13948 (N_13948,N_13737,N_13679);
and U13949 (N_13949,N_13793,N_13654);
or U13950 (N_13950,N_13892,N_13864);
xnor U13951 (N_13951,N_13804,N_13844);
xor U13952 (N_13952,N_13833,N_13825);
and U13953 (N_13953,N_13925,N_13853);
xor U13954 (N_13954,N_13807,N_13872);
nand U13955 (N_13955,N_13917,N_13880);
nand U13956 (N_13956,N_13865,N_13890);
or U13957 (N_13957,N_13826,N_13875);
and U13958 (N_13958,N_13930,N_13944);
nand U13959 (N_13959,N_13881,N_13812);
nor U13960 (N_13960,N_13846,N_13908);
nor U13961 (N_13961,N_13879,N_13888);
nand U13962 (N_13962,N_13911,N_13814);
xnor U13963 (N_13963,N_13909,N_13856);
and U13964 (N_13964,N_13947,N_13946);
xor U13965 (N_13965,N_13855,N_13926);
and U13966 (N_13966,N_13852,N_13802);
xnor U13967 (N_13967,N_13859,N_13941);
or U13968 (N_13968,N_13886,N_13839);
xnor U13969 (N_13969,N_13869,N_13929);
nor U13970 (N_13970,N_13940,N_13893);
xor U13971 (N_13971,N_13948,N_13942);
and U13972 (N_13972,N_13928,N_13830);
xnor U13973 (N_13973,N_13907,N_13897);
nand U13974 (N_13974,N_13836,N_13834);
nor U13975 (N_13975,N_13937,N_13916);
nor U13976 (N_13976,N_13887,N_13906);
nand U13977 (N_13977,N_13843,N_13882);
xor U13978 (N_13978,N_13811,N_13805);
nand U13979 (N_13979,N_13823,N_13813);
and U13980 (N_13980,N_13871,N_13935);
nor U13981 (N_13981,N_13803,N_13854);
xor U13982 (N_13982,N_13857,N_13945);
or U13983 (N_13983,N_13848,N_13847);
nor U13984 (N_13984,N_13806,N_13845);
xor U13985 (N_13985,N_13835,N_13896);
and U13986 (N_13986,N_13933,N_13810);
xor U13987 (N_13987,N_13820,N_13801);
xnor U13988 (N_13988,N_13922,N_13920);
or U13989 (N_13989,N_13943,N_13838);
or U13990 (N_13990,N_13918,N_13894);
nand U13991 (N_13991,N_13824,N_13949);
nand U13992 (N_13992,N_13912,N_13923);
xnor U13993 (N_13993,N_13900,N_13938);
nor U13994 (N_13994,N_13818,N_13841);
nor U13995 (N_13995,N_13858,N_13921);
and U13996 (N_13996,N_13874,N_13876);
and U13997 (N_13997,N_13889,N_13939);
nand U13998 (N_13998,N_13924,N_13800);
xor U13999 (N_13999,N_13808,N_13832);
nand U14000 (N_14000,N_13904,N_13932);
nand U14001 (N_14001,N_13863,N_13870);
or U14002 (N_14002,N_13840,N_13815);
xnor U14003 (N_14003,N_13931,N_13903);
or U14004 (N_14004,N_13919,N_13861);
and U14005 (N_14005,N_13899,N_13868);
xor U14006 (N_14006,N_13884,N_13849);
and U14007 (N_14007,N_13829,N_13913);
or U14008 (N_14008,N_13862,N_13915);
or U14009 (N_14009,N_13850,N_13901);
xor U14010 (N_14010,N_13914,N_13898);
nand U14011 (N_14011,N_13905,N_13831);
nor U14012 (N_14012,N_13895,N_13816);
and U14013 (N_14013,N_13927,N_13883);
nand U14014 (N_14014,N_13821,N_13851);
and U14015 (N_14015,N_13866,N_13936);
nor U14016 (N_14016,N_13891,N_13827);
or U14017 (N_14017,N_13809,N_13934);
nor U14018 (N_14018,N_13877,N_13910);
xnor U14019 (N_14019,N_13819,N_13878);
nor U14020 (N_14020,N_13828,N_13873);
nand U14021 (N_14021,N_13817,N_13867);
or U14022 (N_14022,N_13885,N_13837);
nand U14023 (N_14023,N_13902,N_13860);
or U14024 (N_14024,N_13822,N_13842);
or U14025 (N_14025,N_13826,N_13914);
and U14026 (N_14026,N_13893,N_13840);
or U14027 (N_14027,N_13818,N_13812);
xnor U14028 (N_14028,N_13929,N_13880);
nand U14029 (N_14029,N_13812,N_13869);
xnor U14030 (N_14030,N_13899,N_13833);
nor U14031 (N_14031,N_13913,N_13909);
or U14032 (N_14032,N_13932,N_13840);
xor U14033 (N_14033,N_13833,N_13835);
or U14034 (N_14034,N_13809,N_13850);
or U14035 (N_14035,N_13914,N_13944);
xor U14036 (N_14036,N_13935,N_13919);
or U14037 (N_14037,N_13817,N_13825);
nand U14038 (N_14038,N_13847,N_13854);
nor U14039 (N_14039,N_13903,N_13901);
xnor U14040 (N_14040,N_13925,N_13869);
xor U14041 (N_14041,N_13911,N_13869);
or U14042 (N_14042,N_13877,N_13908);
or U14043 (N_14043,N_13832,N_13814);
xor U14044 (N_14044,N_13847,N_13835);
nand U14045 (N_14045,N_13915,N_13810);
xor U14046 (N_14046,N_13839,N_13854);
or U14047 (N_14047,N_13883,N_13919);
nor U14048 (N_14048,N_13939,N_13907);
and U14049 (N_14049,N_13915,N_13841);
and U14050 (N_14050,N_13899,N_13839);
or U14051 (N_14051,N_13903,N_13865);
nand U14052 (N_14052,N_13813,N_13860);
nand U14053 (N_14053,N_13933,N_13833);
and U14054 (N_14054,N_13928,N_13907);
xor U14055 (N_14055,N_13811,N_13942);
and U14056 (N_14056,N_13849,N_13804);
or U14057 (N_14057,N_13848,N_13896);
and U14058 (N_14058,N_13903,N_13814);
xor U14059 (N_14059,N_13879,N_13814);
and U14060 (N_14060,N_13927,N_13937);
xor U14061 (N_14061,N_13838,N_13870);
and U14062 (N_14062,N_13940,N_13829);
nand U14063 (N_14063,N_13909,N_13807);
or U14064 (N_14064,N_13938,N_13944);
nor U14065 (N_14065,N_13885,N_13946);
nor U14066 (N_14066,N_13834,N_13838);
nor U14067 (N_14067,N_13889,N_13896);
nand U14068 (N_14068,N_13926,N_13927);
or U14069 (N_14069,N_13878,N_13803);
or U14070 (N_14070,N_13856,N_13836);
nor U14071 (N_14071,N_13852,N_13928);
and U14072 (N_14072,N_13840,N_13865);
xnor U14073 (N_14073,N_13836,N_13925);
nor U14074 (N_14074,N_13894,N_13817);
nand U14075 (N_14075,N_13849,N_13937);
nor U14076 (N_14076,N_13928,N_13860);
or U14077 (N_14077,N_13890,N_13934);
xnor U14078 (N_14078,N_13938,N_13857);
and U14079 (N_14079,N_13816,N_13948);
or U14080 (N_14080,N_13815,N_13863);
or U14081 (N_14081,N_13839,N_13859);
or U14082 (N_14082,N_13858,N_13826);
nor U14083 (N_14083,N_13849,N_13814);
and U14084 (N_14084,N_13830,N_13941);
or U14085 (N_14085,N_13839,N_13890);
nand U14086 (N_14086,N_13937,N_13909);
nand U14087 (N_14087,N_13911,N_13864);
nand U14088 (N_14088,N_13928,N_13906);
nand U14089 (N_14089,N_13945,N_13941);
or U14090 (N_14090,N_13825,N_13866);
nor U14091 (N_14091,N_13861,N_13913);
or U14092 (N_14092,N_13896,N_13911);
and U14093 (N_14093,N_13803,N_13932);
or U14094 (N_14094,N_13930,N_13888);
nand U14095 (N_14095,N_13829,N_13848);
nand U14096 (N_14096,N_13878,N_13840);
xor U14097 (N_14097,N_13838,N_13905);
or U14098 (N_14098,N_13804,N_13903);
xnor U14099 (N_14099,N_13848,N_13897);
nand U14100 (N_14100,N_13975,N_13985);
nor U14101 (N_14101,N_13982,N_14078);
or U14102 (N_14102,N_14004,N_14048);
and U14103 (N_14103,N_14038,N_14046);
nor U14104 (N_14104,N_13993,N_14059);
and U14105 (N_14105,N_14085,N_14045);
nand U14106 (N_14106,N_13981,N_13996);
nand U14107 (N_14107,N_14061,N_14033);
nor U14108 (N_14108,N_13995,N_14080);
nand U14109 (N_14109,N_14034,N_14007);
nand U14110 (N_14110,N_13984,N_14006);
or U14111 (N_14111,N_14098,N_13999);
xnor U14112 (N_14112,N_13971,N_14068);
xor U14113 (N_14113,N_13977,N_14073);
nand U14114 (N_14114,N_14064,N_14032);
and U14115 (N_14115,N_14031,N_14057);
nand U14116 (N_14116,N_14077,N_14060);
nor U14117 (N_14117,N_14000,N_14087);
nor U14118 (N_14118,N_13950,N_14089);
nand U14119 (N_14119,N_14018,N_13988);
nor U14120 (N_14120,N_14088,N_14090);
or U14121 (N_14121,N_14039,N_14092);
nor U14122 (N_14122,N_13965,N_14010);
nand U14123 (N_14123,N_13997,N_14044);
or U14124 (N_14124,N_13998,N_14075);
nor U14125 (N_14125,N_13953,N_13974);
nand U14126 (N_14126,N_14015,N_13972);
nand U14127 (N_14127,N_14040,N_14049);
nor U14128 (N_14128,N_14008,N_14097);
nand U14129 (N_14129,N_14047,N_14037);
and U14130 (N_14130,N_14009,N_13964);
and U14131 (N_14131,N_14011,N_13961);
or U14132 (N_14132,N_14093,N_14095);
nor U14133 (N_14133,N_13968,N_13980);
nor U14134 (N_14134,N_13973,N_14016);
xor U14135 (N_14135,N_14072,N_14083);
and U14136 (N_14136,N_13992,N_14074);
xnor U14137 (N_14137,N_13956,N_14017);
and U14138 (N_14138,N_13983,N_13986);
and U14139 (N_14139,N_13991,N_14052);
or U14140 (N_14140,N_14055,N_14099);
or U14141 (N_14141,N_13957,N_14081);
or U14142 (N_14142,N_14028,N_13951);
nand U14143 (N_14143,N_13979,N_13969);
nand U14144 (N_14144,N_14051,N_13960);
and U14145 (N_14145,N_14091,N_13962);
or U14146 (N_14146,N_13955,N_14062);
and U14147 (N_14147,N_14050,N_13994);
nand U14148 (N_14148,N_14013,N_13954);
nand U14149 (N_14149,N_14025,N_14058);
xor U14150 (N_14150,N_14066,N_14019);
or U14151 (N_14151,N_14056,N_14029);
nor U14152 (N_14152,N_14036,N_14021);
or U14153 (N_14153,N_14043,N_14065);
and U14154 (N_14154,N_13970,N_14003);
and U14155 (N_14155,N_13952,N_13978);
xor U14156 (N_14156,N_14035,N_14069);
nor U14157 (N_14157,N_14094,N_14041);
and U14158 (N_14158,N_14071,N_14079);
xnor U14159 (N_14159,N_14024,N_14022);
xnor U14160 (N_14160,N_14053,N_14005);
xnor U14161 (N_14161,N_13987,N_13967);
nand U14162 (N_14162,N_14082,N_14012);
nor U14163 (N_14163,N_14063,N_14076);
and U14164 (N_14164,N_14096,N_14067);
nor U14165 (N_14165,N_14084,N_14030);
nor U14166 (N_14166,N_13958,N_13989);
and U14167 (N_14167,N_13976,N_14014);
nand U14168 (N_14168,N_14086,N_13963);
nor U14169 (N_14169,N_14070,N_14023);
and U14170 (N_14170,N_13966,N_13959);
xnor U14171 (N_14171,N_14001,N_14020);
or U14172 (N_14172,N_14042,N_14026);
or U14173 (N_14173,N_14027,N_14054);
and U14174 (N_14174,N_13990,N_14002);
nor U14175 (N_14175,N_13961,N_14053);
and U14176 (N_14176,N_13950,N_13954);
nor U14177 (N_14177,N_14092,N_14024);
nand U14178 (N_14178,N_14010,N_14087);
and U14179 (N_14179,N_14064,N_14020);
nand U14180 (N_14180,N_14011,N_13959);
xor U14181 (N_14181,N_14044,N_14016);
and U14182 (N_14182,N_14013,N_14032);
and U14183 (N_14183,N_14078,N_14021);
nand U14184 (N_14184,N_14074,N_14044);
nor U14185 (N_14185,N_13999,N_14081);
xnor U14186 (N_14186,N_14023,N_14042);
or U14187 (N_14187,N_13998,N_14050);
nand U14188 (N_14188,N_14050,N_14031);
or U14189 (N_14189,N_13993,N_14050);
or U14190 (N_14190,N_14099,N_13977);
nor U14191 (N_14191,N_14089,N_14076);
and U14192 (N_14192,N_14062,N_14043);
and U14193 (N_14193,N_14099,N_13959);
and U14194 (N_14194,N_14027,N_14009);
and U14195 (N_14195,N_13965,N_14090);
or U14196 (N_14196,N_14001,N_14076);
xnor U14197 (N_14197,N_13950,N_14050);
xnor U14198 (N_14198,N_14083,N_14041);
or U14199 (N_14199,N_14025,N_14098);
xor U14200 (N_14200,N_14038,N_14040);
and U14201 (N_14201,N_14020,N_14008);
xor U14202 (N_14202,N_14054,N_13991);
nor U14203 (N_14203,N_14072,N_13968);
nor U14204 (N_14204,N_13957,N_13959);
or U14205 (N_14205,N_14070,N_14004);
nand U14206 (N_14206,N_14016,N_14026);
xor U14207 (N_14207,N_14069,N_14007);
nand U14208 (N_14208,N_14063,N_13955);
xnor U14209 (N_14209,N_14091,N_13982);
xnor U14210 (N_14210,N_14084,N_14028);
or U14211 (N_14211,N_14061,N_14014);
and U14212 (N_14212,N_14023,N_14097);
or U14213 (N_14213,N_13973,N_14065);
or U14214 (N_14214,N_14020,N_14052);
nor U14215 (N_14215,N_14081,N_14028);
and U14216 (N_14216,N_14044,N_14065);
and U14217 (N_14217,N_14030,N_14019);
nand U14218 (N_14218,N_13995,N_14042);
nor U14219 (N_14219,N_14037,N_14040);
nand U14220 (N_14220,N_13950,N_14087);
xor U14221 (N_14221,N_13951,N_14058);
or U14222 (N_14222,N_13964,N_14021);
nand U14223 (N_14223,N_13988,N_13950);
or U14224 (N_14224,N_14043,N_13988);
nand U14225 (N_14225,N_13960,N_14024);
and U14226 (N_14226,N_14091,N_14031);
or U14227 (N_14227,N_14033,N_14007);
nand U14228 (N_14228,N_14098,N_13954);
or U14229 (N_14229,N_14027,N_13994);
xnor U14230 (N_14230,N_14076,N_13968);
nor U14231 (N_14231,N_13964,N_13962);
and U14232 (N_14232,N_14065,N_13965);
xor U14233 (N_14233,N_13977,N_13967);
xor U14234 (N_14234,N_13978,N_14089);
xnor U14235 (N_14235,N_13954,N_14024);
nor U14236 (N_14236,N_14065,N_13983);
nor U14237 (N_14237,N_13957,N_14041);
and U14238 (N_14238,N_13980,N_14062);
nor U14239 (N_14239,N_14066,N_14068);
and U14240 (N_14240,N_14055,N_14040);
xnor U14241 (N_14241,N_13965,N_14045);
or U14242 (N_14242,N_13982,N_14064);
or U14243 (N_14243,N_13988,N_14063);
xnor U14244 (N_14244,N_14041,N_14022);
or U14245 (N_14245,N_14057,N_14094);
or U14246 (N_14246,N_13953,N_13968);
nand U14247 (N_14247,N_13992,N_13956);
nand U14248 (N_14248,N_14092,N_13998);
xor U14249 (N_14249,N_14091,N_13972);
or U14250 (N_14250,N_14162,N_14101);
xor U14251 (N_14251,N_14241,N_14119);
xnor U14252 (N_14252,N_14249,N_14182);
or U14253 (N_14253,N_14168,N_14247);
and U14254 (N_14254,N_14161,N_14213);
nand U14255 (N_14255,N_14169,N_14136);
nor U14256 (N_14256,N_14235,N_14114);
or U14257 (N_14257,N_14203,N_14180);
nor U14258 (N_14258,N_14166,N_14157);
or U14259 (N_14259,N_14217,N_14199);
and U14260 (N_14260,N_14248,N_14227);
xor U14261 (N_14261,N_14244,N_14100);
xor U14262 (N_14262,N_14155,N_14194);
xor U14263 (N_14263,N_14118,N_14219);
xnor U14264 (N_14264,N_14245,N_14156);
nor U14265 (N_14265,N_14149,N_14193);
or U14266 (N_14266,N_14115,N_14223);
and U14267 (N_14267,N_14145,N_14148);
or U14268 (N_14268,N_14220,N_14186);
nand U14269 (N_14269,N_14122,N_14110);
nor U14270 (N_14270,N_14151,N_14154);
and U14271 (N_14271,N_14230,N_14107);
or U14272 (N_14272,N_14197,N_14196);
nor U14273 (N_14273,N_14132,N_14211);
nand U14274 (N_14274,N_14215,N_14112);
nor U14275 (N_14275,N_14130,N_14127);
nand U14276 (N_14276,N_14187,N_14181);
xnor U14277 (N_14277,N_14147,N_14205);
and U14278 (N_14278,N_14240,N_14189);
xor U14279 (N_14279,N_14228,N_14242);
and U14280 (N_14280,N_14214,N_14200);
xnor U14281 (N_14281,N_14139,N_14212);
or U14282 (N_14282,N_14106,N_14123);
xnor U14283 (N_14283,N_14134,N_14208);
and U14284 (N_14284,N_14108,N_14120);
nor U14285 (N_14285,N_14141,N_14150);
and U14286 (N_14286,N_14216,N_14239);
or U14287 (N_14287,N_14144,N_14138);
nand U14288 (N_14288,N_14229,N_14178);
or U14289 (N_14289,N_14125,N_14175);
nor U14290 (N_14290,N_14137,N_14224);
and U14291 (N_14291,N_14170,N_14143);
xor U14292 (N_14292,N_14204,N_14195);
and U14293 (N_14293,N_14116,N_14103);
nor U14294 (N_14294,N_14124,N_14160);
nand U14295 (N_14295,N_14135,N_14201);
and U14296 (N_14296,N_14206,N_14209);
or U14297 (N_14297,N_14238,N_14218);
and U14298 (N_14298,N_14164,N_14173);
nor U14299 (N_14299,N_14192,N_14163);
or U14300 (N_14300,N_14185,N_14126);
xor U14301 (N_14301,N_14237,N_14222);
or U14302 (N_14302,N_14225,N_14152);
nand U14303 (N_14303,N_14102,N_14128);
or U14304 (N_14304,N_14105,N_14179);
and U14305 (N_14305,N_14231,N_14153);
or U14306 (N_14306,N_14171,N_14188);
nor U14307 (N_14307,N_14165,N_14129);
xor U14308 (N_14308,N_14146,N_14236);
nor U14309 (N_14309,N_14131,N_14117);
nor U14310 (N_14310,N_14172,N_14104);
nand U14311 (N_14311,N_14140,N_14177);
xnor U14312 (N_14312,N_14159,N_14232);
nand U14313 (N_14313,N_14221,N_14207);
and U14314 (N_14314,N_14191,N_14113);
and U14315 (N_14315,N_14167,N_14198);
nor U14316 (N_14316,N_14142,N_14190);
xnor U14317 (N_14317,N_14111,N_14243);
and U14318 (N_14318,N_14246,N_14109);
xnor U14319 (N_14319,N_14183,N_14210);
xnor U14320 (N_14320,N_14184,N_14176);
xnor U14321 (N_14321,N_14202,N_14234);
and U14322 (N_14322,N_14226,N_14121);
or U14323 (N_14323,N_14133,N_14174);
nand U14324 (N_14324,N_14233,N_14158);
nand U14325 (N_14325,N_14206,N_14182);
nor U14326 (N_14326,N_14150,N_14221);
or U14327 (N_14327,N_14238,N_14241);
xor U14328 (N_14328,N_14246,N_14198);
and U14329 (N_14329,N_14239,N_14120);
or U14330 (N_14330,N_14241,N_14235);
and U14331 (N_14331,N_14211,N_14195);
or U14332 (N_14332,N_14175,N_14227);
nor U14333 (N_14333,N_14138,N_14152);
and U14334 (N_14334,N_14191,N_14152);
nor U14335 (N_14335,N_14237,N_14207);
or U14336 (N_14336,N_14178,N_14176);
nand U14337 (N_14337,N_14139,N_14243);
and U14338 (N_14338,N_14192,N_14138);
or U14339 (N_14339,N_14211,N_14227);
nand U14340 (N_14340,N_14172,N_14170);
or U14341 (N_14341,N_14127,N_14111);
or U14342 (N_14342,N_14123,N_14217);
nand U14343 (N_14343,N_14194,N_14158);
or U14344 (N_14344,N_14145,N_14162);
or U14345 (N_14345,N_14137,N_14155);
or U14346 (N_14346,N_14207,N_14205);
nand U14347 (N_14347,N_14211,N_14226);
or U14348 (N_14348,N_14109,N_14134);
nand U14349 (N_14349,N_14215,N_14164);
nor U14350 (N_14350,N_14137,N_14221);
xor U14351 (N_14351,N_14133,N_14218);
and U14352 (N_14352,N_14213,N_14135);
or U14353 (N_14353,N_14176,N_14213);
nor U14354 (N_14354,N_14222,N_14175);
xnor U14355 (N_14355,N_14247,N_14113);
nor U14356 (N_14356,N_14136,N_14230);
and U14357 (N_14357,N_14153,N_14119);
xor U14358 (N_14358,N_14167,N_14175);
xnor U14359 (N_14359,N_14200,N_14137);
xnor U14360 (N_14360,N_14143,N_14211);
and U14361 (N_14361,N_14107,N_14223);
xor U14362 (N_14362,N_14244,N_14131);
or U14363 (N_14363,N_14244,N_14170);
nand U14364 (N_14364,N_14117,N_14129);
nor U14365 (N_14365,N_14203,N_14143);
and U14366 (N_14366,N_14197,N_14244);
nor U14367 (N_14367,N_14125,N_14174);
nand U14368 (N_14368,N_14168,N_14230);
nand U14369 (N_14369,N_14189,N_14226);
or U14370 (N_14370,N_14205,N_14193);
xor U14371 (N_14371,N_14120,N_14147);
xor U14372 (N_14372,N_14243,N_14149);
or U14373 (N_14373,N_14108,N_14129);
nand U14374 (N_14374,N_14161,N_14169);
nand U14375 (N_14375,N_14163,N_14138);
xor U14376 (N_14376,N_14178,N_14187);
nand U14377 (N_14377,N_14120,N_14237);
nand U14378 (N_14378,N_14178,N_14161);
nor U14379 (N_14379,N_14101,N_14203);
nand U14380 (N_14380,N_14160,N_14212);
xor U14381 (N_14381,N_14108,N_14206);
nand U14382 (N_14382,N_14219,N_14185);
nand U14383 (N_14383,N_14226,N_14143);
nand U14384 (N_14384,N_14157,N_14214);
nand U14385 (N_14385,N_14125,N_14230);
or U14386 (N_14386,N_14237,N_14205);
nor U14387 (N_14387,N_14122,N_14133);
nor U14388 (N_14388,N_14190,N_14151);
nor U14389 (N_14389,N_14173,N_14236);
or U14390 (N_14390,N_14115,N_14106);
nor U14391 (N_14391,N_14232,N_14219);
xor U14392 (N_14392,N_14215,N_14106);
nand U14393 (N_14393,N_14206,N_14246);
nand U14394 (N_14394,N_14194,N_14221);
and U14395 (N_14395,N_14155,N_14103);
xnor U14396 (N_14396,N_14177,N_14154);
xnor U14397 (N_14397,N_14193,N_14240);
nor U14398 (N_14398,N_14106,N_14198);
nand U14399 (N_14399,N_14207,N_14151);
or U14400 (N_14400,N_14358,N_14268);
or U14401 (N_14401,N_14364,N_14389);
nand U14402 (N_14402,N_14260,N_14306);
nand U14403 (N_14403,N_14316,N_14394);
nor U14404 (N_14404,N_14393,N_14338);
and U14405 (N_14405,N_14353,N_14309);
xnor U14406 (N_14406,N_14337,N_14387);
nor U14407 (N_14407,N_14279,N_14314);
nor U14408 (N_14408,N_14335,N_14351);
xnor U14409 (N_14409,N_14320,N_14342);
xor U14410 (N_14410,N_14341,N_14304);
or U14411 (N_14411,N_14308,N_14333);
xnor U14412 (N_14412,N_14330,N_14296);
nand U14413 (N_14413,N_14311,N_14383);
nand U14414 (N_14414,N_14332,N_14310);
xor U14415 (N_14415,N_14371,N_14266);
and U14416 (N_14416,N_14328,N_14271);
xor U14417 (N_14417,N_14315,N_14374);
nor U14418 (N_14418,N_14297,N_14360);
xor U14419 (N_14419,N_14323,N_14265);
nand U14420 (N_14420,N_14354,N_14349);
or U14421 (N_14421,N_14388,N_14288);
and U14422 (N_14422,N_14317,N_14272);
nor U14423 (N_14423,N_14299,N_14385);
or U14424 (N_14424,N_14283,N_14390);
nor U14425 (N_14425,N_14380,N_14263);
nand U14426 (N_14426,N_14298,N_14352);
or U14427 (N_14427,N_14340,N_14292);
nor U14428 (N_14428,N_14356,N_14274);
nand U14429 (N_14429,N_14280,N_14348);
nand U14430 (N_14430,N_14258,N_14325);
and U14431 (N_14431,N_14275,N_14350);
nor U14432 (N_14432,N_14397,N_14251);
xor U14433 (N_14433,N_14264,N_14273);
and U14434 (N_14434,N_14285,N_14363);
nor U14435 (N_14435,N_14366,N_14253);
xnor U14436 (N_14436,N_14278,N_14286);
nand U14437 (N_14437,N_14294,N_14329);
and U14438 (N_14438,N_14368,N_14300);
nor U14439 (N_14439,N_14276,N_14321);
or U14440 (N_14440,N_14375,N_14396);
or U14441 (N_14441,N_14290,N_14334);
and U14442 (N_14442,N_14384,N_14324);
nor U14443 (N_14443,N_14399,N_14381);
nand U14444 (N_14444,N_14287,N_14301);
and U14445 (N_14445,N_14250,N_14267);
xnor U14446 (N_14446,N_14269,N_14339);
nand U14447 (N_14447,N_14254,N_14293);
nor U14448 (N_14448,N_14346,N_14391);
nor U14449 (N_14449,N_14367,N_14257);
xnor U14450 (N_14450,N_14365,N_14379);
xor U14451 (N_14451,N_14395,N_14305);
nor U14452 (N_14452,N_14376,N_14319);
nand U14453 (N_14453,N_14262,N_14261);
and U14454 (N_14454,N_14252,N_14284);
xnor U14455 (N_14455,N_14357,N_14303);
nand U14456 (N_14456,N_14256,N_14277);
and U14457 (N_14457,N_14281,N_14386);
and U14458 (N_14458,N_14270,N_14322);
xor U14459 (N_14459,N_14373,N_14345);
or U14460 (N_14460,N_14377,N_14355);
and U14461 (N_14461,N_14259,N_14369);
nor U14462 (N_14462,N_14295,N_14361);
and U14463 (N_14463,N_14382,N_14347);
nor U14464 (N_14464,N_14326,N_14255);
nand U14465 (N_14465,N_14282,N_14359);
xnor U14466 (N_14466,N_14343,N_14398);
or U14467 (N_14467,N_14313,N_14312);
nor U14468 (N_14468,N_14307,N_14331);
nor U14469 (N_14469,N_14372,N_14318);
xor U14470 (N_14470,N_14336,N_14392);
or U14471 (N_14471,N_14291,N_14344);
or U14472 (N_14472,N_14327,N_14362);
or U14473 (N_14473,N_14289,N_14378);
nor U14474 (N_14474,N_14302,N_14370);
nor U14475 (N_14475,N_14370,N_14289);
or U14476 (N_14476,N_14287,N_14334);
nand U14477 (N_14477,N_14317,N_14375);
xor U14478 (N_14478,N_14323,N_14324);
nand U14479 (N_14479,N_14368,N_14274);
nor U14480 (N_14480,N_14341,N_14399);
nand U14481 (N_14481,N_14356,N_14327);
xnor U14482 (N_14482,N_14325,N_14309);
or U14483 (N_14483,N_14283,N_14305);
xnor U14484 (N_14484,N_14328,N_14338);
xor U14485 (N_14485,N_14283,N_14300);
or U14486 (N_14486,N_14291,N_14329);
and U14487 (N_14487,N_14367,N_14397);
or U14488 (N_14488,N_14397,N_14380);
nor U14489 (N_14489,N_14369,N_14266);
xor U14490 (N_14490,N_14360,N_14316);
xor U14491 (N_14491,N_14251,N_14339);
nor U14492 (N_14492,N_14355,N_14255);
xor U14493 (N_14493,N_14267,N_14283);
nand U14494 (N_14494,N_14363,N_14355);
nand U14495 (N_14495,N_14398,N_14364);
and U14496 (N_14496,N_14286,N_14290);
or U14497 (N_14497,N_14372,N_14361);
or U14498 (N_14498,N_14380,N_14339);
nor U14499 (N_14499,N_14274,N_14390);
xnor U14500 (N_14500,N_14306,N_14287);
nor U14501 (N_14501,N_14360,N_14250);
nor U14502 (N_14502,N_14251,N_14285);
and U14503 (N_14503,N_14397,N_14292);
nand U14504 (N_14504,N_14304,N_14361);
or U14505 (N_14505,N_14281,N_14349);
and U14506 (N_14506,N_14283,N_14281);
nand U14507 (N_14507,N_14291,N_14378);
nand U14508 (N_14508,N_14374,N_14258);
nand U14509 (N_14509,N_14320,N_14284);
or U14510 (N_14510,N_14341,N_14370);
and U14511 (N_14511,N_14368,N_14315);
nor U14512 (N_14512,N_14262,N_14364);
or U14513 (N_14513,N_14332,N_14330);
nand U14514 (N_14514,N_14347,N_14348);
or U14515 (N_14515,N_14287,N_14387);
nand U14516 (N_14516,N_14259,N_14311);
or U14517 (N_14517,N_14353,N_14366);
xnor U14518 (N_14518,N_14283,N_14268);
or U14519 (N_14519,N_14268,N_14286);
nand U14520 (N_14520,N_14257,N_14294);
or U14521 (N_14521,N_14269,N_14336);
or U14522 (N_14522,N_14313,N_14274);
nand U14523 (N_14523,N_14253,N_14322);
and U14524 (N_14524,N_14301,N_14390);
nor U14525 (N_14525,N_14328,N_14348);
xor U14526 (N_14526,N_14369,N_14258);
and U14527 (N_14527,N_14382,N_14383);
nand U14528 (N_14528,N_14343,N_14310);
nand U14529 (N_14529,N_14303,N_14273);
nor U14530 (N_14530,N_14268,N_14388);
xor U14531 (N_14531,N_14312,N_14372);
or U14532 (N_14532,N_14252,N_14263);
xor U14533 (N_14533,N_14342,N_14323);
nand U14534 (N_14534,N_14329,N_14365);
and U14535 (N_14535,N_14350,N_14253);
or U14536 (N_14536,N_14281,N_14328);
and U14537 (N_14537,N_14254,N_14370);
nand U14538 (N_14538,N_14387,N_14369);
xor U14539 (N_14539,N_14340,N_14252);
xor U14540 (N_14540,N_14383,N_14263);
or U14541 (N_14541,N_14287,N_14347);
nand U14542 (N_14542,N_14255,N_14399);
nor U14543 (N_14543,N_14390,N_14305);
nor U14544 (N_14544,N_14392,N_14332);
nor U14545 (N_14545,N_14370,N_14342);
xor U14546 (N_14546,N_14271,N_14360);
nor U14547 (N_14547,N_14336,N_14333);
and U14548 (N_14548,N_14346,N_14350);
xor U14549 (N_14549,N_14366,N_14251);
and U14550 (N_14550,N_14527,N_14439);
nand U14551 (N_14551,N_14458,N_14423);
or U14552 (N_14552,N_14414,N_14430);
xnor U14553 (N_14553,N_14406,N_14465);
xor U14554 (N_14554,N_14533,N_14490);
and U14555 (N_14555,N_14456,N_14521);
xor U14556 (N_14556,N_14469,N_14449);
or U14557 (N_14557,N_14511,N_14419);
and U14558 (N_14558,N_14534,N_14532);
nand U14559 (N_14559,N_14546,N_14545);
nand U14560 (N_14560,N_14515,N_14503);
nor U14561 (N_14561,N_14524,N_14452);
or U14562 (N_14562,N_14429,N_14416);
xor U14563 (N_14563,N_14421,N_14445);
nand U14564 (N_14564,N_14529,N_14492);
nand U14565 (N_14565,N_14462,N_14493);
or U14566 (N_14566,N_14468,N_14495);
xor U14567 (N_14567,N_14478,N_14438);
and U14568 (N_14568,N_14473,N_14483);
or U14569 (N_14569,N_14488,N_14505);
nor U14570 (N_14570,N_14442,N_14472);
nor U14571 (N_14571,N_14408,N_14522);
and U14572 (N_14572,N_14513,N_14540);
or U14573 (N_14573,N_14501,N_14497);
xnor U14574 (N_14574,N_14548,N_14507);
nand U14575 (N_14575,N_14502,N_14475);
xnor U14576 (N_14576,N_14436,N_14433);
and U14577 (N_14577,N_14525,N_14494);
nand U14578 (N_14578,N_14415,N_14482);
nor U14579 (N_14579,N_14413,N_14437);
nor U14580 (N_14580,N_14491,N_14451);
nor U14581 (N_14581,N_14435,N_14481);
nor U14582 (N_14582,N_14487,N_14520);
xnor U14583 (N_14583,N_14455,N_14518);
or U14584 (N_14584,N_14538,N_14476);
and U14585 (N_14585,N_14528,N_14454);
and U14586 (N_14586,N_14407,N_14517);
nor U14587 (N_14587,N_14453,N_14508);
and U14588 (N_14588,N_14461,N_14499);
nand U14589 (N_14589,N_14420,N_14542);
and U14590 (N_14590,N_14471,N_14460);
and U14591 (N_14591,N_14530,N_14531);
xor U14592 (N_14592,N_14440,N_14426);
and U14593 (N_14593,N_14411,N_14485);
nand U14594 (N_14594,N_14480,N_14500);
or U14595 (N_14595,N_14410,N_14539);
nor U14596 (N_14596,N_14427,N_14467);
nor U14597 (N_14597,N_14403,N_14510);
nand U14598 (N_14598,N_14523,N_14526);
or U14599 (N_14599,N_14434,N_14459);
nand U14600 (N_14600,N_14448,N_14544);
and U14601 (N_14601,N_14432,N_14409);
and U14602 (N_14602,N_14418,N_14463);
nor U14603 (N_14603,N_14474,N_14541);
and U14604 (N_14604,N_14504,N_14417);
xnor U14605 (N_14605,N_14457,N_14401);
nand U14606 (N_14606,N_14516,N_14484);
or U14607 (N_14607,N_14535,N_14549);
or U14608 (N_14608,N_14498,N_14512);
or U14609 (N_14609,N_14477,N_14470);
xnor U14610 (N_14610,N_14547,N_14543);
xor U14611 (N_14611,N_14514,N_14506);
nor U14612 (N_14612,N_14509,N_14464);
nor U14613 (N_14613,N_14479,N_14447);
and U14614 (N_14614,N_14441,N_14466);
xnor U14615 (N_14615,N_14536,N_14428);
nand U14616 (N_14616,N_14444,N_14446);
or U14617 (N_14617,N_14537,N_14422);
nand U14618 (N_14618,N_14486,N_14519);
xor U14619 (N_14619,N_14489,N_14400);
xor U14620 (N_14620,N_14424,N_14412);
and U14621 (N_14621,N_14443,N_14496);
xnor U14622 (N_14622,N_14450,N_14425);
nand U14623 (N_14623,N_14405,N_14402);
or U14624 (N_14624,N_14431,N_14404);
or U14625 (N_14625,N_14417,N_14410);
or U14626 (N_14626,N_14525,N_14535);
or U14627 (N_14627,N_14503,N_14469);
and U14628 (N_14628,N_14546,N_14430);
or U14629 (N_14629,N_14423,N_14491);
or U14630 (N_14630,N_14406,N_14548);
nand U14631 (N_14631,N_14501,N_14517);
xnor U14632 (N_14632,N_14500,N_14432);
and U14633 (N_14633,N_14440,N_14520);
nor U14634 (N_14634,N_14438,N_14462);
nand U14635 (N_14635,N_14504,N_14517);
xor U14636 (N_14636,N_14501,N_14547);
xnor U14637 (N_14637,N_14423,N_14476);
nand U14638 (N_14638,N_14490,N_14404);
nand U14639 (N_14639,N_14498,N_14490);
xnor U14640 (N_14640,N_14546,N_14429);
nand U14641 (N_14641,N_14488,N_14425);
nor U14642 (N_14642,N_14402,N_14534);
xnor U14643 (N_14643,N_14483,N_14424);
nor U14644 (N_14644,N_14533,N_14420);
and U14645 (N_14645,N_14511,N_14525);
and U14646 (N_14646,N_14413,N_14474);
or U14647 (N_14647,N_14407,N_14529);
nor U14648 (N_14648,N_14437,N_14470);
xor U14649 (N_14649,N_14456,N_14491);
nand U14650 (N_14650,N_14530,N_14448);
or U14651 (N_14651,N_14426,N_14442);
or U14652 (N_14652,N_14488,N_14416);
or U14653 (N_14653,N_14461,N_14443);
nand U14654 (N_14654,N_14528,N_14422);
nor U14655 (N_14655,N_14469,N_14528);
and U14656 (N_14656,N_14540,N_14447);
nor U14657 (N_14657,N_14482,N_14548);
or U14658 (N_14658,N_14525,N_14514);
and U14659 (N_14659,N_14541,N_14539);
nand U14660 (N_14660,N_14526,N_14467);
or U14661 (N_14661,N_14414,N_14545);
nand U14662 (N_14662,N_14490,N_14522);
or U14663 (N_14663,N_14438,N_14514);
xnor U14664 (N_14664,N_14487,N_14491);
or U14665 (N_14665,N_14510,N_14472);
xnor U14666 (N_14666,N_14509,N_14419);
nand U14667 (N_14667,N_14480,N_14423);
xor U14668 (N_14668,N_14502,N_14443);
nor U14669 (N_14669,N_14477,N_14478);
and U14670 (N_14670,N_14410,N_14548);
xnor U14671 (N_14671,N_14539,N_14524);
or U14672 (N_14672,N_14494,N_14421);
xnor U14673 (N_14673,N_14445,N_14496);
nand U14674 (N_14674,N_14522,N_14511);
xor U14675 (N_14675,N_14549,N_14523);
or U14676 (N_14676,N_14548,N_14435);
or U14677 (N_14677,N_14426,N_14520);
xnor U14678 (N_14678,N_14488,N_14500);
xnor U14679 (N_14679,N_14428,N_14480);
and U14680 (N_14680,N_14528,N_14458);
or U14681 (N_14681,N_14527,N_14444);
nor U14682 (N_14682,N_14477,N_14406);
nand U14683 (N_14683,N_14430,N_14465);
nand U14684 (N_14684,N_14523,N_14522);
xor U14685 (N_14685,N_14494,N_14402);
or U14686 (N_14686,N_14486,N_14455);
nand U14687 (N_14687,N_14504,N_14467);
or U14688 (N_14688,N_14495,N_14449);
and U14689 (N_14689,N_14520,N_14461);
or U14690 (N_14690,N_14501,N_14455);
and U14691 (N_14691,N_14535,N_14467);
xor U14692 (N_14692,N_14491,N_14462);
xor U14693 (N_14693,N_14509,N_14510);
xor U14694 (N_14694,N_14503,N_14511);
nand U14695 (N_14695,N_14526,N_14489);
and U14696 (N_14696,N_14524,N_14478);
or U14697 (N_14697,N_14499,N_14531);
or U14698 (N_14698,N_14445,N_14494);
nand U14699 (N_14699,N_14478,N_14450);
or U14700 (N_14700,N_14552,N_14618);
and U14701 (N_14701,N_14615,N_14642);
and U14702 (N_14702,N_14587,N_14652);
or U14703 (N_14703,N_14562,N_14666);
nand U14704 (N_14704,N_14621,N_14609);
or U14705 (N_14705,N_14683,N_14691);
nor U14706 (N_14706,N_14571,N_14688);
xor U14707 (N_14707,N_14566,N_14631);
or U14708 (N_14708,N_14656,N_14603);
and U14709 (N_14709,N_14674,N_14696);
and U14710 (N_14710,N_14561,N_14601);
and U14711 (N_14711,N_14558,N_14675);
and U14712 (N_14712,N_14598,N_14551);
xor U14713 (N_14713,N_14567,N_14677);
and U14714 (N_14714,N_14629,N_14689);
and U14715 (N_14715,N_14625,N_14659);
nand U14716 (N_14716,N_14636,N_14581);
or U14717 (N_14717,N_14678,N_14638);
xor U14718 (N_14718,N_14639,N_14588);
nor U14719 (N_14719,N_14637,N_14654);
xnor U14720 (N_14720,N_14557,N_14590);
xnor U14721 (N_14721,N_14664,N_14597);
xor U14722 (N_14722,N_14679,N_14699);
or U14723 (N_14723,N_14644,N_14628);
and U14724 (N_14724,N_14617,N_14655);
xor U14725 (N_14725,N_14563,N_14694);
nor U14726 (N_14726,N_14661,N_14633);
and U14727 (N_14727,N_14573,N_14667);
and U14728 (N_14728,N_14632,N_14580);
nand U14729 (N_14729,N_14579,N_14649);
or U14730 (N_14730,N_14564,N_14627);
nand U14731 (N_14731,N_14653,N_14616);
nor U14732 (N_14732,N_14589,N_14591);
or U14733 (N_14733,N_14635,N_14550);
nor U14734 (N_14734,N_14612,N_14695);
nor U14735 (N_14735,N_14614,N_14592);
nor U14736 (N_14736,N_14572,N_14555);
xnor U14737 (N_14737,N_14608,N_14575);
nand U14738 (N_14738,N_14693,N_14605);
xor U14739 (N_14739,N_14619,N_14604);
nand U14740 (N_14740,N_14595,N_14553);
nand U14741 (N_14741,N_14669,N_14650);
nor U14742 (N_14742,N_14574,N_14630);
and U14743 (N_14743,N_14682,N_14687);
or U14744 (N_14744,N_14560,N_14576);
nand U14745 (N_14745,N_14570,N_14611);
and U14746 (N_14746,N_14648,N_14554);
xnor U14747 (N_14747,N_14577,N_14586);
and U14748 (N_14748,N_14673,N_14556);
nor U14749 (N_14749,N_14585,N_14643);
and U14750 (N_14750,N_14583,N_14559);
or U14751 (N_14751,N_14657,N_14698);
nor U14752 (N_14752,N_14565,N_14665);
nand U14753 (N_14753,N_14658,N_14602);
nor U14754 (N_14754,N_14641,N_14690);
xor U14755 (N_14755,N_14645,N_14606);
and U14756 (N_14756,N_14697,N_14623);
and U14757 (N_14757,N_14670,N_14626);
or U14758 (N_14758,N_14686,N_14599);
xor U14759 (N_14759,N_14676,N_14578);
or U14760 (N_14760,N_14640,N_14663);
nand U14761 (N_14761,N_14685,N_14672);
xnor U14762 (N_14762,N_14593,N_14634);
or U14763 (N_14763,N_14668,N_14596);
nand U14764 (N_14764,N_14692,N_14582);
nor U14765 (N_14765,N_14620,N_14624);
nor U14766 (N_14766,N_14671,N_14569);
nand U14767 (N_14767,N_14613,N_14681);
nor U14768 (N_14768,N_14680,N_14607);
or U14769 (N_14769,N_14662,N_14568);
nand U14770 (N_14770,N_14660,N_14684);
or U14771 (N_14771,N_14600,N_14646);
and U14772 (N_14772,N_14651,N_14647);
xor U14773 (N_14773,N_14622,N_14584);
xnor U14774 (N_14774,N_14610,N_14594);
and U14775 (N_14775,N_14559,N_14674);
or U14776 (N_14776,N_14571,N_14587);
nand U14777 (N_14777,N_14564,N_14632);
nand U14778 (N_14778,N_14692,N_14627);
xnor U14779 (N_14779,N_14675,N_14640);
and U14780 (N_14780,N_14609,N_14616);
xor U14781 (N_14781,N_14677,N_14581);
xnor U14782 (N_14782,N_14602,N_14616);
nand U14783 (N_14783,N_14613,N_14623);
xnor U14784 (N_14784,N_14598,N_14656);
and U14785 (N_14785,N_14572,N_14668);
nand U14786 (N_14786,N_14674,N_14660);
xnor U14787 (N_14787,N_14559,N_14607);
and U14788 (N_14788,N_14678,N_14585);
and U14789 (N_14789,N_14550,N_14659);
nor U14790 (N_14790,N_14607,N_14599);
and U14791 (N_14791,N_14586,N_14622);
xor U14792 (N_14792,N_14637,N_14661);
and U14793 (N_14793,N_14645,N_14561);
nor U14794 (N_14794,N_14616,N_14684);
xnor U14795 (N_14795,N_14673,N_14550);
nor U14796 (N_14796,N_14647,N_14624);
and U14797 (N_14797,N_14692,N_14687);
nor U14798 (N_14798,N_14668,N_14593);
or U14799 (N_14799,N_14567,N_14648);
and U14800 (N_14800,N_14671,N_14584);
xor U14801 (N_14801,N_14585,N_14667);
and U14802 (N_14802,N_14680,N_14647);
nor U14803 (N_14803,N_14578,N_14606);
or U14804 (N_14804,N_14648,N_14566);
and U14805 (N_14805,N_14597,N_14698);
xor U14806 (N_14806,N_14584,N_14551);
xor U14807 (N_14807,N_14610,N_14593);
and U14808 (N_14808,N_14571,N_14579);
nor U14809 (N_14809,N_14681,N_14586);
and U14810 (N_14810,N_14617,N_14677);
nand U14811 (N_14811,N_14587,N_14662);
and U14812 (N_14812,N_14553,N_14665);
nor U14813 (N_14813,N_14639,N_14665);
nor U14814 (N_14814,N_14596,N_14612);
nand U14815 (N_14815,N_14553,N_14593);
or U14816 (N_14816,N_14643,N_14595);
nand U14817 (N_14817,N_14584,N_14624);
xor U14818 (N_14818,N_14619,N_14570);
or U14819 (N_14819,N_14557,N_14602);
xor U14820 (N_14820,N_14659,N_14645);
nor U14821 (N_14821,N_14663,N_14637);
xor U14822 (N_14822,N_14565,N_14589);
xnor U14823 (N_14823,N_14664,N_14623);
nand U14824 (N_14824,N_14632,N_14667);
nor U14825 (N_14825,N_14559,N_14637);
nor U14826 (N_14826,N_14651,N_14553);
nor U14827 (N_14827,N_14560,N_14655);
nand U14828 (N_14828,N_14650,N_14567);
or U14829 (N_14829,N_14635,N_14626);
and U14830 (N_14830,N_14674,N_14643);
and U14831 (N_14831,N_14665,N_14628);
or U14832 (N_14832,N_14593,N_14608);
nand U14833 (N_14833,N_14615,N_14656);
nand U14834 (N_14834,N_14655,N_14581);
and U14835 (N_14835,N_14670,N_14671);
or U14836 (N_14836,N_14693,N_14618);
nor U14837 (N_14837,N_14688,N_14671);
nor U14838 (N_14838,N_14672,N_14644);
xor U14839 (N_14839,N_14619,N_14586);
nand U14840 (N_14840,N_14682,N_14606);
or U14841 (N_14841,N_14644,N_14665);
and U14842 (N_14842,N_14699,N_14562);
nor U14843 (N_14843,N_14658,N_14652);
or U14844 (N_14844,N_14660,N_14665);
nor U14845 (N_14845,N_14588,N_14592);
nand U14846 (N_14846,N_14607,N_14623);
nand U14847 (N_14847,N_14677,N_14553);
or U14848 (N_14848,N_14656,N_14667);
xor U14849 (N_14849,N_14644,N_14680);
nand U14850 (N_14850,N_14790,N_14832);
or U14851 (N_14851,N_14802,N_14711);
nor U14852 (N_14852,N_14710,N_14743);
xnor U14853 (N_14853,N_14823,N_14846);
nand U14854 (N_14854,N_14749,N_14700);
and U14855 (N_14855,N_14754,N_14767);
nand U14856 (N_14856,N_14764,N_14702);
and U14857 (N_14857,N_14782,N_14740);
xor U14858 (N_14858,N_14715,N_14812);
and U14859 (N_14859,N_14733,N_14789);
xnor U14860 (N_14860,N_14706,N_14713);
xnor U14861 (N_14861,N_14848,N_14744);
and U14862 (N_14862,N_14813,N_14796);
nand U14863 (N_14863,N_14742,N_14801);
xor U14864 (N_14864,N_14709,N_14800);
xnor U14865 (N_14865,N_14772,N_14721);
nor U14866 (N_14866,N_14758,N_14815);
xnor U14867 (N_14867,N_14716,N_14807);
or U14868 (N_14868,N_14818,N_14824);
or U14869 (N_14869,N_14774,N_14842);
xor U14870 (N_14870,N_14745,N_14834);
and U14871 (N_14871,N_14722,N_14791);
or U14872 (N_14872,N_14762,N_14830);
and U14873 (N_14873,N_14819,N_14712);
xor U14874 (N_14874,N_14811,N_14732);
and U14875 (N_14875,N_14746,N_14769);
nor U14876 (N_14876,N_14776,N_14816);
nor U14877 (N_14877,N_14720,N_14844);
and U14878 (N_14878,N_14707,N_14838);
xor U14879 (N_14879,N_14792,N_14755);
nor U14880 (N_14880,N_14752,N_14788);
xnor U14881 (N_14881,N_14831,N_14836);
xnor U14882 (N_14882,N_14747,N_14804);
and U14883 (N_14883,N_14775,N_14741);
or U14884 (N_14884,N_14765,N_14773);
and U14885 (N_14885,N_14717,N_14771);
and U14886 (N_14886,N_14793,N_14703);
nor U14887 (N_14887,N_14817,N_14763);
or U14888 (N_14888,N_14806,N_14794);
or U14889 (N_14889,N_14777,N_14739);
xnor U14890 (N_14890,N_14839,N_14704);
nand U14891 (N_14891,N_14840,N_14843);
nor U14892 (N_14892,N_14829,N_14701);
xnor U14893 (N_14893,N_14736,N_14761);
and U14894 (N_14894,N_14705,N_14833);
and U14895 (N_14895,N_14785,N_14750);
nand U14896 (N_14896,N_14734,N_14735);
or U14897 (N_14897,N_14738,N_14827);
and U14898 (N_14898,N_14726,N_14799);
and U14899 (N_14899,N_14847,N_14759);
and U14900 (N_14900,N_14837,N_14810);
nand U14901 (N_14901,N_14727,N_14748);
or U14902 (N_14902,N_14753,N_14841);
nand U14903 (N_14903,N_14809,N_14786);
nand U14904 (N_14904,N_14768,N_14784);
nor U14905 (N_14905,N_14787,N_14730);
nor U14906 (N_14906,N_14714,N_14825);
or U14907 (N_14907,N_14724,N_14783);
xor U14908 (N_14908,N_14737,N_14820);
xor U14909 (N_14909,N_14756,N_14797);
or U14910 (N_14910,N_14719,N_14731);
and U14911 (N_14911,N_14808,N_14795);
nor U14912 (N_14912,N_14778,N_14828);
nor U14913 (N_14913,N_14781,N_14803);
and U14914 (N_14914,N_14822,N_14849);
nor U14915 (N_14915,N_14729,N_14780);
nor U14916 (N_14916,N_14798,N_14760);
and U14917 (N_14917,N_14728,N_14805);
xor U14918 (N_14918,N_14766,N_14708);
or U14919 (N_14919,N_14751,N_14757);
or U14920 (N_14920,N_14718,N_14725);
nand U14921 (N_14921,N_14770,N_14826);
nor U14922 (N_14922,N_14835,N_14723);
nor U14923 (N_14923,N_14821,N_14814);
and U14924 (N_14924,N_14845,N_14779);
and U14925 (N_14925,N_14781,N_14778);
xor U14926 (N_14926,N_14806,N_14732);
and U14927 (N_14927,N_14729,N_14811);
or U14928 (N_14928,N_14796,N_14799);
and U14929 (N_14929,N_14769,N_14800);
or U14930 (N_14930,N_14838,N_14732);
and U14931 (N_14931,N_14843,N_14816);
nand U14932 (N_14932,N_14835,N_14798);
and U14933 (N_14933,N_14743,N_14793);
or U14934 (N_14934,N_14800,N_14819);
and U14935 (N_14935,N_14717,N_14772);
xnor U14936 (N_14936,N_14820,N_14726);
xor U14937 (N_14937,N_14793,N_14800);
and U14938 (N_14938,N_14704,N_14814);
or U14939 (N_14939,N_14712,N_14784);
nor U14940 (N_14940,N_14731,N_14710);
and U14941 (N_14941,N_14715,N_14831);
or U14942 (N_14942,N_14744,N_14787);
xnor U14943 (N_14943,N_14839,N_14715);
or U14944 (N_14944,N_14770,N_14761);
nand U14945 (N_14945,N_14791,N_14701);
nand U14946 (N_14946,N_14779,N_14758);
and U14947 (N_14947,N_14736,N_14796);
or U14948 (N_14948,N_14727,N_14781);
nor U14949 (N_14949,N_14711,N_14793);
xor U14950 (N_14950,N_14804,N_14828);
or U14951 (N_14951,N_14713,N_14781);
or U14952 (N_14952,N_14807,N_14749);
or U14953 (N_14953,N_14848,N_14766);
nor U14954 (N_14954,N_14758,N_14710);
or U14955 (N_14955,N_14824,N_14833);
nor U14956 (N_14956,N_14817,N_14772);
xor U14957 (N_14957,N_14774,N_14727);
nor U14958 (N_14958,N_14719,N_14832);
nor U14959 (N_14959,N_14712,N_14740);
nand U14960 (N_14960,N_14753,N_14803);
nand U14961 (N_14961,N_14802,N_14760);
nor U14962 (N_14962,N_14796,N_14809);
nand U14963 (N_14963,N_14748,N_14773);
nor U14964 (N_14964,N_14825,N_14719);
nand U14965 (N_14965,N_14790,N_14711);
and U14966 (N_14966,N_14806,N_14799);
nand U14967 (N_14967,N_14813,N_14785);
and U14968 (N_14968,N_14764,N_14716);
nor U14969 (N_14969,N_14825,N_14780);
nand U14970 (N_14970,N_14834,N_14845);
and U14971 (N_14971,N_14715,N_14704);
xnor U14972 (N_14972,N_14733,N_14744);
or U14973 (N_14973,N_14715,N_14769);
nor U14974 (N_14974,N_14758,N_14754);
nor U14975 (N_14975,N_14700,N_14848);
nor U14976 (N_14976,N_14739,N_14751);
nand U14977 (N_14977,N_14700,N_14767);
or U14978 (N_14978,N_14780,N_14760);
nor U14979 (N_14979,N_14722,N_14817);
xnor U14980 (N_14980,N_14710,N_14725);
or U14981 (N_14981,N_14790,N_14723);
nand U14982 (N_14982,N_14725,N_14787);
or U14983 (N_14983,N_14778,N_14800);
nor U14984 (N_14984,N_14706,N_14835);
or U14985 (N_14985,N_14847,N_14746);
nand U14986 (N_14986,N_14713,N_14757);
xnor U14987 (N_14987,N_14734,N_14808);
nor U14988 (N_14988,N_14809,N_14727);
xor U14989 (N_14989,N_14749,N_14801);
nor U14990 (N_14990,N_14785,N_14718);
nand U14991 (N_14991,N_14708,N_14715);
or U14992 (N_14992,N_14703,N_14710);
and U14993 (N_14993,N_14836,N_14705);
or U14994 (N_14994,N_14845,N_14726);
and U14995 (N_14995,N_14816,N_14728);
xor U14996 (N_14996,N_14790,N_14712);
nand U14997 (N_14997,N_14842,N_14738);
and U14998 (N_14998,N_14788,N_14817);
and U14999 (N_14999,N_14769,N_14710);
nor UO_0 (O_0,N_14878,N_14900);
nor UO_1 (O_1,N_14951,N_14963);
nor UO_2 (O_2,N_14898,N_14988);
and UO_3 (O_3,N_14999,N_14907);
xnor UO_4 (O_4,N_14905,N_14984);
or UO_5 (O_5,N_14978,N_14927);
nor UO_6 (O_6,N_14941,N_14889);
nor UO_7 (O_7,N_14993,N_14996);
nand UO_8 (O_8,N_14949,N_14950);
nand UO_9 (O_9,N_14852,N_14880);
nand UO_10 (O_10,N_14961,N_14934);
or UO_11 (O_11,N_14915,N_14892);
nor UO_12 (O_12,N_14863,N_14954);
nor UO_13 (O_13,N_14874,N_14860);
nor UO_14 (O_14,N_14901,N_14980);
xor UO_15 (O_15,N_14896,N_14899);
nor UO_16 (O_16,N_14955,N_14912);
and UO_17 (O_17,N_14973,N_14919);
or UO_18 (O_18,N_14997,N_14937);
xnor UO_19 (O_19,N_14931,N_14855);
nand UO_20 (O_20,N_14903,N_14953);
nand UO_21 (O_21,N_14959,N_14992);
nor UO_22 (O_22,N_14886,N_14872);
nand UO_23 (O_23,N_14853,N_14858);
and UO_24 (O_24,N_14940,N_14917);
xnor UO_25 (O_25,N_14938,N_14987);
nand UO_26 (O_26,N_14936,N_14869);
xor UO_27 (O_27,N_14883,N_14884);
nand UO_28 (O_28,N_14902,N_14876);
or UO_29 (O_29,N_14966,N_14945);
nand UO_30 (O_30,N_14962,N_14910);
nand UO_31 (O_31,N_14995,N_14894);
xnor UO_32 (O_32,N_14879,N_14967);
and UO_33 (O_33,N_14991,N_14908);
nor UO_34 (O_34,N_14911,N_14933);
or UO_35 (O_35,N_14952,N_14969);
xor UO_36 (O_36,N_14965,N_14970);
nor UO_37 (O_37,N_14922,N_14975);
or UO_38 (O_38,N_14890,N_14882);
or UO_39 (O_39,N_14976,N_14971);
nor UO_40 (O_40,N_14923,N_14887);
nor UO_41 (O_41,N_14865,N_14946);
and UO_42 (O_42,N_14918,N_14960);
or UO_43 (O_43,N_14968,N_14928);
nand UO_44 (O_44,N_14875,N_14989);
nor UO_45 (O_45,N_14861,N_14943);
nand UO_46 (O_46,N_14930,N_14870);
or UO_47 (O_47,N_14888,N_14981);
nor UO_48 (O_48,N_14924,N_14998);
nor UO_49 (O_49,N_14885,N_14916);
xnor UO_50 (O_50,N_14921,N_14873);
nand UO_51 (O_51,N_14850,N_14914);
or UO_52 (O_52,N_14926,N_14895);
nand UO_53 (O_53,N_14957,N_14897);
or UO_54 (O_54,N_14944,N_14877);
nor UO_55 (O_55,N_14904,N_14868);
xor UO_56 (O_56,N_14956,N_14851);
nor UO_57 (O_57,N_14866,N_14925);
or UO_58 (O_58,N_14979,N_14986);
nand UO_59 (O_59,N_14909,N_14948);
and UO_60 (O_60,N_14871,N_14862);
nor UO_61 (O_61,N_14854,N_14985);
nand UO_62 (O_62,N_14994,N_14920);
nor UO_63 (O_63,N_14891,N_14935);
xnor UO_64 (O_64,N_14881,N_14939);
and UO_65 (O_65,N_14974,N_14857);
xor UO_66 (O_66,N_14983,N_14942);
or UO_67 (O_67,N_14972,N_14864);
nor UO_68 (O_68,N_14990,N_14977);
nor UO_69 (O_69,N_14964,N_14906);
nand UO_70 (O_70,N_14982,N_14932);
or UO_71 (O_71,N_14958,N_14913);
xor UO_72 (O_72,N_14856,N_14893);
or UO_73 (O_73,N_14929,N_14867);
nand UO_74 (O_74,N_14859,N_14947);
or UO_75 (O_75,N_14868,N_14898);
and UO_76 (O_76,N_14977,N_14880);
nand UO_77 (O_77,N_14905,N_14928);
nor UO_78 (O_78,N_14864,N_14917);
and UO_79 (O_79,N_14934,N_14873);
or UO_80 (O_80,N_14877,N_14975);
xor UO_81 (O_81,N_14981,N_14993);
xor UO_82 (O_82,N_14904,N_14981);
and UO_83 (O_83,N_14883,N_14854);
xor UO_84 (O_84,N_14868,N_14963);
or UO_85 (O_85,N_14907,N_14986);
and UO_86 (O_86,N_14910,N_14868);
nor UO_87 (O_87,N_14885,N_14943);
xor UO_88 (O_88,N_14882,N_14919);
and UO_89 (O_89,N_14890,N_14881);
xor UO_90 (O_90,N_14877,N_14903);
nand UO_91 (O_91,N_14998,N_14921);
or UO_92 (O_92,N_14898,N_14968);
nor UO_93 (O_93,N_14996,N_14897);
nand UO_94 (O_94,N_14908,N_14933);
nand UO_95 (O_95,N_14940,N_14986);
xnor UO_96 (O_96,N_14865,N_14964);
nor UO_97 (O_97,N_14975,N_14945);
nand UO_98 (O_98,N_14857,N_14947);
xnor UO_99 (O_99,N_14856,N_14978);
and UO_100 (O_100,N_14942,N_14868);
xnor UO_101 (O_101,N_14964,N_14873);
nand UO_102 (O_102,N_14906,N_14934);
xor UO_103 (O_103,N_14904,N_14854);
and UO_104 (O_104,N_14981,N_14909);
nor UO_105 (O_105,N_14880,N_14909);
or UO_106 (O_106,N_14886,N_14987);
xnor UO_107 (O_107,N_14863,N_14982);
nor UO_108 (O_108,N_14850,N_14930);
nand UO_109 (O_109,N_14997,N_14962);
xor UO_110 (O_110,N_14935,N_14852);
and UO_111 (O_111,N_14875,N_14871);
nand UO_112 (O_112,N_14926,N_14908);
or UO_113 (O_113,N_14915,N_14890);
and UO_114 (O_114,N_14979,N_14861);
xor UO_115 (O_115,N_14891,N_14983);
or UO_116 (O_116,N_14867,N_14988);
and UO_117 (O_117,N_14895,N_14878);
or UO_118 (O_118,N_14935,N_14893);
and UO_119 (O_119,N_14874,N_14963);
xnor UO_120 (O_120,N_14973,N_14980);
and UO_121 (O_121,N_14968,N_14911);
xor UO_122 (O_122,N_14914,N_14879);
nand UO_123 (O_123,N_14856,N_14891);
nand UO_124 (O_124,N_14901,N_14994);
or UO_125 (O_125,N_14899,N_14953);
nor UO_126 (O_126,N_14933,N_14945);
nand UO_127 (O_127,N_14971,N_14883);
or UO_128 (O_128,N_14890,N_14898);
or UO_129 (O_129,N_14869,N_14985);
and UO_130 (O_130,N_14867,N_14986);
nand UO_131 (O_131,N_14917,N_14997);
nand UO_132 (O_132,N_14994,N_14912);
and UO_133 (O_133,N_14857,N_14907);
nand UO_134 (O_134,N_14942,N_14854);
nor UO_135 (O_135,N_14892,N_14978);
xnor UO_136 (O_136,N_14966,N_14937);
or UO_137 (O_137,N_14850,N_14891);
and UO_138 (O_138,N_14996,N_14952);
nand UO_139 (O_139,N_14999,N_14878);
and UO_140 (O_140,N_14928,N_14991);
xor UO_141 (O_141,N_14921,N_14891);
and UO_142 (O_142,N_14870,N_14980);
or UO_143 (O_143,N_14966,N_14855);
xnor UO_144 (O_144,N_14892,N_14914);
nor UO_145 (O_145,N_14854,N_14874);
or UO_146 (O_146,N_14885,N_14850);
xor UO_147 (O_147,N_14985,N_14993);
and UO_148 (O_148,N_14868,N_14941);
or UO_149 (O_149,N_14952,N_14877);
nor UO_150 (O_150,N_14862,N_14913);
nor UO_151 (O_151,N_14876,N_14925);
nand UO_152 (O_152,N_14994,N_14919);
nand UO_153 (O_153,N_14863,N_14903);
or UO_154 (O_154,N_14926,N_14970);
or UO_155 (O_155,N_14968,N_14887);
nand UO_156 (O_156,N_14875,N_14920);
xor UO_157 (O_157,N_14852,N_14927);
nand UO_158 (O_158,N_14923,N_14914);
xnor UO_159 (O_159,N_14957,N_14960);
nand UO_160 (O_160,N_14892,N_14883);
and UO_161 (O_161,N_14964,N_14978);
or UO_162 (O_162,N_14894,N_14906);
xnor UO_163 (O_163,N_14981,N_14863);
nand UO_164 (O_164,N_14931,N_14960);
and UO_165 (O_165,N_14972,N_14992);
nand UO_166 (O_166,N_14896,N_14922);
nand UO_167 (O_167,N_14977,N_14885);
xnor UO_168 (O_168,N_14998,N_14980);
and UO_169 (O_169,N_14984,N_14891);
and UO_170 (O_170,N_14856,N_14976);
or UO_171 (O_171,N_14894,N_14959);
nor UO_172 (O_172,N_14956,N_14891);
xor UO_173 (O_173,N_14988,N_14876);
or UO_174 (O_174,N_14917,N_14978);
nor UO_175 (O_175,N_14934,N_14889);
nand UO_176 (O_176,N_14851,N_14939);
and UO_177 (O_177,N_14871,N_14859);
xnor UO_178 (O_178,N_14872,N_14942);
nand UO_179 (O_179,N_14871,N_14883);
xor UO_180 (O_180,N_14869,N_14906);
nand UO_181 (O_181,N_14955,N_14943);
xnor UO_182 (O_182,N_14935,N_14926);
nor UO_183 (O_183,N_14968,N_14875);
and UO_184 (O_184,N_14991,N_14929);
xor UO_185 (O_185,N_14991,N_14857);
or UO_186 (O_186,N_14932,N_14995);
nor UO_187 (O_187,N_14934,N_14898);
nor UO_188 (O_188,N_14977,N_14985);
xor UO_189 (O_189,N_14880,N_14989);
xor UO_190 (O_190,N_14927,N_14985);
xnor UO_191 (O_191,N_14936,N_14883);
and UO_192 (O_192,N_14888,N_14924);
nor UO_193 (O_193,N_14897,N_14980);
or UO_194 (O_194,N_14909,N_14941);
nand UO_195 (O_195,N_14955,N_14924);
nor UO_196 (O_196,N_14969,N_14855);
nor UO_197 (O_197,N_14915,N_14965);
xor UO_198 (O_198,N_14916,N_14876);
nor UO_199 (O_199,N_14873,N_14859);
and UO_200 (O_200,N_14928,N_14889);
xnor UO_201 (O_201,N_14957,N_14994);
xor UO_202 (O_202,N_14916,N_14865);
and UO_203 (O_203,N_14880,N_14913);
xnor UO_204 (O_204,N_14957,N_14854);
or UO_205 (O_205,N_14943,N_14904);
or UO_206 (O_206,N_14873,N_14943);
xnor UO_207 (O_207,N_14943,N_14985);
xor UO_208 (O_208,N_14880,N_14988);
xor UO_209 (O_209,N_14910,N_14951);
nor UO_210 (O_210,N_14903,N_14993);
xor UO_211 (O_211,N_14984,N_14909);
xnor UO_212 (O_212,N_14900,N_14874);
or UO_213 (O_213,N_14912,N_14964);
xor UO_214 (O_214,N_14862,N_14915);
and UO_215 (O_215,N_14886,N_14981);
or UO_216 (O_216,N_14855,N_14935);
and UO_217 (O_217,N_14884,N_14854);
and UO_218 (O_218,N_14931,N_14934);
or UO_219 (O_219,N_14874,N_14896);
nand UO_220 (O_220,N_14973,N_14850);
nand UO_221 (O_221,N_14996,N_14989);
nand UO_222 (O_222,N_14902,N_14907);
and UO_223 (O_223,N_14984,N_14907);
or UO_224 (O_224,N_14943,N_14966);
and UO_225 (O_225,N_14971,N_14899);
or UO_226 (O_226,N_14959,N_14900);
or UO_227 (O_227,N_14876,N_14989);
nand UO_228 (O_228,N_14861,N_14970);
nand UO_229 (O_229,N_14992,N_14958);
xnor UO_230 (O_230,N_14992,N_14893);
nand UO_231 (O_231,N_14999,N_14882);
xor UO_232 (O_232,N_14880,N_14889);
or UO_233 (O_233,N_14912,N_14882);
xnor UO_234 (O_234,N_14886,N_14889);
or UO_235 (O_235,N_14968,N_14958);
or UO_236 (O_236,N_14854,N_14851);
nor UO_237 (O_237,N_14992,N_14910);
and UO_238 (O_238,N_14955,N_14882);
nor UO_239 (O_239,N_14977,N_14949);
nand UO_240 (O_240,N_14957,N_14988);
or UO_241 (O_241,N_14855,N_14915);
nand UO_242 (O_242,N_14875,N_14919);
nor UO_243 (O_243,N_14858,N_14889);
or UO_244 (O_244,N_14991,N_14956);
nor UO_245 (O_245,N_14934,N_14913);
nand UO_246 (O_246,N_14889,N_14856);
and UO_247 (O_247,N_14867,N_14938);
nor UO_248 (O_248,N_14964,N_14887);
and UO_249 (O_249,N_14876,N_14986);
nor UO_250 (O_250,N_14962,N_14918);
nor UO_251 (O_251,N_14978,N_14919);
or UO_252 (O_252,N_14946,N_14869);
nor UO_253 (O_253,N_14909,N_14983);
nand UO_254 (O_254,N_14993,N_14923);
nor UO_255 (O_255,N_14997,N_14866);
or UO_256 (O_256,N_14877,N_14886);
xor UO_257 (O_257,N_14863,N_14907);
and UO_258 (O_258,N_14892,N_14975);
or UO_259 (O_259,N_14881,N_14851);
and UO_260 (O_260,N_14983,N_14981);
and UO_261 (O_261,N_14972,N_14862);
nor UO_262 (O_262,N_14936,N_14975);
nor UO_263 (O_263,N_14885,N_14927);
nand UO_264 (O_264,N_14971,N_14993);
nand UO_265 (O_265,N_14913,N_14909);
xnor UO_266 (O_266,N_14966,N_14993);
and UO_267 (O_267,N_14928,N_14945);
xor UO_268 (O_268,N_14873,N_14929);
nor UO_269 (O_269,N_14933,N_14869);
nor UO_270 (O_270,N_14996,N_14885);
or UO_271 (O_271,N_14902,N_14851);
or UO_272 (O_272,N_14952,N_14973);
nand UO_273 (O_273,N_14921,N_14904);
nand UO_274 (O_274,N_14977,N_14855);
xor UO_275 (O_275,N_14855,N_14993);
nand UO_276 (O_276,N_14939,N_14858);
xor UO_277 (O_277,N_14912,N_14982);
nand UO_278 (O_278,N_14869,N_14892);
or UO_279 (O_279,N_14943,N_14880);
nand UO_280 (O_280,N_14904,N_14923);
or UO_281 (O_281,N_14939,N_14934);
nor UO_282 (O_282,N_14975,N_14871);
nor UO_283 (O_283,N_14895,N_14853);
and UO_284 (O_284,N_14896,N_14986);
nor UO_285 (O_285,N_14854,N_14876);
xnor UO_286 (O_286,N_14939,N_14992);
xnor UO_287 (O_287,N_14945,N_14857);
xor UO_288 (O_288,N_14926,N_14955);
xor UO_289 (O_289,N_14894,N_14853);
nand UO_290 (O_290,N_14979,N_14941);
xnor UO_291 (O_291,N_14860,N_14876);
xnor UO_292 (O_292,N_14978,N_14990);
and UO_293 (O_293,N_14854,N_14893);
xnor UO_294 (O_294,N_14874,N_14911);
xor UO_295 (O_295,N_14907,N_14971);
nand UO_296 (O_296,N_14851,N_14862);
nand UO_297 (O_297,N_14883,N_14979);
and UO_298 (O_298,N_14955,N_14992);
or UO_299 (O_299,N_14854,N_14873);
nand UO_300 (O_300,N_14916,N_14948);
or UO_301 (O_301,N_14887,N_14895);
or UO_302 (O_302,N_14892,N_14852);
nand UO_303 (O_303,N_14859,N_14882);
nand UO_304 (O_304,N_14895,N_14894);
nor UO_305 (O_305,N_14924,N_14946);
or UO_306 (O_306,N_14903,N_14852);
or UO_307 (O_307,N_14965,N_14926);
nand UO_308 (O_308,N_14987,N_14856);
or UO_309 (O_309,N_14948,N_14954);
or UO_310 (O_310,N_14886,N_14928);
or UO_311 (O_311,N_14933,N_14893);
xor UO_312 (O_312,N_14933,N_14974);
nor UO_313 (O_313,N_14874,N_14920);
and UO_314 (O_314,N_14931,N_14917);
or UO_315 (O_315,N_14994,N_14974);
and UO_316 (O_316,N_14986,N_14994);
or UO_317 (O_317,N_14886,N_14929);
xnor UO_318 (O_318,N_14962,N_14917);
xor UO_319 (O_319,N_14929,N_14866);
nand UO_320 (O_320,N_14957,N_14859);
or UO_321 (O_321,N_14922,N_14935);
or UO_322 (O_322,N_14951,N_14907);
or UO_323 (O_323,N_14873,N_14979);
and UO_324 (O_324,N_14967,N_14936);
nor UO_325 (O_325,N_14941,N_14958);
nor UO_326 (O_326,N_14885,N_14990);
or UO_327 (O_327,N_14940,N_14901);
and UO_328 (O_328,N_14879,N_14921);
or UO_329 (O_329,N_14869,N_14880);
nand UO_330 (O_330,N_14967,N_14917);
and UO_331 (O_331,N_14996,N_14971);
xor UO_332 (O_332,N_14943,N_14905);
nand UO_333 (O_333,N_14977,N_14936);
nor UO_334 (O_334,N_14927,N_14859);
xnor UO_335 (O_335,N_14993,N_14949);
and UO_336 (O_336,N_14924,N_14970);
nor UO_337 (O_337,N_14854,N_14902);
xnor UO_338 (O_338,N_14921,N_14983);
xnor UO_339 (O_339,N_14913,N_14964);
nor UO_340 (O_340,N_14931,N_14990);
nand UO_341 (O_341,N_14915,N_14894);
xor UO_342 (O_342,N_14873,N_14858);
and UO_343 (O_343,N_14992,N_14936);
nand UO_344 (O_344,N_14923,N_14958);
nand UO_345 (O_345,N_14854,N_14892);
xor UO_346 (O_346,N_14914,N_14896);
nand UO_347 (O_347,N_14968,N_14871);
or UO_348 (O_348,N_14872,N_14978);
or UO_349 (O_349,N_14893,N_14984);
nand UO_350 (O_350,N_14969,N_14947);
nand UO_351 (O_351,N_14986,N_14875);
and UO_352 (O_352,N_14904,N_14880);
or UO_353 (O_353,N_14913,N_14916);
nand UO_354 (O_354,N_14937,N_14887);
and UO_355 (O_355,N_14933,N_14962);
or UO_356 (O_356,N_14890,N_14985);
nand UO_357 (O_357,N_14875,N_14911);
xnor UO_358 (O_358,N_14907,N_14988);
nor UO_359 (O_359,N_14915,N_14959);
xor UO_360 (O_360,N_14947,N_14893);
xnor UO_361 (O_361,N_14864,N_14936);
or UO_362 (O_362,N_14902,N_14893);
nor UO_363 (O_363,N_14954,N_14865);
xnor UO_364 (O_364,N_14983,N_14900);
xnor UO_365 (O_365,N_14998,N_14984);
and UO_366 (O_366,N_14938,N_14976);
xnor UO_367 (O_367,N_14992,N_14853);
nor UO_368 (O_368,N_14953,N_14906);
nor UO_369 (O_369,N_14982,N_14946);
or UO_370 (O_370,N_14954,N_14952);
nor UO_371 (O_371,N_14921,N_14917);
or UO_372 (O_372,N_14925,N_14889);
or UO_373 (O_373,N_14972,N_14976);
nand UO_374 (O_374,N_14982,N_14936);
nand UO_375 (O_375,N_14953,N_14885);
xor UO_376 (O_376,N_14851,N_14927);
or UO_377 (O_377,N_14947,N_14942);
nor UO_378 (O_378,N_14866,N_14909);
nand UO_379 (O_379,N_14905,N_14858);
and UO_380 (O_380,N_14895,N_14919);
nand UO_381 (O_381,N_14984,N_14937);
or UO_382 (O_382,N_14959,N_14877);
and UO_383 (O_383,N_14897,N_14925);
and UO_384 (O_384,N_14963,N_14929);
or UO_385 (O_385,N_14959,N_14972);
xor UO_386 (O_386,N_14958,N_14880);
nand UO_387 (O_387,N_14971,N_14938);
nor UO_388 (O_388,N_14973,N_14886);
and UO_389 (O_389,N_14916,N_14923);
nor UO_390 (O_390,N_14948,N_14962);
or UO_391 (O_391,N_14864,N_14858);
nand UO_392 (O_392,N_14927,N_14944);
xnor UO_393 (O_393,N_14861,N_14974);
nand UO_394 (O_394,N_14862,N_14996);
or UO_395 (O_395,N_14958,N_14904);
nor UO_396 (O_396,N_14950,N_14896);
nand UO_397 (O_397,N_14855,N_14897);
nand UO_398 (O_398,N_14872,N_14975);
xor UO_399 (O_399,N_14909,N_14929);
or UO_400 (O_400,N_14899,N_14928);
or UO_401 (O_401,N_14858,N_14898);
xnor UO_402 (O_402,N_14921,N_14996);
and UO_403 (O_403,N_14883,N_14943);
nor UO_404 (O_404,N_14951,N_14896);
and UO_405 (O_405,N_14908,N_14900);
xnor UO_406 (O_406,N_14963,N_14968);
nor UO_407 (O_407,N_14883,N_14925);
xnor UO_408 (O_408,N_14994,N_14855);
xor UO_409 (O_409,N_14962,N_14981);
nand UO_410 (O_410,N_14985,N_14907);
nand UO_411 (O_411,N_14855,N_14948);
and UO_412 (O_412,N_14896,N_14898);
or UO_413 (O_413,N_14920,N_14982);
xnor UO_414 (O_414,N_14867,N_14918);
and UO_415 (O_415,N_14864,N_14976);
xnor UO_416 (O_416,N_14930,N_14936);
or UO_417 (O_417,N_14974,N_14894);
nand UO_418 (O_418,N_14921,N_14883);
nand UO_419 (O_419,N_14911,N_14854);
nor UO_420 (O_420,N_14912,N_14906);
xnor UO_421 (O_421,N_14908,N_14947);
nand UO_422 (O_422,N_14862,N_14914);
nor UO_423 (O_423,N_14879,N_14894);
nor UO_424 (O_424,N_14880,N_14879);
or UO_425 (O_425,N_14894,N_14992);
nand UO_426 (O_426,N_14967,N_14990);
and UO_427 (O_427,N_14927,N_14918);
xnor UO_428 (O_428,N_14972,N_14950);
nor UO_429 (O_429,N_14994,N_14889);
and UO_430 (O_430,N_14866,N_14891);
or UO_431 (O_431,N_14895,N_14953);
or UO_432 (O_432,N_14859,N_14895);
nand UO_433 (O_433,N_14871,N_14897);
xnor UO_434 (O_434,N_14946,N_14980);
nor UO_435 (O_435,N_14992,N_14914);
nor UO_436 (O_436,N_14963,N_14973);
xor UO_437 (O_437,N_14880,N_14903);
nand UO_438 (O_438,N_14900,N_14996);
nor UO_439 (O_439,N_14927,N_14854);
nor UO_440 (O_440,N_14957,N_14949);
xnor UO_441 (O_441,N_14979,N_14944);
nand UO_442 (O_442,N_14869,N_14950);
nand UO_443 (O_443,N_14900,N_14879);
or UO_444 (O_444,N_14982,N_14985);
or UO_445 (O_445,N_14923,N_14976);
or UO_446 (O_446,N_14977,N_14961);
and UO_447 (O_447,N_14945,N_14953);
and UO_448 (O_448,N_14867,N_14965);
or UO_449 (O_449,N_14939,N_14863);
xor UO_450 (O_450,N_14903,N_14888);
nor UO_451 (O_451,N_14861,N_14972);
xor UO_452 (O_452,N_14864,N_14957);
and UO_453 (O_453,N_14895,N_14976);
xnor UO_454 (O_454,N_14928,N_14907);
nor UO_455 (O_455,N_14968,N_14986);
and UO_456 (O_456,N_14851,N_14867);
or UO_457 (O_457,N_14909,N_14896);
nor UO_458 (O_458,N_14922,N_14909);
and UO_459 (O_459,N_14912,N_14884);
nor UO_460 (O_460,N_14914,N_14858);
nor UO_461 (O_461,N_14888,N_14988);
and UO_462 (O_462,N_14939,N_14903);
nand UO_463 (O_463,N_14925,N_14968);
or UO_464 (O_464,N_14888,N_14969);
xnor UO_465 (O_465,N_14967,N_14974);
nor UO_466 (O_466,N_14907,N_14923);
or UO_467 (O_467,N_14875,N_14892);
or UO_468 (O_468,N_14916,N_14860);
or UO_469 (O_469,N_14969,N_14883);
and UO_470 (O_470,N_14867,N_14896);
and UO_471 (O_471,N_14941,N_14955);
nor UO_472 (O_472,N_14923,N_14929);
xor UO_473 (O_473,N_14912,N_14937);
nand UO_474 (O_474,N_14997,N_14854);
nor UO_475 (O_475,N_14933,N_14999);
and UO_476 (O_476,N_14851,N_14963);
or UO_477 (O_477,N_14922,N_14863);
or UO_478 (O_478,N_14992,N_14908);
nor UO_479 (O_479,N_14878,N_14990);
and UO_480 (O_480,N_14961,N_14974);
or UO_481 (O_481,N_14942,N_14963);
or UO_482 (O_482,N_14974,N_14972);
xor UO_483 (O_483,N_14965,N_14894);
or UO_484 (O_484,N_14982,N_14995);
nand UO_485 (O_485,N_14907,N_14981);
nand UO_486 (O_486,N_14861,N_14866);
and UO_487 (O_487,N_14943,N_14988);
nor UO_488 (O_488,N_14987,N_14970);
nor UO_489 (O_489,N_14944,N_14989);
nor UO_490 (O_490,N_14903,N_14858);
nor UO_491 (O_491,N_14929,N_14948);
nor UO_492 (O_492,N_14978,N_14970);
xnor UO_493 (O_493,N_14871,N_14892);
or UO_494 (O_494,N_14891,N_14962);
and UO_495 (O_495,N_14915,N_14990);
xor UO_496 (O_496,N_14955,N_14938);
nor UO_497 (O_497,N_14995,N_14877);
and UO_498 (O_498,N_14917,N_14876);
nand UO_499 (O_499,N_14872,N_14996);
and UO_500 (O_500,N_14987,N_14931);
or UO_501 (O_501,N_14876,N_14918);
and UO_502 (O_502,N_14896,N_14875);
nor UO_503 (O_503,N_14965,N_14917);
and UO_504 (O_504,N_14870,N_14996);
xor UO_505 (O_505,N_14893,N_14964);
and UO_506 (O_506,N_14915,N_14876);
xnor UO_507 (O_507,N_14998,N_14953);
nand UO_508 (O_508,N_14985,N_14973);
xnor UO_509 (O_509,N_14890,N_14906);
nand UO_510 (O_510,N_14936,N_14889);
nor UO_511 (O_511,N_14913,N_14858);
and UO_512 (O_512,N_14966,N_14958);
or UO_513 (O_513,N_14964,N_14999);
nor UO_514 (O_514,N_14919,N_14893);
nor UO_515 (O_515,N_14894,N_14877);
or UO_516 (O_516,N_14947,N_14894);
nand UO_517 (O_517,N_14948,N_14951);
xor UO_518 (O_518,N_14948,N_14911);
or UO_519 (O_519,N_14907,N_14957);
xnor UO_520 (O_520,N_14981,N_14935);
nand UO_521 (O_521,N_14853,N_14940);
nand UO_522 (O_522,N_14993,N_14872);
or UO_523 (O_523,N_14929,N_14943);
and UO_524 (O_524,N_14859,N_14932);
nand UO_525 (O_525,N_14940,N_14923);
nand UO_526 (O_526,N_14959,N_14999);
nor UO_527 (O_527,N_14973,N_14928);
nand UO_528 (O_528,N_14938,N_14972);
or UO_529 (O_529,N_14963,N_14998);
or UO_530 (O_530,N_14981,N_14953);
nor UO_531 (O_531,N_14880,N_14982);
and UO_532 (O_532,N_14957,N_14932);
and UO_533 (O_533,N_14930,N_14971);
or UO_534 (O_534,N_14954,N_14868);
or UO_535 (O_535,N_14967,N_14873);
xor UO_536 (O_536,N_14928,N_14913);
nor UO_537 (O_537,N_14890,N_14872);
and UO_538 (O_538,N_14960,N_14929);
xor UO_539 (O_539,N_14856,N_14929);
xnor UO_540 (O_540,N_14893,N_14965);
and UO_541 (O_541,N_14859,N_14909);
xor UO_542 (O_542,N_14862,N_14891);
or UO_543 (O_543,N_14946,N_14851);
xnor UO_544 (O_544,N_14915,N_14865);
nand UO_545 (O_545,N_14875,N_14878);
xnor UO_546 (O_546,N_14864,N_14959);
xnor UO_547 (O_547,N_14907,N_14904);
xor UO_548 (O_548,N_14873,N_14956);
xor UO_549 (O_549,N_14851,N_14977);
or UO_550 (O_550,N_14875,N_14982);
nand UO_551 (O_551,N_14988,N_14851);
or UO_552 (O_552,N_14861,N_14855);
or UO_553 (O_553,N_14966,N_14938);
and UO_554 (O_554,N_14932,N_14857);
and UO_555 (O_555,N_14852,N_14992);
xor UO_556 (O_556,N_14904,N_14970);
nor UO_557 (O_557,N_14867,N_14985);
xnor UO_558 (O_558,N_14864,N_14983);
xor UO_559 (O_559,N_14850,N_14857);
xnor UO_560 (O_560,N_14880,N_14885);
xor UO_561 (O_561,N_14888,N_14963);
nor UO_562 (O_562,N_14862,N_14876);
nand UO_563 (O_563,N_14998,N_14905);
xnor UO_564 (O_564,N_14984,N_14942);
or UO_565 (O_565,N_14893,N_14941);
and UO_566 (O_566,N_14905,N_14995);
nor UO_567 (O_567,N_14890,N_14899);
xor UO_568 (O_568,N_14963,N_14904);
xnor UO_569 (O_569,N_14959,N_14880);
xor UO_570 (O_570,N_14990,N_14947);
or UO_571 (O_571,N_14927,N_14926);
or UO_572 (O_572,N_14857,N_14917);
or UO_573 (O_573,N_14960,N_14940);
nand UO_574 (O_574,N_14971,N_14902);
nor UO_575 (O_575,N_14862,N_14859);
nand UO_576 (O_576,N_14998,N_14942);
or UO_577 (O_577,N_14871,N_14960);
and UO_578 (O_578,N_14853,N_14970);
and UO_579 (O_579,N_14881,N_14998);
nor UO_580 (O_580,N_14918,N_14983);
nor UO_581 (O_581,N_14929,N_14885);
nor UO_582 (O_582,N_14913,N_14996);
nand UO_583 (O_583,N_14933,N_14855);
or UO_584 (O_584,N_14916,N_14962);
and UO_585 (O_585,N_14858,N_14881);
or UO_586 (O_586,N_14947,N_14869);
or UO_587 (O_587,N_14988,N_14954);
nor UO_588 (O_588,N_14994,N_14887);
and UO_589 (O_589,N_14854,N_14933);
nor UO_590 (O_590,N_14916,N_14945);
xor UO_591 (O_591,N_14926,N_14853);
nor UO_592 (O_592,N_14859,N_14996);
or UO_593 (O_593,N_14967,N_14973);
or UO_594 (O_594,N_14948,N_14914);
nor UO_595 (O_595,N_14872,N_14958);
and UO_596 (O_596,N_14905,N_14873);
nor UO_597 (O_597,N_14878,N_14876);
nor UO_598 (O_598,N_14956,N_14909);
or UO_599 (O_599,N_14964,N_14968);
xnor UO_600 (O_600,N_14920,N_14989);
nand UO_601 (O_601,N_14860,N_14891);
xor UO_602 (O_602,N_14928,N_14948);
xnor UO_603 (O_603,N_14893,N_14928);
nor UO_604 (O_604,N_14876,N_14947);
nand UO_605 (O_605,N_14996,N_14909);
or UO_606 (O_606,N_14954,N_14858);
nor UO_607 (O_607,N_14963,N_14956);
xnor UO_608 (O_608,N_14919,N_14923);
nand UO_609 (O_609,N_14924,N_14932);
nand UO_610 (O_610,N_14893,N_14914);
nor UO_611 (O_611,N_14863,N_14867);
and UO_612 (O_612,N_14908,N_14982);
or UO_613 (O_613,N_14950,N_14967);
and UO_614 (O_614,N_14884,N_14930);
xor UO_615 (O_615,N_14971,N_14967);
nand UO_616 (O_616,N_14909,N_14927);
and UO_617 (O_617,N_14979,N_14976);
xnor UO_618 (O_618,N_14897,N_14859);
and UO_619 (O_619,N_14934,N_14979);
or UO_620 (O_620,N_14863,N_14947);
nor UO_621 (O_621,N_14950,N_14983);
or UO_622 (O_622,N_14933,N_14991);
nand UO_623 (O_623,N_14891,N_14864);
xnor UO_624 (O_624,N_14980,N_14938);
xnor UO_625 (O_625,N_14887,N_14903);
nand UO_626 (O_626,N_14863,N_14894);
nand UO_627 (O_627,N_14972,N_14966);
nor UO_628 (O_628,N_14971,N_14929);
and UO_629 (O_629,N_14971,N_14903);
xor UO_630 (O_630,N_14958,N_14862);
nor UO_631 (O_631,N_14988,N_14992);
or UO_632 (O_632,N_14892,N_14937);
and UO_633 (O_633,N_14986,N_14982);
and UO_634 (O_634,N_14933,N_14953);
or UO_635 (O_635,N_14981,N_14941);
nor UO_636 (O_636,N_14924,N_14910);
xnor UO_637 (O_637,N_14972,N_14889);
xor UO_638 (O_638,N_14883,N_14951);
and UO_639 (O_639,N_14915,N_14910);
nor UO_640 (O_640,N_14949,N_14964);
or UO_641 (O_641,N_14918,N_14871);
xor UO_642 (O_642,N_14901,N_14974);
or UO_643 (O_643,N_14993,N_14912);
nor UO_644 (O_644,N_14960,N_14994);
and UO_645 (O_645,N_14876,N_14853);
nor UO_646 (O_646,N_14911,N_14940);
nand UO_647 (O_647,N_14942,N_14951);
and UO_648 (O_648,N_14963,N_14859);
and UO_649 (O_649,N_14942,N_14972);
or UO_650 (O_650,N_14862,N_14861);
xor UO_651 (O_651,N_14876,N_14906);
nand UO_652 (O_652,N_14884,N_14915);
or UO_653 (O_653,N_14876,N_14877);
nand UO_654 (O_654,N_14891,N_14942);
or UO_655 (O_655,N_14941,N_14898);
nor UO_656 (O_656,N_14851,N_14959);
xnor UO_657 (O_657,N_14930,N_14861);
nand UO_658 (O_658,N_14979,N_14931);
xnor UO_659 (O_659,N_14963,N_14858);
and UO_660 (O_660,N_14984,N_14904);
nand UO_661 (O_661,N_14944,N_14857);
nor UO_662 (O_662,N_14874,N_14972);
nor UO_663 (O_663,N_14992,N_14904);
nor UO_664 (O_664,N_14995,N_14981);
or UO_665 (O_665,N_14969,N_14990);
nand UO_666 (O_666,N_14952,N_14982);
xor UO_667 (O_667,N_14854,N_14860);
nand UO_668 (O_668,N_14953,N_14880);
nand UO_669 (O_669,N_14990,N_14854);
nand UO_670 (O_670,N_14915,N_14907);
nand UO_671 (O_671,N_14894,N_14916);
nand UO_672 (O_672,N_14979,N_14984);
and UO_673 (O_673,N_14895,N_14955);
nand UO_674 (O_674,N_14874,N_14947);
nand UO_675 (O_675,N_14926,N_14940);
nand UO_676 (O_676,N_14926,N_14915);
xor UO_677 (O_677,N_14893,N_14989);
nor UO_678 (O_678,N_14870,N_14867);
and UO_679 (O_679,N_14886,N_14975);
nor UO_680 (O_680,N_14979,N_14923);
or UO_681 (O_681,N_14903,N_14920);
nand UO_682 (O_682,N_14926,N_14963);
and UO_683 (O_683,N_14859,N_14955);
or UO_684 (O_684,N_14893,N_14954);
nor UO_685 (O_685,N_14989,N_14903);
nand UO_686 (O_686,N_14863,N_14899);
nand UO_687 (O_687,N_14940,N_14962);
and UO_688 (O_688,N_14956,N_14969);
xor UO_689 (O_689,N_14898,N_14916);
xor UO_690 (O_690,N_14995,N_14888);
and UO_691 (O_691,N_14854,N_14962);
xnor UO_692 (O_692,N_14937,N_14954);
or UO_693 (O_693,N_14920,N_14905);
nor UO_694 (O_694,N_14919,N_14914);
xnor UO_695 (O_695,N_14909,N_14861);
and UO_696 (O_696,N_14875,N_14857);
xnor UO_697 (O_697,N_14941,N_14965);
and UO_698 (O_698,N_14900,N_14991);
nand UO_699 (O_699,N_14885,N_14878);
nand UO_700 (O_700,N_14884,N_14996);
and UO_701 (O_701,N_14880,N_14984);
or UO_702 (O_702,N_14967,N_14893);
xor UO_703 (O_703,N_14851,N_14874);
xor UO_704 (O_704,N_14963,N_14876);
nand UO_705 (O_705,N_14895,N_14860);
nand UO_706 (O_706,N_14909,N_14862);
nor UO_707 (O_707,N_14947,N_14860);
nand UO_708 (O_708,N_14906,N_14880);
nand UO_709 (O_709,N_14894,N_14958);
nand UO_710 (O_710,N_14896,N_14968);
or UO_711 (O_711,N_14992,N_14994);
xnor UO_712 (O_712,N_14935,N_14912);
or UO_713 (O_713,N_14913,N_14875);
xnor UO_714 (O_714,N_14929,N_14978);
nor UO_715 (O_715,N_14901,N_14857);
nor UO_716 (O_716,N_14851,N_14955);
nand UO_717 (O_717,N_14914,N_14856);
and UO_718 (O_718,N_14894,N_14988);
or UO_719 (O_719,N_14984,N_14855);
or UO_720 (O_720,N_14924,N_14886);
or UO_721 (O_721,N_14927,N_14891);
nand UO_722 (O_722,N_14921,N_14853);
or UO_723 (O_723,N_14900,N_14961);
xnor UO_724 (O_724,N_14977,N_14971);
xor UO_725 (O_725,N_14985,N_14864);
nor UO_726 (O_726,N_14947,N_14918);
xnor UO_727 (O_727,N_14917,N_14852);
or UO_728 (O_728,N_14865,N_14986);
nor UO_729 (O_729,N_14988,N_14910);
or UO_730 (O_730,N_14908,N_14897);
nor UO_731 (O_731,N_14970,N_14950);
or UO_732 (O_732,N_14899,N_14887);
and UO_733 (O_733,N_14951,N_14923);
and UO_734 (O_734,N_14962,N_14943);
nor UO_735 (O_735,N_14996,N_14945);
nand UO_736 (O_736,N_14987,N_14913);
xnor UO_737 (O_737,N_14896,N_14864);
or UO_738 (O_738,N_14942,N_14911);
and UO_739 (O_739,N_14861,N_14920);
or UO_740 (O_740,N_14929,N_14903);
and UO_741 (O_741,N_14995,N_14946);
or UO_742 (O_742,N_14869,N_14886);
nor UO_743 (O_743,N_14993,N_14889);
or UO_744 (O_744,N_14977,N_14996);
xnor UO_745 (O_745,N_14923,N_14905);
and UO_746 (O_746,N_14971,N_14931);
nand UO_747 (O_747,N_14924,N_14935);
or UO_748 (O_748,N_14894,N_14939);
nor UO_749 (O_749,N_14949,N_14922);
and UO_750 (O_750,N_14903,N_14976);
nand UO_751 (O_751,N_14900,N_14891);
nand UO_752 (O_752,N_14913,N_14936);
nand UO_753 (O_753,N_14965,N_14865);
xor UO_754 (O_754,N_14883,N_14897);
nand UO_755 (O_755,N_14854,N_14930);
and UO_756 (O_756,N_14988,N_14895);
nand UO_757 (O_757,N_14869,N_14887);
nand UO_758 (O_758,N_14907,N_14889);
and UO_759 (O_759,N_14929,N_14858);
xnor UO_760 (O_760,N_14858,N_14906);
nor UO_761 (O_761,N_14897,N_14918);
nor UO_762 (O_762,N_14976,N_14950);
xor UO_763 (O_763,N_14928,N_14917);
xnor UO_764 (O_764,N_14972,N_14920);
and UO_765 (O_765,N_14969,N_14863);
nand UO_766 (O_766,N_14992,N_14951);
nand UO_767 (O_767,N_14886,N_14998);
and UO_768 (O_768,N_14870,N_14874);
and UO_769 (O_769,N_14986,N_14981);
nor UO_770 (O_770,N_14854,N_14888);
xnor UO_771 (O_771,N_14934,N_14947);
nor UO_772 (O_772,N_14968,N_14955);
nor UO_773 (O_773,N_14857,N_14956);
xor UO_774 (O_774,N_14979,N_14851);
nand UO_775 (O_775,N_14856,N_14960);
and UO_776 (O_776,N_14904,N_14991);
or UO_777 (O_777,N_14921,N_14951);
nand UO_778 (O_778,N_14982,N_14931);
xor UO_779 (O_779,N_14869,N_14942);
nor UO_780 (O_780,N_14859,N_14888);
or UO_781 (O_781,N_14931,N_14913);
nand UO_782 (O_782,N_14914,N_14880);
nor UO_783 (O_783,N_14994,N_14876);
nor UO_784 (O_784,N_14950,N_14885);
and UO_785 (O_785,N_14963,N_14966);
nand UO_786 (O_786,N_14882,N_14898);
xor UO_787 (O_787,N_14867,N_14940);
nand UO_788 (O_788,N_14943,N_14881);
and UO_789 (O_789,N_14858,N_14976);
nor UO_790 (O_790,N_14985,N_14992);
or UO_791 (O_791,N_14928,N_14879);
nor UO_792 (O_792,N_14882,N_14939);
nor UO_793 (O_793,N_14899,N_14966);
and UO_794 (O_794,N_14951,N_14913);
or UO_795 (O_795,N_14927,N_14955);
nand UO_796 (O_796,N_14863,N_14980);
nor UO_797 (O_797,N_14909,N_14907);
or UO_798 (O_798,N_14895,N_14992);
nand UO_799 (O_799,N_14950,N_14850);
xor UO_800 (O_800,N_14988,N_14900);
or UO_801 (O_801,N_14936,N_14854);
or UO_802 (O_802,N_14855,N_14945);
or UO_803 (O_803,N_14896,N_14970);
and UO_804 (O_804,N_14965,N_14996);
xor UO_805 (O_805,N_14872,N_14907);
nor UO_806 (O_806,N_14937,N_14933);
and UO_807 (O_807,N_14862,N_14967);
nand UO_808 (O_808,N_14992,N_14983);
xor UO_809 (O_809,N_14945,N_14999);
nor UO_810 (O_810,N_14922,N_14916);
or UO_811 (O_811,N_14882,N_14950);
nand UO_812 (O_812,N_14878,N_14893);
nor UO_813 (O_813,N_14959,N_14927);
and UO_814 (O_814,N_14910,N_14861);
and UO_815 (O_815,N_14933,N_14947);
xor UO_816 (O_816,N_14922,N_14989);
and UO_817 (O_817,N_14944,N_14864);
nor UO_818 (O_818,N_14925,N_14932);
or UO_819 (O_819,N_14872,N_14965);
nand UO_820 (O_820,N_14997,N_14914);
nor UO_821 (O_821,N_14966,N_14871);
xnor UO_822 (O_822,N_14957,N_14917);
and UO_823 (O_823,N_14964,N_14890);
nor UO_824 (O_824,N_14949,N_14868);
and UO_825 (O_825,N_14942,N_14904);
nor UO_826 (O_826,N_14961,N_14903);
xor UO_827 (O_827,N_14931,N_14914);
and UO_828 (O_828,N_14882,N_14960);
or UO_829 (O_829,N_14910,N_14950);
nor UO_830 (O_830,N_14903,N_14927);
or UO_831 (O_831,N_14931,N_14850);
and UO_832 (O_832,N_14899,N_14982);
nand UO_833 (O_833,N_14930,N_14907);
nor UO_834 (O_834,N_14919,N_14928);
xnor UO_835 (O_835,N_14855,N_14989);
or UO_836 (O_836,N_14898,N_14949);
nand UO_837 (O_837,N_14945,N_14889);
and UO_838 (O_838,N_14868,N_14905);
nand UO_839 (O_839,N_14903,N_14900);
nand UO_840 (O_840,N_14973,N_14926);
or UO_841 (O_841,N_14997,N_14987);
xor UO_842 (O_842,N_14980,N_14899);
xnor UO_843 (O_843,N_14989,N_14952);
xnor UO_844 (O_844,N_14884,N_14920);
xor UO_845 (O_845,N_14962,N_14996);
nand UO_846 (O_846,N_14869,N_14937);
or UO_847 (O_847,N_14971,N_14852);
or UO_848 (O_848,N_14878,N_14914);
or UO_849 (O_849,N_14957,N_14979);
and UO_850 (O_850,N_14915,N_14850);
or UO_851 (O_851,N_14927,N_14948);
xnor UO_852 (O_852,N_14873,N_14885);
nand UO_853 (O_853,N_14981,N_14870);
nand UO_854 (O_854,N_14945,N_14939);
xor UO_855 (O_855,N_14939,N_14893);
xor UO_856 (O_856,N_14967,N_14923);
xnor UO_857 (O_857,N_14928,N_14983);
and UO_858 (O_858,N_14915,N_14923);
and UO_859 (O_859,N_14984,N_14881);
nand UO_860 (O_860,N_14939,N_14916);
and UO_861 (O_861,N_14928,N_14993);
and UO_862 (O_862,N_14949,N_14921);
nor UO_863 (O_863,N_14989,N_14871);
nand UO_864 (O_864,N_14922,N_14926);
nand UO_865 (O_865,N_14899,N_14886);
or UO_866 (O_866,N_14867,N_14942);
xor UO_867 (O_867,N_14929,N_14939);
xnor UO_868 (O_868,N_14915,N_14870);
nand UO_869 (O_869,N_14958,N_14907);
and UO_870 (O_870,N_14949,N_14959);
and UO_871 (O_871,N_14958,N_14911);
and UO_872 (O_872,N_14850,N_14985);
and UO_873 (O_873,N_14898,N_14979);
or UO_874 (O_874,N_14991,N_14880);
nand UO_875 (O_875,N_14921,N_14914);
or UO_876 (O_876,N_14914,N_14940);
nand UO_877 (O_877,N_14945,N_14959);
or UO_878 (O_878,N_14904,N_14972);
nand UO_879 (O_879,N_14890,N_14999);
or UO_880 (O_880,N_14950,N_14915);
nor UO_881 (O_881,N_14905,N_14914);
and UO_882 (O_882,N_14996,N_14891);
nand UO_883 (O_883,N_14851,N_14919);
nor UO_884 (O_884,N_14995,N_14859);
or UO_885 (O_885,N_14990,N_14891);
nand UO_886 (O_886,N_14923,N_14982);
or UO_887 (O_887,N_14952,N_14935);
xor UO_888 (O_888,N_14857,N_14876);
and UO_889 (O_889,N_14924,N_14877);
nand UO_890 (O_890,N_14989,N_14869);
xor UO_891 (O_891,N_14921,N_14931);
and UO_892 (O_892,N_14926,N_14856);
nand UO_893 (O_893,N_14954,N_14960);
xor UO_894 (O_894,N_14916,N_14961);
nand UO_895 (O_895,N_14883,N_14905);
and UO_896 (O_896,N_14884,N_14859);
or UO_897 (O_897,N_14950,N_14911);
or UO_898 (O_898,N_14940,N_14948);
nand UO_899 (O_899,N_14968,N_14893);
and UO_900 (O_900,N_14932,N_14918);
nor UO_901 (O_901,N_14964,N_14926);
nor UO_902 (O_902,N_14941,N_14908);
or UO_903 (O_903,N_14905,N_14930);
xor UO_904 (O_904,N_14960,N_14966);
xnor UO_905 (O_905,N_14867,N_14977);
nor UO_906 (O_906,N_14947,N_14954);
and UO_907 (O_907,N_14912,N_14932);
xnor UO_908 (O_908,N_14924,N_14927);
nor UO_909 (O_909,N_14875,N_14958);
nor UO_910 (O_910,N_14880,N_14863);
nand UO_911 (O_911,N_14986,N_14997);
nand UO_912 (O_912,N_14973,N_14959);
and UO_913 (O_913,N_14960,N_14925);
and UO_914 (O_914,N_14944,N_14935);
nor UO_915 (O_915,N_14999,N_14924);
nand UO_916 (O_916,N_14890,N_14967);
xnor UO_917 (O_917,N_14883,N_14850);
or UO_918 (O_918,N_14868,N_14980);
or UO_919 (O_919,N_14924,N_14905);
and UO_920 (O_920,N_14907,N_14921);
or UO_921 (O_921,N_14907,N_14931);
or UO_922 (O_922,N_14916,N_14942);
xor UO_923 (O_923,N_14960,N_14851);
or UO_924 (O_924,N_14972,N_14855);
xor UO_925 (O_925,N_14918,N_14981);
or UO_926 (O_926,N_14949,N_14901);
and UO_927 (O_927,N_14870,N_14903);
nor UO_928 (O_928,N_14885,N_14988);
nor UO_929 (O_929,N_14928,N_14940);
xnor UO_930 (O_930,N_14864,N_14908);
nand UO_931 (O_931,N_14869,N_14979);
nor UO_932 (O_932,N_14960,N_14874);
and UO_933 (O_933,N_14945,N_14912);
and UO_934 (O_934,N_14893,N_14921);
and UO_935 (O_935,N_14881,N_14912);
and UO_936 (O_936,N_14978,N_14896);
nand UO_937 (O_937,N_14914,N_14937);
and UO_938 (O_938,N_14899,N_14990);
nand UO_939 (O_939,N_14934,N_14936);
or UO_940 (O_940,N_14995,N_14886);
xnor UO_941 (O_941,N_14869,N_14968);
nand UO_942 (O_942,N_14931,N_14955);
nand UO_943 (O_943,N_14944,N_14881);
nand UO_944 (O_944,N_14910,N_14975);
xnor UO_945 (O_945,N_14907,N_14989);
xor UO_946 (O_946,N_14986,N_14862);
xor UO_947 (O_947,N_14869,N_14956);
and UO_948 (O_948,N_14982,N_14856);
or UO_949 (O_949,N_14925,N_14896);
and UO_950 (O_950,N_14854,N_14929);
and UO_951 (O_951,N_14913,N_14933);
and UO_952 (O_952,N_14874,N_14923);
nand UO_953 (O_953,N_14993,N_14942);
xor UO_954 (O_954,N_14892,N_14991);
nand UO_955 (O_955,N_14986,N_14996);
and UO_956 (O_956,N_14867,N_14979);
xnor UO_957 (O_957,N_14910,N_14982);
nand UO_958 (O_958,N_14855,N_14979);
and UO_959 (O_959,N_14870,N_14918);
or UO_960 (O_960,N_14920,N_14882);
or UO_961 (O_961,N_14955,N_14888);
nor UO_962 (O_962,N_14949,N_14968);
xor UO_963 (O_963,N_14896,N_14919);
nor UO_964 (O_964,N_14982,N_14869);
xnor UO_965 (O_965,N_14917,N_14977);
xor UO_966 (O_966,N_14908,N_14994);
xor UO_967 (O_967,N_14879,N_14990);
nand UO_968 (O_968,N_14965,N_14964);
and UO_969 (O_969,N_14864,N_14955);
and UO_970 (O_970,N_14964,N_14904);
and UO_971 (O_971,N_14872,N_14976);
nor UO_972 (O_972,N_14981,N_14976);
and UO_973 (O_973,N_14974,N_14885);
xnor UO_974 (O_974,N_14872,N_14982);
and UO_975 (O_975,N_14907,N_14851);
nor UO_976 (O_976,N_14887,N_14874);
nor UO_977 (O_977,N_14861,N_14877);
nor UO_978 (O_978,N_14907,N_14861);
or UO_979 (O_979,N_14881,N_14862);
xnor UO_980 (O_980,N_14877,N_14935);
and UO_981 (O_981,N_14941,N_14934);
nor UO_982 (O_982,N_14894,N_14933);
or UO_983 (O_983,N_14993,N_14934);
and UO_984 (O_984,N_14881,N_14855);
or UO_985 (O_985,N_14914,N_14894);
nor UO_986 (O_986,N_14908,N_14934);
nand UO_987 (O_987,N_14965,N_14945);
nand UO_988 (O_988,N_14930,N_14888);
or UO_989 (O_989,N_14951,N_14936);
nor UO_990 (O_990,N_14995,N_14962);
or UO_991 (O_991,N_14929,N_14892);
xnor UO_992 (O_992,N_14966,N_14953);
and UO_993 (O_993,N_14980,N_14969);
xor UO_994 (O_994,N_14903,N_14914);
xor UO_995 (O_995,N_14962,N_14850);
xnor UO_996 (O_996,N_14971,N_14920);
or UO_997 (O_997,N_14857,N_14893);
nor UO_998 (O_998,N_14926,N_14952);
or UO_999 (O_999,N_14991,N_14985);
or UO_1000 (O_1000,N_14943,N_14859);
nor UO_1001 (O_1001,N_14908,N_14937);
and UO_1002 (O_1002,N_14987,N_14980);
nand UO_1003 (O_1003,N_14940,N_14882);
xnor UO_1004 (O_1004,N_14913,N_14895);
xor UO_1005 (O_1005,N_14982,N_14928);
or UO_1006 (O_1006,N_14957,N_14853);
nor UO_1007 (O_1007,N_14950,N_14956);
or UO_1008 (O_1008,N_14914,N_14917);
and UO_1009 (O_1009,N_14870,N_14973);
or UO_1010 (O_1010,N_14850,N_14960);
and UO_1011 (O_1011,N_14970,N_14916);
xnor UO_1012 (O_1012,N_14962,N_14977);
or UO_1013 (O_1013,N_14850,N_14920);
and UO_1014 (O_1014,N_14957,N_14911);
nor UO_1015 (O_1015,N_14972,N_14993);
and UO_1016 (O_1016,N_14888,N_14934);
or UO_1017 (O_1017,N_14905,N_14989);
nand UO_1018 (O_1018,N_14859,N_14982);
and UO_1019 (O_1019,N_14922,N_14924);
nand UO_1020 (O_1020,N_14964,N_14894);
xnor UO_1021 (O_1021,N_14877,N_14901);
xnor UO_1022 (O_1022,N_14941,N_14929);
and UO_1023 (O_1023,N_14946,N_14905);
nor UO_1024 (O_1024,N_14916,N_14971);
or UO_1025 (O_1025,N_14886,N_14922);
nor UO_1026 (O_1026,N_14924,N_14934);
nand UO_1027 (O_1027,N_14937,N_14999);
or UO_1028 (O_1028,N_14898,N_14855);
and UO_1029 (O_1029,N_14987,N_14972);
xor UO_1030 (O_1030,N_14882,N_14957);
or UO_1031 (O_1031,N_14851,N_14893);
and UO_1032 (O_1032,N_14923,N_14970);
nor UO_1033 (O_1033,N_14901,N_14871);
nor UO_1034 (O_1034,N_14877,N_14987);
and UO_1035 (O_1035,N_14953,N_14938);
nor UO_1036 (O_1036,N_14964,N_14924);
nor UO_1037 (O_1037,N_14966,N_14873);
nand UO_1038 (O_1038,N_14886,N_14923);
or UO_1039 (O_1039,N_14980,N_14930);
and UO_1040 (O_1040,N_14929,N_14966);
xnor UO_1041 (O_1041,N_14971,N_14874);
and UO_1042 (O_1042,N_14987,N_14995);
nand UO_1043 (O_1043,N_14960,N_14932);
xor UO_1044 (O_1044,N_14956,N_14932);
nor UO_1045 (O_1045,N_14944,N_14977);
or UO_1046 (O_1046,N_14856,N_14981);
and UO_1047 (O_1047,N_14856,N_14988);
nand UO_1048 (O_1048,N_14898,N_14913);
nor UO_1049 (O_1049,N_14923,N_14926);
nor UO_1050 (O_1050,N_14907,N_14916);
nand UO_1051 (O_1051,N_14976,N_14881);
and UO_1052 (O_1052,N_14933,N_14899);
nor UO_1053 (O_1053,N_14916,N_14918);
xnor UO_1054 (O_1054,N_14909,N_14930);
or UO_1055 (O_1055,N_14941,N_14971);
or UO_1056 (O_1056,N_14962,N_14955);
and UO_1057 (O_1057,N_14877,N_14945);
nor UO_1058 (O_1058,N_14943,N_14906);
nand UO_1059 (O_1059,N_14942,N_14879);
nand UO_1060 (O_1060,N_14921,N_14930);
xor UO_1061 (O_1061,N_14984,N_14890);
xor UO_1062 (O_1062,N_14916,N_14879);
or UO_1063 (O_1063,N_14941,N_14976);
nor UO_1064 (O_1064,N_14885,N_14937);
and UO_1065 (O_1065,N_14959,N_14899);
and UO_1066 (O_1066,N_14953,N_14886);
and UO_1067 (O_1067,N_14909,N_14904);
nor UO_1068 (O_1068,N_14874,N_14973);
nor UO_1069 (O_1069,N_14985,N_14999);
nand UO_1070 (O_1070,N_14917,N_14986);
and UO_1071 (O_1071,N_14955,N_14947);
nor UO_1072 (O_1072,N_14999,N_14966);
or UO_1073 (O_1073,N_14931,N_14866);
and UO_1074 (O_1074,N_14937,N_14929);
or UO_1075 (O_1075,N_14915,N_14871);
nor UO_1076 (O_1076,N_14994,N_14918);
or UO_1077 (O_1077,N_14980,N_14924);
nand UO_1078 (O_1078,N_14909,N_14882);
and UO_1079 (O_1079,N_14868,N_14866);
nand UO_1080 (O_1080,N_14989,N_14933);
nand UO_1081 (O_1081,N_14861,N_14879);
nand UO_1082 (O_1082,N_14912,N_14856);
nand UO_1083 (O_1083,N_14884,N_14946);
nor UO_1084 (O_1084,N_14879,N_14884);
nor UO_1085 (O_1085,N_14920,N_14943);
nand UO_1086 (O_1086,N_14912,N_14957);
nand UO_1087 (O_1087,N_14990,N_14876);
or UO_1088 (O_1088,N_14925,N_14906);
xor UO_1089 (O_1089,N_14964,N_14972);
and UO_1090 (O_1090,N_14926,N_14974);
and UO_1091 (O_1091,N_14957,N_14978);
and UO_1092 (O_1092,N_14976,N_14988);
or UO_1093 (O_1093,N_14865,N_14918);
nor UO_1094 (O_1094,N_14946,N_14895);
and UO_1095 (O_1095,N_14915,N_14918);
xnor UO_1096 (O_1096,N_14900,N_14870);
nand UO_1097 (O_1097,N_14890,N_14861);
xor UO_1098 (O_1098,N_14899,N_14879);
nor UO_1099 (O_1099,N_14994,N_14929);
xnor UO_1100 (O_1100,N_14981,N_14857);
xor UO_1101 (O_1101,N_14983,N_14986);
xnor UO_1102 (O_1102,N_14928,N_14875);
and UO_1103 (O_1103,N_14883,N_14976);
nand UO_1104 (O_1104,N_14870,N_14880);
nand UO_1105 (O_1105,N_14933,N_14977);
nand UO_1106 (O_1106,N_14895,N_14982);
or UO_1107 (O_1107,N_14907,N_14899);
nor UO_1108 (O_1108,N_14972,N_14948);
nor UO_1109 (O_1109,N_14909,N_14958);
xor UO_1110 (O_1110,N_14878,N_14997);
nand UO_1111 (O_1111,N_14979,N_14969);
nand UO_1112 (O_1112,N_14921,N_14888);
nor UO_1113 (O_1113,N_14986,N_14926);
xnor UO_1114 (O_1114,N_14992,N_14998);
nand UO_1115 (O_1115,N_14956,N_14945);
and UO_1116 (O_1116,N_14980,N_14921);
xor UO_1117 (O_1117,N_14983,N_14937);
xor UO_1118 (O_1118,N_14995,N_14876);
nor UO_1119 (O_1119,N_14924,N_14869);
nor UO_1120 (O_1120,N_14885,N_14963);
and UO_1121 (O_1121,N_14956,N_14988);
xnor UO_1122 (O_1122,N_14896,N_14911);
nor UO_1123 (O_1123,N_14880,N_14854);
nand UO_1124 (O_1124,N_14976,N_14992);
and UO_1125 (O_1125,N_14981,N_14967);
nand UO_1126 (O_1126,N_14956,N_14923);
xnor UO_1127 (O_1127,N_14918,N_14989);
nor UO_1128 (O_1128,N_14953,N_14939);
or UO_1129 (O_1129,N_14932,N_14916);
nor UO_1130 (O_1130,N_14874,N_14981);
nand UO_1131 (O_1131,N_14879,N_14956);
and UO_1132 (O_1132,N_14875,N_14932);
nor UO_1133 (O_1133,N_14988,N_14872);
and UO_1134 (O_1134,N_14932,N_14931);
and UO_1135 (O_1135,N_14884,N_14871);
or UO_1136 (O_1136,N_14910,N_14850);
or UO_1137 (O_1137,N_14959,N_14910);
nand UO_1138 (O_1138,N_14873,N_14997);
and UO_1139 (O_1139,N_14952,N_14906);
or UO_1140 (O_1140,N_14894,N_14860);
xor UO_1141 (O_1141,N_14921,N_14862);
xor UO_1142 (O_1142,N_14968,N_14996);
or UO_1143 (O_1143,N_14989,N_14940);
nand UO_1144 (O_1144,N_14862,N_14957);
and UO_1145 (O_1145,N_14924,N_14975);
nor UO_1146 (O_1146,N_14986,N_14951);
and UO_1147 (O_1147,N_14850,N_14937);
nand UO_1148 (O_1148,N_14938,N_14911);
nor UO_1149 (O_1149,N_14877,N_14873);
and UO_1150 (O_1150,N_14924,N_14978);
nand UO_1151 (O_1151,N_14901,N_14892);
nand UO_1152 (O_1152,N_14973,N_14880);
and UO_1153 (O_1153,N_14862,N_14956);
xor UO_1154 (O_1154,N_14932,N_14967);
nor UO_1155 (O_1155,N_14872,N_14947);
nand UO_1156 (O_1156,N_14953,N_14904);
or UO_1157 (O_1157,N_14881,N_14875);
or UO_1158 (O_1158,N_14994,N_14910);
nand UO_1159 (O_1159,N_14966,N_14927);
and UO_1160 (O_1160,N_14896,N_14865);
nand UO_1161 (O_1161,N_14852,N_14923);
or UO_1162 (O_1162,N_14966,N_14931);
or UO_1163 (O_1163,N_14913,N_14859);
xor UO_1164 (O_1164,N_14875,N_14851);
or UO_1165 (O_1165,N_14949,N_14979);
nand UO_1166 (O_1166,N_14882,N_14887);
nand UO_1167 (O_1167,N_14994,N_14941);
nand UO_1168 (O_1168,N_14902,N_14898);
nand UO_1169 (O_1169,N_14971,N_14851);
nor UO_1170 (O_1170,N_14997,N_14896);
and UO_1171 (O_1171,N_14961,N_14925);
or UO_1172 (O_1172,N_14897,N_14854);
nor UO_1173 (O_1173,N_14910,N_14961);
xnor UO_1174 (O_1174,N_14918,N_14904);
and UO_1175 (O_1175,N_14853,N_14914);
nand UO_1176 (O_1176,N_14889,N_14943);
xor UO_1177 (O_1177,N_14993,N_14991);
nor UO_1178 (O_1178,N_14892,N_14958);
xnor UO_1179 (O_1179,N_14875,N_14893);
or UO_1180 (O_1180,N_14946,N_14920);
or UO_1181 (O_1181,N_14938,N_14948);
or UO_1182 (O_1182,N_14873,N_14925);
and UO_1183 (O_1183,N_14953,N_14868);
or UO_1184 (O_1184,N_14968,N_14974);
nand UO_1185 (O_1185,N_14852,N_14967);
nand UO_1186 (O_1186,N_14950,N_14889);
nor UO_1187 (O_1187,N_14948,N_14939);
nor UO_1188 (O_1188,N_14931,N_14874);
xor UO_1189 (O_1189,N_14937,N_14938);
nand UO_1190 (O_1190,N_14989,N_14968);
xnor UO_1191 (O_1191,N_14851,N_14952);
nand UO_1192 (O_1192,N_14902,N_14952);
nor UO_1193 (O_1193,N_14977,N_14928);
nor UO_1194 (O_1194,N_14965,N_14892);
and UO_1195 (O_1195,N_14854,N_14863);
nand UO_1196 (O_1196,N_14881,N_14866);
xor UO_1197 (O_1197,N_14976,N_14885);
xnor UO_1198 (O_1198,N_14858,N_14899);
nand UO_1199 (O_1199,N_14866,N_14984);
nor UO_1200 (O_1200,N_14985,N_14915);
nor UO_1201 (O_1201,N_14901,N_14921);
and UO_1202 (O_1202,N_14979,N_14936);
nor UO_1203 (O_1203,N_14860,N_14954);
xor UO_1204 (O_1204,N_14972,N_14900);
xor UO_1205 (O_1205,N_14943,N_14999);
nand UO_1206 (O_1206,N_14870,N_14865);
and UO_1207 (O_1207,N_14878,N_14880);
nand UO_1208 (O_1208,N_14920,N_14954);
nand UO_1209 (O_1209,N_14892,N_14916);
and UO_1210 (O_1210,N_14857,N_14862);
or UO_1211 (O_1211,N_14880,N_14896);
xnor UO_1212 (O_1212,N_14874,N_14881);
or UO_1213 (O_1213,N_14918,N_14973);
xnor UO_1214 (O_1214,N_14924,N_14853);
or UO_1215 (O_1215,N_14999,N_14902);
xor UO_1216 (O_1216,N_14954,N_14976);
nand UO_1217 (O_1217,N_14885,N_14975);
or UO_1218 (O_1218,N_14867,N_14971);
or UO_1219 (O_1219,N_14934,N_14890);
and UO_1220 (O_1220,N_14854,N_14910);
or UO_1221 (O_1221,N_14951,N_14984);
xnor UO_1222 (O_1222,N_14998,N_14878);
or UO_1223 (O_1223,N_14947,N_14960);
xor UO_1224 (O_1224,N_14879,N_14925);
nor UO_1225 (O_1225,N_14903,N_14968);
and UO_1226 (O_1226,N_14906,N_14947);
and UO_1227 (O_1227,N_14989,N_14971);
xnor UO_1228 (O_1228,N_14903,N_14985);
xor UO_1229 (O_1229,N_14958,N_14982);
or UO_1230 (O_1230,N_14904,N_14945);
xor UO_1231 (O_1231,N_14983,N_14931);
nor UO_1232 (O_1232,N_14994,N_14984);
and UO_1233 (O_1233,N_14923,N_14935);
nand UO_1234 (O_1234,N_14912,N_14874);
xnor UO_1235 (O_1235,N_14913,N_14943);
nor UO_1236 (O_1236,N_14874,N_14897);
or UO_1237 (O_1237,N_14850,N_14925);
nand UO_1238 (O_1238,N_14979,N_14878);
and UO_1239 (O_1239,N_14860,N_14865);
nand UO_1240 (O_1240,N_14899,N_14900);
and UO_1241 (O_1241,N_14935,N_14906);
or UO_1242 (O_1242,N_14880,N_14980);
nand UO_1243 (O_1243,N_14978,N_14966);
nand UO_1244 (O_1244,N_14987,N_14928);
and UO_1245 (O_1245,N_14963,N_14856);
nand UO_1246 (O_1246,N_14929,N_14953);
nand UO_1247 (O_1247,N_14887,N_14877);
nand UO_1248 (O_1248,N_14918,N_14941);
nor UO_1249 (O_1249,N_14972,N_14933);
nor UO_1250 (O_1250,N_14878,N_14899);
nand UO_1251 (O_1251,N_14990,N_14919);
nand UO_1252 (O_1252,N_14852,N_14939);
nand UO_1253 (O_1253,N_14894,N_14884);
nor UO_1254 (O_1254,N_14910,N_14869);
and UO_1255 (O_1255,N_14900,N_14888);
nor UO_1256 (O_1256,N_14923,N_14955);
nor UO_1257 (O_1257,N_14916,N_14931);
xor UO_1258 (O_1258,N_14892,N_14853);
nand UO_1259 (O_1259,N_14911,N_14993);
nor UO_1260 (O_1260,N_14899,N_14956);
nor UO_1261 (O_1261,N_14875,N_14943);
nand UO_1262 (O_1262,N_14963,N_14866);
and UO_1263 (O_1263,N_14975,N_14964);
or UO_1264 (O_1264,N_14916,N_14969);
nor UO_1265 (O_1265,N_14970,N_14925);
nand UO_1266 (O_1266,N_14902,N_14935);
and UO_1267 (O_1267,N_14986,N_14964);
nor UO_1268 (O_1268,N_14879,N_14973);
xnor UO_1269 (O_1269,N_14991,N_14953);
nor UO_1270 (O_1270,N_14982,N_14934);
nor UO_1271 (O_1271,N_14916,N_14908);
or UO_1272 (O_1272,N_14887,N_14926);
and UO_1273 (O_1273,N_14884,N_14865);
nand UO_1274 (O_1274,N_14860,N_14862);
nor UO_1275 (O_1275,N_14933,N_14878);
xnor UO_1276 (O_1276,N_14927,N_14915);
or UO_1277 (O_1277,N_14913,N_14981);
xnor UO_1278 (O_1278,N_14921,N_14995);
nor UO_1279 (O_1279,N_14865,N_14866);
and UO_1280 (O_1280,N_14875,N_14895);
nand UO_1281 (O_1281,N_14851,N_14903);
or UO_1282 (O_1282,N_14892,N_14996);
xor UO_1283 (O_1283,N_14923,N_14894);
nor UO_1284 (O_1284,N_14932,N_14952);
xnor UO_1285 (O_1285,N_14982,N_14956);
xor UO_1286 (O_1286,N_14891,N_14933);
nor UO_1287 (O_1287,N_14933,N_14950);
nor UO_1288 (O_1288,N_14944,N_14904);
and UO_1289 (O_1289,N_14852,N_14898);
and UO_1290 (O_1290,N_14983,N_14881);
or UO_1291 (O_1291,N_14905,N_14967);
nand UO_1292 (O_1292,N_14996,N_14867);
nand UO_1293 (O_1293,N_14941,N_14951);
nand UO_1294 (O_1294,N_14851,N_14870);
xnor UO_1295 (O_1295,N_14999,N_14946);
and UO_1296 (O_1296,N_14875,N_14909);
xnor UO_1297 (O_1297,N_14884,N_14972);
nand UO_1298 (O_1298,N_14927,N_14958);
nand UO_1299 (O_1299,N_14999,N_14913);
nand UO_1300 (O_1300,N_14853,N_14945);
and UO_1301 (O_1301,N_14888,N_14998);
xor UO_1302 (O_1302,N_14901,N_14928);
and UO_1303 (O_1303,N_14958,N_14854);
nor UO_1304 (O_1304,N_14895,N_14863);
nor UO_1305 (O_1305,N_14897,N_14975);
xor UO_1306 (O_1306,N_14853,N_14880);
nor UO_1307 (O_1307,N_14934,N_14975);
or UO_1308 (O_1308,N_14985,N_14877);
xnor UO_1309 (O_1309,N_14858,N_14988);
or UO_1310 (O_1310,N_14957,N_14855);
or UO_1311 (O_1311,N_14851,N_14876);
nor UO_1312 (O_1312,N_14880,N_14933);
or UO_1313 (O_1313,N_14914,N_14960);
nor UO_1314 (O_1314,N_14887,N_14971);
or UO_1315 (O_1315,N_14922,N_14979);
xnor UO_1316 (O_1316,N_14896,N_14938);
and UO_1317 (O_1317,N_14936,N_14918);
or UO_1318 (O_1318,N_14897,N_14959);
nand UO_1319 (O_1319,N_14960,N_14985);
nand UO_1320 (O_1320,N_14910,N_14934);
nor UO_1321 (O_1321,N_14947,N_14882);
nor UO_1322 (O_1322,N_14865,N_14897);
or UO_1323 (O_1323,N_14919,N_14890);
nor UO_1324 (O_1324,N_14911,N_14853);
nand UO_1325 (O_1325,N_14969,N_14925);
nand UO_1326 (O_1326,N_14869,N_14877);
or UO_1327 (O_1327,N_14910,N_14867);
or UO_1328 (O_1328,N_14863,N_14996);
xnor UO_1329 (O_1329,N_14945,N_14958);
or UO_1330 (O_1330,N_14874,N_14959);
nand UO_1331 (O_1331,N_14868,N_14957);
nor UO_1332 (O_1332,N_14900,N_14939);
nand UO_1333 (O_1333,N_14959,N_14868);
nor UO_1334 (O_1334,N_14946,N_14901);
nand UO_1335 (O_1335,N_14883,N_14964);
nand UO_1336 (O_1336,N_14851,N_14973);
or UO_1337 (O_1337,N_14851,N_14852);
or UO_1338 (O_1338,N_14953,N_14905);
and UO_1339 (O_1339,N_14971,N_14922);
xnor UO_1340 (O_1340,N_14913,N_14937);
or UO_1341 (O_1341,N_14892,N_14855);
xnor UO_1342 (O_1342,N_14861,N_14896);
and UO_1343 (O_1343,N_14920,N_14964);
or UO_1344 (O_1344,N_14975,N_14980);
or UO_1345 (O_1345,N_14997,N_14875);
xnor UO_1346 (O_1346,N_14934,N_14950);
xnor UO_1347 (O_1347,N_14919,N_14974);
nand UO_1348 (O_1348,N_14977,N_14914);
nand UO_1349 (O_1349,N_14983,N_14960);
and UO_1350 (O_1350,N_14956,N_14985);
xnor UO_1351 (O_1351,N_14957,N_14935);
xor UO_1352 (O_1352,N_14926,N_14882);
nor UO_1353 (O_1353,N_14989,N_14975);
nor UO_1354 (O_1354,N_14911,N_14892);
and UO_1355 (O_1355,N_14874,N_14905);
and UO_1356 (O_1356,N_14941,N_14996);
nand UO_1357 (O_1357,N_14861,N_14955);
xor UO_1358 (O_1358,N_14918,N_14949);
and UO_1359 (O_1359,N_14981,N_14916);
or UO_1360 (O_1360,N_14908,N_14878);
xnor UO_1361 (O_1361,N_14947,N_14962);
and UO_1362 (O_1362,N_14886,N_14861);
xnor UO_1363 (O_1363,N_14967,N_14875);
nand UO_1364 (O_1364,N_14901,N_14998);
and UO_1365 (O_1365,N_14998,N_14932);
nand UO_1366 (O_1366,N_14921,N_14953);
and UO_1367 (O_1367,N_14908,N_14868);
xnor UO_1368 (O_1368,N_14944,N_14903);
xor UO_1369 (O_1369,N_14939,N_14859);
xnor UO_1370 (O_1370,N_14881,N_14867);
or UO_1371 (O_1371,N_14978,N_14911);
nand UO_1372 (O_1372,N_14870,N_14855);
and UO_1373 (O_1373,N_14963,N_14864);
and UO_1374 (O_1374,N_14905,N_14991);
xnor UO_1375 (O_1375,N_14905,N_14981);
nor UO_1376 (O_1376,N_14952,N_14915);
or UO_1377 (O_1377,N_14944,N_14917);
nor UO_1378 (O_1378,N_14860,N_14922);
nand UO_1379 (O_1379,N_14893,N_14882);
and UO_1380 (O_1380,N_14974,N_14886);
nor UO_1381 (O_1381,N_14949,N_14944);
and UO_1382 (O_1382,N_14869,N_14998);
nor UO_1383 (O_1383,N_14878,N_14929);
nand UO_1384 (O_1384,N_14998,N_14999);
xor UO_1385 (O_1385,N_14948,N_14993);
nor UO_1386 (O_1386,N_14939,N_14932);
and UO_1387 (O_1387,N_14897,N_14877);
nand UO_1388 (O_1388,N_14948,N_14973);
nand UO_1389 (O_1389,N_14925,N_14885);
nand UO_1390 (O_1390,N_14877,N_14858);
and UO_1391 (O_1391,N_14957,N_14925);
and UO_1392 (O_1392,N_14996,N_14938);
and UO_1393 (O_1393,N_14911,N_14882);
nand UO_1394 (O_1394,N_14888,N_14899);
nor UO_1395 (O_1395,N_14995,N_14986);
nor UO_1396 (O_1396,N_14968,N_14908);
nand UO_1397 (O_1397,N_14878,N_14984);
or UO_1398 (O_1398,N_14985,N_14892);
or UO_1399 (O_1399,N_14865,N_14977);
and UO_1400 (O_1400,N_14854,N_14944);
and UO_1401 (O_1401,N_14881,N_14887);
and UO_1402 (O_1402,N_14967,N_14993);
nor UO_1403 (O_1403,N_14990,N_14855);
nor UO_1404 (O_1404,N_14954,N_14886);
xor UO_1405 (O_1405,N_14961,N_14952);
nor UO_1406 (O_1406,N_14922,N_14878);
and UO_1407 (O_1407,N_14858,N_14910);
or UO_1408 (O_1408,N_14987,N_14954);
or UO_1409 (O_1409,N_14916,N_14874);
nor UO_1410 (O_1410,N_14993,N_14856);
nand UO_1411 (O_1411,N_14859,N_14869);
or UO_1412 (O_1412,N_14871,N_14887);
nor UO_1413 (O_1413,N_14862,N_14951);
nor UO_1414 (O_1414,N_14956,N_14877);
nor UO_1415 (O_1415,N_14923,N_14995);
or UO_1416 (O_1416,N_14871,N_14951);
nor UO_1417 (O_1417,N_14859,N_14962);
xnor UO_1418 (O_1418,N_14971,N_14940);
nand UO_1419 (O_1419,N_14946,N_14940);
or UO_1420 (O_1420,N_14872,N_14884);
or UO_1421 (O_1421,N_14929,N_14874);
nand UO_1422 (O_1422,N_14922,N_14932);
and UO_1423 (O_1423,N_14855,N_14851);
nand UO_1424 (O_1424,N_14862,N_14948);
nand UO_1425 (O_1425,N_14857,N_14937);
nor UO_1426 (O_1426,N_14932,N_14906);
xor UO_1427 (O_1427,N_14880,N_14932);
nor UO_1428 (O_1428,N_14978,N_14851);
or UO_1429 (O_1429,N_14950,N_14923);
xnor UO_1430 (O_1430,N_14879,N_14947);
and UO_1431 (O_1431,N_14860,N_14936);
and UO_1432 (O_1432,N_14868,N_14962);
and UO_1433 (O_1433,N_14851,N_14894);
nor UO_1434 (O_1434,N_14971,N_14882);
or UO_1435 (O_1435,N_14893,N_14911);
and UO_1436 (O_1436,N_14854,N_14998);
or UO_1437 (O_1437,N_14956,N_14993);
nand UO_1438 (O_1438,N_14909,N_14876);
nand UO_1439 (O_1439,N_14981,N_14893);
and UO_1440 (O_1440,N_14916,N_14903);
and UO_1441 (O_1441,N_14924,N_14858);
nor UO_1442 (O_1442,N_14912,N_14930);
nor UO_1443 (O_1443,N_14989,N_14976);
or UO_1444 (O_1444,N_14897,N_14960);
and UO_1445 (O_1445,N_14863,N_14953);
nor UO_1446 (O_1446,N_14974,N_14957);
xnor UO_1447 (O_1447,N_14922,N_14929);
nor UO_1448 (O_1448,N_14968,N_14941);
or UO_1449 (O_1449,N_14957,N_14890);
nand UO_1450 (O_1450,N_14906,N_14966);
and UO_1451 (O_1451,N_14967,N_14970);
or UO_1452 (O_1452,N_14860,N_14956);
and UO_1453 (O_1453,N_14954,N_14983);
or UO_1454 (O_1454,N_14922,N_14883);
xnor UO_1455 (O_1455,N_14957,N_14863);
and UO_1456 (O_1456,N_14911,N_14903);
or UO_1457 (O_1457,N_14948,N_14921);
and UO_1458 (O_1458,N_14910,N_14880);
nand UO_1459 (O_1459,N_14851,N_14891);
or UO_1460 (O_1460,N_14982,N_14909);
nand UO_1461 (O_1461,N_14941,N_14858);
or UO_1462 (O_1462,N_14958,N_14920);
xnor UO_1463 (O_1463,N_14872,N_14936);
nand UO_1464 (O_1464,N_14976,N_14911);
xnor UO_1465 (O_1465,N_14999,N_14983);
nor UO_1466 (O_1466,N_14907,N_14942);
and UO_1467 (O_1467,N_14922,N_14867);
nor UO_1468 (O_1468,N_14903,N_14901);
and UO_1469 (O_1469,N_14860,N_14902);
nand UO_1470 (O_1470,N_14998,N_14892);
or UO_1471 (O_1471,N_14865,N_14858);
nand UO_1472 (O_1472,N_14960,N_14965);
nor UO_1473 (O_1473,N_14943,N_14960);
or UO_1474 (O_1474,N_14910,N_14957);
nand UO_1475 (O_1475,N_14877,N_14933);
and UO_1476 (O_1476,N_14983,N_14879);
nor UO_1477 (O_1477,N_14908,N_14953);
nor UO_1478 (O_1478,N_14877,N_14997);
nor UO_1479 (O_1479,N_14974,N_14978);
and UO_1480 (O_1480,N_14913,N_14957);
xor UO_1481 (O_1481,N_14974,N_14940);
nand UO_1482 (O_1482,N_14962,N_14896);
and UO_1483 (O_1483,N_14994,N_14907);
and UO_1484 (O_1484,N_14908,N_14877);
nor UO_1485 (O_1485,N_14959,N_14860);
or UO_1486 (O_1486,N_14965,N_14929);
nand UO_1487 (O_1487,N_14880,N_14893);
or UO_1488 (O_1488,N_14919,N_14918);
or UO_1489 (O_1489,N_14876,N_14911);
xnor UO_1490 (O_1490,N_14870,N_14963);
and UO_1491 (O_1491,N_14879,N_14980);
nor UO_1492 (O_1492,N_14907,N_14943);
and UO_1493 (O_1493,N_14866,N_14956);
nor UO_1494 (O_1494,N_14959,N_14962);
xnor UO_1495 (O_1495,N_14997,N_14952);
or UO_1496 (O_1496,N_14979,N_14906);
or UO_1497 (O_1497,N_14992,N_14882);
nor UO_1498 (O_1498,N_14953,N_14964);
nand UO_1499 (O_1499,N_14875,N_14916);
nor UO_1500 (O_1500,N_14892,N_14968);
xor UO_1501 (O_1501,N_14919,N_14929);
and UO_1502 (O_1502,N_14981,N_14947);
or UO_1503 (O_1503,N_14988,N_14915);
or UO_1504 (O_1504,N_14946,N_14852);
xor UO_1505 (O_1505,N_14950,N_14855);
nand UO_1506 (O_1506,N_14852,N_14921);
nor UO_1507 (O_1507,N_14993,N_14907);
and UO_1508 (O_1508,N_14927,N_14880);
or UO_1509 (O_1509,N_14914,N_14864);
or UO_1510 (O_1510,N_14982,N_14915);
or UO_1511 (O_1511,N_14994,N_14959);
or UO_1512 (O_1512,N_14895,N_14876);
and UO_1513 (O_1513,N_14999,N_14949);
and UO_1514 (O_1514,N_14941,N_14928);
or UO_1515 (O_1515,N_14893,N_14948);
nand UO_1516 (O_1516,N_14976,N_14865);
xnor UO_1517 (O_1517,N_14877,N_14972);
xnor UO_1518 (O_1518,N_14859,N_14904);
xor UO_1519 (O_1519,N_14872,N_14879);
nand UO_1520 (O_1520,N_14860,N_14886);
nor UO_1521 (O_1521,N_14986,N_14942);
or UO_1522 (O_1522,N_14996,N_14854);
and UO_1523 (O_1523,N_14970,N_14930);
nand UO_1524 (O_1524,N_14890,N_14955);
nand UO_1525 (O_1525,N_14938,N_14964);
xor UO_1526 (O_1526,N_14886,N_14927);
and UO_1527 (O_1527,N_14984,N_14897);
and UO_1528 (O_1528,N_14880,N_14924);
or UO_1529 (O_1529,N_14885,N_14960);
nand UO_1530 (O_1530,N_14938,N_14952);
nor UO_1531 (O_1531,N_14979,N_14930);
xor UO_1532 (O_1532,N_14918,N_14952);
nand UO_1533 (O_1533,N_14955,N_14961);
nand UO_1534 (O_1534,N_14943,N_14939);
nor UO_1535 (O_1535,N_14958,N_14997);
nand UO_1536 (O_1536,N_14878,N_14991);
nand UO_1537 (O_1537,N_14890,N_14970);
nor UO_1538 (O_1538,N_14917,N_14873);
nor UO_1539 (O_1539,N_14876,N_14937);
or UO_1540 (O_1540,N_14949,N_14935);
nand UO_1541 (O_1541,N_14870,N_14947);
xor UO_1542 (O_1542,N_14873,N_14880);
nor UO_1543 (O_1543,N_14859,N_14863);
or UO_1544 (O_1544,N_14964,N_14942);
or UO_1545 (O_1545,N_14925,N_14909);
or UO_1546 (O_1546,N_14991,N_14965);
nor UO_1547 (O_1547,N_14921,N_14969);
and UO_1548 (O_1548,N_14906,N_14892);
nand UO_1549 (O_1549,N_14936,N_14956);
nor UO_1550 (O_1550,N_14988,N_14924);
or UO_1551 (O_1551,N_14953,N_14917);
or UO_1552 (O_1552,N_14914,N_14982);
nor UO_1553 (O_1553,N_14851,N_14974);
and UO_1554 (O_1554,N_14999,N_14871);
nand UO_1555 (O_1555,N_14854,N_14914);
nor UO_1556 (O_1556,N_14902,N_14981);
nand UO_1557 (O_1557,N_14943,N_14942);
or UO_1558 (O_1558,N_14947,N_14987);
nor UO_1559 (O_1559,N_14935,N_14864);
xor UO_1560 (O_1560,N_14880,N_14921);
nor UO_1561 (O_1561,N_14866,N_14901);
xnor UO_1562 (O_1562,N_14948,N_14942);
or UO_1563 (O_1563,N_14892,N_14950);
nand UO_1564 (O_1564,N_14910,N_14895);
xor UO_1565 (O_1565,N_14955,N_14995);
and UO_1566 (O_1566,N_14990,N_14984);
or UO_1567 (O_1567,N_14935,N_14921);
xnor UO_1568 (O_1568,N_14851,N_14934);
xnor UO_1569 (O_1569,N_14965,N_14940);
and UO_1570 (O_1570,N_14850,N_14867);
and UO_1571 (O_1571,N_14894,N_14943);
or UO_1572 (O_1572,N_14930,N_14924);
xnor UO_1573 (O_1573,N_14929,N_14902);
nor UO_1574 (O_1574,N_14884,N_14869);
xnor UO_1575 (O_1575,N_14852,N_14983);
nor UO_1576 (O_1576,N_14967,N_14980);
nor UO_1577 (O_1577,N_14907,N_14933);
xnor UO_1578 (O_1578,N_14976,N_14867);
nand UO_1579 (O_1579,N_14959,N_14998);
nor UO_1580 (O_1580,N_14951,N_14972);
nand UO_1581 (O_1581,N_14964,N_14866);
and UO_1582 (O_1582,N_14889,N_14906);
and UO_1583 (O_1583,N_14853,N_14901);
nor UO_1584 (O_1584,N_14944,N_14874);
nor UO_1585 (O_1585,N_14924,N_14928);
xor UO_1586 (O_1586,N_14955,N_14932);
xor UO_1587 (O_1587,N_14905,N_14898);
nor UO_1588 (O_1588,N_14907,N_14940);
nand UO_1589 (O_1589,N_14896,N_14952);
nor UO_1590 (O_1590,N_14973,N_14960);
nand UO_1591 (O_1591,N_14887,N_14875);
or UO_1592 (O_1592,N_14951,N_14889);
or UO_1593 (O_1593,N_14880,N_14883);
nand UO_1594 (O_1594,N_14965,N_14857);
nand UO_1595 (O_1595,N_14918,N_14928);
nor UO_1596 (O_1596,N_14857,N_14856);
xor UO_1597 (O_1597,N_14917,N_14903);
nand UO_1598 (O_1598,N_14918,N_14997);
or UO_1599 (O_1599,N_14970,N_14857);
xor UO_1600 (O_1600,N_14953,N_14876);
nand UO_1601 (O_1601,N_14880,N_14998);
nand UO_1602 (O_1602,N_14895,N_14862);
xnor UO_1603 (O_1603,N_14905,N_14926);
xor UO_1604 (O_1604,N_14902,N_14863);
nand UO_1605 (O_1605,N_14938,N_14851);
nand UO_1606 (O_1606,N_14897,N_14998);
or UO_1607 (O_1607,N_14871,N_14936);
nand UO_1608 (O_1608,N_14911,N_14884);
or UO_1609 (O_1609,N_14939,N_14888);
xor UO_1610 (O_1610,N_14999,N_14892);
and UO_1611 (O_1611,N_14993,N_14861);
nand UO_1612 (O_1612,N_14877,N_14902);
nor UO_1613 (O_1613,N_14942,N_14952);
or UO_1614 (O_1614,N_14906,N_14857);
and UO_1615 (O_1615,N_14867,N_14895);
nor UO_1616 (O_1616,N_14852,N_14874);
or UO_1617 (O_1617,N_14906,N_14973);
nor UO_1618 (O_1618,N_14896,N_14934);
and UO_1619 (O_1619,N_14927,N_14887);
or UO_1620 (O_1620,N_14914,N_14995);
nor UO_1621 (O_1621,N_14966,N_14991);
nor UO_1622 (O_1622,N_14939,N_14989);
xor UO_1623 (O_1623,N_14987,N_14918);
or UO_1624 (O_1624,N_14967,N_14882);
or UO_1625 (O_1625,N_14992,N_14927);
xor UO_1626 (O_1626,N_14887,N_14863);
xnor UO_1627 (O_1627,N_14953,N_14852);
nor UO_1628 (O_1628,N_14880,N_14920);
nand UO_1629 (O_1629,N_14929,N_14931);
and UO_1630 (O_1630,N_14948,N_14991);
xor UO_1631 (O_1631,N_14928,N_14954);
and UO_1632 (O_1632,N_14971,N_14984);
nor UO_1633 (O_1633,N_14953,N_14894);
or UO_1634 (O_1634,N_14899,N_14913);
nor UO_1635 (O_1635,N_14965,N_14931);
or UO_1636 (O_1636,N_14959,N_14852);
nand UO_1637 (O_1637,N_14882,N_14894);
nand UO_1638 (O_1638,N_14938,N_14918);
and UO_1639 (O_1639,N_14900,N_14960);
and UO_1640 (O_1640,N_14974,N_14912);
and UO_1641 (O_1641,N_14978,N_14850);
and UO_1642 (O_1642,N_14967,N_14870);
xor UO_1643 (O_1643,N_14981,N_14978);
xor UO_1644 (O_1644,N_14870,N_14945);
nand UO_1645 (O_1645,N_14931,N_14906);
nor UO_1646 (O_1646,N_14886,N_14911);
xor UO_1647 (O_1647,N_14898,N_14966);
nor UO_1648 (O_1648,N_14985,N_14886);
and UO_1649 (O_1649,N_14932,N_14873);
or UO_1650 (O_1650,N_14873,N_14931);
nand UO_1651 (O_1651,N_14979,N_14932);
nand UO_1652 (O_1652,N_14928,N_14906);
and UO_1653 (O_1653,N_14853,N_14890);
nand UO_1654 (O_1654,N_14905,N_14872);
nand UO_1655 (O_1655,N_14885,N_14945);
and UO_1656 (O_1656,N_14981,N_14862);
xnor UO_1657 (O_1657,N_14945,N_14909);
xor UO_1658 (O_1658,N_14974,N_14950);
xor UO_1659 (O_1659,N_14971,N_14872);
nand UO_1660 (O_1660,N_14902,N_14905);
nor UO_1661 (O_1661,N_14921,N_14964);
nand UO_1662 (O_1662,N_14954,N_14855);
xnor UO_1663 (O_1663,N_14881,N_14923);
nor UO_1664 (O_1664,N_14857,N_14943);
xor UO_1665 (O_1665,N_14924,N_14987);
or UO_1666 (O_1666,N_14853,N_14961);
xor UO_1667 (O_1667,N_14939,N_14862);
nor UO_1668 (O_1668,N_14931,N_14872);
and UO_1669 (O_1669,N_14968,N_14975);
xor UO_1670 (O_1670,N_14925,N_14956);
or UO_1671 (O_1671,N_14909,N_14952);
and UO_1672 (O_1672,N_14945,N_14983);
nor UO_1673 (O_1673,N_14874,N_14967);
nor UO_1674 (O_1674,N_14887,N_14909);
xor UO_1675 (O_1675,N_14961,N_14931);
or UO_1676 (O_1676,N_14928,N_14852);
nand UO_1677 (O_1677,N_14850,N_14964);
nor UO_1678 (O_1678,N_14895,N_14987);
nor UO_1679 (O_1679,N_14996,N_14959);
nand UO_1680 (O_1680,N_14951,N_14970);
or UO_1681 (O_1681,N_14927,N_14912);
and UO_1682 (O_1682,N_14928,N_14876);
nand UO_1683 (O_1683,N_14940,N_14892);
and UO_1684 (O_1684,N_14979,N_14983);
nor UO_1685 (O_1685,N_14929,N_14987);
nor UO_1686 (O_1686,N_14922,N_14898);
or UO_1687 (O_1687,N_14892,N_14907);
nor UO_1688 (O_1688,N_14917,N_14988);
and UO_1689 (O_1689,N_14872,N_14951);
nor UO_1690 (O_1690,N_14887,N_14914);
xor UO_1691 (O_1691,N_14871,N_14911);
or UO_1692 (O_1692,N_14887,N_14907);
nand UO_1693 (O_1693,N_14898,N_14879);
nand UO_1694 (O_1694,N_14850,N_14989);
xnor UO_1695 (O_1695,N_14901,N_14937);
nand UO_1696 (O_1696,N_14893,N_14970);
or UO_1697 (O_1697,N_14898,N_14992);
xnor UO_1698 (O_1698,N_14915,N_14983);
nor UO_1699 (O_1699,N_14936,N_14944);
or UO_1700 (O_1700,N_14868,N_14960);
or UO_1701 (O_1701,N_14933,N_14866);
nor UO_1702 (O_1702,N_14950,N_14930);
or UO_1703 (O_1703,N_14997,N_14975);
nand UO_1704 (O_1704,N_14969,N_14882);
nand UO_1705 (O_1705,N_14924,N_14873);
or UO_1706 (O_1706,N_14989,N_14881);
and UO_1707 (O_1707,N_14892,N_14941);
and UO_1708 (O_1708,N_14885,N_14931);
xnor UO_1709 (O_1709,N_14916,N_14960);
or UO_1710 (O_1710,N_14883,N_14981);
nand UO_1711 (O_1711,N_14879,N_14999);
xnor UO_1712 (O_1712,N_14985,N_14882);
nand UO_1713 (O_1713,N_14940,N_14850);
nor UO_1714 (O_1714,N_14856,N_14937);
nor UO_1715 (O_1715,N_14899,N_14942);
and UO_1716 (O_1716,N_14988,N_14919);
nor UO_1717 (O_1717,N_14940,N_14891);
xnor UO_1718 (O_1718,N_14884,N_14980);
nor UO_1719 (O_1719,N_14941,N_14867);
or UO_1720 (O_1720,N_14916,N_14984);
and UO_1721 (O_1721,N_14853,N_14874);
and UO_1722 (O_1722,N_14866,N_14902);
and UO_1723 (O_1723,N_14927,N_14981);
or UO_1724 (O_1724,N_14962,N_14956);
or UO_1725 (O_1725,N_14894,N_14926);
nor UO_1726 (O_1726,N_14940,N_14958);
nor UO_1727 (O_1727,N_14878,N_14870);
or UO_1728 (O_1728,N_14979,N_14958);
and UO_1729 (O_1729,N_14910,N_14928);
xnor UO_1730 (O_1730,N_14978,N_14986);
and UO_1731 (O_1731,N_14963,N_14910);
xnor UO_1732 (O_1732,N_14969,N_14856);
nand UO_1733 (O_1733,N_14859,N_14965);
nand UO_1734 (O_1734,N_14890,N_14950);
nand UO_1735 (O_1735,N_14990,N_14858);
or UO_1736 (O_1736,N_14865,N_14863);
xnor UO_1737 (O_1737,N_14946,N_14948);
and UO_1738 (O_1738,N_14991,N_14972);
or UO_1739 (O_1739,N_14923,N_14902);
nor UO_1740 (O_1740,N_14876,N_14901);
and UO_1741 (O_1741,N_14895,N_14952);
xnor UO_1742 (O_1742,N_14923,N_14920);
xnor UO_1743 (O_1743,N_14909,N_14855);
xor UO_1744 (O_1744,N_14964,N_14884);
and UO_1745 (O_1745,N_14987,N_14894);
xor UO_1746 (O_1746,N_14959,N_14963);
nand UO_1747 (O_1747,N_14856,N_14888);
nor UO_1748 (O_1748,N_14969,N_14928);
nor UO_1749 (O_1749,N_14896,N_14903);
or UO_1750 (O_1750,N_14998,N_14861);
and UO_1751 (O_1751,N_14899,N_14909);
and UO_1752 (O_1752,N_14930,N_14961);
or UO_1753 (O_1753,N_14911,N_14936);
or UO_1754 (O_1754,N_14943,N_14950);
and UO_1755 (O_1755,N_14901,N_14908);
nand UO_1756 (O_1756,N_14916,N_14869);
and UO_1757 (O_1757,N_14883,N_14910);
nand UO_1758 (O_1758,N_14965,N_14982);
nand UO_1759 (O_1759,N_14968,N_14960);
or UO_1760 (O_1760,N_14942,N_14985);
and UO_1761 (O_1761,N_14905,N_14994);
nand UO_1762 (O_1762,N_14969,N_14937);
and UO_1763 (O_1763,N_14901,N_14941);
nand UO_1764 (O_1764,N_14999,N_14888);
nor UO_1765 (O_1765,N_14892,N_14851);
or UO_1766 (O_1766,N_14909,N_14891);
and UO_1767 (O_1767,N_14991,N_14939);
and UO_1768 (O_1768,N_14873,N_14899);
or UO_1769 (O_1769,N_14989,N_14947);
or UO_1770 (O_1770,N_14971,N_14905);
and UO_1771 (O_1771,N_14978,N_14932);
and UO_1772 (O_1772,N_14970,N_14920);
nand UO_1773 (O_1773,N_14998,N_14988);
nor UO_1774 (O_1774,N_14997,N_14980);
nor UO_1775 (O_1775,N_14859,N_14902);
or UO_1776 (O_1776,N_14911,N_14894);
and UO_1777 (O_1777,N_14852,N_14954);
nor UO_1778 (O_1778,N_14913,N_14890);
or UO_1779 (O_1779,N_14961,N_14933);
nor UO_1780 (O_1780,N_14982,N_14981);
or UO_1781 (O_1781,N_14917,N_14868);
or UO_1782 (O_1782,N_14983,N_14955);
nor UO_1783 (O_1783,N_14910,N_14997);
and UO_1784 (O_1784,N_14999,N_14954);
or UO_1785 (O_1785,N_14975,N_14970);
and UO_1786 (O_1786,N_14922,N_14948);
and UO_1787 (O_1787,N_14907,N_14959);
and UO_1788 (O_1788,N_14990,N_14971);
nand UO_1789 (O_1789,N_14991,N_14866);
xnor UO_1790 (O_1790,N_14873,N_14995);
or UO_1791 (O_1791,N_14973,N_14907);
and UO_1792 (O_1792,N_14991,N_14943);
xnor UO_1793 (O_1793,N_14940,N_14851);
nor UO_1794 (O_1794,N_14880,N_14866);
nor UO_1795 (O_1795,N_14870,N_14997);
nand UO_1796 (O_1796,N_14920,N_14898);
nor UO_1797 (O_1797,N_14985,N_14933);
or UO_1798 (O_1798,N_14901,N_14939);
nand UO_1799 (O_1799,N_14965,N_14916);
xnor UO_1800 (O_1800,N_14978,N_14922);
and UO_1801 (O_1801,N_14941,N_14998);
and UO_1802 (O_1802,N_14897,N_14852);
xor UO_1803 (O_1803,N_14957,N_14914);
xor UO_1804 (O_1804,N_14885,N_14939);
nor UO_1805 (O_1805,N_14870,N_14964);
xor UO_1806 (O_1806,N_14915,N_14935);
nand UO_1807 (O_1807,N_14858,N_14987);
or UO_1808 (O_1808,N_14990,N_14942);
or UO_1809 (O_1809,N_14910,N_14918);
and UO_1810 (O_1810,N_14924,N_14972);
nor UO_1811 (O_1811,N_14911,N_14914);
xor UO_1812 (O_1812,N_14895,N_14954);
nand UO_1813 (O_1813,N_14864,N_14853);
nor UO_1814 (O_1814,N_14998,N_14906);
xnor UO_1815 (O_1815,N_14977,N_14972);
xnor UO_1816 (O_1816,N_14866,N_14996);
xnor UO_1817 (O_1817,N_14875,N_14883);
nand UO_1818 (O_1818,N_14878,N_14949);
nand UO_1819 (O_1819,N_14920,N_14940);
and UO_1820 (O_1820,N_14924,N_14923);
and UO_1821 (O_1821,N_14969,N_14870);
and UO_1822 (O_1822,N_14926,N_14931);
or UO_1823 (O_1823,N_14852,N_14931);
xor UO_1824 (O_1824,N_14967,N_14933);
and UO_1825 (O_1825,N_14969,N_14919);
nand UO_1826 (O_1826,N_14982,N_14865);
and UO_1827 (O_1827,N_14898,N_14899);
nand UO_1828 (O_1828,N_14957,N_14941);
or UO_1829 (O_1829,N_14867,N_14983);
and UO_1830 (O_1830,N_14937,N_14947);
nor UO_1831 (O_1831,N_14913,N_14949);
or UO_1832 (O_1832,N_14964,N_14980);
nand UO_1833 (O_1833,N_14995,N_14937);
or UO_1834 (O_1834,N_14978,N_14886);
xnor UO_1835 (O_1835,N_14956,N_14905);
nand UO_1836 (O_1836,N_14903,N_14886);
nor UO_1837 (O_1837,N_14955,N_14893);
or UO_1838 (O_1838,N_14911,N_14908);
or UO_1839 (O_1839,N_14919,N_14985);
or UO_1840 (O_1840,N_14958,N_14976);
nand UO_1841 (O_1841,N_14866,N_14864);
nand UO_1842 (O_1842,N_14896,N_14947);
xor UO_1843 (O_1843,N_14932,N_14966);
or UO_1844 (O_1844,N_14894,N_14956);
nor UO_1845 (O_1845,N_14881,N_14872);
nor UO_1846 (O_1846,N_14886,N_14859);
nor UO_1847 (O_1847,N_14989,N_14860);
nor UO_1848 (O_1848,N_14915,N_14925);
nand UO_1849 (O_1849,N_14877,N_14917);
nand UO_1850 (O_1850,N_14865,N_14951);
or UO_1851 (O_1851,N_14969,N_14962);
xnor UO_1852 (O_1852,N_14927,N_14908);
and UO_1853 (O_1853,N_14880,N_14887);
xnor UO_1854 (O_1854,N_14937,N_14858);
and UO_1855 (O_1855,N_14882,N_14852);
xnor UO_1856 (O_1856,N_14999,N_14856);
and UO_1857 (O_1857,N_14870,N_14864);
nor UO_1858 (O_1858,N_14941,N_14896);
xnor UO_1859 (O_1859,N_14987,N_14853);
nand UO_1860 (O_1860,N_14914,N_14956);
and UO_1861 (O_1861,N_14981,N_14899);
nor UO_1862 (O_1862,N_14999,N_14904);
xnor UO_1863 (O_1863,N_14927,N_14923);
and UO_1864 (O_1864,N_14970,N_14897);
nand UO_1865 (O_1865,N_14914,N_14961);
nor UO_1866 (O_1866,N_14895,N_14971);
xor UO_1867 (O_1867,N_14925,N_14990);
or UO_1868 (O_1868,N_14998,N_14875);
xnor UO_1869 (O_1869,N_14982,N_14901);
nor UO_1870 (O_1870,N_14880,N_14983);
xnor UO_1871 (O_1871,N_14923,N_14941);
nand UO_1872 (O_1872,N_14899,N_14931);
xor UO_1873 (O_1873,N_14924,N_14859);
xor UO_1874 (O_1874,N_14863,N_14877);
nor UO_1875 (O_1875,N_14999,N_14960);
or UO_1876 (O_1876,N_14992,N_14872);
nor UO_1877 (O_1877,N_14993,N_14984);
nor UO_1878 (O_1878,N_14916,N_14882);
nor UO_1879 (O_1879,N_14893,N_14897);
xnor UO_1880 (O_1880,N_14969,N_14972);
nor UO_1881 (O_1881,N_14949,N_14989);
nand UO_1882 (O_1882,N_14977,N_14950);
or UO_1883 (O_1883,N_14979,N_14902);
xnor UO_1884 (O_1884,N_14977,N_14923);
xor UO_1885 (O_1885,N_14954,N_14978);
or UO_1886 (O_1886,N_14919,N_14900);
nand UO_1887 (O_1887,N_14988,N_14897);
or UO_1888 (O_1888,N_14990,N_14886);
or UO_1889 (O_1889,N_14904,N_14989);
xnor UO_1890 (O_1890,N_14964,N_14927);
nor UO_1891 (O_1891,N_14851,N_14926);
nor UO_1892 (O_1892,N_14964,N_14889);
or UO_1893 (O_1893,N_14998,N_14950);
or UO_1894 (O_1894,N_14975,N_14898);
nand UO_1895 (O_1895,N_14902,N_14950);
nor UO_1896 (O_1896,N_14863,N_14951);
and UO_1897 (O_1897,N_14881,N_14999);
nor UO_1898 (O_1898,N_14969,N_14940);
xnor UO_1899 (O_1899,N_14870,N_14992);
xor UO_1900 (O_1900,N_14932,N_14876);
or UO_1901 (O_1901,N_14855,N_14917);
xnor UO_1902 (O_1902,N_14911,N_14860);
nand UO_1903 (O_1903,N_14929,N_14972);
nor UO_1904 (O_1904,N_14942,N_14991);
nand UO_1905 (O_1905,N_14955,N_14891);
and UO_1906 (O_1906,N_14978,N_14865);
nand UO_1907 (O_1907,N_14978,N_14983);
nand UO_1908 (O_1908,N_14909,N_14910);
xor UO_1909 (O_1909,N_14862,N_14928);
xor UO_1910 (O_1910,N_14988,N_14973);
nor UO_1911 (O_1911,N_14873,N_14865);
or UO_1912 (O_1912,N_14862,N_14933);
xor UO_1913 (O_1913,N_14963,N_14869);
nand UO_1914 (O_1914,N_14930,N_14999);
nor UO_1915 (O_1915,N_14963,N_14907);
nand UO_1916 (O_1916,N_14882,N_14958);
xnor UO_1917 (O_1917,N_14997,N_14922);
xnor UO_1918 (O_1918,N_14873,N_14850);
xnor UO_1919 (O_1919,N_14918,N_14900);
nand UO_1920 (O_1920,N_14944,N_14992);
nor UO_1921 (O_1921,N_14859,N_14933);
nand UO_1922 (O_1922,N_14976,N_14977);
nor UO_1923 (O_1923,N_14909,N_14888);
nand UO_1924 (O_1924,N_14877,N_14918);
nand UO_1925 (O_1925,N_14951,N_14945);
and UO_1926 (O_1926,N_14965,N_14909);
xor UO_1927 (O_1927,N_14917,N_14862);
or UO_1928 (O_1928,N_14992,N_14901);
and UO_1929 (O_1929,N_14933,N_14923);
or UO_1930 (O_1930,N_14889,N_14922);
nor UO_1931 (O_1931,N_14853,N_14878);
nand UO_1932 (O_1932,N_14906,N_14987);
or UO_1933 (O_1933,N_14964,N_14984);
xor UO_1934 (O_1934,N_14895,N_14981);
or UO_1935 (O_1935,N_14880,N_14867);
and UO_1936 (O_1936,N_14888,N_14954);
nor UO_1937 (O_1937,N_14851,N_14904);
and UO_1938 (O_1938,N_14976,N_14879);
and UO_1939 (O_1939,N_14993,N_14878);
nor UO_1940 (O_1940,N_14924,N_14968);
and UO_1941 (O_1941,N_14871,N_14948);
or UO_1942 (O_1942,N_14900,N_14886);
xor UO_1943 (O_1943,N_14897,N_14964);
xor UO_1944 (O_1944,N_14907,N_14935);
and UO_1945 (O_1945,N_14943,N_14870);
nand UO_1946 (O_1946,N_14954,N_14894);
and UO_1947 (O_1947,N_14950,N_14859);
or UO_1948 (O_1948,N_14926,N_14983);
nor UO_1949 (O_1949,N_14949,N_14865);
nand UO_1950 (O_1950,N_14867,N_14951);
nand UO_1951 (O_1951,N_14923,N_14882);
nor UO_1952 (O_1952,N_14946,N_14997);
or UO_1953 (O_1953,N_14995,N_14908);
or UO_1954 (O_1954,N_14861,N_14901);
nand UO_1955 (O_1955,N_14999,N_14936);
or UO_1956 (O_1956,N_14890,N_14889);
xor UO_1957 (O_1957,N_14871,N_14930);
nor UO_1958 (O_1958,N_14971,N_14850);
nand UO_1959 (O_1959,N_14983,N_14952);
or UO_1960 (O_1960,N_14869,N_14957);
and UO_1961 (O_1961,N_14917,N_14938);
and UO_1962 (O_1962,N_14905,N_14966);
or UO_1963 (O_1963,N_14872,N_14977);
xnor UO_1964 (O_1964,N_14946,N_14913);
or UO_1965 (O_1965,N_14938,N_14968);
xor UO_1966 (O_1966,N_14915,N_14924);
and UO_1967 (O_1967,N_14895,N_14935);
and UO_1968 (O_1968,N_14893,N_14901);
xor UO_1969 (O_1969,N_14981,N_14930);
nand UO_1970 (O_1970,N_14898,N_14900);
and UO_1971 (O_1971,N_14930,N_14976);
and UO_1972 (O_1972,N_14954,N_14866);
nor UO_1973 (O_1973,N_14925,N_14894);
xor UO_1974 (O_1974,N_14924,N_14967);
or UO_1975 (O_1975,N_14951,N_14925);
and UO_1976 (O_1976,N_14867,N_14860);
and UO_1977 (O_1977,N_14960,N_14854);
or UO_1978 (O_1978,N_14912,N_14965);
xor UO_1979 (O_1979,N_14998,N_14926);
xor UO_1980 (O_1980,N_14936,N_14978);
and UO_1981 (O_1981,N_14938,N_14960);
nor UO_1982 (O_1982,N_14924,N_14984);
xor UO_1983 (O_1983,N_14856,N_14870);
or UO_1984 (O_1984,N_14928,N_14909);
and UO_1985 (O_1985,N_14905,N_14888);
and UO_1986 (O_1986,N_14928,N_14868);
and UO_1987 (O_1987,N_14981,N_14897);
or UO_1988 (O_1988,N_14945,N_14874);
and UO_1989 (O_1989,N_14957,N_14909);
xor UO_1990 (O_1990,N_14945,N_14898);
nand UO_1991 (O_1991,N_14899,N_14906);
xnor UO_1992 (O_1992,N_14933,N_14865);
and UO_1993 (O_1993,N_14952,N_14933);
xnor UO_1994 (O_1994,N_14945,N_14908);
nor UO_1995 (O_1995,N_14887,N_14967);
nand UO_1996 (O_1996,N_14867,N_14904);
xor UO_1997 (O_1997,N_14878,N_14911);
or UO_1998 (O_1998,N_14855,N_14918);
nor UO_1999 (O_1999,N_14916,N_14912);
endmodule