module basic_500_3000_500_6_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_234,In_32);
and U1 (N_1,In_307,In_300);
and U2 (N_2,In_382,In_355);
and U3 (N_3,In_36,In_44);
nor U4 (N_4,In_365,In_281);
nand U5 (N_5,In_453,In_169);
nor U6 (N_6,In_127,In_384);
nand U7 (N_7,In_261,In_470);
and U8 (N_8,In_130,In_323);
nand U9 (N_9,In_478,In_195);
nor U10 (N_10,In_396,In_487);
or U11 (N_11,In_143,In_97);
nand U12 (N_12,In_499,In_353);
nor U13 (N_13,In_344,In_229);
or U14 (N_14,In_406,In_188);
and U15 (N_15,In_171,In_274);
and U16 (N_16,In_456,In_479);
or U17 (N_17,In_463,In_179);
or U18 (N_18,In_400,In_175);
nand U19 (N_19,In_40,In_139);
nand U20 (N_20,In_318,In_420);
nor U21 (N_21,In_118,In_152);
nor U22 (N_22,In_245,In_460);
nand U23 (N_23,In_391,In_451);
nand U24 (N_24,In_23,In_297);
or U25 (N_25,In_96,In_208);
or U26 (N_26,In_220,In_122);
nor U27 (N_27,In_256,In_452);
nand U28 (N_28,In_407,In_393);
nor U29 (N_29,In_343,In_54);
or U30 (N_30,In_434,In_81);
xnor U31 (N_31,In_136,In_285);
or U32 (N_32,In_277,In_445);
or U33 (N_33,In_295,In_93);
and U34 (N_34,In_283,In_103);
nand U35 (N_35,In_123,In_383);
or U36 (N_36,In_217,In_207);
and U37 (N_37,In_429,In_278);
and U38 (N_38,In_158,In_153);
nor U39 (N_39,In_101,In_498);
nor U40 (N_40,In_329,In_259);
nand U41 (N_41,In_430,In_227);
and U42 (N_42,In_338,In_233);
or U43 (N_43,In_141,In_110);
nand U44 (N_44,In_161,In_174);
or U45 (N_45,In_299,In_155);
and U46 (N_46,In_399,In_372);
or U47 (N_47,In_120,In_409);
xnor U48 (N_48,In_362,In_66);
nor U49 (N_49,In_346,In_380);
nand U50 (N_50,In_211,In_405);
nand U51 (N_51,In_45,In_444);
and U52 (N_52,In_13,In_454);
nor U53 (N_53,In_337,In_388);
nand U54 (N_54,In_25,In_48);
or U55 (N_55,In_417,In_342);
or U56 (N_56,In_176,In_357);
nand U57 (N_57,In_328,In_241);
or U58 (N_58,In_270,In_92);
nand U59 (N_59,In_128,In_121);
and U60 (N_60,In_472,In_116);
nand U61 (N_61,In_293,In_30);
nand U62 (N_62,In_288,In_154);
and U63 (N_63,In_77,In_471);
and U64 (N_64,In_401,In_126);
nor U65 (N_65,In_332,In_247);
and U66 (N_66,In_1,In_68);
and U67 (N_67,In_351,In_137);
or U68 (N_68,In_19,In_146);
nor U69 (N_69,In_0,In_482);
nand U70 (N_70,In_381,In_199);
or U71 (N_71,In_273,In_361);
or U72 (N_72,In_100,In_63);
or U73 (N_73,In_474,In_2);
or U74 (N_74,In_115,In_484);
or U75 (N_75,In_99,In_242);
and U76 (N_76,In_119,In_157);
or U77 (N_77,In_373,In_201);
and U78 (N_78,In_258,In_308);
or U79 (N_79,In_431,In_87);
and U80 (N_80,In_62,In_438);
and U81 (N_81,In_240,In_186);
nand U82 (N_82,In_184,In_348);
or U83 (N_83,In_224,In_8);
or U84 (N_84,In_398,In_10);
nor U85 (N_85,In_330,In_428);
and U86 (N_86,In_282,In_410);
nor U87 (N_87,In_422,In_341);
nand U88 (N_88,In_279,In_483);
or U89 (N_89,In_271,In_289);
and U90 (N_90,In_378,In_440);
and U91 (N_91,In_53,In_339);
nand U92 (N_92,In_39,In_156);
nand U93 (N_93,In_491,In_371);
or U94 (N_94,In_243,In_73);
or U95 (N_95,In_497,In_476);
nor U96 (N_96,In_395,In_272);
nor U97 (N_97,In_38,In_57);
or U98 (N_98,In_284,In_369);
and U99 (N_99,In_26,In_427);
and U100 (N_100,In_455,In_166);
and U101 (N_101,In_292,In_244);
nand U102 (N_102,In_345,In_140);
nand U103 (N_103,In_204,In_206);
nor U104 (N_104,In_350,In_263);
nor U105 (N_105,In_327,In_102);
nand U106 (N_106,In_11,In_433);
nor U107 (N_107,In_88,In_90);
or U108 (N_108,In_210,In_200);
or U109 (N_109,In_326,In_34);
nand U110 (N_110,In_192,In_370);
nor U111 (N_111,In_402,In_82);
nand U112 (N_112,In_219,In_173);
nand U113 (N_113,In_182,In_276);
or U114 (N_114,In_132,In_55);
and U115 (N_115,In_397,In_421);
or U116 (N_116,In_253,In_251);
or U117 (N_117,In_58,In_449);
or U118 (N_118,In_91,In_333);
nand U119 (N_119,In_213,In_321);
nor U120 (N_120,In_22,In_267);
nor U121 (N_121,In_481,In_492);
nor U122 (N_122,In_203,In_108);
or U123 (N_123,In_309,In_266);
and U124 (N_124,In_84,In_368);
nor U125 (N_125,In_262,In_390);
or U126 (N_126,In_467,In_113);
nor U127 (N_127,In_469,In_67);
and U128 (N_128,In_79,In_360);
nand U129 (N_129,In_458,In_268);
and U130 (N_130,In_107,In_163);
and U131 (N_131,In_43,In_86);
nand U132 (N_132,In_59,In_56);
nor U133 (N_133,In_376,In_95);
and U134 (N_134,In_112,In_74);
nor U135 (N_135,In_144,In_159);
or U136 (N_136,In_49,In_218);
or U137 (N_137,In_425,In_117);
and U138 (N_138,In_465,In_486);
or U139 (N_139,In_435,In_183);
or U140 (N_140,In_364,In_291);
nor U141 (N_141,In_94,In_457);
nor U142 (N_142,In_109,In_215);
or U143 (N_143,In_387,In_489);
nand U144 (N_144,In_28,In_172);
and U145 (N_145,In_269,In_7);
or U146 (N_146,In_325,In_488);
nand U147 (N_147,In_237,In_15);
or U148 (N_148,In_375,In_314);
nor U149 (N_149,In_374,In_89);
nand U150 (N_150,In_287,In_131);
and U151 (N_151,In_392,In_441);
nor U152 (N_152,In_302,In_104);
or U153 (N_153,In_347,In_177);
and U154 (N_154,In_459,In_150);
nor U155 (N_155,In_490,In_65);
nand U156 (N_156,In_443,In_47);
and U157 (N_157,In_191,In_187);
and U158 (N_158,In_304,In_496);
and U159 (N_159,In_138,In_423);
nor U160 (N_160,In_209,In_27);
or U161 (N_161,In_148,In_125);
nor U162 (N_162,In_14,In_411);
and U163 (N_163,In_305,In_35);
nor U164 (N_164,In_151,In_301);
nand U165 (N_165,In_389,In_167);
and U166 (N_166,In_133,In_322);
and U167 (N_167,In_303,In_290);
nand U168 (N_168,In_260,In_31);
nor U169 (N_169,In_468,In_228);
nor U170 (N_170,In_239,In_439);
and U171 (N_171,In_466,In_358);
and U172 (N_172,In_377,In_248);
nand U173 (N_173,In_356,In_462);
and U174 (N_174,In_394,In_379);
nand U175 (N_175,In_16,In_60);
and U176 (N_176,In_20,In_147);
xor U177 (N_177,In_464,In_250);
or U178 (N_178,In_331,In_76);
and U179 (N_179,In_461,In_419);
or U180 (N_180,In_72,In_349);
nor U181 (N_181,In_29,In_178);
and U182 (N_182,In_216,In_414);
and U183 (N_183,In_42,In_316);
and U184 (N_184,In_189,In_142);
nor U185 (N_185,In_426,In_75);
nand U186 (N_186,In_46,In_418);
or U187 (N_187,In_145,In_315);
nor U188 (N_188,In_223,In_231);
and U189 (N_189,In_447,In_286);
nor U190 (N_190,In_298,In_185);
nand U191 (N_191,In_225,In_311);
and U192 (N_192,In_5,In_106);
or U193 (N_193,In_275,In_352);
and U194 (N_194,In_129,In_181);
nor U195 (N_195,In_164,In_255);
nor U196 (N_196,In_437,In_124);
or U197 (N_197,In_485,In_264);
nor U198 (N_198,In_236,In_312);
nor U199 (N_199,In_385,In_69);
and U200 (N_200,In_111,In_359);
or U201 (N_201,In_162,In_98);
nor U202 (N_202,In_12,In_412);
nand U203 (N_203,In_477,In_252);
nor U204 (N_204,In_473,In_50);
nor U205 (N_205,In_408,In_70);
nand U206 (N_206,In_340,In_37);
nand U207 (N_207,In_17,In_80);
or U208 (N_208,In_18,In_202);
nand U209 (N_209,In_403,In_436);
nor U210 (N_210,In_190,In_114);
nor U211 (N_211,In_9,In_363);
or U212 (N_212,In_212,In_180);
nand U213 (N_213,In_249,In_85);
nand U214 (N_214,In_366,In_222);
and U215 (N_215,In_221,In_24);
nor U216 (N_216,In_257,In_165);
or U217 (N_217,In_51,In_254);
or U218 (N_218,In_230,In_196);
nand U219 (N_219,In_306,In_442);
or U220 (N_220,In_367,In_493);
and U221 (N_221,In_448,In_480);
or U222 (N_222,In_280,In_194);
nor U223 (N_223,In_238,In_386);
nand U224 (N_224,In_41,In_6);
nand U225 (N_225,In_170,In_416);
and U226 (N_226,In_83,In_294);
and U227 (N_227,In_324,In_475);
or U228 (N_228,In_71,In_334);
and U229 (N_229,In_317,In_235);
nand U230 (N_230,In_446,In_52);
and U231 (N_231,In_160,In_64);
and U232 (N_232,In_354,In_21);
or U233 (N_233,In_197,In_3);
and U234 (N_234,In_336,In_320);
and U235 (N_235,In_413,In_424);
or U236 (N_236,In_246,In_135);
nor U237 (N_237,In_4,In_33);
or U238 (N_238,In_265,In_313);
or U239 (N_239,In_198,In_78);
nor U240 (N_240,In_319,In_494);
or U241 (N_241,In_226,In_134);
or U242 (N_242,In_149,In_495);
nor U243 (N_243,In_205,In_296);
or U244 (N_244,In_404,In_415);
and U245 (N_245,In_232,In_105);
and U246 (N_246,In_193,In_214);
nand U247 (N_247,In_432,In_61);
or U248 (N_248,In_310,In_450);
or U249 (N_249,In_168,In_335);
nor U250 (N_250,In_348,In_386);
or U251 (N_251,In_497,In_33);
or U252 (N_252,In_206,In_464);
or U253 (N_253,In_358,In_291);
nor U254 (N_254,In_313,In_21);
nand U255 (N_255,In_468,In_203);
nand U256 (N_256,In_292,In_448);
and U257 (N_257,In_84,In_47);
or U258 (N_258,In_411,In_164);
nor U259 (N_259,In_360,In_4);
nor U260 (N_260,In_258,In_65);
nand U261 (N_261,In_375,In_426);
nand U262 (N_262,In_21,In_77);
and U263 (N_263,In_469,In_60);
nand U264 (N_264,In_132,In_343);
or U265 (N_265,In_251,In_234);
or U266 (N_266,In_230,In_306);
and U267 (N_267,In_362,In_493);
nand U268 (N_268,In_246,In_380);
nand U269 (N_269,In_279,In_11);
nand U270 (N_270,In_289,In_346);
or U271 (N_271,In_44,In_282);
nor U272 (N_272,In_231,In_492);
nor U273 (N_273,In_309,In_317);
nor U274 (N_274,In_56,In_97);
nor U275 (N_275,In_5,In_166);
nand U276 (N_276,In_439,In_271);
and U277 (N_277,In_98,In_317);
and U278 (N_278,In_468,In_440);
nand U279 (N_279,In_361,In_142);
nor U280 (N_280,In_310,In_300);
and U281 (N_281,In_393,In_259);
or U282 (N_282,In_183,In_322);
nor U283 (N_283,In_210,In_389);
nand U284 (N_284,In_409,In_363);
nand U285 (N_285,In_112,In_228);
nand U286 (N_286,In_45,In_254);
or U287 (N_287,In_79,In_480);
and U288 (N_288,In_397,In_197);
nand U289 (N_289,In_62,In_55);
nor U290 (N_290,In_235,In_52);
and U291 (N_291,In_404,In_467);
or U292 (N_292,In_303,In_443);
nor U293 (N_293,In_326,In_192);
nand U294 (N_294,In_157,In_495);
and U295 (N_295,In_19,In_412);
nand U296 (N_296,In_29,In_59);
nor U297 (N_297,In_424,In_415);
nand U298 (N_298,In_240,In_112);
or U299 (N_299,In_469,In_193);
and U300 (N_300,In_398,In_126);
or U301 (N_301,In_322,In_1);
nand U302 (N_302,In_26,In_364);
nor U303 (N_303,In_15,In_279);
nand U304 (N_304,In_253,In_454);
nand U305 (N_305,In_445,In_105);
and U306 (N_306,In_59,In_319);
or U307 (N_307,In_308,In_180);
xor U308 (N_308,In_95,In_208);
or U309 (N_309,In_312,In_132);
nor U310 (N_310,In_321,In_441);
and U311 (N_311,In_408,In_358);
nand U312 (N_312,In_280,In_248);
nor U313 (N_313,In_378,In_102);
and U314 (N_314,In_442,In_223);
nand U315 (N_315,In_9,In_7);
nand U316 (N_316,In_98,In_197);
and U317 (N_317,In_42,In_78);
and U318 (N_318,In_281,In_369);
or U319 (N_319,In_468,In_59);
nor U320 (N_320,In_294,In_487);
nand U321 (N_321,In_414,In_260);
nand U322 (N_322,In_30,In_257);
nor U323 (N_323,In_44,In_131);
and U324 (N_324,In_52,In_34);
and U325 (N_325,In_404,In_16);
nand U326 (N_326,In_446,In_458);
nor U327 (N_327,In_197,In_114);
or U328 (N_328,In_221,In_19);
and U329 (N_329,In_425,In_165);
nor U330 (N_330,In_440,In_382);
or U331 (N_331,In_348,In_61);
nor U332 (N_332,In_459,In_320);
nand U333 (N_333,In_467,In_442);
and U334 (N_334,In_287,In_292);
or U335 (N_335,In_77,In_467);
and U336 (N_336,In_225,In_60);
nor U337 (N_337,In_447,In_143);
nor U338 (N_338,In_177,In_166);
and U339 (N_339,In_434,In_171);
or U340 (N_340,In_257,In_408);
nor U341 (N_341,In_316,In_467);
nor U342 (N_342,In_438,In_157);
nand U343 (N_343,In_43,In_409);
nor U344 (N_344,In_125,In_329);
xnor U345 (N_345,In_320,In_283);
and U346 (N_346,In_284,In_438);
nand U347 (N_347,In_13,In_48);
or U348 (N_348,In_25,In_267);
nand U349 (N_349,In_175,In_247);
and U350 (N_350,In_336,In_319);
or U351 (N_351,In_250,In_160);
and U352 (N_352,In_22,In_89);
or U353 (N_353,In_317,In_465);
and U354 (N_354,In_301,In_186);
nand U355 (N_355,In_16,In_67);
nand U356 (N_356,In_51,In_94);
nor U357 (N_357,In_465,In_403);
and U358 (N_358,In_229,In_166);
or U359 (N_359,In_451,In_431);
and U360 (N_360,In_25,In_57);
nand U361 (N_361,In_282,In_231);
and U362 (N_362,In_305,In_194);
nor U363 (N_363,In_93,In_298);
nor U364 (N_364,In_459,In_371);
nor U365 (N_365,In_64,In_49);
or U366 (N_366,In_223,In_199);
nand U367 (N_367,In_295,In_225);
and U368 (N_368,In_151,In_209);
and U369 (N_369,In_18,In_62);
and U370 (N_370,In_297,In_150);
and U371 (N_371,In_133,In_363);
or U372 (N_372,In_281,In_77);
or U373 (N_373,In_71,In_110);
nor U374 (N_374,In_149,In_0);
or U375 (N_375,In_257,In_205);
nand U376 (N_376,In_126,In_344);
nand U377 (N_377,In_308,In_202);
and U378 (N_378,In_489,In_113);
or U379 (N_379,In_303,In_366);
nor U380 (N_380,In_252,In_8);
or U381 (N_381,In_300,In_36);
nand U382 (N_382,In_363,In_281);
or U383 (N_383,In_253,In_60);
nor U384 (N_384,In_156,In_412);
nor U385 (N_385,In_286,In_467);
or U386 (N_386,In_485,In_405);
or U387 (N_387,In_37,In_230);
nand U388 (N_388,In_65,In_395);
and U389 (N_389,In_290,In_142);
or U390 (N_390,In_457,In_204);
nor U391 (N_391,In_310,In_46);
or U392 (N_392,In_356,In_282);
nor U393 (N_393,In_172,In_191);
or U394 (N_394,In_185,In_309);
and U395 (N_395,In_492,In_488);
or U396 (N_396,In_18,In_107);
nor U397 (N_397,In_125,In_330);
or U398 (N_398,In_227,In_38);
nand U399 (N_399,In_290,In_413);
or U400 (N_400,In_128,In_22);
nor U401 (N_401,In_198,In_318);
or U402 (N_402,In_461,In_412);
and U403 (N_403,In_320,In_400);
or U404 (N_404,In_146,In_211);
nand U405 (N_405,In_60,In_398);
nand U406 (N_406,In_405,In_406);
and U407 (N_407,In_234,In_296);
or U408 (N_408,In_198,In_427);
or U409 (N_409,In_164,In_129);
and U410 (N_410,In_102,In_268);
or U411 (N_411,In_344,In_57);
and U412 (N_412,In_371,In_227);
and U413 (N_413,In_206,In_144);
nand U414 (N_414,In_256,In_434);
and U415 (N_415,In_93,In_15);
and U416 (N_416,In_225,In_237);
nor U417 (N_417,In_154,In_65);
or U418 (N_418,In_447,In_303);
nor U419 (N_419,In_249,In_353);
nor U420 (N_420,In_96,In_452);
nor U421 (N_421,In_341,In_15);
nand U422 (N_422,In_110,In_360);
nor U423 (N_423,In_412,In_370);
nor U424 (N_424,In_457,In_165);
nor U425 (N_425,In_223,In_406);
or U426 (N_426,In_360,In_365);
and U427 (N_427,In_176,In_8);
and U428 (N_428,In_264,In_338);
and U429 (N_429,In_299,In_151);
nand U430 (N_430,In_480,In_357);
and U431 (N_431,In_417,In_293);
or U432 (N_432,In_452,In_355);
and U433 (N_433,In_360,In_447);
nor U434 (N_434,In_435,In_150);
or U435 (N_435,In_178,In_271);
and U436 (N_436,In_385,In_130);
and U437 (N_437,In_16,In_15);
and U438 (N_438,In_258,In_334);
nor U439 (N_439,In_208,In_103);
nor U440 (N_440,In_439,In_205);
and U441 (N_441,In_107,In_337);
nor U442 (N_442,In_416,In_246);
xnor U443 (N_443,In_195,In_446);
and U444 (N_444,In_227,In_191);
or U445 (N_445,In_280,In_335);
or U446 (N_446,In_483,In_12);
or U447 (N_447,In_231,In_102);
or U448 (N_448,In_73,In_47);
or U449 (N_449,In_242,In_155);
xor U450 (N_450,In_9,In_298);
nor U451 (N_451,In_365,In_379);
nand U452 (N_452,In_426,In_149);
and U453 (N_453,In_455,In_228);
nand U454 (N_454,In_345,In_184);
nor U455 (N_455,In_489,In_134);
nand U456 (N_456,In_476,In_147);
nor U457 (N_457,In_445,In_457);
and U458 (N_458,In_214,In_211);
or U459 (N_459,In_304,In_449);
nand U460 (N_460,In_74,In_376);
nor U461 (N_461,In_466,In_278);
or U462 (N_462,In_265,In_139);
nand U463 (N_463,In_73,In_300);
nand U464 (N_464,In_186,In_428);
or U465 (N_465,In_270,In_285);
or U466 (N_466,In_277,In_43);
nand U467 (N_467,In_192,In_327);
and U468 (N_468,In_433,In_113);
and U469 (N_469,In_77,In_197);
or U470 (N_470,In_217,In_320);
nor U471 (N_471,In_160,In_364);
or U472 (N_472,In_244,In_282);
or U473 (N_473,In_495,In_406);
nand U474 (N_474,In_443,In_199);
or U475 (N_475,In_402,In_384);
nor U476 (N_476,In_295,In_208);
nor U477 (N_477,In_324,In_347);
and U478 (N_478,In_421,In_38);
and U479 (N_479,In_4,In_234);
and U480 (N_480,In_55,In_66);
or U481 (N_481,In_488,In_494);
and U482 (N_482,In_462,In_304);
nor U483 (N_483,In_38,In_327);
or U484 (N_484,In_110,In_349);
and U485 (N_485,In_85,In_21);
nor U486 (N_486,In_16,In_129);
or U487 (N_487,In_207,In_392);
or U488 (N_488,In_216,In_171);
nor U489 (N_489,In_495,In_128);
nor U490 (N_490,In_350,In_101);
and U491 (N_491,In_366,In_460);
xor U492 (N_492,In_133,In_47);
and U493 (N_493,In_261,In_298);
or U494 (N_494,In_411,In_388);
or U495 (N_495,In_291,In_246);
and U496 (N_496,In_437,In_54);
or U497 (N_497,In_186,In_257);
nand U498 (N_498,In_88,In_454);
and U499 (N_499,In_129,In_249);
nor U500 (N_500,N_209,N_38);
or U501 (N_501,N_473,N_314);
and U502 (N_502,N_238,N_324);
nor U503 (N_503,N_213,N_273);
nor U504 (N_504,N_239,N_150);
or U505 (N_505,N_437,N_191);
nand U506 (N_506,N_403,N_155);
nand U507 (N_507,N_463,N_454);
or U508 (N_508,N_84,N_296);
nand U509 (N_509,N_249,N_250);
nor U510 (N_510,N_363,N_115);
and U511 (N_511,N_147,N_307);
or U512 (N_512,N_393,N_383);
nor U513 (N_513,N_75,N_428);
and U514 (N_514,N_472,N_65);
nor U515 (N_515,N_110,N_76);
nor U516 (N_516,N_229,N_398);
and U517 (N_517,N_64,N_104);
nand U518 (N_518,N_341,N_60);
nor U519 (N_519,N_465,N_170);
xnor U520 (N_520,N_163,N_3);
or U521 (N_521,N_448,N_466);
nor U522 (N_522,N_282,N_156);
nor U523 (N_523,N_131,N_424);
and U524 (N_524,N_72,N_486);
or U525 (N_525,N_196,N_280);
nand U526 (N_526,N_235,N_475);
and U527 (N_527,N_369,N_234);
and U528 (N_528,N_322,N_43);
or U529 (N_529,N_237,N_417);
nor U530 (N_530,N_259,N_394);
xor U531 (N_531,N_294,N_88);
xor U532 (N_532,N_297,N_230);
or U533 (N_533,N_87,N_160);
or U534 (N_534,N_491,N_105);
and U535 (N_535,N_327,N_34);
nor U536 (N_536,N_246,N_21);
and U537 (N_537,N_86,N_319);
nand U538 (N_538,N_128,N_182);
or U539 (N_539,N_467,N_165);
or U540 (N_540,N_323,N_379);
and U541 (N_541,N_114,N_14);
and U542 (N_542,N_103,N_0);
nand U543 (N_543,N_208,N_42);
nor U544 (N_544,N_415,N_405);
or U545 (N_545,N_357,N_350);
nor U546 (N_546,N_412,N_74);
and U547 (N_547,N_248,N_312);
or U548 (N_548,N_227,N_495);
and U549 (N_549,N_427,N_13);
and U550 (N_550,N_391,N_429);
nand U551 (N_551,N_149,N_68);
nor U552 (N_552,N_171,N_489);
nand U553 (N_553,N_245,N_377);
nor U554 (N_554,N_140,N_387);
nand U555 (N_555,N_175,N_368);
nor U556 (N_556,N_49,N_58);
nor U557 (N_557,N_308,N_356);
nand U558 (N_558,N_422,N_57);
nand U559 (N_559,N_108,N_203);
and U560 (N_560,N_301,N_287);
nand U561 (N_561,N_216,N_173);
and U562 (N_562,N_404,N_425);
nand U563 (N_563,N_482,N_284);
nor U564 (N_564,N_408,N_347);
and U565 (N_565,N_263,N_77);
or U566 (N_566,N_154,N_265);
nor U567 (N_567,N_82,N_158);
nand U568 (N_568,N_221,N_313);
nand U569 (N_569,N_143,N_26);
or U570 (N_570,N_242,N_286);
nor U571 (N_571,N_325,N_195);
and U572 (N_572,N_252,N_185);
nand U573 (N_573,N_63,N_254);
or U574 (N_574,N_348,N_7);
or U575 (N_575,N_447,N_187);
nand U576 (N_576,N_397,N_219);
xnor U577 (N_577,N_93,N_362);
or U578 (N_578,N_90,N_339);
and U579 (N_579,N_304,N_6);
nor U580 (N_580,N_162,N_32);
nand U581 (N_581,N_410,N_126);
and U582 (N_582,N_8,N_469);
nand U583 (N_583,N_376,N_320);
and U584 (N_584,N_92,N_443);
and U585 (N_585,N_207,N_311);
nor U586 (N_586,N_251,N_416);
and U587 (N_587,N_27,N_285);
or U588 (N_588,N_420,N_373);
or U589 (N_589,N_25,N_176);
or U590 (N_590,N_432,N_266);
nand U591 (N_591,N_204,N_29);
nand U592 (N_592,N_371,N_241);
nand U593 (N_593,N_134,N_497);
and U594 (N_594,N_411,N_271);
nand U595 (N_595,N_5,N_326);
and U596 (N_596,N_35,N_381);
or U597 (N_597,N_70,N_228);
or U598 (N_598,N_192,N_402);
and U599 (N_599,N_139,N_66);
or U600 (N_600,N_351,N_464);
and U601 (N_601,N_189,N_396);
or U602 (N_602,N_374,N_123);
or U603 (N_603,N_161,N_215);
nor U604 (N_604,N_107,N_353);
and U605 (N_605,N_364,N_367);
and U606 (N_606,N_361,N_109);
or U607 (N_607,N_119,N_168);
or U608 (N_608,N_352,N_380);
or U609 (N_609,N_132,N_283);
nor U610 (N_610,N_253,N_205);
or U611 (N_611,N_455,N_372);
and U612 (N_612,N_384,N_481);
nand U613 (N_613,N_336,N_337);
nor U614 (N_614,N_11,N_55);
nand U615 (N_615,N_487,N_181);
and U616 (N_616,N_483,N_124);
or U617 (N_617,N_365,N_264);
or U618 (N_618,N_51,N_122);
xor U619 (N_619,N_257,N_413);
and U620 (N_620,N_133,N_426);
nor U621 (N_621,N_153,N_40);
or U622 (N_622,N_389,N_210);
or U623 (N_623,N_444,N_125);
or U624 (N_624,N_378,N_451);
nor U625 (N_625,N_449,N_19);
or U626 (N_626,N_97,N_438);
nor U627 (N_627,N_91,N_340);
nand U628 (N_628,N_401,N_180);
xor U629 (N_629,N_95,N_261);
or U630 (N_630,N_256,N_288);
and U631 (N_631,N_289,N_30);
and U632 (N_632,N_355,N_130);
or U633 (N_633,N_146,N_16);
or U634 (N_634,N_36,N_79);
nand U635 (N_635,N_354,N_421);
nand U636 (N_636,N_435,N_338);
or U637 (N_637,N_233,N_275);
nor U638 (N_638,N_419,N_20);
nand U639 (N_639,N_277,N_118);
nand U640 (N_640,N_111,N_452);
or U641 (N_641,N_329,N_212);
nand U642 (N_642,N_445,N_144);
nor U643 (N_643,N_59,N_492);
nand U644 (N_644,N_223,N_12);
nand U645 (N_645,N_457,N_85);
nor U646 (N_646,N_71,N_267);
or U647 (N_647,N_499,N_1);
or U648 (N_648,N_117,N_247);
nor U649 (N_649,N_194,N_61);
nand U650 (N_650,N_120,N_330);
nand U651 (N_651,N_346,N_260);
or U652 (N_652,N_459,N_344);
or U653 (N_653,N_106,N_262);
nand U654 (N_654,N_164,N_218);
and U655 (N_655,N_231,N_332);
or U656 (N_656,N_167,N_309);
or U657 (N_657,N_136,N_485);
and U658 (N_658,N_9,N_81);
and U659 (N_659,N_148,N_206);
nand U660 (N_660,N_98,N_243);
nor U661 (N_661,N_101,N_96);
or U662 (N_662,N_47,N_484);
nand U663 (N_663,N_453,N_462);
and U664 (N_664,N_349,N_39);
or U665 (N_665,N_102,N_135);
nand U666 (N_666,N_15,N_423);
nand U667 (N_667,N_56,N_138);
and U668 (N_668,N_166,N_80);
and U669 (N_669,N_310,N_183);
nand U670 (N_670,N_222,N_316);
nand U671 (N_671,N_331,N_343);
and U672 (N_672,N_468,N_434);
nor U673 (N_673,N_184,N_33);
nor U674 (N_674,N_201,N_305);
nor U675 (N_675,N_112,N_461);
or U676 (N_676,N_137,N_386);
nor U677 (N_677,N_23,N_290);
nand U678 (N_678,N_99,N_450);
nand U679 (N_679,N_276,N_214);
nor U680 (N_680,N_78,N_236);
or U681 (N_681,N_306,N_244);
nor U682 (N_682,N_129,N_441);
nand U683 (N_683,N_18,N_198);
and U684 (N_684,N_50,N_360);
or U685 (N_685,N_328,N_400);
or U686 (N_686,N_321,N_113);
or U687 (N_687,N_159,N_281);
nor U688 (N_688,N_226,N_358);
nor U689 (N_689,N_177,N_318);
or U690 (N_690,N_479,N_295);
nand U691 (N_691,N_291,N_232);
nor U692 (N_692,N_480,N_334);
and U693 (N_693,N_269,N_498);
or U694 (N_694,N_279,N_493);
nand U695 (N_695,N_460,N_418);
or U696 (N_696,N_414,N_151);
nor U697 (N_697,N_385,N_470);
nand U698 (N_698,N_220,N_54);
nor U699 (N_699,N_217,N_24);
and U700 (N_700,N_258,N_382);
or U701 (N_701,N_458,N_433);
or U702 (N_702,N_145,N_188);
or U703 (N_703,N_157,N_240);
nor U704 (N_704,N_292,N_293);
and U705 (N_705,N_268,N_496);
or U706 (N_706,N_333,N_442);
or U707 (N_707,N_89,N_52);
nor U708 (N_708,N_45,N_4);
and U709 (N_709,N_69,N_28);
nor U710 (N_710,N_22,N_17);
and U711 (N_711,N_395,N_174);
nor U712 (N_712,N_488,N_127);
and U713 (N_713,N_270,N_37);
nand U714 (N_714,N_62,N_366);
or U715 (N_715,N_67,N_299);
nor U716 (N_716,N_169,N_478);
nor U717 (N_717,N_141,N_83);
or U718 (N_718,N_121,N_390);
and U719 (N_719,N_456,N_202);
nor U720 (N_720,N_359,N_199);
nor U721 (N_721,N_490,N_494);
and U722 (N_722,N_300,N_477);
nand U723 (N_723,N_116,N_388);
nand U724 (N_724,N_152,N_431);
and U725 (N_725,N_474,N_409);
nand U726 (N_726,N_193,N_446);
and U727 (N_727,N_439,N_53);
nor U728 (N_728,N_46,N_100);
nand U729 (N_729,N_178,N_370);
xor U730 (N_730,N_200,N_476);
and U731 (N_731,N_436,N_41);
nor U732 (N_732,N_211,N_335);
and U733 (N_733,N_302,N_399);
nand U734 (N_734,N_255,N_406);
and U735 (N_735,N_392,N_94);
or U736 (N_736,N_44,N_303);
nand U737 (N_737,N_2,N_430);
nand U738 (N_738,N_224,N_407);
nor U739 (N_739,N_274,N_272);
nand U740 (N_740,N_48,N_197);
or U741 (N_741,N_10,N_342);
and U742 (N_742,N_142,N_315);
and U743 (N_743,N_225,N_317);
and U744 (N_744,N_172,N_73);
and U745 (N_745,N_440,N_179);
nand U746 (N_746,N_186,N_278);
and U747 (N_747,N_190,N_31);
nand U748 (N_748,N_345,N_471);
nand U749 (N_749,N_298,N_375);
nor U750 (N_750,N_137,N_161);
and U751 (N_751,N_451,N_402);
nor U752 (N_752,N_112,N_366);
or U753 (N_753,N_151,N_277);
nand U754 (N_754,N_313,N_372);
nor U755 (N_755,N_59,N_496);
and U756 (N_756,N_192,N_191);
or U757 (N_757,N_200,N_89);
and U758 (N_758,N_170,N_71);
nor U759 (N_759,N_445,N_216);
or U760 (N_760,N_285,N_165);
nand U761 (N_761,N_170,N_155);
or U762 (N_762,N_206,N_236);
or U763 (N_763,N_351,N_357);
nand U764 (N_764,N_381,N_345);
nor U765 (N_765,N_416,N_410);
nand U766 (N_766,N_320,N_452);
nand U767 (N_767,N_143,N_317);
nand U768 (N_768,N_266,N_478);
and U769 (N_769,N_293,N_273);
nor U770 (N_770,N_178,N_420);
nor U771 (N_771,N_16,N_459);
and U772 (N_772,N_115,N_442);
or U773 (N_773,N_10,N_432);
and U774 (N_774,N_405,N_5);
nor U775 (N_775,N_459,N_145);
or U776 (N_776,N_334,N_83);
nor U777 (N_777,N_448,N_355);
nand U778 (N_778,N_478,N_254);
nand U779 (N_779,N_390,N_319);
xnor U780 (N_780,N_244,N_419);
nor U781 (N_781,N_438,N_266);
nor U782 (N_782,N_326,N_379);
nor U783 (N_783,N_259,N_390);
nand U784 (N_784,N_478,N_357);
nand U785 (N_785,N_464,N_342);
or U786 (N_786,N_173,N_244);
nor U787 (N_787,N_118,N_350);
nor U788 (N_788,N_181,N_236);
and U789 (N_789,N_181,N_306);
nor U790 (N_790,N_192,N_461);
nand U791 (N_791,N_3,N_51);
nand U792 (N_792,N_388,N_480);
nor U793 (N_793,N_445,N_463);
and U794 (N_794,N_394,N_377);
nor U795 (N_795,N_291,N_126);
or U796 (N_796,N_120,N_170);
nor U797 (N_797,N_239,N_79);
nand U798 (N_798,N_277,N_120);
or U799 (N_799,N_329,N_84);
nor U800 (N_800,N_7,N_184);
nand U801 (N_801,N_9,N_245);
and U802 (N_802,N_260,N_212);
nor U803 (N_803,N_199,N_312);
nor U804 (N_804,N_439,N_54);
nand U805 (N_805,N_81,N_283);
and U806 (N_806,N_389,N_330);
nor U807 (N_807,N_465,N_250);
nor U808 (N_808,N_27,N_371);
or U809 (N_809,N_419,N_339);
or U810 (N_810,N_262,N_94);
nand U811 (N_811,N_278,N_2);
nand U812 (N_812,N_226,N_491);
nand U813 (N_813,N_436,N_447);
and U814 (N_814,N_351,N_172);
and U815 (N_815,N_126,N_242);
nor U816 (N_816,N_465,N_498);
nand U817 (N_817,N_499,N_27);
and U818 (N_818,N_113,N_481);
nand U819 (N_819,N_154,N_89);
and U820 (N_820,N_204,N_52);
nor U821 (N_821,N_94,N_422);
nor U822 (N_822,N_458,N_482);
nor U823 (N_823,N_430,N_288);
or U824 (N_824,N_202,N_120);
nor U825 (N_825,N_250,N_345);
or U826 (N_826,N_330,N_204);
nand U827 (N_827,N_370,N_334);
or U828 (N_828,N_421,N_162);
and U829 (N_829,N_496,N_266);
or U830 (N_830,N_41,N_112);
or U831 (N_831,N_473,N_170);
or U832 (N_832,N_56,N_86);
or U833 (N_833,N_341,N_346);
and U834 (N_834,N_191,N_21);
or U835 (N_835,N_462,N_374);
or U836 (N_836,N_277,N_191);
nor U837 (N_837,N_491,N_33);
and U838 (N_838,N_479,N_38);
and U839 (N_839,N_367,N_295);
nand U840 (N_840,N_90,N_419);
nor U841 (N_841,N_94,N_159);
nand U842 (N_842,N_369,N_372);
xor U843 (N_843,N_272,N_26);
or U844 (N_844,N_116,N_72);
nand U845 (N_845,N_243,N_186);
nand U846 (N_846,N_468,N_266);
nor U847 (N_847,N_38,N_370);
or U848 (N_848,N_117,N_480);
nand U849 (N_849,N_257,N_32);
nand U850 (N_850,N_216,N_371);
and U851 (N_851,N_46,N_326);
or U852 (N_852,N_30,N_63);
and U853 (N_853,N_429,N_332);
or U854 (N_854,N_189,N_79);
nor U855 (N_855,N_11,N_124);
or U856 (N_856,N_242,N_484);
and U857 (N_857,N_95,N_275);
or U858 (N_858,N_182,N_480);
nor U859 (N_859,N_134,N_165);
xnor U860 (N_860,N_334,N_46);
and U861 (N_861,N_173,N_405);
or U862 (N_862,N_308,N_197);
or U863 (N_863,N_182,N_367);
nor U864 (N_864,N_439,N_377);
nand U865 (N_865,N_246,N_205);
or U866 (N_866,N_132,N_468);
nor U867 (N_867,N_345,N_348);
nor U868 (N_868,N_103,N_347);
nand U869 (N_869,N_326,N_461);
and U870 (N_870,N_482,N_258);
nor U871 (N_871,N_243,N_278);
nor U872 (N_872,N_270,N_128);
nand U873 (N_873,N_224,N_393);
nor U874 (N_874,N_103,N_408);
or U875 (N_875,N_381,N_108);
nand U876 (N_876,N_192,N_295);
or U877 (N_877,N_91,N_176);
and U878 (N_878,N_218,N_202);
or U879 (N_879,N_475,N_297);
and U880 (N_880,N_423,N_272);
nand U881 (N_881,N_476,N_169);
nor U882 (N_882,N_153,N_14);
and U883 (N_883,N_244,N_282);
and U884 (N_884,N_252,N_194);
or U885 (N_885,N_305,N_327);
and U886 (N_886,N_455,N_269);
nor U887 (N_887,N_85,N_476);
or U888 (N_888,N_82,N_40);
or U889 (N_889,N_389,N_227);
nor U890 (N_890,N_242,N_95);
or U891 (N_891,N_305,N_452);
and U892 (N_892,N_131,N_329);
nand U893 (N_893,N_401,N_359);
and U894 (N_894,N_413,N_248);
or U895 (N_895,N_56,N_334);
nand U896 (N_896,N_5,N_18);
nand U897 (N_897,N_445,N_103);
or U898 (N_898,N_210,N_216);
nor U899 (N_899,N_55,N_273);
nor U900 (N_900,N_371,N_221);
and U901 (N_901,N_303,N_253);
or U902 (N_902,N_468,N_72);
and U903 (N_903,N_162,N_442);
and U904 (N_904,N_397,N_351);
nand U905 (N_905,N_342,N_222);
or U906 (N_906,N_127,N_276);
nand U907 (N_907,N_284,N_443);
and U908 (N_908,N_463,N_91);
nor U909 (N_909,N_110,N_235);
or U910 (N_910,N_41,N_162);
and U911 (N_911,N_477,N_182);
nor U912 (N_912,N_78,N_220);
nor U913 (N_913,N_116,N_356);
and U914 (N_914,N_458,N_435);
nor U915 (N_915,N_201,N_441);
nand U916 (N_916,N_219,N_301);
or U917 (N_917,N_131,N_330);
nor U918 (N_918,N_135,N_163);
and U919 (N_919,N_87,N_463);
and U920 (N_920,N_278,N_449);
and U921 (N_921,N_346,N_60);
and U922 (N_922,N_249,N_296);
nor U923 (N_923,N_291,N_50);
or U924 (N_924,N_273,N_151);
nand U925 (N_925,N_404,N_280);
nor U926 (N_926,N_78,N_229);
and U927 (N_927,N_228,N_260);
nor U928 (N_928,N_31,N_326);
nand U929 (N_929,N_167,N_428);
or U930 (N_930,N_153,N_457);
nand U931 (N_931,N_191,N_454);
or U932 (N_932,N_212,N_276);
and U933 (N_933,N_483,N_64);
and U934 (N_934,N_242,N_24);
nor U935 (N_935,N_14,N_497);
or U936 (N_936,N_209,N_156);
and U937 (N_937,N_424,N_292);
or U938 (N_938,N_341,N_55);
nand U939 (N_939,N_342,N_30);
and U940 (N_940,N_28,N_498);
or U941 (N_941,N_3,N_119);
or U942 (N_942,N_174,N_375);
xnor U943 (N_943,N_455,N_141);
nand U944 (N_944,N_318,N_60);
or U945 (N_945,N_59,N_157);
xnor U946 (N_946,N_47,N_307);
and U947 (N_947,N_423,N_213);
and U948 (N_948,N_208,N_339);
nand U949 (N_949,N_133,N_106);
nand U950 (N_950,N_61,N_45);
and U951 (N_951,N_199,N_399);
or U952 (N_952,N_17,N_316);
nand U953 (N_953,N_157,N_497);
nor U954 (N_954,N_333,N_108);
nand U955 (N_955,N_497,N_443);
nand U956 (N_956,N_334,N_256);
nor U957 (N_957,N_441,N_310);
nor U958 (N_958,N_107,N_417);
and U959 (N_959,N_352,N_307);
or U960 (N_960,N_495,N_49);
nand U961 (N_961,N_280,N_347);
nand U962 (N_962,N_335,N_76);
and U963 (N_963,N_50,N_460);
nand U964 (N_964,N_298,N_283);
and U965 (N_965,N_327,N_250);
nor U966 (N_966,N_289,N_229);
or U967 (N_967,N_468,N_355);
and U968 (N_968,N_61,N_329);
or U969 (N_969,N_83,N_379);
nor U970 (N_970,N_67,N_390);
or U971 (N_971,N_88,N_170);
nor U972 (N_972,N_222,N_79);
and U973 (N_973,N_199,N_206);
or U974 (N_974,N_123,N_434);
nor U975 (N_975,N_178,N_484);
nand U976 (N_976,N_177,N_208);
nand U977 (N_977,N_327,N_259);
and U978 (N_978,N_140,N_237);
xnor U979 (N_979,N_240,N_97);
and U980 (N_980,N_258,N_386);
or U981 (N_981,N_418,N_314);
nand U982 (N_982,N_129,N_383);
and U983 (N_983,N_94,N_69);
nand U984 (N_984,N_37,N_296);
and U985 (N_985,N_229,N_179);
or U986 (N_986,N_454,N_464);
nor U987 (N_987,N_263,N_389);
or U988 (N_988,N_118,N_87);
nand U989 (N_989,N_123,N_184);
nand U990 (N_990,N_373,N_334);
and U991 (N_991,N_85,N_10);
nand U992 (N_992,N_357,N_340);
nor U993 (N_993,N_324,N_26);
nand U994 (N_994,N_87,N_206);
or U995 (N_995,N_176,N_238);
nor U996 (N_996,N_322,N_113);
nor U997 (N_997,N_36,N_84);
nor U998 (N_998,N_327,N_202);
or U999 (N_999,N_211,N_131);
nor U1000 (N_1000,N_564,N_739);
and U1001 (N_1001,N_525,N_507);
and U1002 (N_1002,N_946,N_968);
or U1003 (N_1003,N_956,N_963);
and U1004 (N_1004,N_897,N_930);
or U1005 (N_1005,N_642,N_686);
nor U1006 (N_1006,N_588,N_785);
nand U1007 (N_1007,N_694,N_817);
and U1008 (N_1008,N_703,N_548);
nand U1009 (N_1009,N_974,N_699);
nor U1010 (N_1010,N_800,N_528);
nor U1011 (N_1011,N_945,N_854);
nor U1012 (N_1012,N_631,N_611);
nand U1013 (N_1013,N_531,N_584);
and U1014 (N_1014,N_766,N_894);
nand U1015 (N_1015,N_558,N_644);
nand U1016 (N_1016,N_562,N_934);
and U1017 (N_1017,N_598,N_695);
and U1018 (N_1018,N_753,N_794);
and U1019 (N_1019,N_761,N_841);
and U1020 (N_1020,N_704,N_986);
nand U1021 (N_1021,N_574,N_778);
nor U1022 (N_1022,N_876,N_690);
or U1023 (N_1023,N_955,N_745);
nor U1024 (N_1024,N_554,N_937);
nor U1025 (N_1025,N_655,N_594);
and U1026 (N_1026,N_881,N_685);
nand U1027 (N_1027,N_616,N_688);
nand U1028 (N_1028,N_799,N_786);
or U1029 (N_1029,N_816,N_541);
nor U1030 (N_1030,N_676,N_991);
and U1031 (N_1031,N_681,N_669);
and U1032 (N_1032,N_994,N_770);
nor U1033 (N_1033,N_902,N_600);
nor U1034 (N_1034,N_896,N_579);
nand U1035 (N_1035,N_793,N_901);
nand U1036 (N_1036,N_749,N_863);
nand U1037 (N_1037,N_743,N_877);
and U1038 (N_1038,N_936,N_552);
and U1039 (N_1039,N_540,N_519);
nor U1040 (N_1040,N_625,N_737);
nor U1041 (N_1041,N_859,N_965);
nand U1042 (N_1042,N_849,N_708);
nand U1043 (N_1043,N_995,N_972);
or U1044 (N_1044,N_866,N_914);
or U1045 (N_1045,N_890,N_728);
and U1046 (N_1046,N_730,N_673);
and U1047 (N_1047,N_647,N_510);
nor U1048 (N_1048,N_501,N_821);
or U1049 (N_1049,N_858,N_813);
nor U1050 (N_1050,N_707,N_668);
or U1051 (N_1051,N_561,N_944);
nor U1052 (N_1052,N_735,N_885);
or U1053 (N_1053,N_533,N_651);
or U1054 (N_1054,N_763,N_582);
and U1055 (N_1055,N_522,N_978);
or U1056 (N_1056,N_768,N_626);
and U1057 (N_1057,N_727,N_933);
nand U1058 (N_1058,N_526,N_609);
or U1059 (N_1059,N_776,N_575);
nand U1060 (N_1060,N_537,N_736);
and U1061 (N_1061,N_912,N_523);
nor U1062 (N_1062,N_790,N_569);
or U1063 (N_1063,N_840,N_857);
or U1064 (N_1064,N_604,N_970);
and U1065 (N_1065,N_880,N_976);
or U1066 (N_1066,N_649,N_867);
nand U1067 (N_1067,N_764,N_532);
or U1068 (N_1068,N_572,N_715);
nand U1069 (N_1069,N_678,N_920);
and U1070 (N_1070,N_536,N_516);
nor U1071 (N_1071,N_985,N_560);
and U1072 (N_1072,N_789,N_629);
or U1073 (N_1073,N_882,N_843);
or U1074 (N_1074,N_787,N_940);
nand U1075 (N_1075,N_658,N_862);
or U1076 (N_1076,N_634,N_839);
and U1077 (N_1077,N_636,N_871);
and U1078 (N_1078,N_621,N_975);
or U1079 (N_1079,N_734,N_996);
and U1080 (N_1080,N_928,N_701);
or U1081 (N_1081,N_723,N_827);
and U1082 (N_1082,N_815,N_774);
or U1083 (N_1083,N_557,N_587);
and U1084 (N_1084,N_846,N_689);
nand U1085 (N_1085,N_622,N_812);
or U1086 (N_1086,N_771,N_993);
and U1087 (N_1087,N_853,N_795);
nor U1088 (N_1088,N_726,N_779);
and U1089 (N_1089,N_830,N_889);
nor U1090 (N_1090,N_508,N_610);
or U1091 (N_1091,N_578,N_665);
and U1092 (N_1092,N_635,N_529);
nor U1093 (N_1093,N_987,N_534);
nor U1094 (N_1094,N_545,N_868);
or U1095 (N_1095,N_500,N_645);
nand U1096 (N_1096,N_856,N_580);
nor U1097 (N_1097,N_744,N_538);
and U1098 (N_1098,N_513,N_576);
and U1099 (N_1099,N_746,N_973);
and U1100 (N_1100,N_801,N_627);
nor U1101 (N_1101,N_939,N_718);
and U1102 (N_1102,N_721,N_884);
and U1103 (N_1103,N_667,N_542);
nor U1104 (N_1104,N_742,N_664);
nor U1105 (N_1105,N_630,N_589);
or U1106 (N_1106,N_691,N_546);
or U1107 (N_1107,N_819,N_765);
nand U1108 (N_1108,N_504,N_696);
or U1109 (N_1109,N_679,N_767);
nor U1110 (N_1110,N_581,N_731);
nand U1111 (N_1111,N_879,N_961);
nand U1112 (N_1112,N_949,N_924);
nor U1113 (N_1113,N_848,N_603);
or U1114 (N_1114,N_942,N_663);
nor U1115 (N_1115,N_977,N_543);
or U1116 (N_1116,N_938,N_873);
nand U1117 (N_1117,N_711,N_989);
nor U1118 (N_1118,N_814,N_806);
nand U1119 (N_1119,N_754,N_878);
or U1120 (N_1120,N_820,N_583);
and U1121 (N_1121,N_913,N_652);
nand U1122 (N_1122,N_818,N_633);
or U1123 (N_1123,N_666,N_967);
and U1124 (N_1124,N_998,N_653);
and U1125 (N_1125,N_577,N_568);
nand U1126 (N_1126,N_670,N_953);
and U1127 (N_1127,N_599,N_788);
or U1128 (N_1128,N_810,N_671);
nor U1129 (N_1129,N_521,N_792);
or U1130 (N_1130,N_809,N_729);
xnor U1131 (N_1131,N_672,N_505);
nor U1132 (N_1132,N_960,N_803);
and U1133 (N_1133,N_834,N_674);
or U1134 (N_1134,N_722,N_719);
or U1135 (N_1135,N_926,N_916);
or U1136 (N_1136,N_586,N_962);
nand U1137 (N_1137,N_907,N_826);
or U1138 (N_1138,N_808,N_844);
nor U1139 (N_1139,N_905,N_733);
nand U1140 (N_1140,N_931,N_682);
and U1141 (N_1141,N_798,N_898);
nor U1142 (N_1142,N_511,N_999);
and U1143 (N_1143,N_888,N_551);
or U1144 (N_1144,N_796,N_782);
nand U1145 (N_1145,N_908,N_656);
nor U1146 (N_1146,N_822,N_570);
and U1147 (N_1147,N_615,N_646);
or U1148 (N_1148,N_693,N_851);
nand U1149 (N_1149,N_850,N_716);
nor U1150 (N_1150,N_904,N_966);
nor U1151 (N_1151,N_592,N_791);
nand U1152 (N_1152,N_982,N_654);
nor U1153 (N_1153,N_947,N_911);
or U1154 (N_1154,N_825,N_984);
or U1155 (N_1155,N_662,N_772);
and U1156 (N_1156,N_958,N_864);
nor U1157 (N_1157,N_832,N_530);
or U1158 (N_1158,N_648,N_698);
nor U1159 (N_1159,N_833,N_502);
nand U1160 (N_1160,N_874,N_969);
nand U1161 (N_1161,N_520,N_650);
or U1162 (N_1162,N_917,N_556);
nand U1163 (N_1163,N_837,N_855);
or U1164 (N_1164,N_811,N_614);
nor U1165 (N_1165,N_619,N_971);
nand U1166 (N_1166,N_952,N_712);
and U1167 (N_1167,N_524,N_758);
nand U1168 (N_1168,N_724,N_935);
nor U1169 (N_1169,N_738,N_983);
and U1170 (N_1170,N_829,N_892);
and U1171 (N_1171,N_802,N_607);
nand U1172 (N_1172,N_943,N_845);
or U1173 (N_1173,N_680,N_677);
nor U1174 (N_1174,N_515,N_852);
and U1175 (N_1175,N_612,N_957);
and U1176 (N_1176,N_988,N_608);
nor U1177 (N_1177,N_567,N_748);
and U1178 (N_1178,N_573,N_591);
or U1179 (N_1179,N_784,N_509);
nand U1180 (N_1180,N_835,N_517);
nor U1181 (N_1181,N_838,N_613);
and U1182 (N_1182,N_828,N_700);
nor U1183 (N_1183,N_948,N_807);
or U1184 (N_1184,N_997,N_883);
and U1185 (N_1185,N_891,N_929);
or U1186 (N_1186,N_563,N_797);
nor U1187 (N_1187,N_714,N_675);
or U1188 (N_1188,N_842,N_954);
nor U1189 (N_1189,N_660,N_623);
and U1190 (N_1190,N_659,N_941);
nand U1191 (N_1191,N_910,N_593);
nor U1192 (N_1192,N_628,N_595);
and U1193 (N_1193,N_893,N_951);
and U1194 (N_1194,N_661,N_773);
nor U1195 (N_1195,N_585,N_950);
nor U1196 (N_1196,N_717,N_602);
and U1197 (N_1197,N_550,N_597);
and U1198 (N_1198,N_702,N_705);
nand U1199 (N_1199,N_847,N_692);
and U1200 (N_1200,N_747,N_709);
and U1201 (N_1201,N_909,N_861);
and U1202 (N_1202,N_566,N_555);
nor U1203 (N_1203,N_918,N_506);
or U1204 (N_1204,N_710,N_870);
nand U1205 (N_1205,N_922,N_990);
nor U1206 (N_1206,N_601,N_915);
and U1207 (N_1207,N_887,N_606);
nand U1208 (N_1208,N_759,N_544);
nor U1209 (N_1209,N_756,N_777);
or U1210 (N_1210,N_921,N_637);
and U1211 (N_1211,N_618,N_643);
and U1212 (N_1212,N_869,N_539);
nand U1213 (N_1213,N_617,N_518);
or U1214 (N_1214,N_751,N_605);
nor U1215 (N_1215,N_639,N_804);
nand U1216 (N_1216,N_684,N_527);
and U1217 (N_1217,N_780,N_981);
nand U1218 (N_1218,N_725,N_836);
or U1219 (N_1219,N_865,N_872);
nand U1220 (N_1220,N_927,N_762);
and U1221 (N_1221,N_752,N_620);
nor U1222 (N_1222,N_740,N_683);
nand U1223 (N_1223,N_755,N_657);
nor U1224 (N_1224,N_706,N_980);
and U1225 (N_1225,N_632,N_805);
or U1226 (N_1226,N_959,N_624);
nor U1227 (N_1227,N_823,N_553);
and U1228 (N_1228,N_596,N_783);
nand U1229 (N_1229,N_923,N_906);
nand U1230 (N_1230,N_741,N_775);
nand U1231 (N_1231,N_590,N_875);
or U1232 (N_1232,N_886,N_769);
and U1233 (N_1233,N_559,N_899);
nor U1234 (N_1234,N_697,N_760);
nand U1235 (N_1235,N_992,N_979);
or U1236 (N_1236,N_903,N_514);
and U1237 (N_1237,N_565,N_687);
nor U1238 (N_1238,N_964,N_831);
nor U1239 (N_1239,N_781,N_919);
and U1240 (N_1240,N_571,N_932);
or U1241 (N_1241,N_503,N_732);
and U1242 (N_1242,N_860,N_549);
and U1243 (N_1243,N_720,N_900);
xnor U1244 (N_1244,N_512,N_535);
or U1245 (N_1245,N_750,N_641);
nor U1246 (N_1246,N_895,N_638);
and U1247 (N_1247,N_547,N_640);
nor U1248 (N_1248,N_713,N_757);
nor U1249 (N_1249,N_824,N_925);
or U1250 (N_1250,N_951,N_914);
nand U1251 (N_1251,N_637,N_641);
or U1252 (N_1252,N_518,N_520);
nand U1253 (N_1253,N_810,N_984);
or U1254 (N_1254,N_751,N_565);
nand U1255 (N_1255,N_764,N_595);
nor U1256 (N_1256,N_712,N_927);
or U1257 (N_1257,N_757,N_636);
nand U1258 (N_1258,N_531,N_966);
nand U1259 (N_1259,N_653,N_660);
or U1260 (N_1260,N_522,N_642);
nor U1261 (N_1261,N_965,N_864);
or U1262 (N_1262,N_870,N_689);
nor U1263 (N_1263,N_971,N_569);
or U1264 (N_1264,N_985,N_944);
nor U1265 (N_1265,N_923,N_879);
or U1266 (N_1266,N_742,N_905);
nor U1267 (N_1267,N_507,N_688);
nand U1268 (N_1268,N_536,N_634);
nor U1269 (N_1269,N_768,N_558);
nor U1270 (N_1270,N_749,N_880);
nor U1271 (N_1271,N_799,N_974);
and U1272 (N_1272,N_757,N_542);
nor U1273 (N_1273,N_951,N_675);
nand U1274 (N_1274,N_568,N_559);
and U1275 (N_1275,N_633,N_692);
and U1276 (N_1276,N_732,N_816);
or U1277 (N_1277,N_895,N_657);
and U1278 (N_1278,N_629,N_966);
and U1279 (N_1279,N_864,N_555);
nor U1280 (N_1280,N_926,N_750);
or U1281 (N_1281,N_726,N_811);
nor U1282 (N_1282,N_831,N_647);
nand U1283 (N_1283,N_734,N_982);
nand U1284 (N_1284,N_914,N_625);
xnor U1285 (N_1285,N_866,N_740);
nand U1286 (N_1286,N_724,N_603);
or U1287 (N_1287,N_528,N_526);
or U1288 (N_1288,N_840,N_535);
or U1289 (N_1289,N_722,N_942);
and U1290 (N_1290,N_602,N_973);
or U1291 (N_1291,N_507,N_984);
or U1292 (N_1292,N_764,N_893);
nor U1293 (N_1293,N_529,N_643);
and U1294 (N_1294,N_584,N_533);
nand U1295 (N_1295,N_642,N_785);
nor U1296 (N_1296,N_903,N_727);
nor U1297 (N_1297,N_787,N_605);
and U1298 (N_1298,N_524,N_602);
nor U1299 (N_1299,N_919,N_531);
and U1300 (N_1300,N_780,N_681);
and U1301 (N_1301,N_999,N_690);
and U1302 (N_1302,N_745,N_792);
or U1303 (N_1303,N_560,N_641);
or U1304 (N_1304,N_670,N_697);
nor U1305 (N_1305,N_696,N_555);
nand U1306 (N_1306,N_885,N_584);
or U1307 (N_1307,N_547,N_626);
nand U1308 (N_1308,N_921,N_762);
and U1309 (N_1309,N_985,N_759);
nor U1310 (N_1310,N_893,N_856);
or U1311 (N_1311,N_585,N_703);
nor U1312 (N_1312,N_671,N_946);
or U1313 (N_1313,N_715,N_874);
nand U1314 (N_1314,N_798,N_705);
nor U1315 (N_1315,N_660,N_787);
or U1316 (N_1316,N_805,N_651);
nand U1317 (N_1317,N_563,N_729);
or U1318 (N_1318,N_544,N_806);
or U1319 (N_1319,N_782,N_870);
nand U1320 (N_1320,N_660,N_845);
nor U1321 (N_1321,N_856,N_763);
and U1322 (N_1322,N_659,N_814);
and U1323 (N_1323,N_878,N_857);
and U1324 (N_1324,N_867,N_927);
nand U1325 (N_1325,N_663,N_521);
and U1326 (N_1326,N_574,N_568);
or U1327 (N_1327,N_851,N_922);
nand U1328 (N_1328,N_712,N_766);
or U1329 (N_1329,N_780,N_701);
nand U1330 (N_1330,N_700,N_892);
and U1331 (N_1331,N_698,N_927);
or U1332 (N_1332,N_673,N_539);
nand U1333 (N_1333,N_518,N_849);
nand U1334 (N_1334,N_874,N_981);
nand U1335 (N_1335,N_978,N_776);
or U1336 (N_1336,N_826,N_853);
or U1337 (N_1337,N_575,N_712);
nand U1338 (N_1338,N_649,N_964);
and U1339 (N_1339,N_930,N_980);
and U1340 (N_1340,N_695,N_897);
nor U1341 (N_1341,N_745,N_922);
and U1342 (N_1342,N_983,N_726);
nand U1343 (N_1343,N_945,N_676);
or U1344 (N_1344,N_931,N_517);
xnor U1345 (N_1345,N_960,N_567);
nor U1346 (N_1346,N_759,N_785);
nand U1347 (N_1347,N_878,N_938);
nand U1348 (N_1348,N_825,N_965);
or U1349 (N_1349,N_724,N_912);
or U1350 (N_1350,N_687,N_992);
and U1351 (N_1351,N_814,N_585);
nand U1352 (N_1352,N_503,N_658);
nand U1353 (N_1353,N_874,N_506);
nand U1354 (N_1354,N_812,N_814);
nor U1355 (N_1355,N_888,N_751);
nor U1356 (N_1356,N_706,N_749);
or U1357 (N_1357,N_969,N_721);
nor U1358 (N_1358,N_520,N_952);
and U1359 (N_1359,N_716,N_860);
nand U1360 (N_1360,N_630,N_893);
and U1361 (N_1361,N_615,N_881);
and U1362 (N_1362,N_730,N_529);
or U1363 (N_1363,N_881,N_876);
and U1364 (N_1364,N_669,N_667);
nor U1365 (N_1365,N_806,N_789);
or U1366 (N_1366,N_613,N_500);
and U1367 (N_1367,N_821,N_705);
nand U1368 (N_1368,N_577,N_666);
nand U1369 (N_1369,N_976,N_763);
nand U1370 (N_1370,N_961,N_842);
nor U1371 (N_1371,N_970,N_927);
nor U1372 (N_1372,N_677,N_815);
or U1373 (N_1373,N_587,N_530);
or U1374 (N_1374,N_731,N_545);
and U1375 (N_1375,N_521,N_720);
nand U1376 (N_1376,N_675,N_660);
nand U1377 (N_1377,N_815,N_941);
and U1378 (N_1378,N_621,N_578);
and U1379 (N_1379,N_607,N_801);
or U1380 (N_1380,N_636,N_690);
nand U1381 (N_1381,N_721,N_795);
or U1382 (N_1382,N_752,N_532);
nor U1383 (N_1383,N_530,N_711);
nor U1384 (N_1384,N_850,N_899);
nand U1385 (N_1385,N_673,N_982);
nor U1386 (N_1386,N_701,N_531);
nand U1387 (N_1387,N_869,N_606);
nand U1388 (N_1388,N_692,N_989);
nand U1389 (N_1389,N_501,N_773);
and U1390 (N_1390,N_605,N_931);
or U1391 (N_1391,N_584,N_834);
and U1392 (N_1392,N_889,N_948);
or U1393 (N_1393,N_890,N_836);
or U1394 (N_1394,N_892,N_510);
or U1395 (N_1395,N_808,N_797);
or U1396 (N_1396,N_671,N_956);
and U1397 (N_1397,N_653,N_617);
xnor U1398 (N_1398,N_751,N_718);
nor U1399 (N_1399,N_519,N_760);
nor U1400 (N_1400,N_837,N_608);
nand U1401 (N_1401,N_598,N_641);
nand U1402 (N_1402,N_941,N_764);
nand U1403 (N_1403,N_744,N_903);
nand U1404 (N_1404,N_661,N_987);
and U1405 (N_1405,N_652,N_621);
nand U1406 (N_1406,N_624,N_974);
nand U1407 (N_1407,N_761,N_971);
or U1408 (N_1408,N_724,N_949);
nand U1409 (N_1409,N_901,N_874);
nor U1410 (N_1410,N_693,N_724);
nor U1411 (N_1411,N_689,N_852);
nor U1412 (N_1412,N_972,N_593);
and U1413 (N_1413,N_599,N_781);
xor U1414 (N_1414,N_652,N_849);
nand U1415 (N_1415,N_986,N_822);
or U1416 (N_1416,N_969,N_981);
nand U1417 (N_1417,N_797,N_513);
and U1418 (N_1418,N_834,N_835);
or U1419 (N_1419,N_702,N_680);
or U1420 (N_1420,N_592,N_715);
and U1421 (N_1421,N_500,N_840);
nor U1422 (N_1422,N_993,N_766);
nand U1423 (N_1423,N_551,N_654);
or U1424 (N_1424,N_770,N_673);
or U1425 (N_1425,N_633,N_842);
or U1426 (N_1426,N_595,N_686);
nor U1427 (N_1427,N_664,N_914);
nand U1428 (N_1428,N_574,N_892);
nor U1429 (N_1429,N_881,N_671);
and U1430 (N_1430,N_548,N_754);
and U1431 (N_1431,N_837,N_800);
xor U1432 (N_1432,N_753,N_538);
nor U1433 (N_1433,N_753,N_638);
and U1434 (N_1434,N_833,N_972);
and U1435 (N_1435,N_674,N_802);
xor U1436 (N_1436,N_928,N_716);
and U1437 (N_1437,N_608,N_797);
nor U1438 (N_1438,N_574,N_572);
and U1439 (N_1439,N_732,N_578);
nor U1440 (N_1440,N_864,N_962);
nor U1441 (N_1441,N_644,N_574);
nor U1442 (N_1442,N_999,N_651);
nor U1443 (N_1443,N_681,N_989);
and U1444 (N_1444,N_691,N_952);
or U1445 (N_1445,N_804,N_572);
and U1446 (N_1446,N_555,N_528);
xnor U1447 (N_1447,N_951,N_854);
and U1448 (N_1448,N_950,N_602);
or U1449 (N_1449,N_576,N_528);
or U1450 (N_1450,N_579,N_613);
or U1451 (N_1451,N_981,N_675);
nor U1452 (N_1452,N_661,N_702);
or U1453 (N_1453,N_705,N_611);
nor U1454 (N_1454,N_973,N_982);
or U1455 (N_1455,N_783,N_665);
and U1456 (N_1456,N_827,N_877);
nor U1457 (N_1457,N_842,N_505);
or U1458 (N_1458,N_736,N_675);
and U1459 (N_1459,N_957,N_959);
nand U1460 (N_1460,N_960,N_847);
and U1461 (N_1461,N_520,N_547);
nand U1462 (N_1462,N_618,N_994);
and U1463 (N_1463,N_741,N_586);
nor U1464 (N_1464,N_835,N_750);
or U1465 (N_1465,N_522,N_872);
nor U1466 (N_1466,N_932,N_631);
nor U1467 (N_1467,N_579,N_602);
and U1468 (N_1468,N_956,N_860);
nand U1469 (N_1469,N_686,N_908);
nand U1470 (N_1470,N_937,N_974);
and U1471 (N_1471,N_971,N_638);
nor U1472 (N_1472,N_951,N_516);
nor U1473 (N_1473,N_921,N_880);
or U1474 (N_1474,N_627,N_945);
nand U1475 (N_1475,N_575,N_535);
nor U1476 (N_1476,N_761,N_910);
or U1477 (N_1477,N_531,N_963);
or U1478 (N_1478,N_779,N_822);
nor U1479 (N_1479,N_699,N_842);
and U1480 (N_1480,N_509,N_741);
nor U1481 (N_1481,N_573,N_598);
and U1482 (N_1482,N_725,N_570);
nor U1483 (N_1483,N_568,N_884);
nor U1484 (N_1484,N_969,N_791);
nand U1485 (N_1485,N_684,N_727);
or U1486 (N_1486,N_980,N_912);
nor U1487 (N_1487,N_564,N_507);
or U1488 (N_1488,N_619,N_988);
nor U1489 (N_1489,N_609,N_901);
or U1490 (N_1490,N_711,N_699);
nor U1491 (N_1491,N_664,N_735);
or U1492 (N_1492,N_539,N_681);
or U1493 (N_1493,N_900,N_822);
and U1494 (N_1494,N_501,N_681);
nor U1495 (N_1495,N_702,N_791);
nand U1496 (N_1496,N_961,N_691);
nor U1497 (N_1497,N_821,N_552);
and U1498 (N_1498,N_673,N_607);
and U1499 (N_1499,N_610,N_694);
and U1500 (N_1500,N_1045,N_1134);
and U1501 (N_1501,N_1067,N_1430);
nor U1502 (N_1502,N_1065,N_1253);
nor U1503 (N_1503,N_1431,N_1017);
or U1504 (N_1504,N_1244,N_1285);
or U1505 (N_1505,N_1393,N_1129);
nor U1506 (N_1506,N_1101,N_1457);
and U1507 (N_1507,N_1131,N_1441);
nor U1508 (N_1508,N_1432,N_1102);
and U1509 (N_1509,N_1236,N_1080);
and U1510 (N_1510,N_1235,N_1185);
nand U1511 (N_1511,N_1190,N_1212);
nand U1512 (N_1512,N_1445,N_1480);
nor U1513 (N_1513,N_1455,N_1448);
or U1514 (N_1514,N_1085,N_1366);
nand U1515 (N_1515,N_1155,N_1382);
or U1516 (N_1516,N_1268,N_1088);
and U1517 (N_1517,N_1002,N_1196);
and U1518 (N_1518,N_1453,N_1215);
nand U1519 (N_1519,N_1343,N_1136);
or U1520 (N_1520,N_1380,N_1043);
and U1521 (N_1521,N_1114,N_1429);
or U1522 (N_1522,N_1158,N_1025);
and U1523 (N_1523,N_1014,N_1274);
and U1524 (N_1524,N_1009,N_1118);
and U1525 (N_1525,N_1006,N_1409);
and U1526 (N_1526,N_1095,N_1223);
or U1527 (N_1527,N_1449,N_1394);
nand U1528 (N_1528,N_1228,N_1444);
nor U1529 (N_1529,N_1027,N_1159);
nand U1530 (N_1530,N_1010,N_1066);
nor U1531 (N_1531,N_1309,N_1093);
nand U1532 (N_1532,N_1142,N_1301);
and U1533 (N_1533,N_1036,N_1075);
and U1534 (N_1534,N_1367,N_1479);
and U1535 (N_1535,N_1054,N_1051);
nand U1536 (N_1536,N_1202,N_1355);
and U1537 (N_1537,N_1466,N_1205);
nand U1538 (N_1538,N_1099,N_1057);
nor U1539 (N_1539,N_1345,N_1385);
and U1540 (N_1540,N_1378,N_1069);
or U1541 (N_1541,N_1061,N_1071);
nand U1542 (N_1542,N_1214,N_1074);
xnor U1543 (N_1543,N_1091,N_1259);
nor U1544 (N_1544,N_1348,N_1217);
nand U1545 (N_1545,N_1277,N_1260);
or U1546 (N_1546,N_1022,N_1225);
and U1547 (N_1547,N_1387,N_1470);
nor U1548 (N_1548,N_1276,N_1181);
or U1549 (N_1549,N_1497,N_1331);
nor U1550 (N_1550,N_1172,N_1433);
nand U1551 (N_1551,N_1216,N_1314);
nand U1552 (N_1552,N_1306,N_1398);
and U1553 (N_1553,N_1100,N_1210);
nor U1554 (N_1554,N_1330,N_1384);
or U1555 (N_1555,N_1334,N_1462);
or U1556 (N_1556,N_1186,N_1126);
nand U1557 (N_1557,N_1255,N_1180);
nand U1558 (N_1558,N_1411,N_1233);
nand U1559 (N_1559,N_1220,N_1239);
and U1560 (N_1560,N_1089,N_1325);
nor U1561 (N_1561,N_1272,N_1287);
or U1562 (N_1562,N_1403,N_1408);
and U1563 (N_1563,N_1068,N_1351);
or U1564 (N_1564,N_1019,N_1293);
and U1565 (N_1565,N_1153,N_1034);
and U1566 (N_1566,N_1229,N_1486);
nand U1567 (N_1567,N_1324,N_1204);
and U1568 (N_1568,N_1464,N_1015);
nand U1569 (N_1569,N_1033,N_1224);
nand U1570 (N_1570,N_1168,N_1283);
nand U1571 (N_1571,N_1278,N_1371);
nand U1572 (N_1572,N_1249,N_1284);
or U1573 (N_1573,N_1289,N_1127);
and U1574 (N_1574,N_1468,N_1439);
or U1575 (N_1575,N_1044,N_1389);
or U1576 (N_1576,N_1148,N_1428);
nor U1577 (N_1577,N_1157,N_1340);
and U1578 (N_1578,N_1230,N_1182);
and U1579 (N_1579,N_1177,N_1245);
nand U1580 (N_1580,N_1046,N_1011);
and U1581 (N_1581,N_1417,N_1405);
nand U1582 (N_1582,N_1476,N_1161);
or U1583 (N_1583,N_1474,N_1262);
or U1584 (N_1584,N_1116,N_1307);
nor U1585 (N_1585,N_1218,N_1333);
nand U1586 (N_1586,N_1248,N_1492);
nor U1587 (N_1587,N_1195,N_1193);
and U1588 (N_1588,N_1243,N_1156);
or U1589 (N_1589,N_1146,N_1339);
nor U1590 (N_1590,N_1421,N_1087);
or U1591 (N_1591,N_1499,N_1108);
nand U1592 (N_1592,N_1013,N_1247);
nor U1593 (N_1593,N_1179,N_1377);
or U1594 (N_1594,N_1008,N_1083);
and U1595 (N_1595,N_1113,N_1053);
nor U1596 (N_1596,N_1124,N_1270);
or U1597 (N_1597,N_1496,N_1016);
or U1598 (N_1598,N_1313,N_1420);
and U1599 (N_1599,N_1232,N_1381);
nor U1600 (N_1600,N_1438,N_1332);
or U1601 (N_1601,N_1375,N_1026);
or U1602 (N_1602,N_1240,N_1483);
or U1603 (N_1603,N_1425,N_1359);
nor U1604 (N_1604,N_1299,N_1471);
nand U1605 (N_1605,N_1227,N_1110);
and U1606 (N_1606,N_1165,N_1327);
nand U1607 (N_1607,N_1077,N_1163);
nand U1608 (N_1608,N_1261,N_1335);
nand U1609 (N_1609,N_1374,N_1213);
or U1610 (N_1610,N_1388,N_1115);
nand U1611 (N_1611,N_1047,N_1317);
or U1612 (N_1612,N_1279,N_1312);
and U1613 (N_1613,N_1282,N_1450);
nand U1614 (N_1614,N_1275,N_1092);
or U1615 (N_1615,N_1437,N_1297);
nor U1616 (N_1616,N_1201,N_1139);
nand U1617 (N_1617,N_1020,N_1004);
nor U1618 (N_1618,N_1104,N_1487);
nor U1619 (N_1619,N_1086,N_1198);
or U1620 (N_1620,N_1484,N_1251);
and U1621 (N_1621,N_1003,N_1234);
or U1622 (N_1622,N_1176,N_1356);
nor U1623 (N_1623,N_1197,N_1132);
nor U1624 (N_1624,N_1137,N_1117);
nand U1625 (N_1625,N_1064,N_1296);
or U1626 (N_1626,N_1273,N_1167);
nand U1627 (N_1627,N_1434,N_1338);
nand U1628 (N_1628,N_1370,N_1029);
nor U1629 (N_1629,N_1191,N_1467);
nor U1630 (N_1630,N_1458,N_1291);
nand U1631 (N_1631,N_1125,N_1424);
nor U1632 (N_1632,N_1265,N_1000);
or U1633 (N_1633,N_1368,N_1138);
and U1634 (N_1634,N_1012,N_1469);
or U1635 (N_1635,N_1485,N_1264);
nor U1636 (N_1636,N_1373,N_1226);
or U1637 (N_1637,N_1475,N_1414);
nor U1638 (N_1638,N_1362,N_1030);
or U1639 (N_1639,N_1070,N_1342);
nor U1640 (N_1640,N_1473,N_1059);
or U1641 (N_1641,N_1040,N_1256);
nor U1642 (N_1642,N_1222,N_1081);
nor U1643 (N_1643,N_1105,N_1446);
nor U1644 (N_1644,N_1308,N_1250);
and U1645 (N_1645,N_1426,N_1038);
or U1646 (N_1646,N_1147,N_1018);
or U1647 (N_1647,N_1488,N_1358);
or U1648 (N_1648,N_1401,N_1060);
nand U1649 (N_1649,N_1383,N_1252);
nand U1650 (N_1650,N_1454,N_1001);
nand U1651 (N_1651,N_1058,N_1231);
and U1652 (N_1652,N_1072,N_1035);
and U1653 (N_1653,N_1318,N_1328);
nand U1654 (N_1654,N_1322,N_1295);
nor U1655 (N_1655,N_1143,N_1007);
or U1656 (N_1656,N_1112,N_1052);
nand U1657 (N_1657,N_1173,N_1491);
nor U1658 (N_1658,N_1106,N_1365);
or U1659 (N_1659,N_1315,N_1149);
nor U1660 (N_1660,N_1406,N_1412);
and U1661 (N_1661,N_1094,N_1402);
nand U1662 (N_1662,N_1397,N_1290);
and U1663 (N_1663,N_1478,N_1311);
or U1664 (N_1664,N_1152,N_1489);
xor U1665 (N_1665,N_1140,N_1258);
and U1666 (N_1666,N_1498,N_1336);
or U1667 (N_1667,N_1456,N_1145);
nor U1668 (N_1668,N_1109,N_1344);
or U1669 (N_1669,N_1031,N_1178);
or U1670 (N_1670,N_1292,N_1271);
or U1671 (N_1671,N_1465,N_1305);
nand U1672 (N_1672,N_1329,N_1376);
or U1673 (N_1673,N_1407,N_1347);
nor U1674 (N_1674,N_1481,N_1495);
nand U1675 (N_1675,N_1286,N_1039);
nand U1676 (N_1676,N_1133,N_1281);
and U1677 (N_1677,N_1372,N_1396);
or U1678 (N_1678,N_1169,N_1410);
nor U1679 (N_1679,N_1360,N_1219);
nor U1680 (N_1680,N_1392,N_1390);
nor U1681 (N_1681,N_1056,N_1097);
nor U1682 (N_1682,N_1354,N_1207);
nand U1683 (N_1683,N_1206,N_1404);
nor U1684 (N_1684,N_1337,N_1144);
nor U1685 (N_1685,N_1310,N_1280);
nor U1686 (N_1686,N_1341,N_1269);
and U1687 (N_1687,N_1451,N_1440);
nand U1688 (N_1688,N_1078,N_1084);
nand U1689 (N_1689,N_1111,N_1416);
and U1690 (N_1690,N_1288,N_1494);
nor U1691 (N_1691,N_1493,N_1399);
nor U1692 (N_1692,N_1427,N_1023);
nor U1693 (N_1693,N_1461,N_1150);
or U1694 (N_1694,N_1005,N_1452);
nor U1695 (N_1695,N_1203,N_1184);
or U1696 (N_1696,N_1418,N_1237);
nor U1697 (N_1697,N_1119,N_1141);
nand U1698 (N_1698,N_1208,N_1443);
or U1699 (N_1699,N_1049,N_1175);
nand U1700 (N_1700,N_1135,N_1189);
nand U1701 (N_1701,N_1364,N_1257);
nor U1702 (N_1702,N_1246,N_1096);
or U1703 (N_1703,N_1188,N_1166);
or U1704 (N_1704,N_1160,N_1221);
or U1705 (N_1705,N_1363,N_1042);
and U1706 (N_1706,N_1082,N_1170);
and U1707 (N_1707,N_1357,N_1041);
nand U1708 (N_1708,N_1028,N_1266);
nand U1709 (N_1709,N_1321,N_1164);
or U1710 (N_1710,N_1200,N_1482);
nor U1711 (N_1711,N_1346,N_1199);
and U1712 (N_1712,N_1120,N_1459);
nand U1713 (N_1713,N_1422,N_1294);
or U1714 (N_1714,N_1128,N_1103);
and U1715 (N_1715,N_1162,N_1263);
or U1716 (N_1716,N_1187,N_1021);
nor U1717 (N_1717,N_1123,N_1151);
and U1718 (N_1718,N_1242,N_1415);
and U1719 (N_1719,N_1463,N_1037);
nand U1720 (N_1720,N_1316,N_1154);
nor U1721 (N_1721,N_1032,N_1209);
nand U1722 (N_1722,N_1395,N_1379);
xor U1723 (N_1723,N_1076,N_1098);
nand U1724 (N_1724,N_1107,N_1300);
nand U1725 (N_1725,N_1254,N_1460);
and U1726 (N_1726,N_1211,N_1369);
nor U1727 (N_1727,N_1024,N_1062);
nand U1728 (N_1728,N_1436,N_1423);
nor U1729 (N_1729,N_1194,N_1241);
or U1730 (N_1730,N_1063,N_1349);
nand U1731 (N_1731,N_1319,N_1386);
or U1732 (N_1732,N_1419,N_1490);
or U1733 (N_1733,N_1400,N_1320);
nor U1734 (N_1734,N_1353,N_1238);
and U1735 (N_1735,N_1447,N_1361);
nor U1736 (N_1736,N_1323,N_1050);
nand U1737 (N_1737,N_1174,N_1304);
nand U1738 (N_1738,N_1413,N_1192);
nor U1739 (N_1739,N_1391,N_1352);
nand U1740 (N_1740,N_1267,N_1090);
and U1741 (N_1741,N_1472,N_1055);
or U1742 (N_1742,N_1326,N_1079);
and U1743 (N_1743,N_1442,N_1350);
and U1744 (N_1744,N_1048,N_1435);
nand U1745 (N_1745,N_1298,N_1121);
nand U1746 (N_1746,N_1122,N_1303);
or U1747 (N_1747,N_1477,N_1302);
or U1748 (N_1748,N_1130,N_1073);
and U1749 (N_1749,N_1183,N_1171);
or U1750 (N_1750,N_1285,N_1306);
nor U1751 (N_1751,N_1268,N_1026);
nand U1752 (N_1752,N_1388,N_1226);
or U1753 (N_1753,N_1475,N_1105);
and U1754 (N_1754,N_1046,N_1073);
or U1755 (N_1755,N_1257,N_1494);
nor U1756 (N_1756,N_1006,N_1394);
nor U1757 (N_1757,N_1292,N_1006);
and U1758 (N_1758,N_1284,N_1348);
nor U1759 (N_1759,N_1437,N_1354);
nor U1760 (N_1760,N_1168,N_1243);
nor U1761 (N_1761,N_1332,N_1106);
nor U1762 (N_1762,N_1114,N_1407);
or U1763 (N_1763,N_1340,N_1468);
nand U1764 (N_1764,N_1159,N_1197);
or U1765 (N_1765,N_1156,N_1059);
and U1766 (N_1766,N_1381,N_1141);
nand U1767 (N_1767,N_1111,N_1479);
or U1768 (N_1768,N_1021,N_1216);
nor U1769 (N_1769,N_1086,N_1184);
or U1770 (N_1770,N_1399,N_1108);
nand U1771 (N_1771,N_1137,N_1118);
or U1772 (N_1772,N_1401,N_1435);
xnor U1773 (N_1773,N_1360,N_1026);
or U1774 (N_1774,N_1467,N_1209);
or U1775 (N_1775,N_1378,N_1366);
or U1776 (N_1776,N_1401,N_1135);
nor U1777 (N_1777,N_1397,N_1056);
and U1778 (N_1778,N_1313,N_1298);
and U1779 (N_1779,N_1394,N_1331);
nand U1780 (N_1780,N_1428,N_1139);
nor U1781 (N_1781,N_1180,N_1015);
or U1782 (N_1782,N_1197,N_1413);
or U1783 (N_1783,N_1375,N_1157);
and U1784 (N_1784,N_1151,N_1192);
or U1785 (N_1785,N_1184,N_1071);
nand U1786 (N_1786,N_1476,N_1120);
or U1787 (N_1787,N_1481,N_1298);
nand U1788 (N_1788,N_1258,N_1283);
nand U1789 (N_1789,N_1171,N_1004);
nand U1790 (N_1790,N_1331,N_1104);
or U1791 (N_1791,N_1138,N_1213);
and U1792 (N_1792,N_1341,N_1298);
and U1793 (N_1793,N_1015,N_1354);
nand U1794 (N_1794,N_1010,N_1168);
nor U1795 (N_1795,N_1215,N_1245);
and U1796 (N_1796,N_1161,N_1176);
nor U1797 (N_1797,N_1408,N_1198);
and U1798 (N_1798,N_1150,N_1076);
and U1799 (N_1799,N_1331,N_1080);
nor U1800 (N_1800,N_1411,N_1123);
and U1801 (N_1801,N_1262,N_1022);
nand U1802 (N_1802,N_1158,N_1127);
or U1803 (N_1803,N_1105,N_1411);
and U1804 (N_1804,N_1362,N_1463);
or U1805 (N_1805,N_1072,N_1239);
and U1806 (N_1806,N_1296,N_1137);
or U1807 (N_1807,N_1181,N_1216);
nand U1808 (N_1808,N_1343,N_1356);
and U1809 (N_1809,N_1457,N_1433);
nor U1810 (N_1810,N_1224,N_1284);
and U1811 (N_1811,N_1475,N_1288);
nand U1812 (N_1812,N_1339,N_1298);
and U1813 (N_1813,N_1317,N_1039);
nand U1814 (N_1814,N_1027,N_1008);
nand U1815 (N_1815,N_1180,N_1468);
nor U1816 (N_1816,N_1171,N_1058);
nor U1817 (N_1817,N_1052,N_1280);
or U1818 (N_1818,N_1238,N_1462);
nor U1819 (N_1819,N_1025,N_1026);
nor U1820 (N_1820,N_1381,N_1280);
and U1821 (N_1821,N_1273,N_1058);
nand U1822 (N_1822,N_1141,N_1104);
or U1823 (N_1823,N_1086,N_1423);
nand U1824 (N_1824,N_1171,N_1436);
xor U1825 (N_1825,N_1217,N_1388);
and U1826 (N_1826,N_1165,N_1352);
and U1827 (N_1827,N_1070,N_1176);
nand U1828 (N_1828,N_1498,N_1372);
nand U1829 (N_1829,N_1087,N_1001);
and U1830 (N_1830,N_1453,N_1176);
nand U1831 (N_1831,N_1455,N_1280);
and U1832 (N_1832,N_1169,N_1468);
or U1833 (N_1833,N_1012,N_1158);
and U1834 (N_1834,N_1161,N_1061);
or U1835 (N_1835,N_1161,N_1314);
or U1836 (N_1836,N_1476,N_1350);
or U1837 (N_1837,N_1334,N_1307);
and U1838 (N_1838,N_1491,N_1299);
and U1839 (N_1839,N_1303,N_1149);
nand U1840 (N_1840,N_1166,N_1232);
nand U1841 (N_1841,N_1223,N_1138);
or U1842 (N_1842,N_1184,N_1034);
nand U1843 (N_1843,N_1008,N_1473);
or U1844 (N_1844,N_1041,N_1129);
nand U1845 (N_1845,N_1131,N_1470);
xor U1846 (N_1846,N_1073,N_1307);
nor U1847 (N_1847,N_1134,N_1320);
and U1848 (N_1848,N_1399,N_1092);
or U1849 (N_1849,N_1191,N_1170);
nor U1850 (N_1850,N_1131,N_1270);
and U1851 (N_1851,N_1037,N_1105);
nand U1852 (N_1852,N_1077,N_1256);
nor U1853 (N_1853,N_1245,N_1041);
nor U1854 (N_1854,N_1230,N_1276);
nand U1855 (N_1855,N_1057,N_1395);
nand U1856 (N_1856,N_1167,N_1379);
nor U1857 (N_1857,N_1024,N_1254);
nand U1858 (N_1858,N_1430,N_1457);
and U1859 (N_1859,N_1272,N_1122);
nor U1860 (N_1860,N_1250,N_1026);
nor U1861 (N_1861,N_1127,N_1369);
and U1862 (N_1862,N_1270,N_1447);
or U1863 (N_1863,N_1125,N_1052);
nor U1864 (N_1864,N_1135,N_1134);
nor U1865 (N_1865,N_1001,N_1123);
or U1866 (N_1866,N_1305,N_1271);
nor U1867 (N_1867,N_1164,N_1435);
nor U1868 (N_1868,N_1354,N_1095);
and U1869 (N_1869,N_1480,N_1274);
nand U1870 (N_1870,N_1347,N_1074);
or U1871 (N_1871,N_1050,N_1228);
and U1872 (N_1872,N_1320,N_1356);
nand U1873 (N_1873,N_1230,N_1250);
or U1874 (N_1874,N_1233,N_1116);
and U1875 (N_1875,N_1350,N_1334);
and U1876 (N_1876,N_1322,N_1485);
nor U1877 (N_1877,N_1076,N_1024);
or U1878 (N_1878,N_1477,N_1099);
nand U1879 (N_1879,N_1225,N_1050);
or U1880 (N_1880,N_1251,N_1322);
nand U1881 (N_1881,N_1152,N_1395);
nand U1882 (N_1882,N_1147,N_1210);
and U1883 (N_1883,N_1356,N_1148);
or U1884 (N_1884,N_1045,N_1443);
nor U1885 (N_1885,N_1125,N_1113);
nand U1886 (N_1886,N_1075,N_1247);
and U1887 (N_1887,N_1268,N_1064);
nor U1888 (N_1888,N_1371,N_1188);
nand U1889 (N_1889,N_1496,N_1263);
and U1890 (N_1890,N_1245,N_1263);
and U1891 (N_1891,N_1067,N_1300);
and U1892 (N_1892,N_1085,N_1438);
nand U1893 (N_1893,N_1185,N_1438);
or U1894 (N_1894,N_1357,N_1101);
and U1895 (N_1895,N_1091,N_1402);
nand U1896 (N_1896,N_1239,N_1224);
nor U1897 (N_1897,N_1382,N_1120);
nor U1898 (N_1898,N_1486,N_1324);
nand U1899 (N_1899,N_1263,N_1033);
or U1900 (N_1900,N_1173,N_1158);
or U1901 (N_1901,N_1067,N_1220);
and U1902 (N_1902,N_1391,N_1251);
nor U1903 (N_1903,N_1271,N_1079);
or U1904 (N_1904,N_1066,N_1130);
nand U1905 (N_1905,N_1458,N_1000);
and U1906 (N_1906,N_1468,N_1301);
and U1907 (N_1907,N_1463,N_1364);
or U1908 (N_1908,N_1056,N_1118);
nand U1909 (N_1909,N_1452,N_1044);
or U1910 (N_1910,N_1499,N_1112);
or U1911 (N_1911,N_1088,N_1242);
and U1912 (N_1912,N_1148,N_1225);
or U1913 (N_1913,N_1243,N_1468);
and U1914 (N_1914,N_1181,N_1359);
nand U1915 (N_1915,N_1256,N_1228);
nand U1916 (N_1916,N_1230,N_1151);
or U1917 (N_1917,N_1030,N_1208);
and U1918 (N_1918,N_1246,N_1440);
nor U1919 (N_1919,N_1261,N_1476);
or U1920 (N_1920,N_1019,N_1341);
nand U1921 (N_1921,N_1331,N_1379);
and U1922 (N_1922,N_1166,N_1248);
nand U1923 (N_1923,N_1408,N_1345);
nand U1924 (N_1924,N_1217,N_1443);
nor U1925 (N_1925,N_1499,N_1198);
nor U1926 (N_1926,N_1113,N_1337);
and U1927 (N_1927,N_1373,N_1009);
nor U1928 (N_1928,N_1382,N_1261);
or U1929 (N_1929,N_1429,N_1349);
and U1930 (N_1930,N_1072,N_1410);
nand U1931 (N_1931,N_1078,N_1284);
nor U1932 (N_1932,N_1161,N_1403);
and U1933 (N_1933,N_1322,N_1000);
xnor U1934 (N_1934,N_1179,N_1387);
or U1935 (N_1935,N_1401,N_1115);
nand U1936 (N_1936,N_1313,N_1035);
and U1937 (N_1937,N_1042,N_1262);
nand U1938 (N_1938,N_1455,N_1422);
nor U1939 (N_1939,N_1345,N_1132);
or U1940 (N_1940,N_1307,N_1452);
and U1941 (N_1941,N_1025,N_1138);
nor U1942 (N_1942,N_1079,N_1076);
or U1943 (N_1943,N_1456,N_1186);
or U1944 (N_1944,N_1170,N_1221);
nor U1945 (N_1945,N_1265,N_1081);
or U1946 (N_1946,N_1408,N_1006);
nand U1947 (N_1947,N_1256,N_1039);
nand U1948 (N_1948,N_1187,N_1257);
or U1949 (N_1949,N_1436,N_1025);
nor U1950 (N_1950,N_1168,N_1334);
and U1951 (N_1951,N_1041,N_1375);
nand U1952 (N_1952,N_1496,N_1253);
or U1953 (N_1953,N_1290,N_1057);
nor U1954 (N_1954,N_1128,N_1056);
and U1955 (N_1955,N_1286,N_1326);
and U1956 (N_1956,N_1048,N_1273);
nand U1957 (N_1957,N_1035,N_1414);
and U1958 (N_1958,N_1373,N_1098);
nand U1959 (N_1959,N_1423,N_1208);
xor U1960 (N_1960,N_1387,N_1039);
or U1961 (N_1961,N_1179,N_1335);
and U1962 (N_1962,N_1417,N_1152);
nand U1963 (N_1963,N_1025,N_1081);
nand U1964 (N_1964,N_1018,N_1179);
nor U1965 (N_1965,N_1427,N_1214);
nand U1966 (N_1966,N_1168,N_1388);
nand U1967 (N_1967,N_1145,N_1347);
nor U1968 (N_1968,N_1367,N_1344);
or U1969 (N_1969,N_1336,N_1348);
nor U1970 (N_1970,N_1069,N_1290);
nor U1971 (N_1971,N_1494,N_1076);
nor U1972 (N_1972,N_1176,N_1058);
and U1973 (N_1973,N_1189,N_1137);
nand U1974 (N_1974,N_1176,N_1193);
nand U1975 (N_1975,N_1297,N_1047);
or U1976 (N_1976,N_1200,N_1214);
and U1977 (N_1977,N_1178,N_1066);
or U1978 (N_1978,N_1191,N_1433);
nor U1979 (N_1979,N_1317,N_1266);
or U1980 (N_1980,N_1283,N_1170);
nand U1981 (N_1981,N_1131,N_1392);
nand U1982 (N_1982,N_1170,N_1486);
nor U1983 (N_1983,N_1000,N_1406);
nor U1984 (N_1984,N_1067,N_1383);
and U1985 (N_1985,N_1402,N_1258);
nor U1986 (N_1986,N_1186,N_1341);
nor U1987 (N_1987,N_1145,N_1019);
and U1988 (N_1988,N_1006,N_1092);
nand U1989 (N_1989,N_1364,N_1170);
or U1990 (N_1990,N_1294,N_1112);
or U1991 (N_1991,N_1410,N_1490);
nor U1992 (N_1992,N_1415,N_1440);
and U1993 (N_1993,N_1322,N_1011);
and U1994 (N_1994,N_1285,N_1119);
or U1995 (N_1995,N_1225,N_1267);
or U1996 (N_1996,N_1495,N_1296);
and U1997 (N_1997,N_1353,N_1336);
or U1998 (N_1998,N_1165,N_1116);
and U1999 (N_1999,N_1300,N_1333);
and U2000 (N_2000,N_1631,N_1775);
nor U2001 (N_2001,N_1820,N_1831);
or U2002 (N_2002,N_1748,N_1567);
or U2003 (N_2003,N_1997,N_1500);
nor U2004 (N_2004,N_1896,N_1787);
and U2005 (N_2005,N_1734,N_1880);
or U2006 (N_2006,N_1900,N_1566);
and U2007 (N_2007,N_1797,N_1601);
and U2008 (N_2008,N_1784,N_1619);
or U2009 (N_2009,N_1836,N_1942);
nor U2010 (N_2010,N_1966,N_1668);
and U2011 (N_2011,N_1945,N_1865);
nor U2012 (N_2012,N_1955,N_1649);
nand U2013 (N_2013,N_1569,N_1572);
nand U2014 (N_2014,N_1749,N_1573);
nor U2015 (N_2015,N_1730,N_1981);
or U2016 (N_2016,N_1946,N_1646);
nand U2017 (N_2017,N_1916,N_1765);
or U2018 (N_2018,N_1568,N_1724);
nand U2019 (N_2019,N_1701,N_1881);
nor U2020 (N_2020,N_1590,N_1764);
nor U2021 (N_2021,N_1517,N_1920);
or U2022 (N_2022,N_1848,N_1849);
nor U2023 (N_2023,N_1729,N_1698);
and U2024 (N_2024,N_1737,N_1702);
and U2025 (N_2025,N_1598,N_1963);
nor U2026 (N_2026,N_1885,N_1861);
nand U2027 (N_2027,N_1659,N_1661);
and U2028 (N_2028,N_1531,N_1964);
nor U2029 (N_2029,N_1965,N_1754);
nand U2030 (N_2030,N_1697,N_1663);
nand U2031 (N_2031,N_1851,N_1662);
or U2032 (N_2032,N_1871,N_1632);
or U2033 (N_2033,N_1579,N_1687);
and U2034 (N_2034,N_1793,N_1919);
nand U2035 (N_2035,N_1895,N_1984);
nand U2036 (N_2036,N_1758,N_1656);
and U2037 (N_2037,N_1892,N_1975);
nand U2038 (N_2038,N_1888,N_1961);
nor U2039 (N_2039,N_1636,N_1533);
nor U2040 (N_2040,N_1501,N_1766);
and U2041 (N_2041,N_1671,N_1937);
nor U2042 (N_2042,N_1982,N_1915);
or U2043 (N_2043,N_1586,N_1930);
and U2044 (N_2044,N_1527,N_1771);
nor U2045 (N_2045,N_1655,N_1824);
or U2046 (N_2046,N_1773,N_1794);
nor U2047 (N_2047,N_1875,N_1745);
or U2048 (N_2048,N_1544,N_1582);
nand U2049 (N_2049,N_1968,N_1502);
nand U2050 (N_2050,N_1938,N_1746);
and U2051 (N_2051,N_1805,N_1756);
or U2052 (N_2052,N_1577,N_1912);
or U2053 (N_2053,N_1904,N_1578);
nand U2054 (N_2054,N_1508,N_1782);
nand U2055 (N_2055,N_1560,N_1506);
or U2056 (N_2056,N_1750,N_1647);
nor U2057 (N_2057,N_1948,N_1600);
nor U2058 (N_2058,N_1993,N_1684);
nand U2059 (N_2059,N_1715,N_1813);
and U2060 (N_2060,N_1726,N_1798);
nor U2061 (N_2061,N_1792,N_1922);
nor U2062 (N_2062,N_1595,N_1510);
and U2063 (N_2063,N_1858,N_1516);
and U2064 (N_2064,N_1983,N_1676);
nor U2065 (N_2065,N_1806,N_1640);
and U2066 (N_2066,N_1995,N_1905);
nor U2067 (N_2067,N_1908,N_1882);
or U2068 (N_2068,N_1866,N_1914);
nand U2069 (N_2069,N_1906,N_1974);
nor U2070 (N_2070,N_1776,N_1522);
and U2071 (N_2071,N_1725,N_1518);
nand U2072 (N_2072,N_1665,N_1845);
or U2073 (N_2073,N_1755,N_1509);
nor U2074 (N_2074,N_1700,N_1778);
or U2075 (N_2075,N_1587,N_1760);
nand U2076 (N_2076,N_1580,N_1648);
nor U2077 (N_2077,N_1660,N_1657);
and U2078 (N_2078,N_1543,N_1802);
or U2079 (N_2079,N_1901,N_1690);
and U2080 (N_2080,N_1694,N_1538);
nand U2081 (N_2081,N_1996,N_1633);
nor U2082 (N_2082,N_1923,N_1894);
nand U2083 (N_2083,N_1994,N_1583);
or U2084 (N_2084,N_1615,N_1673);
nand U2085 (N_2085,N_1744,N_1635);
and U2086 (N_2086,N_1859,N_1712);
nor U2087 (N_2087,N_1971,N_1856);
nand U2088 (N_2088,N_1772,N_1986);
nor U2089 (N_2089,N_1591,N_1514);
nor U2090 (N_2090,N_1990,N_1747);
or U2091 (N_2091,N_1988,N_1785);
nand U2092 (N_2092,N_1989,N_1622);
or U2093 (N_2093,N_1650,N_1852);
nand U2094 (N_2094,N_1672,N_1571);
nor U2095 (N_2095,N_1829,N_1556);
or U2096 (N_2096,N_1873,N_1952);
or U2097 (N_2097,N_1770,N_1999);
nor U2098 (N_2098,N_1523,N_1709);
and U2099 (N_2099,N_1774,N_1921);
nor U2100 (N_2100,N_1821,N_1722);
or U2101 (N_2101,N_1530,N_1757);
or U2102 (N_2102,N_1616,N_1847);
nor U2103 (N_2103,N_1638,N_1608);
or U2104 (N_2104,N_1675,N_1887);
or U2105 (N_2105,N_1507,N_1628);
and U2106 (N_2106,N_1515,N_1819);
and U2107 (N_2107,N_1614,N_1740);
or U2108 (N_2108,N_1893,N_1738);
nand U2109 (N_2109,N_1877,N_1960);
nor U2110 (N_2110,N_1947,N_1634);
or U2111 (N_2111,N_1874,N_1827);
nand U2112 (N_2112,N_1727,N_1951);
and U2113 (N_2113,N_1529,N_1547);
and U2114 (N_2114,N_1610,N_1644);
and U2115 (N_2115,N_1759,N_1589);
or U2116 (N_2116,N_1789,N_1941);
nor U2117 (N_2117,N_1899,N_1599);
or U2118 (N_2118,N_1826,N_1867);
nand U2119 (N_2119,N_1584,N_1788);
nand U2120 (N_2120,N_1557,N_1933);
or U2121 (N_2121,N_1537,N_1605);
nor U2122 (N_2122,N_1504,N_1574);
nor U2123 (N_2123,N_1979,N_1607);
and U2124 (N_2124,N_1843,N_1695);
and U2125 (N_2125,N_1670,N_1932);
and U2126 (N_2126,N_1811,N_1884);
nand U2127 (N_2127,N_1623,N_1834);
or U2128 (N_2128,N_1751,N_1783);
nand U2129 (N_2129,N_1817,N_1704);
nand U2130 (N_2130,N_1553,N_1611);
and U2131 (N_2131,N_1597,N_1588);
nor U2132 (N_2132,N_1902,N_1521);
nand U2133 (N_2133,N_1559,N_1909);
and U2134 (N_2134,N_1763,N_1535);
or U2135 (N_2135,N_1546,N_1864);
or U2136 (N_2136,N_1511,N_1689);
nor U2137 (N_2137,N_1762,N_1603);
nor U2138 (N_2138,N_1703,N_1682);
nand U2139 (N_2139,N_1850,N_1713);
nor U2140 (N_2140,N_1918,N_1736);
or U2141 (N_2141,N_1863,N_1780);
nor U2142 (N_2142,N_1627,N_1653);
nor U2143 (N_2143,N_1869,N_1854);
nand U2144 (N_2144,N_1645,N_1562);
or U2145 (N_2145,N_1803,N_1739);
and U2146 (N_2146,N_1526,N_1609);
nor U2147 (N_2147,N_1800,N_1998);
and U2148 (N_2148,N_1534,N_1992);
nor U2149 (N_2149,N_1666,N_1679);
nand U2150 (N_2150,N_1621,N_1718);
nand U2151 (N_2151,N_1801,N_1812);
nor U2152 (N_2152,N_1551,N_1719);
or U2153 (N_2153,N_1927,N_1924);
or U2154 (N_2154,N_1565,N_1853);
or U2155 (N_2155,N_1620,N_1541);
nor U2156 (N_2156,N_1716,N_1624);
xnor U2157 (N_2157,N_1711,N_1618);
or U2158 (N_2158,N_1581,N_1561);
nor U2159 (N_2159,N_1870,N_1779);
and U2160 (N_2160,N_1532,N_1804);
and U2161 (N_2161,N_1691,N_1707);
nor U2162 (N_2162,N_1939,N_1987);
nand U2163 (N_2163,N_1536,N_1807);
and U2164 (N_2164,N_1903,N_1911);
nand U2165 (N_2165,N_1957,N_1596);
nor U2166 (N_2166,N_1652,N_1592);
or U2167 (N_2167,N_1625,N_1575);
or U2168 (N_2168,N_1825,N_1838);
nor U2169 (N_2169,N_1976,N_1554);
and U2170 (N_2170,N_1814,N_1723);
nor U2171 (N_2171,N_1769,N_1639);
nand U2172 (N_2172,N_1664,N_1910);
nor U2173 (N_2173,N_1889,N_1768);
or U2174 (N_2174,N_1855,N_1970);
nand U2175 (N_2175,N_1777,N_1753);
and U2176 (N_2176,N_1934,N_1860);
nand U2177 (N_2177,N_1840,N_1897);
nor U2178 (N_2178,N_1710,N_1637);
and U2179 (N_2179,N_1728,N_1823);
and U2180 (N_2180,N_1956,N_1962);
nand U2181 (N_2181,N_1721,N_1630);
and U2182 (N_2182,N_1809,N_1949);
and U2183 (N_2183,N_1642,N_1503);
and U2184 (N_2184,N_1980,N_1810);
nand U2185 (N_2185,N_1604,N_1545);
nand U2186 (N_2186,N_1626,N_1576);
nand U2187 (N_2187,N_1818,N_1958);
and U2188 (N_2188,N_1542,N_1950);
and U2189 (N_2189,N_1525,N_1972);
xor U2190 (N_2190,N_1594,N_1841);
nor U2191 (N_2191,N_1549,N_1886);
nand U2192 (N_2192,N_1752,N_1844);
or U2193 (N_2193,N_1781,N_1693);
nand U2194 (N_2194,N_1907,N_1686);
or U2195 (N_2195,N_1846,N_1935);
nor U2196 (N_2196,N_1548,N_1822);
nand U2197 (N_2197,N_1761,N_1735);
and U2198 (N_2198,N_1786,N_1868);
or U2199 (N_2199,N_1977,N_1519);
or U2200 (N_2200,N_1943,N_1732);
and U2201 (N_2201,N_1688,N_1931);
and U2202 (N_2202,N_1641,N_1832);
and U2203 (N_2203,N_1940,N_1883);
nor U2204 (N_2204,N_1528,N_1513);
and U2205 (N_2205,N_1898,N_1552);
or U2206 (N_2206,N_1555,N_1925);
or U2207 (N_2207,N_1917,N_1696);
and U2208 (N_2208,N_1606,N_1862);
nor U2209 (N_2209,N_1959,N_1558);
nand U2210 (N_2210,N_1717,N_1651);
nor U2211 (N_2211,N_1563,N_1683);
nand U2212 (N_2212,N_1954,N_1678);
nor U2213 (N_2213,N_1731,N_1808);
and U2214 (N_2214,N_1878,N_1767);
or U2215 (N_2215,N_1602,N_1570);
or U2216 (N_2216,N_1944,N_1505);
nand U2217 (N_2217,N_1512,N_1973);
and U2218 (N_2218,N_1828,N_1699);
and U2219 (N_2219,N_1706,N_1833);
or U2220 (N_2220,N_1643,N_1978);
nand U2221 (N_2221,N_1742,N_1692);
nand U2222 (N_2222,N_1879,N_1926);
and U2223 (N_2223,N_1585,N_1658);
or U2224 (N_2224,N_1654,N_1876);
nand U2225 (N_2225,N_1796,N_1837);
and U2226 (N_2226,N_1791,N_1795);
nand U2227 (N_2227,N_1815,N_1593);
or U2228 (N_2228,N_1857,N_1991);
nor U2229 (N_2229,N_1685,N_1677);
nand U2230 (N_2230,N_1936,N_1799);
nand U2231 (N_2231,N_1667,N_1613);
and U2232 (N_2232,N_1669,N_1520);
nand U2233 (N_2233,N_1612,N_1629);
nor U2234 (N_2234,N_1872,N_1953);
and U2235 (N_2235,N_1830,N_1720);
and U2236 (N_2236,N_1839,N_1835);
or U2237 (N_2237,N_1524,N_1680);
or U2238 (N_2238,N_1550,N_1705);
nor U2239 (N_2239,N_1617,N_1708);
or U2240 (N_2240,N_1539,N_1842);
or U2241 (N_2241,N_1969,N_1674);
nand U2242 (N_2242,N_1741,N_1928);
or U2243 (N_2243,N_1564,N_1790);
nand U2244 (N_2244,N_1540,N_1891);
and U2245 (N_2245,N_1816,N_1681);
nand U2246 (N_2246,N_1929,N_1714);
nand U2247 (N_2247,N_1733,N_1743);
and U2248 (N_2248,N_1913,N_1890);
or U2249 (N_2249,N_1967,N_1985);
nor U2250 (N_2250,N_1676,N_1896);
nand U2251 (N_2251,N_1873,N_1823);
or U2252 (N_2252,N_1583,N_1565);
and U2253 (N_2253,N_1671,N_1564);
or U2254 (N_2254,N_1964,N_1560);
or U2255 (N_2255,N_1959,N_1529);
and U2256 (N_2256,N_1937,N_1537);
and U2257 (N_2257,N_1950,N_1641);
and U2258 (N_2258,N_1826,N_1871);
nor U2259 (N_2259,N_1918,N_1863);
nor U2260 (N_2260,N_1576,N_1690);
or U2261 (N_2261,N_1751,N_1780);
nand U2262 (N_2262,N_1750,N_1588);
nand U2263 (N_2263,N_1688,N_1714);
nor U2264 (N_2264,N_1672,N_1900);
nand U2265 (N_2265,N_1677,N_1638);
xor U2266 (N_2266,N_1526,N_1819);
or U2267 (N_2267,N_1901,N_1859);
nand U2268 (N_2268,N_1954,N_1512);
nand U2269 (N_2269,N_1546,N_1876);
or U2270 (N_2270,N_1672,N_1761);
or U2271 (N_2271,N_1555,N_1631);
and U2272 (N_2272,N_1777,N_1936);
nor U2273 (N_2273,N_1899,N_1582);
or U2274 (N_2274,N_1982,N_1676);
xor U2275 (N_2275,N_1873,N_1940);
nor U2276 (N_2276,N_1832,N_1561);
or U2277 (N_2277,N_1523,N_1804);
nand U2278 (N_2278,N_1785,N_1843);
nand U2279 (N_2279,N_1912,N_1952);
and U2280 (N_2280,N_1641,N_1853);
nand U2281 (N_2281,N_1572,N_1516);
nor U2282 (N_2282,N_1544,N_1699);
or U2283 (N_2283,N_1815,N_1964);
and U2284 (N_2284,N_1759,N_1816);
and U2285 (N_2285,N_1954,N_1888);
nand U2286 (N_2286,N_1914,N_1870);
or U2287 (N_2287,N_1518,N_1522);
nor U2288 (N_2288,N_1672,N_1754);
and U2289 (N_2289,N_1822,N_1636);
and U2290 (N_2290,N_1853,N_1667);
or U2291 (N_2291,N_1964,N_1580);
nor U2292 (N_2292,N_1617,N_1621);
nor U2293 (N_2293,N_1652,N_1779);
and U2294 (N_2294,N_1704,N_1546);
nand U2295 (N_2295,N_1842,N_1913);
nor U2296 (N_2296,N_1739,N_1697);
or U2297 (N_2297,N_1793,N_1613);
or U2298 (N_2298,N_1608,N_1597);
nor U2299 (N_2299,N_1673,N_1787);
nand U2300 (N_2300,N_1802,N_1663);
nor U2301 (N_2301,N_1966,N_1839);
and U2302 (N_2302,N_1587,N_1885);
nand U2303 (N_2303,N_1592,N_1964);
or U2304 (N_2304,N_1753,N_1919);
and U2305 (N_2305,N_1668,N_1817);
nor U2306 (N_2306,N_1665,N_1978);
and U2307 (N_2307,N_1510,N_1813);
and U2308 (N_2308,N_1853,N_1770);
or U2309 (N_2309,N_1688,N_1905);
and U2310 (N_2310,N_1994,N_1959);
nand U2311 (N_2311,N_1933,N_1658);
or U2312 (N_2312,N_1761,N_1924);
nand U2313 (N_2313,N_1726,N_1532);
nand U2314 (N_2314,N_1782,N_1833);
nor U2315 (N_2315,N_1791,N_1969);
and U2316 (N_2316,N_1671,N_1805);
nand U2317 (N_2317,N_1547,N_1749);
or U2318 (N_2318,N_1907,N_1634);
or U2319 (N_2319,N_1839,N_1937);
nand U2320 (N_2320,N_1706,N_1857);
nand U2321 (N_2321,N_1858,N_1761);
or U2322 (N_2322,N_1787,N_1685);
nor U2323 (N_2323,N_1800,N_1764);
nand U2324 (N_2324,N_1955,N_1743);
and U2325 (N_2325,N_1631,N_1921);
nand U2326 (N_2326,N_1781,N_1994);
nor U2327 (N_2327,N_1980,N_1716);
and U2328 (N_2328,N_1826,N_1640);
nor U2329 (N_2329,N_1514,N_1638);
or U2330 (N_2330,N_1762,N_1862);
or U2331 (N_2331,N_1555,N_1599);
or U2332 (N_2332,N_1698,N_1846);
nor U2333 (N_2333,N_1793,N_1973);
nor U2334 (N_2334,N_1776,N_1595);
or U2335 (N_2335,N_1805,N_1859);
nor U2336 (N_2336,N_1892,N_1570);
nor U2337 (N_2337,N_1613,N_1809);
nand U2338 (N_2338,N_1905,N_1650);
nor U2339 (N_2339,N_1717,N_1732);
and U2340 (N_2340,N_1778,N_1587);
or U2341 (N_2341,N_1567,N_1881);
or U2342 (N_2342,N_1737,N_1907);
nor U2343 (N_2343,N_1949,N_1946);
nand U2344 (N_2344,N_1709,N_1916);
and U2345 (N_2345,N_1679,N_1915);
and U2346 (N_2346,N_1803,N_1876);
or U2347 (N_2347,N_1840,N_1641);
and U2348 (N_2348,N_1708,N_1725);
or U2349 (N_2349,N_1746,N_1563);
nand U2350 (N_2350,N_1578,N_1866);
nand U2351 (N_2351,N_1922,N_1833);
nor U2352 (N_2352,N_1933,N_1911);
nor U2353 (N_2353,N_1890,N_1561);
nand U2354 (N_2354,N_1659,N_1730);
and U2355 (N_2355,N_1738,N_1588);
and U2356 (N_2356,N_1640,N_1754);
or U2357 (N_2357,N_1690,N_1808);
and U2358 (N_2358,N_1618,N_1623);
or U2359 (N_2359,N_1742,N_1655);
nor U2360 (N_2360,N_1662,N_1595);
nand U2361 (N_2361,N_1990,N_1942);
nand U2362 (N_2362,N_1704,N_1589);
and U2363 (N_2363,N_1935,N_1600);
nand U2364 (N_2364,N_1953,N_1795);
and U2365 (N_2365,N_1740,N_1785);
or U2366 (N_2366,N_1774,N_1597);
or U2367 (N_2367,N_1740,N_1562);
and U2368 (N_2368,N_1596,N_1946);
nor U2369 (N_2369,N_1843,N_1802);
nand U2370 (N_2370,N_1557,N_1873);
xnor U2371 (N_2371,N_1870,N_1941);
and U2372 (N_2372,N_1706,N_1703);
nand U2373 (N_2373,N_1614,N_1871);
nand U2374 (N_2374,N_1547,N_1549);
or U2375 (N_2375,N_1706,N_1627);
and U2376 (N_2376,N_1961,N_1958);
nand U2377 (N_2377,N_1525,N_1500);
nand U2378 (N_2378,N_1976,N_1706);
nor U2379 (N_2379,N_1768,N_1965);
or U2380 (N_2380,N_1819,N_1931);
and U2381 (N_2381,N_1629,N_1893);
nand U2382 (N_2382,N_1758,N_1541);
or U2383 (N_2383,N_1827,N_1650);
or U2384 (N_2384,N_1836,N_1819);
nor U2385 (N_2385,N_1936,N_1835);
nand U2386 (N_2386,N_1676,N_1644);
or U2387 (N_2387,N_1732,N_1568);
or U2388 (N_2388,N_1980,N_1970);
or U2389 (N_2389,N_1610,N_1616);
nand U2390 (N_2390,N_1579,N_1958);
and U2391 (N_2391,N_1514,N_1801);
nand U2392 (N_2392,N_1656,N_1625);
and U2393 (N_2393,N_1634,N_1540);
nand U2394 (N_2394,N_1906,N_1606);
or U2395 (N_2395,N_1519,N_1866);
nand U2396 (N_2396,N_1513,N_1730);
or U2397 (N_2397,N_1504,N_1975);
nand U2398 (N_2398,N_1887,N_1831);
nand U2399 (N_2399,N_1643,N_1987);
nand U2400 (N_2400,N_1670,N_1560);
and U2401 (N_2401,N_1517,N_1852);
nand U2402 (N_2402,N_1588,N_1996);
or U2403 (N_2403,N_1758,N_1819);
nand U2404 (N_2404,N_1898,N_1731);
nor U2405 (N_2405,N_1787,N_1947);
or U2406 (N_2406,N_1689,N_1997);
nand U2407 (N_2407,N_1612,N_1671);
or U2408 (N_2408,N_1815,N_1664);
nand U2409 (N_2409,N_1650,N_1944);
nand U2410 (N_2410,N_1544,N_1810);
nand U2411 (N_2411,N_1888,N_1959);
xor U2412 (N_2412,N_1591,N_1648);
nor U2413 (N_2413,N_1584,N_1688);
nand U2414 (N_2414,N_1557,N_1885);
nor U2415 (N_2415,N_1986,N_1787);
nor U2416 (N_2416,N_1864,N_1678);
and U2417 (N_2417,N_1840,N_1956);
or U2418 (N_2418,N_1943,N_1617);
and U2419 (N_2419,N_1744,N_1736);
and U2420 (N_2420,N_1978,N_1585);
and U2421 (N_2421,N_1651,N_1995);
nor U2422 (N_2422,N_1894,N_1893);
or U2423 (N_2423,N_1973,N_1759);
or U2424 (N_2424,N_1668,N_1538);
nor U2425 (N_2425,N_1797,N_1648);
and U2426 (N_2426,N_1647,N_1753);
and U2427 (N_2427,N_1822,N_1623);
nand U2428 (N_2428,N_1951,N_1965);
nor U2429 (N_2429,N_1846,N_1869);
or U2430 (N_2430,N_1697,N_1807);
and U2431 (N_2431,N_1601,N_1519);
and U2432 (N_2432,N_1865,N_1719);
or U2433 (N_2433,N_1777,N_1705);
nor U2434 (N_2434,N_1872,N_1938);
nor U2435 (N_2435,N_1789,N_1622);
or U2436 (N_2436,N_1653,N_1841);
or U2437 (N_2437,N_1990,N_1672);
and U2438 (N_2438,N_1587,N_1838);
or U2439 (N_2439,N_1786,N_1777);
and U2440 (N_2440,N_1750,N_1504);
nor U2441 (N_2441,N_1933,N_1543);
nand U2442 (N_2442,N_1961,N_1984);
nand U2443 (N_2443,N_1903,N_1718);
and U2444 (N_2444,N_1826,N_1702);
nand U2445 (N_2445,N_1616,N_1652);
and U2446 (N_2446,N_1792,N_1627);
and U2447 (N_2447,N_1805,N_1629);
nor U2448 (N_2448,N_1647,N_1901);
or U2449 (N_2449,N_1626,N_1881);
nor U2450 (N_2450,N_1956,N_1630);
and U2451 (N_2451,N_1967,N_1842);
nor U2452 (N_2452,N_1744,N_1689);
nand U2453 (N_2453,N_1830,N_1816);
nand U2454 (N_2454,N_1631,N_1566);
and U2455 (N_2455,N_1644,N_1890);
xnor U2456 (N_2456,N_1776,N_1502);
or U2457 (N_2457,N_1737,N_1739);
nand U2458 (N_2458,N_1806,N_1524);
and U2459 (N_2459,N_1521,N_1616);
nand U2460 (N_2460,N_1759,N_1768);
or U2461 (N_2461,N_1751,N_1743);
nor U2462 (N_2462,N_1996,N_1699);
or U2463 (N_2463,N_1548,N_1830);
nor U2464 (N_2464,N_1786,N_1701);
or U2465 (N_2465,N_1841,N_1711);
and U2466 (N_2466,N_1679,N_1975);
nor U2467 (N_2467,N_1835,N_1916);
nor U2468 (N_2468,N_1967,N_1765);
nor U2469 (N_2469,N_1582,N_1505);
or U2470 (N_2470,N_1618,N_1967);
nor U2471 (N_2471,N_1543,N_1553);
or U2472 (N_2472,N_1918,N_1778);
nand U2473 (N_2473,N_1881,N_1884);
xnor U2474 (N_2474,N_1729,N_1511);
nand U2475 (N_2475,N_1818,N_1880);
nor U2476 (N_2476,N_1721,N_1759);
nor U2477 (N_2477,N_1781,N_1719);
nand U2478 (N_2478,N_1700,N_1544);
nand U2479 (N_2479,N_1770,N_1633);
nor U2480 (N_2480,N_1853,N_1630);
or U2481 (N_2481,N_1898,N_1800);
nand U2482 (N_2482,N_1542,N_1837);
xnor U2483 (N_2483,N_1670,N_1919);
nor U2484 (N_2484,N_1511,N_1653);
and U2485 (N_2485,N_1955,N_1742);
and U2486 (N_2486,N_1719,N_1633);
nor U2487 (N_2487,N_1581,N_1830);
nand U2488 (N_2488,N_1672,N_1512);
and U2489 (N_2489,N_1685,N_1533);
or U2490 (N_2490,N_1623,N_1767);
nor U2491 (N_2491,N_1742,N_1930);
and U2492 (N_2492,N_1671,N_1753);
nand U2493 (N_2493,N_1544,N_1761);
or U2494 (N_2494,N_1591,N_1663);
nand U2495 (N_2495,N_1699,N_1805);
nor U2496 (N_2496,N_1710,N_1969);
nor U2497 (N_2497,N_1789,N_1649);
or U2498 (N_2498,N_1871,N_1709);
or U2499 (N_2499,N_1899,N_1561);
or U2500 (N_2500,N_2116,N_2310);
or U2501 (N_2501,N_2115,N_2060);
or U2502 (N_2502,N_2236,N_2367);
nor U2503 (N_2503,N_2037,N_2247);
nor U2504 (N_2504,N_2369,N_2129);
nand U2505 (N_2505,N_2487,N_2462);
xnor U2506 (N_2506,N_2222,N_2305);
nor U2507 (N_2507,N_2112,N_2482);
or U2508 (N_2508,N_2296,N_2049);
or U2509 (N_2509,N_2366,N_2011);
nor U2510 (N_2510,N_2139,N_2051);
nand U2511 (N_2511,N_2337,N_2355);
nor U2512 (N_2512,N_2365,N_2014);
and U2513 (N_2513,N_2055,N_2453);
and U2514 (N_2514,N_2145,N_2403);
and U2515 (N_2515,N_2009,N_2321);
or U2516 (N_2516,N_2467,N_2298);
and U2517 (N_2517,N_2007,N_2344);
nor U2518 (N_2518,N_2108,N_2197);
and U2519 (N_2519,N_2074,N_2183);
nor U2520 (N_2520,N_2226,N_2280);
nand U2521 (N_2521,N_2312,N_2345);
and U2522 (N_2522,N_2036,N_2028);
or U2523 (N_2523,N_2152,N_2488);
or U2524 (N_2524,N_2350,N_2335);
nor U2525 (N_2525,N_2282,N_2422);
nor U2526 (N_2526,N_2044,N_2409);
and U2527 (N_2527,N_2429,N_2072);
nand U2528 (N_2528,N_2299,N_2033);
and U2529 (N_2529,N_2228,N_2277);
nor U2530 (N_2530,N_2489,N_2245);
and U2531 (N_2531,N_2180,N_2319);
nand U2532 (N_2532,N_2320,N_2169);
or U2533 (N_2533,N_2221,N_2030);
nor U2534 (N_2534,N_2091,N_2371);
and U2535 (N_2535,N_2040,N_2132);
and U2536 (N_2536,N_2164,N_2410);
or U2537 (N_2537,N_2414,N_2356);
nor U2538 (N_2538,N_2032,N_2271);
xnor U2539 (N_2539,N_2084,N_2288);
or U2540 (N_2540,N_2459,N_2000);
and U2541 (N_2541,N_2497,N_2433);
nor U2542 (N_2542,N_2437,N_2346);
or U2543 (N_2543,N_2292,N_2441);
nand U2544 (N_2544,N_2024,N_2191);
nor U2545 (N_2545,N_2223,N_2151);
nand U2546 (N_2546,N_2383,N_2390);
and U2547 (N_2547,N_2008,N_2498);
nand U2548 (N_2548,N_2456,N_2318);
nand U2549 (N_2549,N_2465,N_2314);
nor U2550 (N_2550,N_2206,N_2176);
and U2551 (N_2551,N_2067,N_2159);
and U2552 (N_2552,N_2449,N_2316);
or U2553 (N_2553,N_2405,N_2034);
nor U2554 (N_2554,N_2411,N_2499);
nor U2555 (N_2555,N_2094,N_2204);
and U2556 (N_2556,N_2017,N_2170);
or U2557 (N_2557,N_2003,N_2266);
or U2558 (N_2558,N_2158,N_2398);
and U2559 (N_2559,N_2098,N_2363);
nor U2560 (N_2560,N_2246,N_2184);
nor U2561 (N_2561,N_2291,N_2047);
and U2562 (N_2562,N_2218,N_2205);
and U2563 (N_2563,N_2395,N_2278);
nor U2564 (N_2564,N_2311,N_2479);
nand U2565 (N_2565,N_2481,N_2454);
and U2566 (N_2566,N_2105,N_2213);
or U2567 (N_2567,N_2069,N_2207);
nand U2568 (N_2568,N_2270,N_2334);
nor U2569 (N_2569,N_2463,N_2294);
and U2570 (N_2570,N_2201,N_2285);
nor U2571 (N_2571,N_2413,N_2096);
nor U2572 (N_2572,N_2234,N_2438);
nand U2573 (N_2573,N_2153,N_2005);
nor U2574 (N_2574,N_2124,N_2351);
or U2575 (N_2575,N_2147,N_2202);
and U2576 (N_2576,N_2235,N_2066);
nor U2577 (N_2577,N_2090,N_2237);
and U2578 (N_2578,N_2231,N_2377);
nand U2579 (N_2579,N_2308,N_2391);
xnor U2580 (N_2580,N_2160,N_2379);
nand U2581 (N_2581,N_2209,N_2070);
nand U2582 (N_2582,N_2293,N_2386);
or U2583 (N_2583,N_2196,N_2327);
or U2584 (N_2584,N_2466,N_2264);
and U2585 (N_2585,N_2303,N_2250);
or U2586 (N_2586,N_2057,N_2156);
nor U2587 (N_2587,N_2172,N_2342);
or U2588 (N_2588,N_2210,N_2200);
nor U2589 (N_2589,N_2135,N_2330);
nor U2590 (N_2590,N_2217,N_2452);
and U2591 (N_2591,N_2439,N_2179);
or U2592 (N_2592,N_2307,N_2127);
nor U2593 (N_2593,N_2100,N_2042);
nand U2594 (N_2594,N_2381,N_2259);
nor U2595 (N_2595,N_2078,N_2050);
nor U2596 (N_2596,N_2103,N_2167);
nor U2597 (N_2597,N_2265,N_2359);
nand U2598 (N_2598,N_2415,N_2473);
or U2599 (N_2599,N_2374,N_2175);
nand U2600 (N_2600,N_2338,N_2400);
and U2601 (N_2601,N_2136,N_2494);
nand U2602 (N_2602,N_2284,N_2232);
and U2603 (N_2603,N_2333,N_2272);
and U2604 (N_2604,N_2412,N_2064);
and U2605 (N_2605,N_2077,N_2370);
nor U2606 (N_2606,N_2325,N_2181);
or U2607 (N_2607,N_2140,N_2087);
and U2608 (N_2608,N_2029,N_2276);
or U2609 (N_2609,N_2483,N_2323);
nand U2610 (N_2610,N_2297,N_2134);
nand U2611 (N_2611,N_2031,N_2387);
nand U2612 (N_2612,N_2025,N_2171);
and U2613 (N_2613,N_2089,N_2052);
and U2614 (N_2614,N_2262,N_2464);
or U2615 (N_2615,N_2404,N_2239);
or U2616 (N_2616,N_2434,N_2068);
nand U2617 (N_2617,N_2469,N_2058);
or U2618 (N_2618,N_2336,N_2255);
nand U2619 (N_2619,N_2023,N_2130);
and U2620 (N_2620,N_2418,N_2062);
nor U2621 (N_2621,N_2249,N_2475);
nor U2622 (N_2622,N_2182,N_2461);
or U2623 (N_2623,N_2491,N_2476);
and U2624 (N_2624,N_2406,N_2106);
or U2625 (N_2625,N_2486,N_2141);
nand U2626 (N_2626,N_2382,N_2079);
and U2627 (N_2627,N_2065,N_2004);
nor U2628 (N_2628,N_2195,N_2021);
nand U2629 (N_2629,N_2286,N_2485);
nand U2630 (N_2630,N_2394,N_2402);
nor U2631 (N_2631,N_2053,N_2093);
and U2632 (N_2632,N_2484,N_2086);
and U2633 (N_2633,N_2080,N_2443);
nand U2634 (N_2634,N_2426,N_2375);
or U2635 (N_2635,N_2309,N_2424);
or U2636 (N_2636,N_2144,N_2243);
nand U2637 (N_2637,N_2177,N_2254);
nor U2638 (N_2638,N_2161,N_2117);
or U2639 (N_2639,N_2348,N_2347);
nand U2640 (N_2640,N_2211,N_2075);
nor U2641 (N_2641,N_2146,N_2378);
nor U2642 (N_2642,N_2421,N_2107);
or U2643 (N_2643,N_2490,N_2353);
nor U2644 (N_2644,N_2142,N_2263);
and U2645 (N_2645,N_2495,N_2315);
nor U2646 (N_2646,N_2155,N_2471);
nor U2647 (N_2647,N_2099,N_2267);
or U2648 (N_2648,N_2457,N_2419);
or U2649 (N_2649,N_2339,N_2396);
nand U2650 (N_2650,N_2214,N_2193);
nand U2651 (N_2651,N_2240,N_2474);
nor U2652 (N_2652,N_2341,N_2428);
nor U2653 (N_2653,N_2046,N_2258);
and U2654 (N_2654,N_2137,N_2372);
nand U2655 (N_2655,N_2198,N_2120);
xnor U2656 (N_2656,N_2219,N_2477);
and U2657 (N_2657,N_2361,N_2445);
nor U2658 (N_2658,N_2492,N_2302);
or U2659 (N_2659,N_2056,N_2442);
nand U2660 (N_2660,N_2216,N_2225);
nand U2661 (N_2661,N_2328,N_2480);
nor U2662 (N_2662,N_2111,N_2451);
nand U2663 (N_2663,N_2352,N_2035);
nor U2664 (N_2664,N_2331,N_2446);
nor U2665 (N_2665,N_2012,N_2455);
or U2666 (N_2666,N_2189,N_2038);
and U2667 (N_2667,N_2432,N_2119);
nand U2668 (N_2668,N_2022,N_2229);
nand U2669 (N_2669,N_2110,N_2054);
nor U2670 (N_2670,N_2076,N_2283);
nor U2671 (N_2671,N_2427,N_2041);
or U2672 (N_2672,N_2397,N_2138);
nor U2673 (N_2673,N_2496,N_2244);
or U2674 (N_2674,N_2043,N_2125);
and U2675 (N_2675,N_2015,N_2408);
nand U2676 (N_2676,N_2450,N_2287);
or U2677 (N_2677,N_2006,N_2185);
nor U2678 (N_2678,N_2083,N_2092);
and U2679 (N_2679,N_2118,N_2256);
nand U2680 (N_2680,N_2121,N_2238);
nor U2681 (N_2681,N_2313,N_2300);
and U2682 (N_2682,N_2039,N_2131);
or U2683 (N_2683,N_2447,N_2261);
nand U2684 (N_2684,N_2220,N_2349);
nand U2685 (N_2685,N_2279,N_2324);
nand U2686 (N_2686,N_2393,N_2368);
and U2687 (N_2687,N_2085,N_2045);
nor U2688 (N_2688,N_2149,N_2002);
and U2689 (N_2689,N_2001,N_2020);
and U2690 (N_2690,N_2174,N_2304);
nor U2691 (N_2691,N_2097,N_2326);
and U2692 (N_2692,N_2444,N_2269);
xnor U2693 (N_2693,N_2260,N_2088);
and U2694 (N_2694,N_2026,N_2194);
and U2695 (N_2695,N_2157,N_2010);
and U2696 (N_2696,N_2436,N_2357);
or U2697 (N_2697,N_2212,N_2373);
nand U2698 (N_2698,N_2163,N_2448);
or U2699 (N_2699,N_2203,N_2364);
and U2700 (N_2700,N_2102,N_2224);
and U2701 (N_2701,N_2248,N_2317);
or U2702 (N_2702,N_2168,N_2425);
nor U2703 (N_2703,N_2407,N_2460);
nor U2704 (N_2704,N_2019,N_2470);
nand U2705 (N_2705,N_2430,N_2376);
and U2706 (N_2706,N_2192,N_2478);
nand U2707 (N_2707,N_2027,N_2362);
nand U2708 (N_2708,N_2230,N_2186);
nor U2709 (N_2709,N_2241,N_2389);
and U2710 (N_2710,N_2431,N_2178);
nand U2711 (N_2711,N_2360,N_2128);
nor U2712 (N_2712,N_2190,N_2468);
nand U2713 (N_2713,N_2329,N_2187);
nor U2714 (N_2714,N_2275,N_2281);
and U2715 (N_2715,N_2013,N_2435);
nor U2716 (N_2716,N_2257,N_2401);
nor U2717 (N_2717,N_2332,N_2122);
nor U2718 (N_2718,N_2143,N_2289);
nand U2719 (N_2719,N_2420,N_2458);
nand U2720 (N_2720,N_2472,N_2399);
nand U2721 (N_2721,N_2252,N_2380);
nor U2722 (N_2722,N_2301,N_2150);
and U2723 (N_2723,N_2104,N_2188);
nor U2724 (N_2724,N_2173,N_2071);
nand U2725 (N_2725,N_2126,N_2388);
nand U2726 (N_2726,N_2416,N_2162);
or U2727 (N_2727,N_2208,N_2295);
nor U2728 (N_2728,N_2081,N_2016);
or U2729 (N_2729,N_2423,N_2154);
nor U2730 (N_2730,N_2113,N_2440);
nand U2731 (N_2731,N_2322,N_2215);
nor U2732 (N_2732,N_2384,N_2340);
or U2733 (N_2733,N_2306,N_2148);
nor U2734 (N_2734,N_2199,N_2227);
and U2735 (N_2735,N_2385,N_2417);
or U2736 (N_2736,N_2082,N_2343);
nand U2737 (N_2737,N_2123,N_2233);
nor U2738 (N_2738,N_2392,N_2274);
or U2739 (N_2739,N_2063,N_2109);
nand U2740 (N_2740,N_2358,N_2165);
or U2741 (N_2741,N_2048,N_2354);
nor U2742 (N_2742,N_2242,N_2166);
or U2743 (N_2743,N_2493,N_2073);
and U2744 (N_2744,N_2114,N_2101);
xor U2745 (N_2745,N_2095,N_2268);
nor U2746 (N_2746,N_2133,N_2251);
and U2747 (N_2747,N_2018,N_2061);
and U2748 (N_2748,N_2253,N_2290);
nand U2749 (N_2749,N_2273,N_2059);
nand U2750 (N_2750,N_2267,N_2346);
or U2751 (N_2751,N_2308,N_2493);
nor U2752 (N_2752,N_2022,N_2234);
nand U2753 (N_2753,N_2433,N_2161);
nor U2754 (N_2754,N_2394,N_2491);
and U2755 (N_2755,N_2336,N_2436);
nor U2756 (N_2756,N_2164,N_2303);
nor U2757 (N_2757,N_2369,N_2053);
nand U2758 (N_2758,N_2419,N_2105);
nor U2759 (N_2759,N_2222,N_2199);
nor U2760 (N_2760,N_2465,N_2240);
or U2761 (N_2761,N_2280,N_2246);
nand U2762 (N_2762,N_2148,N_2404);
and U2763 (N_2763,N_2471,N_2357);
or U2764 (N_2764,N_2138,N_2328);
nand U2765 (N_2765,N_2398,N_2058);
and U2766 (N_2766,N_2182,N_2395);
nor U2767 (N_2767,N_2189,N_2281);
or U2768 (N_2768,N_2413,N_2012);
nor U2769 (N_2769,N_2407,N_2327);
or U2770 (N_2770,N_2414,N_2243);
nand U2771 (N_2771,N_2310,N_2009);
or U2772 (N_2772,N_2180,N_2350);
or U2773 (N_2773,N_2098,N_2194);
or U2774 (N_2774,N_2288,N_2204);
and U2775 (N_2775,N_2483,N_2055);
nor U2776 (N_2776,N_2022,N_2394);
nor U2777 (N_2777,N_2458,N_2028);
and U2778 (N_2778,N_2040,N_2116);
nand U2779 (N_2779,N_2460,N_2445);
nor U2780 (N_2780,N_2127,N_2457);
nand U2781 (N_2781,N_2221,N_2409);
nor U2782 (N_2782,N_2291,N_2221);
and U2783 (N_2783,N_2423,N_2347);
nor U2784 (N_2784,N_2100,N_2135);
and U2785 (N_2785,N_2164,N_2268);
nor U2786 (N_2786,N_2044,N_2165);
nor U2787 (N_2787,N_2466,N_2313);
or U2788 (N_2788,N_2195,N_2459);
nand U2789 (N_2789,N_2151,N_2076);
nand U2790 (N_2790,N_2296,N_2418);
nor U2791 (N_2791,N_2080,N_2478);
or U2792 (N_2792,N_2443,N_2449);
or U2793 (N_2793,N_2467,N_2492);
or U2794 (N_2794,N_2253,N_2368);
or U2795 (N_2795,N_2137,N_2367);
or U2796 (N_2796,N_2027,N_2467);
and U2797 (N_2797,N_2354,N_2285);
nand U2798 (N_2798,N_2144,N_2386);
and U2799 (N_2799,N_2415,N_2049);
or U2800 (N_2800,N_2468,N_2109);
nand U2801 (N_2801,N_2053,N_2332);
or U2802 (N_2802,N_2451,N_2268);
or U2803 (N_2803,N_2187,N_2312);
and U2804 (N_2804,N_2177,N_2112);
and U2805 (N_2805,N_2369,N_2381);
or U2806 (N_2806,N_2308,N_2172);
and U2807 (N_2807,N_2289,N_2043);
nor U2808 (N_2808,N_2212,N_2278);
and U2809 (N_2809,N_2273,N_2280);
nor U2810 (N_2810,N_2353,N_2304);
and U2811 (N_2811,N_2346,N_2397);
nand U2812 (N_2812,N_2371,N_2292);
and U2813 (N_2813,N_2118,N_2020);
nor U2814 (N_2814,N_2109,N_2249);
or U2815 (N_2815,N_2124,N_2116);
nand U2816 (N_2816,N_2209,N_2360);
or U2817 (N_2817,N_2352,N_2275);
nand U2818 (N_2818,N_2382,N_2303);
and U2819 (N_2819,N_2068,N_2364);
and U2820 (N_2820,N_2496,N_2377);
nor U2821 (N_2821,N_2053,N_2071);
and U2822 (N_2822,N_2270,N_2006);
nand U2823 (N_2823,N_2055,N_2058);
nand U2824 (N_2824,N_2383,N_2336);
and U2825 (N_2825,N_2274,N_2378);
and U2826 (N_2826,N_2291,N_2364);
nor U2827 (N_2827,N_2369,N_2385);
and U2828 (N_2828,N_2418,N_2457);
and U2829 (N_2829,N_2286,N_2408);
nand U2830 (N_2830,N_2136,N_2296);
and U2831 (N_2831,N_2301,N_2393);
or U2832 (N_2832,N_2331,N_2461);
nor U2833 (N_2833,N_2191,N_2154);
nor U2834 (N_2834,N_2314,N_2442);
or U2835 (N_2835,N_2073,N_2343);
nor U2836 (N_2836,N_2318,N_2174);
or U2837 (N_2837,N_2043,N_2483);
nand U2838 (N_2838,N_2077,N_2408);
or U2839 (N_2839,N_2075,N_2082);
nand U2840 (N_2840,N_2232,N_2423);
nor U2841 (N_2841,N_2422,N_2057);
and U2842 (N_2842,N_2179,N_2288);
nand U2843 (N_2843,N_2143,N_2141);
nand U2844 (N_2844,N_2009,N_2151);
nor U2845 (N_2845,N_2187,N_2101);
nand U2846 (N_2846,N_2027,N_2447);
nor U2847 (N_2847,N_2022,N_2404);
nor U2848 (N_2848,N_2236,N_2262);
nor U2849 (N_2849,N_2384,N_2215);
and U2850 (N_2850,N_2420,N_2494);
nor U2851 (N_2851,N_2251,N_2088);
and U2852 (N_2852,N_2456,N_2201);
and U2853 (N_2853,N_2260,N_2046);
nand U2854 (N_2854,N_2434,N_2116);
and U2855 (N_2855,N_2095,N_2078);
and U2856 (N_2856,N_2358,N_2159);
or U2857 (N_2857,N_2026,N_2394);
nor U2858 (N_2858,N_2102,N_2219);
and U2859 (N_2859,N_2037,N_2255);
and U2860 (N_2860,N_2397,N_2070);
nor U2861 (N_2861,N_2263,N_2027);
nor U2862 (N_2862,N_2241,N_2084);
and U2863 (N_2863,N_2194,N_2071);
nand U2864 (N_2864,N_2434,N_2122);
nand U2865 (N_2865,N_2031,N_2144);
and U2866 (N_2866,N_2431,N_2227);
nor U2867 (N_2867,N_2421,N_2372);
nor U2868 (N_2868,N_2084,N_2078);
nand U2869 (N_2869,N_2189,N_2262);
or U2870 (N_2870,N_2361,N_2469);
and U2871 (N_2871,N_2144,N_2435);
and U2872 (N_2872,N_2417,N_2331);
nand U2873 (N_2873,N_2236,N_2429);
and U2874 (N_2874,N_2227,N_2384);
and U2875 (N_2875,N_2060,N_2180);
nand U2876 (N_2876,N_2296,N_2001);
or U2877 (N_2877,N_2240,N_2163);
xnor U2878 (N_2878,N_2038,N_2073);
nand U2879 (N_2879,N_2308,N_2468);
nand U2880 (N_2880,N_2030,N_2104);
and U2881 (N_2881,N_2078,N_2167);
or U2882 (N_2882,N_2495,N_2346);
or U2883 (N_2883,N_2183,N_2039);
nand U2884 (N_2884,N_2154,N_2248);
and U2885 (N_2885,N_2389,N_2273);
nor U2886 (N_2886,N_2467,N_2132);
nand U2887 (N_2887,N_2295,N_2407);
nand U2888 (N_2888,N_2432,N_2053);
or U2889 (N_2889,N_2107,N_2415);
or U2890 (N_2890,N_2349,N_2306);
nor U2891 (N_2891,N_2279,N_2448);
nand U2892 (N_2892,N_2064,N_2156);
nand U2893 (N_2893,N_2357,N_2297);
xor U2894 (N_2894,N_2194,N_2021);
nor U2895 (N_2895,N_2078,N_2003);
nor U2896 (N_2896,N_2408,N_2129);
or U2897 (N_2897,N_2051,N_2123);
and U2898 (N_2898,N_2495,N_2267);
nand U2899 (N_2899,N_2068,N_2079);
nor U2900 (N_2900,N_2067,N_2231);
or U2901 (N_2901,N_2424,N_2441);
nor U2902 (N_2902,N_2456,N_2223);
and U2903 (N_2903,N_2167,N_2267);
nor U2904 (N_2904,N_2375,N_2085);
nand U2905 (N_2905,N_2483,N_2112);
or U2906 (N_2906,N_2068,N_2104);
nor U2907 (N_2907,N_2042,N_2499);
nand U2908 (N_2908,N_2432,N_2200);
nand U2909 (N_2909,N_2408,N_2375);
nor U2910 (N_2910,N_2215,N_2439);
and U2911 (N_2911,N_2463,N_2004);
and U2912 (N_2912,N_2151,N_2496);
nand U2913 (N_2913,N_2024,N_2456);
and U2914 (N_2914,N_2123,N_2388);
or U2915 (N_2915,N_2121,N_2397);
and U2916 (N_2916,N_2007,N_2330);
and U2917 (N_2917,N_2254,N_2357);
nor U2918 (N_2918,N_2031,N_2322);
and U2919 (N_2919,N_2391,N_2182);
nor U2920 (N_2920,N_2462,N_2121);
and U2921 (N_2921,N_2021,N_2312);
nand U2922 (N_2922,N_2379,N_2048);
or U2923 (N_2923,N_2270,N_2017);
nor U2924 (N_2924,N_2157,N_2144);
nand U2925 (N_2925,N_2012,N_2017);
or U2926 (N_2926,N_2025,N_2182);
or U2927 (N_2927,N_2039,N_2114);
nor U2928 (N_2928,N_2010,N_2174);
and U2929 (N_2929,N_2417,N_2144);
or U2930 (N_2930,N_2347,N_2167);
nand U2931 (N_2931,N_2421,N_2090);
or U2932 (N_2932,N_2243,N_2240);
nor U2933 (N_2933,N_2312,N_2318);
or U2934 (N_2934,N_2422,N_2335);
nand U2935 (N_2935,N_2231,N_2044);
nand U2936 (N_2936,N_2416,N_2465);
nor U2937 (N_2937,N_2106,N_2299);
nor U2938 (N_2938,N_2044,N_2170);
xnor U2939 (N_2939,N_2162,N_2451);
or U2940 (N_2940,N_2095,N_2054);
or U2941 (N_2941,N_2202,N_2001);
nor U2942 (N_2942,N_2486,N_2162);
and U2943 (N_2943,N_2446,N_2476);
and U2944 (N_2944,N_2225,N_2274);
nor U2945 (N_2945,N_2218,N_2144);
or U2946 (N_2946,N_2293,N_2337);
and U2947 (N_2947,N_2349,N_2333);
nand U2948 (N_2948,N_2029,N_2173);
and U2949 (N_2949,N_2315,N_2332);
nand U2950 (N_2950,N_2017,N_2059);
and U2951 (N_2951,N_2228,N_2288);
nor U2952 (N_2952,N_2494,N_2197);
nand U2953 (N_2953,N_2068,N_2403);
or U2954 (N_2954,N_2141,N_2431);
xor U2955 (N_2955,N_2465,N_2334);
and U2956 (N_2956,N_2281,N_2483);
nand U2957 (N_2957,N_2138,N_2189);
and U2958 (N_2958,N_2201,N_2323);
or U2959 (N_2959,N_2262,N_2461);
or U2960 (N_2960,N_2074,N_2032);
nand U2961 (N_2961,N_2464,N_2116);
nor U2962 (N_2962,N_2032,N_2292);
nor U2963 (N_2963,N_2448,N_2245);
and U2964 (N_2964,N_2176,N_2455);
nor U2965 (N_2965,N_2091,N_2461);
nand U2966 (N_2966,N_2177,N_2409);
nand U2967 (N_2967,N_2455,N_2407);
and U2968 (N_2968,N_2495,N_2106);
or U2969 (N_2969,N_2041,N_2491);
and U2970 (N_2970,N_2002,N_2185);
and U2971 (N_2971,N_2273,N_2257);
nand U2972 (N_2972,N_2095,N_2213);
nor U2973 (N_2973,N_2035,N_2298);
or U2974 (N_2974,N_2417,N_2164);
xnor U2975 (N_2975,N_2263,N_2083);
nand U2976 (N_2976,N_2485,N_2104);
nand U2977 (N_2977,N_2248,N_2489);
or U2978 (N_2978,N_2340,N_2284);
nor U2979 (N_2979,N_2107,N_2184);
or U2980 (N_2980,N_2286,N_2185);
xor U2981 (N_2981,N_2411,N_2047);
and U2982 (N_2982,N_2374,N_2327);
or U2983 (N_2983,N_2144,N_2158);
and U2984 (N_2984,N_2083,N_2292);
and U2985 (N_2985,N_2293,N_2363);
or U2986 (N_2986,N_2339,N_2161);
nand U2987 (N_2987,N_2248,N_2419);
nor U2988 (N_2988,N_2356,N_2134);
nand U2989 (N_2989,N_2061,N_2373);
xnor U2990 (N_2990,N_2152,N_2485);
or U2991 (N_2991,N_2324,N_2250);
and U2992 (N_2992,N_2214,N_2099);
or U2993 (N_2993,N_2182,N_2332);
nor U2994 (N_2994,N_2308,N_2009);
and U2995 (N_2995,N_2419,N_2232);
xnor U2996 (N_2996,N_2360,N_2469);
or U2997 (N_2997,N_2190,N_2297);
and U2998 (N_2998,N_2381,N_2183);
nor U2999 (N_2999,N_2264,N_2192);
nor UO_0 (O_0,N_2589,N_2724);
nor UO_1 (O_1,N_2790,N_2794);
or UO_2 (O_2,N_2690,N_2560);
or UO_3 (O_3,N_2674,N_2538);
nand UO_4 (O_4,N_2519,N_2749);
or UO_5 (O_5,N_2872,N_2715);
and UO_6 (O_6,N_2796,N_2681);
and UO_7 (O_7,N_2533,N_2734);
nand UO_8 (O_8,N_2858,N_2532);
and UO_9 (O_9,N_2844,N_2861);
nand UO_10 (O_10,N_2615,N_2798);
nor UO_11 (O_11,N_2856,N_2626);
and UO_12 (O_12,N_2832,N_2647);
and UO_13 (O_13,N_2879,N_2621);
nor UO_14 (O_14,N_2812,N_2608);
and UO_15 (O_15,N_2933,N_2887);
or UO_16 (O_16,N_2962,N_2731);
nor UO_17 (O_17,N_2574,N_2946);
nor UO_18 (O_18,N_2776,N_2722);
or UO_19 (O_19,N_2509,N_2991);
or UO_20 (O_20,N_2646,N_2859);
nor UO_21 (O_21,N_2765,N_2529);
and UO_22 (O_22,N_2865,N_2912);
nor UO_23 (O_23,N_2837,N_2672);
nor UO_24 (O_24,N_2809,N_2632);
or UO_25 (O_25,N_2683,N_2945);
nand UO_26 (O_26,N_2652,N_2886);
xor UO_27 (O_27,N_2738,N_2575);
nand UO_28 (O_28,N_2829,N_2642);
and UO_29 (O_29,N_2736,N_2663);
or UO_30 (O_30,N_2511,N_2508);
or UO_31 (O_31,N_2673,N_2970);
nand UO_32 (O_32,N_2655,N_2782);
nor UO_33 (O_33,N_2956,N_2935);
and UO_34 (O_34,N_2840,N_2685);
and UO_35 (O_35,N_2635,N_2803);
or UO_36 (O_36,N_2843,N_2506);
nor UO_37 (O_37,N_2781,N_2658);
xor UO_38 (O_38,N_2791,N_2526);
and UO_39 (O_39,N_2855,N_2628);
nand UO_40 (O_40,N_2810,N_2593);
nor UO_41 (O_41,N_2762,N_2750);
and UO_42 (O_42,N_2889,N_2664);
nor UO_43 (O_43,N_2540,N_2634);
nand UO_44 (O_44,N_2727,N_2691);
nor UO_45 (O_45,N_2981,N_2878);
nand UO_46 (O_46,N_2815,N_2542);
and UO_47 (O_47,N_2573,N_2600);
and UO_48 (O_48,N_2666,N_2951);
and UO_49 (O_49,N_2982,N_2813);
nor UO_50 (O_50,N_2641,N_2607);
nand UO_51 (O_51,N_2637,N_2692);
nor UO_52 (O_52,N_2612,N_2898);
and UO_53 (O_53,N_2834,N_2741);
nor UO_54 (O_54,N_2960,N_2597);
nand UO_55 (O_55,N_2839,N_2604);
and UO_56 (O_56,N_2622,N_2869);
and UO_57 (O_57,N_2548,N_2842);
nor UO_58 (O_58,N_2943,N_2989);
or UO_59 (O_59,N_2510,N_2742);
nor UO_60 (O_60,N_2871,N_2884);
nand UO_61 (O_61,N_2702,N_2732);
nand UO_62 (O_62,N_2903,N_2936);
and UO_63 (O_63,N_2712,N_2649);
and UO_64 (O_64,N_2864,N_2866);
or UO_65 (O_65,N_2583,N_2805);
or UO_66 (O_66,N_2789,N_2890);
nand UO_67 (O_67,N_2678,N_2831);
and UO_68 (O_68,N_2667,N_2881);
or UO_69 (O_69,N_2932,N_2979);
or UO_70 (O_70,N_2744,N_2701);
nor UO_71 (O_71,N_2971,N_2894);
nor UO_72 (O_72,N_2984,N_2916);
nand UO_73 (O_73,N_2908,N_2630);
or UO_74 (O_74,N_2562,N_2696);
nand UO_75 (O_75,N_2503,N_2747);
nand UO_76 (O_76,N_2917,N_2523);
or UO_77 (O_77,N_2624,N_2759);
nor UO_78 (O_78,N_2975,N_2687);
and UO_79 (O_79,N_2717,N_2949);
nor UO_80 (O_80,N_2910,N_2950);
and UO_81 (O_81,N_2927,N_2870);
or UO_82 (O_82,N_2850,N_2911);
and UO_83 (O_83,N_2594,N_2543);
or UO_84 (O_84,N_2801,N_2901);
nand UO_85 (O_85,N_2785,N_2814);
nor UO_86 (O_86,N_2918,N_2558);
nor UO_87 (O_87,N_2599,N_2768);
and UO_88 (O_88,N_2826,N_2955);
or UO_89 (O_89,N_2693,N_2671);
nor UO_90 (O_90,N_2883,N_2587);
xor UO_91 (O_91,N_2576,N_2660);
nor UO_92 (O_92,N_2899,N_2877);
or UO_93 (O_93,N_2875,N_2958);
nand UO_94 (O_94,N_2553,N_2645);
nand UO_95 (O_95,N_2857,N_2686);
nor UO_96 (O_96,N_2682,N_2760);
and UO_97 (O_97,N_2662,N_2797);
nand UO_98 (O_98,N_2851,N_2852);
or UO_99 (O_99,N_2627,N_2518);
and UO_100 (O_100,N_2816,N_2515);
nor UO_101 (O_101,N_2751,N_2728);
nand UO_102 (O_102,N_2570,N_2688);
nand UO_103 (O_103,N_2720,N_2601);
nand UO_104 (O_104,N_2923,N_2572);
or UO_105 (O_105,N_2948,N_2530);
nand UO_106 (O_106,N_2648,N_2522);
or UO_107 (O_107,N_2609,N_2500);
xor UO_108 (O_108,N_2983,N_2555);
or UO_109 (O_109,N_2920,N_2788);
nand UO_110 (O_110,N_2939,N_2959);
and UO_111 (O_111,N_2610,N_2885);
or UO_112 (O_112,N_2703,N_2915);
nor UO_113 (O_113,N_2531,N_2528);
and UO_114 (O_114,N_2643,N_2748);
nor UO_115 (O_115,N_2714,N_2656);
and UO_116 (O_116,N_2502,N_2501);
nand UO_117 (O_117,N_2629,N_2633);
or UO_118 (O_118,N_2735,N_2675);
nor UO_119 (O_119,N_2819,N_2631);
and UO_120 (O_120,N_2704,N_2778);
and UO_121 (O_121,N_2998,N_2914);
and UO_122 (O_122,N_2824,N_2811);
nor UO_123 (O_123,N_2694,N_2669);
nand UO_124 (O_124,N_2758,N_2513);
nor UO_125 (O_125,N_2930,N_2623);
nor UO_126 (O_126,N_2677,N_2584);
nand UO_127 (O_127,N_2854,N_2756);
nand UO_128 (O_128,N_2964,N_2900);
nor UO_129 (O_129,N_2755,N_2557);
or UO_130 (O_130,N_2638,N_2980);
nand UO_131 (O_131,N_2567,N_2876);
and UO_132 (O_132,N_2947,N_2992);
nand UO_133 (O_133,N_2718,N_2619);
nand UO_134 (O_134,N_2963,N_2716);
nor UO_135 (O_135,N_2569,N_2772);
nand UO_136 (O_136,N_2568,N_2783);
or UO_137 (O_137,N_2670,N_2746);
and UO_138 (O_138,N_2591,N_2867);
nor UO_139 (O_139,N_2639,N_2954);
and UO_140 (O_140,N_2986,N_2792);
or UO_141 (O_141,N_2953,N_2997);
nor UO_142 (O_142,N_2689,N_2541);
or UO_143 (O_143,N_2577,N_2882);
nand UO_144 (O_144,N_2547,N_2723);
nor UO_145 (O_145,N_2713,N_2896);
nor UO_146 (O_146,N_2521,N_2551);
and UO_147 (O_147,N_2895,N_2769);
and UO_148 (O_148,N_2847,N_2868);
and UO_149 (O_149,N_2525,N_2514);
nor UO_150 (O_150,N_2793,N_2880);
and UO_151 (O_151,N_2988,N_2775);
nor UO_152 (O_152,N_2873,N_2761);
nor UO_153 (O_153,N_2517,N_2725);
nand UO_154 (O_154,N_2990,N_2684);
nor UO_155 (O_155,N_2544,N_2657);
and UO_156 (O_156,N_2773,N_2611);
and UO_157 (O_157,N_2770,N_2679);
and UO_158 (O_158,N_2571,N_2640);
and UO_159 (O_159,N_2780,N_2994);
nor UO_160 (O_160,N_2730,N_2737);
and UO_161 (O_161,N_2897,N_2937);
or UO_162 (O_162,N_2919,N_2905);
or UO_163 (O_163,N_2833,N_2706);
and UO_164 (O_164,N_2974,N_2556);
nor UO_165 (O_165,N_2996,N_2743);
nand UO_166 (O_166,N_2973,N_2563);
nor UO_167 (O_167,N_2565,N_2554);
nand UO_168 (O_168,N_2764,N_2733);
nor UO_169 (O_169,N_2680,N_2605);
nor UO_170 (O_170,N_2707,N_2938);
nand UO_171 (O_171,N_2698,N_2729);
nor UO_172 (O_172,N_2695,N_2891);
or UO_173 (O_173,N_2754,N_2827);
nand UO_174 (O_174,N_2952,N_2838);
or UO_175 (O_175,N_2863,N_2676);
or UO_176 (O_176,N_2926,N_2909);
nand UO_177 (O_177,N_2820,N_2752);
nor UO_178 (O_178,N_2825,N_2512);
nand UO_179 (O_179,N_2699,N_2786);
or UO_180 (O_180,N_2505,N_2545);
nand UO_181 (O_181,N_2830,N_2957);
and UO_182 (O_182,N_2836,N_2705);
or UO_183 (O_183,N_2590,N_2617);
nor UO_184 (O_184,N_2665,N_2507);
nand UO_185 (O_185,N_2976,N_2807);
or UO_186 (O_186,N_2766,N_2993);
nand UO_187 (O_187,N_2596,N_2921);
and UO_188 (O_188,N_2902,N_2804);
or UO_189 (O_189,N_2579,N_2828);
and UO_190 (O_190,N_2893,N_2636);
or UO_191 (O_191,N_2941,N_2874);
nor UO_192 (O_192,N_2653,N_2549);
nand UO_193 (O_193,N_2802,N_2862);
and UO_194 (O_194,N_2806,N_2823);
nand UO_195 (O_195,N_2739,N_2922);
or UO_196 (O_196,N_2771,N_2582);
nor UO_197 (O_197,N_2931,N_2967);
nand UO_198 (O_198,N_2595,N_2753);
and UO_199 (O_199,N_2940,N_2625);
or UO_200 (O_200,N_2711,N_2561);
and UO_201 (O_201,N_2566,N_2841);
nand UO_202 (O_202,N_2821,N_2559);
and UO_203 (O_203,N_2977,N_2659);
or UO_204 (O_204,N_2613,N_2846);
or UO_205 (O_205,N_2944,N_2999);
nor UO_206 (O_206,N_2777,N_2925);
and UO_207 (O_207,N_2904,N_2961);
or UO_208 (O_208,N_2740,N_2602);
or UO_209 (O_209,N_2709,N_2787);
nor UO_210 (O_210,N_2985,N_2907);
nor UO_211 (O_211,N_2580,N_2520);
nand UO_212 (O_212,N_2592,N_2767);
and UO_213 (O_213,N_2795,N_2719);
nand UO_214 (O_214,N_2585,N_2848);
and UO_215 (O_215,N_2661,N_2668);
nor UO_216 (O_216,N_2757,N_2697);
or UO_217 (O_217,N_2799,N_2708);
and UO_218 (O_218,N_2987,N_2535);
nor UO_219 (O_219,N_2618,N_2906);
nand UO_220 (O_220,N_2995,N_2721);
nor UO_221 (O_221,N_2534,N_2539);
nand UO_222 (O_222,N_2537,N_2784);
or UO_223 (O_223,N_2800,N_2774);
or UO_224 (O_224,N_2527,N_2892);
or UO_225 (O_225,N_2745,N_2966);
nand UO_226 (O_226,N_2928,N_2516);
nand UO_227 (O_227,N_2654,N_2835);
nor UO_228 (O_228,N_2578,N_2651);
and UO_229 (O_229,N_2845,N_2614);
and UO_230 (O_230,N_2924,N_2969);
and UO_231 (O_231,N_2588,N_2888);
or UO_232 (O_232,N_2606,N_2552);
or UO_233 (O_233,N_2808,N_2536);
nor UO_234 (O_234,N_2849,N_2934);
xnor UO_235 (O_235,N_2913,N_2603);
or UO_236 (O_236,N_2644,N_2817);
or UO_237 (O_237,N_2929,N_2504);
nor UO_238 (O_238,N_2598,N_2564);
nor UO_239 (O_239,N_2763,N_2581);
or UO_240 (O_240,N_2650,N_2700);
and UO_241 (O_241,N_2860,N_2978);
nand UO_242 (O_242,N_2550,N_2779);
nand UO_243 (O_243,N_2965,N_2853);
and UO_244 (O_244,N_2586,N_2972);
nand UO_245 (O_245,N_2616,N_2620);
or UO_246 (O_246,N_2546,N_2726);
or UO_247 (O_247,N_2822,N_2710);
and UO_248 (O_248,N_2818,N_2942);
or UO_249 (O_249,N_2524,N_2968);
nor UO_250 (O_250,N_2600,N_2714);
and UO_251 (O_251,N_2508,N_2518);
nand UO_252 (O_252,N_2947,N_2834);
or UO_253 (O_253,N_2539,N_2891);
and UO_254 (O_254,N_2666,N_2736);
and UO_255 (O_255,N_2955,N_2964);
or UO_256 (O_256,N_2859,N_2987);
nand UO_257 (O_257,N_2545,N_2787);
and UO_258 (O_258,N_2725,N_2750);
or UO_259 (O_259,N_2608,N_2681);
nor UO_260 (O_260,N_2525,N_2821);
and UO_261 (O_261,N_2898,N_2674);
and UO_262 (O_262,N_2816,N_2598);
or UO_263 (O_263,N_2730,N_2556);
nor UO_264 (O_264,N_2938,N_2808);
and UO_265 (O_265,N_2791,N_2830);
and UO_266 (O_266,N_2947,N_2572);
nand UO_267 (O_267,N_2699,N_2834);
and UO_268 (O_268,N_2848,N_2651);
or UO_269 (O_269,N_2720,N_2873);
or UO_270 (O_270,N_2817,N_2917);
and UO_271 (O_271,N_2528,N_2865);
nand UO_272 (O_272,N_2572,N_2709);
nand UO_273 (O_273,N_2597,N_2653);
and UO_274 (O_274,N_2542,N_2649);
nand UO_275 (O_275,N_2906,N_2847);
or UO_276 (O_276,N_2752,N_2883);
and UO_277 (O_277,N_2676,N_2597);
nand UO_278 (O_278,N_2603,N_2632);
nand UO_279 (O_279,N_2500,N_2989);
or UO_280 (O_280,N_2673,N_2986);
and UO_281 (O_281,N_2794,N_2896);
and UO_282 (O_282,N_2756,N_2652);
nor UO_283 (O_283,N_2546,N_2571);
nand UO_284 (O_284,N_2912,N_2888);
and UO_285 (O_285,N_2817,N_2658);
or UO_286 (O_286,N_2964,N_2796);
nand UO_287 (O_287,N_2691,N_2603);
and UO_288 (O_288,N_2621,N_2651);
nand UO_289 (O_289,N_2988,N_2684);
nand UO_290 (O_290,N_2535,N_2995);
nand UO_291 (O_291,N_2629,N_2711);
nand UO_292 (O_292,N_2778,N_2647);
or UO_293 (O_293,N_2616,N_2570);
nand UO_294 (O_294,N_2778,N_2694);
or UO_295 (O_295,N_2603,N_2666);
nor UO_296 (O_296,N_2666,N_2694);
and UO_297 (O_297,N_2805,N_2897);
or UO_298 (O_298,N_2758,N_2663);
nor UO_299 (O_299,N_2988,N_2899);
and UO_300 (O_300,N_2868,N_2660);
nand UO_301 (O_301,N_2590,N_2975);
nand UO_302 (O_302,N_2938,N_2704);
nor UO_303 (O_303,N_2860,N_2812);
nand UO_304 (O_304,N_2727,N_2931);
nor UO_305 (O_305,N_2659,N_2957);
and UO_306 (O_306,N_2794,N_2874);
nand UO_307 (O_307,N_2920,N_2576);
or UO_308 (O_308,N_2854,N_2836);
or UO_309 (O_309,N_2886,N_2827);
nand UO_310 (O_310,N_2562,N_2576);
or UO_311 (O_311,N_2576,N_2522);
or UO_312 (O_312,N_2813,N_2796);
or UO_313 (O_313,N_2530,N_2985);
xnor UO_314 (O_314,N_2701,N_2945);
nand UO_315 (O_315,N_2840,N_2512);
nor UO_316 (O_316,N_2572,N_2784);
and UO_317 (O_317,N_2751,N_2834);
and UO_318 (O_318,N_2990,N_2863);
and UO_319 (O_319,N_2825,N_2820);
and UO_320 (O_320,N_2642,N_2889);
or UO_321 (O_321,N_2626,N_2904);
and UO_322 (O_322,N_2687,N_2554);
or UO_323 (O_323,N_2934,N_2988);
nor UO_324 (O_324,N_2745,N_2583);
nand UO_325 (O_325,N_2660,N_2596);
and UO_326 (O_326,N_2815,N_2710);
nor UO_327 (O_327,N_2804,N_2944);
nand UO_328 (O_328,N_2739,N_2808);
nand UO_329 (O_329,N_2724,N_2532);
or UO_330 (O_330,N_2614,N_2781);
nand UO_331 (O_331,N_2815,N_2603);
nand UO_332 (O_332,N_2694,N_2931);
nor UO_333 (O_333,N_2504,N_2551);
nor UO_334 (O_334,N_2999,N_2749);
nor UO_335 (O_335,N_2549,N_2606);
nor UO_336 (O_336,N_2964,N_2601);
and UO_337 (O_337,N_2621,N_2725);
nor UO_338 (O_338,N_2615,N_2838);
or UO_339 (O_339,N_2634,N_2672);
nand UO_340 (O_340,N_2706,N_2993);
nor UO_341 (O_341,N_2939,N_2890);
and UO_342 (O_342,N_2748,N_2505);
or UO_343 (O_343,N_2539,N_2904);
nor UO_344 (O_344,N_2950,N_2947);
nand UO_345 (O_345,N_2569,N_2702);
nand UO_346 (O_346,N_2586,N_2572);
and UO_347 (O_347,N_2723,N_2885);
nand UO_348 (O_348,N_2640,N_2664);
nand UO_349 (O_349,N_2851,N_2800);
nor UO_350 (O_350,N_2815,N_2514);
and UO_351 (O_351,N_2642,N_2883);
nor UO_352 (O_352,N_2823,N_2959);
and UO_353 (O_353,N_2959,N_2973);
or UO_354 (O_354,N_2550,N_2545);
nor UO_355 (O_355,N_2697,N_2835);
nand UO_356 (O_356,N_2633,N_2869);
xor UO_357 (O_357,N_2842,N_2623);
and UO_358 (O_358,N_2901,N_2953);
and UO_359 (O_359,N_2944,N_2595);
and UO_360 (O_360,N_2905,N_2555);
and UO_361 (O_361,N_2794,N_2574);
or UO_362 (O_362,N_2866,N_2730);
nor UO_363 (O_363,N_2633,N_2808);
or UO_364 (O_364,N_2883,N_2502);
nor UO_365 (O_365,N_2522,N_2721);
or UO_366 (O_366,N_2793,N_2968);
nor UO_367 (O_367,N_2977,N_2945);
and UO_368 (O_368,N_2901,N_2828);
nand UO_369 (O_369,N_2769,N_2942);
or UO_370 (O_370,N_2514,N_2540);
or UO_371 (O_371,N_2815,N_2927);
nand UO_372 (O_372,N_2676,N_2953);
and UO_373 (O_373,N_2892,N_2654);
nor UO_374 (O_374,N_2596,N_2987);
or UO_375 (O_375,N_2584,N_2900);
nor UO_376 (O_376,N_2971,N_2989);
nor UO_377 (O_377,N_2509,N_2724);
xor UO_378 (O_378,N_2626,N_2519);
nand UO_379 (O_379,N_2986,N_2637);
or UO_380 (O_380,N_2965,N_2810);
and UO_381 (O_381,N_2600,N_2817);
and UO_382 (O_382,N_2776,N_2740);
nor UO_383 (O_383,N_2711,N_2603);
and UO_384 (O_384,N_2939,N_2582);
and UO_385 (O_385,N_2942,N_2924);
and UO_386 (O_386,N_2604,N_2858);
and UO_387 (O_387,N_2595,N_2622);
nor UO_388 (O_388,N_2786,N_2777);
and UO_389 (O_389,N_2842,N_2927);
or UO_390 (O_390,N_2946,N_2604);
nor UO_391 (O_391,N_2901,N_2544);
nor UO_392 (O_392,N_2848,N_2963);
nor UO_393 (O_393,N_2993,N_2533);
nor UO_394 (O_394,N_2565,N_2814);
nand UO_395 (O_395,N_2868,N_2899);
nor UO_396 (O_396,N_2851,N_2764);
or UO_397 (O_397,N_2818,N_2707);
nor UO_398 (O_398,N_2747,N_2803);
nand UO_399 (O_399,N_2791,N_2567);
or UO_400 (O_400,N_2541,N_2721);
or UO_401 (O_401,N_2585,N_2713);
and UO_402 (O_402,N_2906,N_2596);
and UO_403 (O_403,N_2750,N_2635);
nor UO_404 (O_404,N_2621,N_2602);
nand UO_405 (O_405,N_2665,N_2842);
or UO_406 (O_406,N_2706,N_2787);
and UO_407 (O_407,N_2814,N_2800);
or UO_408 (O_408,N_2629,N_2909);
nand UO_409 (O_409,N_2920,N_2750);
and UO_410 (O_410,N_2897,N_2978);
or UO_411 (O_411,N_2690,N_2523);
nand UO_412 (O_412,N_2940,N_2788);
and UO_413 (O_413,N_2708,N_2979);
nor UO_414 (O_414,N_2882,N_2808);
nand UO_415 (O_415,N_2907,N_2698);
nand UO_416 (O_416,N_2540,N_2650);
and UO_417 (O_417,N_2552,N_2572);
nor UO_418 (O_418,N_2811,N_2910);
nor UO_419 (O_419,N_2753,N_2555);
or UO_420 (O_420,N_2961,N_2965);
and UO_421 (O_421,N_2697,N_2993);
nand UO_422 (O_422,N_2811,N_2684);
or UO_423 (O_423,N_2695,N_2843);
nor UO_424 (O_424,N_2737,N_2551);
nor UO_425 (O_425,N_2959,N_2521);
or UO_426 (O_426,N_2658,N_2771);
nor UO_427 (O_427,N_2689,N_2858);
nand UO_428 (O_428,N_2584,N_2833);
and UO_429 (O_429,N_2579,N_2799);
and UO_430 (O_430,N_2860,N_2641);
and UO_431 (O_431,N_2573,N_2556);
and UO_432 (O_432,N_2508,N_2643);
nand UO_433 (O_433,N_2985,N_2500);
nand UO_434 (O_434,N_2809,N_2703);
and UO_435 (O_435,N_2523,N_2995);
nand UO_436 (O_436,N_2767,N_2891);
or UO_437 (O_437,N_2890,N_2610);
nand UO_438 (O_438,N_2555,N_2848);
nand UO_439 (O_439,N_2889,N_2505);
nor UO_440 (O_440,N_2600,N_2665);
and UO_441 (O_441,N_2959,N_2966);
and UO_442 (O_442,N_2906,N_2857);
or UO_443 (O_443,N_2744,N_2933);
or UO_444 (O_444,N_2746,N_2919);
nand UO_445 (O_445,N_2612,N_2704);
or UO_446 (O_446,N_2903,N_2931);
nor UO_447 (O_447,N_2857,N_2592);
nand UO_448 (O_448,N_2861,N_2800);
and UO_449 (O_449,N_2658,N_2795);
nand UO_450 (O_450,N_2914,N_2712);
nand UO_451 (O_451,N_2847,N_2754);
or UO_452 (O_452,N_2536,N_2936);
or UO_453 (O_453,N_2899,N_2701);
nand UO_454 (O_454,N_2809,N_2782);
nor UO_455 (O_455,N_2622,N_2978);
nand UO_456 (O_456,N_2533,N_2932);
nor UO_457 (O_457,N_2978,N_2678);
nor UO_458 (O_458,N_2988,N_2619);
nand UO_459 (O_459,N_2955,N_2525);
or UO_460 (O_460,N_2855,N_2919);
nand UO_461 (O_461,N_2657,N_2849);
nor UO_462 (O_462,N_2917,N_2689);
or UO_463 (O_463,N_2998,N_2994);
and UO_464 (O_464,N_2589,N_2955);
and UO_465 (O_465,N_2958,N_2647);
nand UO_466 (O_466,N_2990,N_2769);
nand UO_467 (O_467,N_2532,N_2667);
or UO_468 (O_468,N_2568,N_2616);
nand UO_469 (O_469,N_2596,N_2951);
nand UO_470 (O_470,N_2907,N_2505);
nand UO_471 (O_471,N_2584,N_2762);
nor UO_472 (O_472,N_2691,N_2830);
nor UO_473 (O_473,N_2941,N_2592);
nor UO_474 (O_474,N_2798,N_2868);
nor UO_475 (O_475,N_2618,N_2898);
nor UO_476 (O_476,N_2673,N_2661);
nand UO_477 (O_477,N_2910,N_2772);
and UO_478 (O_478,N_2782,N_2653);
or UO_479 (O_479,N_2678,N_2766);
nor UO_480 (O_480,N_2683,N_2654);
and UO_481 (O_481,N_2916,N_2847);
or UO_482 (O_482,N_2739,N_2798);
and UO_483 (O_483,N_2741,N_2761);
nand UO_484 (O_484,N_2818,N_2577);
nand UO_485 (O_485,N_2759,N_2720);
or UO_486 (O_486,N_2658,N_2676);
nand UO_487 (O_487,N_2894,N_2844);
or UO_488 (O_488,N_2983,N_2775);
or UO_489 (O_489,N_2607,N_2642);
nand UO_490 (O_490,N_2781,N_2909);
and UO_491 (O_491,N_2749,N_2635);
and UO_492 (O_492,N_2811,N_2904);
xnor UO_493 (O_493,N_2541,N_2804);
and UO_494 (O_494,N_2764,N_2517);
nor UO_495 (O_495,N_2580,N_2783);
nand UO_496 (O_496,N_2698,N_2664);
and UO_497 (O_497,N_2730,N_2523);
or UO_498 (O_498,N_2503,N_2850);
nor UO_499 (O_499,N_2914,N_2738);
endmodule