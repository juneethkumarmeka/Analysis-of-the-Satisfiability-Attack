module basic_500_3000_500_30_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_227,In_288);
nand U1 (N_1,In_387,In_317);
nand U2 (N_2,In_302,In_70);
and U3 (N_3,In_419,In_282);
and U4 (N_4,In_161,In_328);
or U5 (N_5,In_254,In_231);
nand U6 (N_6,In_379,In_154);
nand U7 (N_7,In_285,In_475);
or U8 (N_8,In_408,In_239);
nand U9 (N_9,In_406,In_412);
or U10 (N_10,In_76,In_458);
nor U11 (N_11,In_382,In_436);
nand U12 (N_12,In_341,In_6);
nand U13 (N_13,In_293,In_314);
nor U14 (N_14,In_391,In_281);
nand U15 (N_15,In_264,In_85);
nor U16 (N_16,In_10,In_483);
nand U17 (N_17,In_35,In_452);
or U18 (N_18,In_273,In_93);
nor U19 (N_19,In_144,In_332);
nor U20 (N_20,In_389,In_4);
nor U21 (N_21,In_178,In_68);
and U22 (N_22,In_245,In_411);
or U23 (N_23,In_40,In_476);
nor U24 (N_24,In_43,In_467);
nor U25 (N_25,In_474,In_418);
or U26 (N_26,In_397,In_185);
or U27 (N_27,In_278,In_12);
or U28 (N_28,In_200,In_63);
or U29 (N_29,In_335,In_9);
or U30 (N_30,In_343,In_41);
and U31 (N_31,In_140,In_148);
nand U32 (N_32,In_420,In_191);
and U33 (N_33,In_102,In_289);
and U34 (N_34,In_143,In_162);
xnor U35 (N_35,In_109,In_434);
nand U36 (N_36,In_182,In_498);
and U37 (N_37,In_244,In_295);
and U38 (N_38,In_131,In_84);
and U39 (N_39,In_189,In_401);
xnor U40 (N_40,In_253,In_303);
nor U41 (N_41,In_318,In_426);
xor U42 (N_42,In_250,In_230);
nand U43 (N_43,In_168,In_356);
nor U44 (N_44,In_75,In_274);
xnor U45 (N_45,In_47,In_352);
nand U46 (N_46,In_67,In_79);
nand U47 (N_47,In_0,In_66);
nand U48 (N_48,In_380,In_181);
and U49 (N_49,In_369,In_284);
or U50 (N_50,In_374,In_243);
nand U51 (N_51,In_27,In_17);
and U52 (N_52,In_429,In_410);
or U53 (N_53,In_431,In_54);
xor U54 (N_54,In_271,In_370);
nand U55 (N_55,In_204,In_398);
nand U56 (N_56,In_486,In_351);
and U57 (N_57,In_188,In_394);
nand U58 (N_58,In_116,In_409);
nand U59 (N_59,In_252,In_355);
nand U60 (N_60,In_172,In_174);
xnor U61 (N_61,In_457,In_215);
xor U62 (N_62,In_350,In_173);
nand U63 (N_63,In_153,In_44);
nor U64 (N_64,In_122,In_320);
nand U65 (N_65,In_150,In_488);
nand U66 (N_66,In_163,In_312);
nor U67 (N_67,In_495,In_141);
nor U68 (N_68,In_92,In_390);
or U69 (N_69,In_91,In_404);
or U70 (N_70,In_211,In_497);
xor U71 (N_71,In_334,In_199);
nand U72 (N_72,In_269,In_489);
or U73 (N_73,In_459,In_177);
and U74 (N_74,In_158,In_145);
xor U75 (N_75,In_104,In_340);
nand U76 (N_76,In_18,In_449);
and U77 (N_77,In_11,In_265);
and U78 (N_78,In_78,In_106);
xor U79 (N_79,In_367,In_45);
and U80 (N_80,In_325,In_267);
or U81 (N_81,In_399,In_442);
nor U82 (N_82,In_258,In_219);
xor U83 (N_83,In_86,In_167);
nand U84 (N_84,In_16,In_236);
or U85 (N_85,In_415,In_324);
nor U86 (N_86,In_443,In_218);
or U87 (N_87,In_99,In_127);
nand U88 (N_88,In_151,In_448);
and U89 (N_89,In_377,In_105);
or U90 (N_90,In_111,In_201);
or U91 (N_91,In_330,In_220);
nand U92 (N_92,In_217,In_248);
xnor U93 (N_93,In_383,In_3);
or U94 (N_94,In_301,In_71);
nand U95 (N_95,In_89,In_19);
or U96 (N_96,In_465,In_364);
and U97 (N_97,In_451,In_316);
nand U98 (N_98,In_128,In_95);
nand U99 (N_99,In_88,In_49);
and U100 (N_100,N_39,N_75);
or U101 (N_101,In_171,N_48);
or U102 (N_102,In_428,N_69);
nor U103 (N_103,In_247,In_469);
xnor U104 (N_104,In_202,N_11);
nor U105 (N_105,N_15,In_31);
or U106 (N_106,In_292,In_493);
and U107 (N_107,In_462,In_494);
nor U108 (N_108,In_22,In_8);
nand U109 (N_109,In_195,In_242);
and U110 (N_110,In_338,In_26);
nand U111 (N_111,In_251,N_83);
nand U112 (N_112,In_138,In_107);
nor U113 (N_113,In_139,In_414);
nand U114 (N_114,In_132,In_296);
nor U115 (N_115,In_56,In_310);
or U116 (N_116,N_37,In_405);
nand U117 (N_117,N_61,In_179);
xnor U118 (N_118,In_36,In_372);
xnor U119 (N_119,N_23,In_87);
nand U120 (N_120,In_280,In_490);
and U121 (N_121,In_433,In_413);
nand U122 (N_122,In_214,In_37);
nand U123 (N_123,N_85,N_96);
or U124 (N_124,In_226,In_129);
nand U125 (N_125,In_55,N_20);
or U126 (N_126,In_463,In_363);
nor U127 (N_127,In_297,In_479);
nand U128 (N_128,In_357,N_82);
or U129 (N_129,In_376,In_42);
nand U130 (N_130,In_20,In_427);
xnor U131 (N_131,In_206,In_275);
nand U132 (N_132,In_50,In_216);
nand U133 (N_133,In_208,In_445);
xor U134 (N_134,In_72,In_361);
and U135 (N_135,In_237,In_435);
and U136 (N_136,In_64,N_57);
nor U137 (N_137,In_198,In_329);
nor U138 (N_138,In_194,In_80);
xor U139 (N_139,N_92,N_51);
nor U140 (N_140,In_395,In_120);
and U141 (N_141,In_203,In_183);
nand U142 (N_142,In_306,In_94);
or U143 (N_143,N_58,In_403);
nor U144 (N_144,In_438,N_7);
and U145 (N_145,In_101,In_126);
nand U146 (N_146,In_470,In_437);
nor U147 (N_147,In_155,In_260);
nand U148 (N_148,In_59,In_473);
or U149 (N_149,In_117,In_118);
or U150 (N_150,N_98,In_491);
or U151 (N_151,In_15,In_1);
or U152 (N_152,In_464,N_81);
and U153 (N_153,In_147,In_108);
and U154 (N_154,In_366,In_441);
or U155 (N_155,In_146,In_2);
nor U156 (N_156,In_480,In_98);
nand U157 (N_157,In_279,N_68);
and U158 (N_158,In_133,In_222);
nor U159 (N_159,In_453,N_18);
and U160 (N_160,In_57,N_19);
or U161 (N_161,In_400,N_26);
xnor U162 (N_162,N_66,In_190);
nand U163 (N_163,In_307,In_160);
and U164 (N_164,In_196,In_234);
or U165 (N_165,In_184,In_136);
nand U166 (N_166,In_384,In_23);
nor U167 (N_167,In_205,In_209);
xor U168 (N_168,N_31,N_74);
xor U169 (N_169,N_53,N_73);
and U170 (N_170,N_3,In_299);
or U171 (N_171,In_378,N_50);
xnor U172 (N_172,In_112,N_71);
and U173 (N_173,In_322,In_485);
nor U174 (N_174,In_487,In_38);
nand U175 (N_175,In_455,In_197);
or U176 (N_176,N_62,In_450);
and U177 (N_177,In_142,In_347);
and U178 (N_178,N_29,N_87);
nand U179 (N_179,In_353,In_333);
and U180 (N_180,In_482,In_32);
or U181 (N_181,N_80,In_33);
nor U182 (N_182,In_61,In_373);
nand U183 (N_183,In_21,In_466);
or U184 (N_184,In_261,N_45);
or U185 (N_185,In_327,In_149);
xnor U186 (N_186,In_124,In_298);
nor U187 (N_187,In_375,N_97);
and U188 (N_188,N_42,In_348);
xor U189 (N_189,N_0,In_423);
nor U190 (N_190,In_152,In_477);
xnor U191 (N_191,In_283,N_94);
and U192 (N_192,N_12,In_51);
nand U193 (N_193,In_319,In_481);
nor U194 (N_194,In_439,In_305);
and U195 (N_195,In_342,In_263);
and U196 (N_196,In_424,In_321);
or U197 (N_197,In_225,In_125);
nand U198 (N_198,In_192,N_22);
nand U199 (N_199,In_461,N_78);
and U200 (N_200,N_171,N_28);
and U201 (N_201,N_137,N_138);
and U202 (N_202,In_157,N_161);
or U203 (N_203,In_58,In_268);
or U204 (N_204,N_167,In_193);
xor U205 (N_205,In_7,N_179);
nand U206 (N_206,In_468,In_444);
xnor U207 (N_207,N_123,In_331);
nand U208 (N_208,N_155,In_416);
nand U209 (N_209,N_139,N_115);
nor U210 (N_210,N_157,N_84);
xnor U211 (N_211,N_165,N_111);
or U212 (N_212,N_63,N_191);
or U213 (N_213,In_393,In_187);
and U214 (N_214,N_76,N_33);
nor U215 (N_215,In_5,In_421);
and U216 (N_216,In_121,N_177);
nand U217 (N_217,In_287,N_89);
xnor U218 (N_218,In_48,In_381);
xor U219 (N_219,In_270,N_113);
xnor U220 (N_220,In_235,In_100);
xor U221 (N_221,N_106,In_169);
or U222 (N_222,In_300,N_35);
or U223 (N_223,N_112,In_53);
xor U224 (N_224,N_178,In_336);
and U225 (N_225,N_166,In_304);
nand U226 (N_226,In_447,In_210);
nor U227 (N_227,N_194,In_308);
xnor U228 (N_228,In_240,N_176);
nor U229 (N_229,In_326,N_55);
nor U230 (N_230,N_143,In_103);
nand U231 (N_231,In_432,N_70);
xnor U232 (N_232,In_176,N_175);
and U233 (N_233,N_180,In_484);
nor U234 (N_234,In_256,N_192);
xor U235 (N_235,In_170,In_337);
nand U236 (N_236,In_460,In_186);
xor U237 (N_237,N_56,In_25);
xnor U238 (N_238,In_119,N_126);
nor U239 (N_239,N_118,In_266);
or U240 (N_240,N_150,In_262);
xor U241 (N_241,In_496,N_135);
nand U242 (N_242,In_456,N_41);
nand U243 (N_243,N_93,N_117);
or U244 (N_244,In_478,In_135);
xnor U245 (N_245,N_122,In_96);
nand U246 (N_246,In_472,N_181);
or U247 (N_247,In_30,N_145);
nor U248 (N_248,In_315,N_114);
or U249 (N_249,N_148,In_29);
nand U250 (N_250,N_64,N_1);
nor U251 (N_251,In_46,In_24);
or U252 (N_252,In_229,In_123);
nor U253 (N_253,In_471,N_65);
xnor U254 (N_254,In_83,N_59);
and U255 (N_255,N_173,N_125);
nor U256 (N_256,N_134,N_199);
nor U257 (N_257,In_39,In_407);
nand U258 (N_258,N_27,N_189);
nand U259 (N_259,N_103,N_49);
and U260 (N_260,In_349,In_224);
nand U261 (N_261,N_116,N_152);
and U262 (N_262,N_174,N_140);
nor U263 (N_263,In_228,In_14);
and U264 (N_264,N_153,N_119);
nor U265 (N_265,N_154,N_13);
nor U266 (N_266,N_34,In_417);
and U267 (N_267,In_392,In_346);
and U268 (N_268,In_388,In_354);
or U269 (N_269,In_74,N_130);
nor U270 (N_270,N_5,In_81);
nor U271 (N_271,N_185,N_162);
nand U272 (N_272,In_277,N_133);
nand U273 (N_273,In_232,N_44);
nor U274 (N_274,In_77,In_60);
or U275 (N_275,In_82,In_402);
xnor U276 (N_276,N_186,N_43);
and U277 (N_277,In_255,N_38);
nand U278 (N_278,In_156,N_110);
and U279 (N_279,N_88,N_188);
nor U280 (N_280,In_238,N_77);
and U281 (N_281,In_276,N_91);
xor U282 (N_282,In_241,In_257);
and U283 (N_283,N_159,In_52);
nor U284 (N_284,N_100,In_115);
nor U285 (N_285,In_164,N_101);
nor U286 (N_286,N_169,In_113);
and U287 (N_287,In_290,N_46);
nand U288 (N_288,N_30,In_362);
and U289 (N_289,N_149,N_156);
or U290 (N_290,N_86,N_24);
nand U291 (N_291,N_54,N_6);
xor U292 (N_292,In_440,N_32);
or U293 (N_293,In_359,N_136);
xnor U294 (N_294,N_109,In_358);
or U295 (N_295,In_365,In_213);
xnor U296 (N_296,In_175,In_249);
or U297 (N_297,N_170,In_212);
and U298 (N_298,N_163,In_386);
and U299 (N_299,In_309,In_34);
xnor U300 (N_300,In_499,N_9);
and U301 (N_301,In_294,In_286);
and U302 (N_302,In_385,N_21);
nor U303 (N_303,N_265,N_240);
or U304 (N_304,N_259,N_221);
nor U305 (N_305,N_235,In_166);
nand U306 (N_306,N_284,N_231);
nand U307 (N_307,N_209,N_296);
or U308 (N_308,N_60,In_492);
and U309 (N_309,N_280,N_232);
nand U310 (N_310,In_137,In_114);
and U311 (N_311,N_246,In_207);
and U312 (N_312,N_214,N_252);
nor U313 (N_313,N_187,N_40);
xnor U314 (N_314,In_313,In_259);
nor U315 (N_315,N_146,N_295);
and U316 (N_316,N_241,N_297);
and U317 (N_317,N_213,N_274);
or U318 (N_318,N_285,N_105);
and U319 (N_319,In_272,N_142);
and U320 (N_320,N_218,N_8);
or U321 (N_321,N_144,In_344);
xnor U322 (N_322,N_128,N_190);
or U323 (N_323,N_263,N_2);
nand U324 (N_324,N_104,N_129);
nor U325 (N_325,N_283,In_97);
and U326 (N_326,In_345,N_196);
nand U327 (N_327,In_323,N_262);
nor U328 (N_328,N_10,N_248);
nand U329 (N_329,In_69,N_256);
nor U330 (N_330,N_36,N_212);
and U331 (N_331,N_224,N_230);
nand U332 (N_332,N_127,N_16);
or U333 (N_333,N_108,N_238);
nor U334 (N_334,N_184,N_267);
nand U335 (N_335,N_233,N_251);
xnor U336 (N_336,In_360,N_299);
nor U337 (N_337,N_239,N_247);
or U338 (N_338,N_286,N_271);
nand U339 (N_339,N_226,N_195);
or U340 (N_340,N_216,N_273);
nor U341 (N_341,N_183,N_225);
or U342 (N_342,N_206,N_253);
and U343 (N_343,N_107,N_260);
nand U344 (N_344,In_90,N_287);
nor U345 (N_345,N_282,N_25);
nor U346 (N_346,N_298,N_268);
nor U347 (N_347,N_215,N_14);
or U348 (N_348,N_281,N_168);
nor U349 (N_349,N_264,N_227);
xnor U350 (N_350,N_229,N_269);
xor U351 (N_351,N_52,N_121);
nand U352 (N_352,N_254,N_270);
and U353 (N_353,In_430,N_131);
and U354 (N_354,N_160,In_246);
xor U355 (N_355,N_291,N_234);
and U356 (N_356,N_292,N_289);
nor U357 (N_357,In_396,N_200);
xnor U358 (N_358,N_147,N_204);
nor U359 (N_359,N_197,N_210);
or U360 (N_360,N_237,N_205);
or U361 (N_361,N_249,N_250);
nor U362 (N_362,N_72,In_368);
or U363 (N_363,In_221,N_67);
or U364 (N_364,N_47,In_446);
and U365 (N_365,N_79,In_180);
nand U366 (N_366,N_294,N_277);
nor U367 (N_367,N_293,N_228);
or U368 (N_368,In_311,N_151);
nor U369 (N_369,N_258,N_95);
nand U370 (N_370,N_244,N_290);
and U371 (N_371,N_198,N_261);
nor U372 (N_372,In_13,N_202);
nand U373 (N_373,N_245,N_164);
or U374 (N_374,N_203,N_217);
nand U375 (N_375,N_207,N_211);
nor U376 (N_376,N_172,In_223);
nand U377 (N_377,N_255,N_266);
nor U378 (N_378,N_193,N_288);
xor U379 (N_379,N_102,In_425);
nor U380 (N_380,In_165,In_28);
or U381 (N_381,N_132,In_62);
nor U382 (N_382,N_219,N_242);
and U383 (N_383,In_454,N_275);
nand U384 (N_384,N_120,In_130);
or U385 (N_385,N_223,In_291);
nor U386 (N_386,In_73,N_201);
nand U387 (N_387,In_371,In_339);
and U388 (N_388,N_182,N_257);
or U389 (N_389,N_272,N_236);
or U390 (N_390,N_17,N_276);
and U391 (N_391,N_124,In_134);
nor U392 (N_392,In_65,N_243);
or U393 (N_393,N_141,In_110);
nor U394 (N_394,N_208,N_90);
or U395 (N_395,In_422,In_159);
and U396 (N_396,N_158,In_233);
or U397 (N_397,N_278,N_99);
or U398 (N_398,N_4,N_220);
nand U399 (N_399,N_222,N_279);
nor U400 (N_400,N_308,N_350);
and U401 (N_401,N_364,N_322);
nand U402 (N_402,N_368,N_343);
xor U403 (N_403,N_396,N_359);
nand U404 (N_404,N_319,N_315);
or U405 (N_405,N_313,N_326);
or U406 (N_406,N_339,N_345);
and U407 (N_407,N_321,N_344);
nand U408 (N_408,N_328,N_318);
nor U409 (N_409,N_306,N_391);
or U410 (N_410,N_395,N_361);
nand U411 (N_411,N_314,N_370);
nor U412 (N_412,N_378,N_338);
nor U413 (N_413,N_300,N_332);
nand U414 (N_414,N_336,N_385);
and U415 (N_415,N_355,N_360);
or U416 (N_416,N_354,N_374);
nor U417 (N_417,N_312,N_311);
nor U418 (N_418,N_329,N_358);
and U419 (N_419,N_324,N_399);
nand U420 (N_420,N_335,N_356);
xor U421 (N_421,N_301,N_390);
or U422 (N_422,N_352,N_382);
or U423 (N_423,N_383,N_353);
and U424 (N_424,N_310,N_376);
nand U425 (N_425,N_375,N_317);
nor U426 (N_426,N_365,N_386);
nand U427 (N_427,N_346,N_337);
or U428 (N_428,N_340,N_398);
and U429 (N_429,N_362,N_381);
nor U430 (N_430,N_397,N_347);
nor U431 (N_431,N_357,N_351);
or U432 (N_432,N_342,N_325);
and U433 (N_433,N_348,N_333);
xnor U434 (N_434,N_303,N_330);
nor U435 (N_435,N_371,N_389);
or U436 (N_436,N_373,N_393);
nor U437 (N_437,N_394,N_349);
nor U438 (N_438,N_384,N_302);
or U439 (N_439,N_392,N_341);
or U440 (N_440,N_380,N_307);
nand U441 (N_441,N_327,N_334);
and U442 (N_442,N_304,N_323);
nor U443 (N_443,N_320,N_309);
or U444 (N_444,N_305,N_379);
and U445 (N_445,N_387,N_366);
and U446 (N_446,N_316,N_377);
and U447 (N_447,N_369,N_331);
nand U448 (N_448,N_367,N_363);
nor U449 (N_449,N_388,N_372);
nand U450 (N_450,N_349,N_304);
and U451 (N_451,N_344,N_347);
nand U452 (N_452,N_309,N_385);
or U453 (N_453,N_300,N_353);
nor U454 (N_454,N_302,N_393);
or U455 (N_455,N_342,N_397);
nor U456 (N_456,N_305,N_383);
and U457 (N_457,N_389,N_344);
or U458 (N_458,N_336,N_377);
xor U459 (N_459,N_384,N_392);
nand U460 (N_460,N_397,N_329);
nand U461 (N_461,N_372,N_383);
nor U462 (N_462,N_378,N_315);
nor U463 (N_463,N_321,N_329);
or U464 (N_464,N_350,N_338);
and U465 (N_465,N_324,N_312);
or U466 (N_466,N_306,N_368);
xor U467 (N_467,N_347,N_384);
or U468 (N_468,N_321,N_312);
nand U469 (N_469,N_301,N_311);
and U470 (N_470,N_347,N_398);
and U471 (N_471,N_385,N_325);
nand U472 (N_472,N_375,N_329);
or U473 (N_473,N_376,N_305);
and U474 (N_474,N_328,N_320);
nand U475 (N_475,N_322,N_317);
or U476 (N_476,N_384,N_307);
nand U477 (N_477,N_349,N_369);
nand U478 (N_478,N_300,N_325);
or U479 (N_479,N_363,N_364);
and U480 (N_480,N_393,N_381);
and U481 (N_481,N_361,N_379);
or U482 (N_482,N_388,N_382);
nand U483 (N_483,N_326,N_345);
nor U484 (N_484,N_347,N_368);
nor U485 (N_485,N_373,N_339);
nor U486 (N_486,N_372,N_308);
or U487 (N_487,N_386,N_356);
nor U488 (N_488,N_376,N_341);
nor U489 (N_489,N_325,N_364);
nor U490 (N_490,N_326,N_384);
nor U491 (N_491,N_347,N_355);
nand U492 (N_492,N_349,N_372);
and U493 (N_493,N_319,N_392);
and U494 (N_494,N_395,N_359);
and U495 (N_495,N_303,N_304);
and U496 (N_496,N_307,N_360);
nand U497 (N_497,N_392,N_305);
nand U498 (N_498,N_386,N_395);
xnor U499 (N_499,N_358,N_383);
and U500 (N_500,N_440,N_421);
or U501 (N_501,N_449,N_447);
nor U502 (N_502,N_487,N_419);
or U503 (N_503,N_460,N_415);
nand U504 (N_504,N_491,N_438);
and U505 (N_505,N_401,N_418);
and U506 (N_506,N_467,N_482);
or U507 (N_507,N_479,N_422);
and U508 (N_508,N_426,N_472);
nand U509 (N_509,N_427,N_442);
and U510 (N_510,N_490,N_425);
or U511 (N_511,N_474,N_454);
or U512 (N_512,N_402,N_469);
nand U513 (N_513,N_408,N_478);
or U514 (N_514,N_455,N_448);
or U515 (N_515,N_488,N_473);
and U516 (N_516,N_461,N_452);
nor U517 (N_517,N_429,N_471);
xnor U518 (N_518,N_434,N_497);
nand U519 (N_519,N_458,N_468);
and U520 (N_520,N_420,N_405);
or U521 (N_521,N_494,N_499);
or U522 (N_522,N_485,N_476);
or U523 (N_523,N_495,N_466);
nand U524 (N_524,N_465,N_430);
nor U525 (N_525,N_498,N_481);
nor U526 (N_526,N_456,N_496);
xnor U527 (N_527,N_489,N_424);
nor U528 (N_528,N_428,N_444);
nand U529 (N_529,N_431,N_470);
and U530 (N_530,N_411,N_450);
nor U531 (N_531,N_493,N_423);
xor U532 (N_532,N_483,N_404);
xor U533 (N_533,N_486,N_441);
nand U534 (N_534,N_451,N_492);
and U535 (N_535,N_453,N_417);
nor U536 (N_536,N_412,N_435);
xor U537 (N_537,N_410,N_436);
nor U538 (N_538,N_459,N_484);
or U539 (N_539,N_439,N_480);
xor U540 (N_540,N_437,N_403);
nor U541 (N_541,N_409,N_446);
nand U542 (N_542,N_416,N_413);
or U543 (N_543,N_463,N_462);
and U544 (N_544,N_464,N_445);
nor U545 (N_545,N_443,N_407);
nand U546 (N_546,N_477,N_433);
and U547 (N_547,N_406,N_457);
xor U548 (N_548,N_432,N_414);
nand U549 (N_549,N_400,N_475);
xor U550 (N_550,N_460,N_448);
xor U551 (N_551,N_478,N_495);
nor U552 (N_552,N_448,N_435);
nand U553 (N_553,N_443,N_451);
and U554 (N_554,N_420,N_423);
nand U555 (N_555,N_405,N_431);
nand U556 (N_556,N_432,N_455);
nor U557 (N_557,N_421,N_456);
or U558 (N_558,N_472,N_452);
and U559 (N_559,N_440,N_484);
nor U560 (N_560,N_403,N_499);
xor U561 (N_561,N_457,N_436);
nor U562 (N_562,N_453,N_466);
nor U563 (N_563,N_451,N_415);
nor U564 (N_564,N_447,N_417);
xnor U565 (N_565,N_453,N_487);
and U566 (N_566,N_467,N_401);
nor U567 (N_567,N_408,N_430);
or U568 (N_568,N_424,N_446);
and U569 (N_569,N_489,N_453);
or U570 (N_570,N_417,N_408);
and U571 (N_571,N_433,N_466);
nor U572 (N_572,N_436,N_447);
or U573 (N_573,N_462,N_400);
nor U574 (N_574,N_407,N_401);
nand U575 (N_575,N_419,N_408);
xor U576 (N_576,N_489,N_434);
nand U577 (N_577,N_436,N_439);
nand U578 (N_578,N_476,N_431);
nand U579 (N_579,N_419,N_409);
nand U580 (N_580,N_425,N_488);
and U581 (N_581,N_410,N_495);
nand U582 (N_582,N_456,N_499);
nand U583 (N_583,N_432,N_451);
and U584 (N_584,N_439,N_400);
nand U585 (N_585,N_435,N_463);
nor U586 (N_586,N_418,N_422);
nor U587 (N_587,N_402,N_414);
nand U588 (N_588,N_439,N_458);
and U589 (N_589,N_465,N_426);
nor U590 (N_590,N_433,N_413);
or U591 (N_591,N_471,N_435);
and U592 (N_592,N_428,N_437);
or U593 (N_593,N_414,N_428);
or U594 (N_594,N_442,N_484);
nor U595 (N_595,N_475,N_482);
nor U596 (N_596,N_425,N_456);
nor U597 (N_597,N_429,N_482);
nand U598 (N_598,N_464,N_400);
nand U599 (N_599,N_446,N_494);
or U600 (N_600,N_584,N_513);
and U601 (N_601,N_539,N_535);
or U602 (N_602,N_547,N_598);
nor U603 (N_603,N_529,N_596);
or U604 (N_604,N_577,N_533);
or U605 (N_605,N_579,N_543);
xor U606 (N_606,N_521,N_595);
and U607 (N_607,N_585,N_545);
nand U608 (N_608,N_518,N_553);
nor U609 (N_609,N_567,N_537);
xor U610 (N_610,N_532,N_519);
xor U611 (N_611,N_597,N_527);
nand U612 (N_612,N_528,N_504);
xor U613 (N_613,N_560,N_536);
xnor U614 (N_614,N_572,N_549);
nor U615 (N_615,N_542,N_509);
and U616 (N_616,N_599,N_505);
nor U617 (N_617,N_561,N_557);
and U618 (N_618,N_569,N_586);
and U619 (N_619,N_524,N_566);
xor U620 (N_620,N_574,N_588);
nor U621 (N_621,N_501,N_568);
xor U622 (N_622,N_573,N_514);
and U623 (N_623,N_523,N_548);
and U624 (N_624,N_525,N_530);
xor U625 (N_625,N_503,N_551);
and U626 (N_626,N_531,N_565);
nor U627 (N_627,N_555,N_550);
and U628 (N_628,N_590,N_500);
nor U629 (N_629,N_512,N_582);
nor U630 (N_630,N_517,N_559);
nor U631 (N_631,N_575,N_516);
nor U632 (N_632,N_578,N_563);
xor U633 (N_633,N_538,N_592);
nand U634 (N_634,N_508,N_507);
or U635 (N_635,N_581,N_540);
or U636 (N_636,N_583,N_526);
xor U637 (N_637,N_554,N_546);
and U638 (N_638,N_544,N_580);
nor U639 (N_639,N_564,N_589);
nand U640 (N_640,N_576,N_570);
or U641 (N_641,N_591,N_534);
and U642 (N_642,N_522,N_587);
nand U643 (N_643,N_510,N_511);
nand U644 (N_644,N_520,N_556);
or U645 (N_645,N_558,N_552);
nor U646 (N_646,N_571,N_562);
and U647 (N_647,N_594,N_515);
or U648 (N_648,N_593,N_506);
nand U649 (N_649,N_541,N_502);
or U650 (N_650,N_567,N_528);
xor U651 (N_651,N_525,N_520);
and U652 (N_652,N_573,N_533);
xor U653 (N_653,N_512,N_594);
nand U654 (N_654,N_593,N_524);
nand U655 (N_655,N_592,N_542);
xor U656 (N_656,N_592,N_590);
or U657 (N_657,N_500,N_525);
nor U658 (N_658,N_536,N_565);
nor U659 (N_659,N_508,N_556);
nand U660 (N_660,N_589,N_510);
nand U661 (N_661,N_535,N_529);
or U662 (N_662,N_501,N_583);
nor U663 (N_663,N_513,N_561);
xor U664 (N_664,N_574,N_521);
and U665 (N_665,N_556,N_511);
and U666 (N_666,N_569,N_547);
or U667 (N_667,N_578,N_535);
and U668 (N_668,N_576,N_531);
or U669 (N_669,N_531,N_549);
or U670 (N_670,N_583,N_588);
xor U671 (N_671,N_525,N_532);
nand U672 (N_672,N_593,N_530);
and U673 (N_673,N_518,N_547);
and U674 (N_674,N_563,N_589);
nand U675 (N_675,N_542,N_518);
or U676 (N_676,N_550,N_557);
nor U677 (N_677,N_594,N_520);
or U678 (N_678,N_525,N_526);
nand U679 (N_679,N_560,N_521);
and U680 (N_680,N_504,N_583);
or U681 (N_681,N_531,N_550);
and U682 (N_682,N_550,N_590);
nand U683 (N_683,N_500,N_598);
and U684 (N_684,N_540,N_514);
nor U685 (N_685,N_589,N_565);
nand U686 (N_686,N_525,N_597);
nor U687 (N_687,N_564,N_508);
nor U688 (N_688,N_524,N_532);
or U689 (N_689,N_544,N_530);
nand U690 (N_690,N_529,N_560);
and U691 (N_691,N_553,N_596);
or U692 (N_692,N_503,N_539);
nand U693 (N_693,N_596,N_570);
and U694 (N_694,N_525,N_513);
and U695 (N_695,N_564,N_538);
and U696 (N_696,N_507,N_575);
or U697 (N_697,N_546,N_577);
and U698 (N_698,N_501,N_527);
and U699 (N_699,N_560,N_558);
nand U700 (N_700,N_655,N_609);
nor U701 (N_701,N_615,N_683);
xnor U702 (N_702,N_633,N_664);
and U703 (N_703,N_602,N_674);
nor U704 (N_704,N_624,N_698);
or U705 (N_705,N_623,N_662);
or U706 (N_706,N_616,N_657);
and U707 (N_707,N_671,N_600);
nand U708 (N_708,N_634,N_647);
xor U709 (N_709,N_693,N_682);
or U710 (N_710,N_640,N_601);
nor U711 (N_711,N_644,N_638);
or U712 (N_712,N_653,N_686);
and U713 (N_713,N_688,N_617);
nor U714 (N_714,N_668,N_670);
nor U715 (N_715,N_630,N_656);
and U716 (N_716,N_680,N_677);
or U717 (N_717,N_666,N_676);
or U718 (N_718,N_611,N_635);
nand U719 (N_719,N_607,N_672);
or U720 (N_720,N_694,N_675);
nor U721 (N_721,N_667,N_603);
nand U722 (N_722,N_649,N_663);
or U723 (N_723,N_641,N_687);
and U724 (N_724,N_637,N_643);
xor U725 (N_725,N_625,N_695);
or U726 (N_726,N_678,N_652);
xnor U727 (N_727,N_669,N_689);
or U728 (N_728,N_650,N_604);
nand U729 (N_729,N_626,N_605);
nand U730 (N_730,N_692,N_679);
nand U731 (N_731,N_651,N_632);
and U732 (N_732,N_654,N_629);
nand U733 (N_733,N_620,N_681);
nand U734 (N_734,N_665,N_646);
nor U735 (N_735,N_613,N_685);
nand U736 (N_736,N_661,N_610);
or U737 (N_737,N_673,N_639);
and U738 (N_738,N_696,N_627);
nor U739 (N_739,N_645,N_606);
nor U740 (N_740,N_660,N_658);
or U741 (N_741,N_648,N_622);
and U742 (N_742,N_636,N_614);
nor U743 (N_743,N_628,N_690);
nand U744 (N_744,N_619,N_618);
nand U745 (N_745,N_697,N_612);
or U746 (N_746,N_691,N_659);
nand U747 (N_747,N_621,N_684);
nor U748 (N_748,N_608,N_642);
nor U749 (N_749,N_631,N_699);
nand U750 (N_750,N_644,N_673);
and U751 (N_751,N_697,N_692);
nor U752 (N_752,N_670,N_640);
or U753 (N_753,N_625,N_699);
nor U754 (N_754,N_680,N_629);
or U755 (N_755,N_665,N_648);
or U756 (N_756,N_615,N_666);
nand U757 (N_757,N_613,N_640);
xnor U758 (N_758,N_667,N_690);
nand U759 (N_759,N_648,N_608);
nor U760 (N_760,N_620,N_699);
nor U761 (N_761,N_646,N_615);
nor U762 (N_762,N_688,N_663);
and U763 (N_763,N_629,N_651);
and U764 (N_764,N_672,N_641);
nand U765 (N_765,N_697,N_627);
nor U766 (N_766,N_643,N_680);
xor U767 (N_767,N_662,N_605);
nand U768 (N_768,N_648,N_691);
nor U769 (N_769,N_658,N_681);
nor U770 (N_770,N_644,N_667);
and U771 (N_771,N_608,N_609);
nand U772 (N_772,N_638,N_620);
nor U773 (N_773,N_624,N_683);
and U774 (N_774,N_683,N_652);
or U775 (N_775,N_695,N_630);
and U776 (N_776,N_607,N_635);
and U777 (N_777,N_692,N_655);
or U778 (N_778,N_666,N_616);
or U779 (N_779,N_677,N_629);
and U780 (N_780,N_666,N_652);
nor U781 (N_781,N_612,N_683);
or U782 (N_782,N_653,N_641);
or U783 (N_783,N_666,N_669);
xor U784 (N_784,N_653,N_642);
or U785 (N_785,N_631,N_629);
or U786 (N_786,N_697,N_678);
nand U787 (N_787,N_613,N_633);
nand U788 (N_788,N_625,N_694);
xor U789 (N_789,N_648,N_641);
and U790 (N_790,N_688,N_675);
and U791 (N_791,N_626,N_642);
or U792 (N_792,N_659,N_652);
nor U793 (N_793,N_672,N_694);
and U794 (N_794,N_663,N_631);
or U795 (N_795,N_643,N_666);
nand U796 (N_796,N_684,N_603);
nor U797 (N_797,N_671,N_619);
and U798 (N_798,N_648,N_609);
and U799 (N_799,N_641,N_699);
or U800 (N_800,N_796,N_754);
nand U801 (N_801,N_744,N_745);
nor U802 (N_802,N_757,N_721);
xor U803 (N_803,N_789,N_761);
and U804 (N_804,N_788,N_722);
xor U805 (N_805,N_792,N_784);
and U806 (N_806,N_791,N_758);
nor U807 (N_807,N_783,N_785);
or U808 (N_808,N_762,N_768);
nand U809 (N_809,N_797,N_713);
or U810 (N_810,N_795,N_719);
and U811 (N_811,N_759,N_769);
or U812 (N_812,N_772,N_787);
nor U813 (N_813,N_782,N_732);
xor U814 (N_814,N_790,N_794);
or U815 (N_815,N_741,N_798);
and U816 (N_816,N_776,N_771);
nand U817 (N_817,N_710,N_726);
or U818 (N_818,N_730,N_767);
nand U819 (N_819,N_786,N_764);
nor U820 (N_820,N_712,N_755);
nor U821 (N_821,N_748,N_766);
nor U822 (N_822,N_773,N_704);
and U823 (N_823,N_746,N_747);
or U824 (N_824,N_735,N_715);
or U825 (N_825,N_717,N_777);
nor U826 (N_826,N_774,N_750);
nand U827 (N_827,N_793,N_749);
nand U828 (N_828,N_725,N_753);
or U829 (N_829,N_763,N_703);
nand U830 (N_830,N_765,N_724);
nor U831 (N_831,N_702,N_728);
xor U832 (N_832,N_736,N_700);
and U833 (N_833,N_711,N_734);
xor U834 (N_834,N_729,N_760);
or U835 (N_835,N_723,N_707);
or U836 (N_836,N_737,N_701);
and U837 (N_837,N_752,N_756);
nor U838 (N_838,N_720,N_743);
xor U839 (N_839,N_727,N_714);
or U840 (N_840,N_716,N_751);
nand U841 (N_841,N_731,N_718);
nand U842 (N_842,N_708,N_778);
nor U843 (N_843,N_705,N_739);
xnor U844 (N_844,N_742,N_799);
and U845 (N_845,N_706,N_780);
or U846 (N_846,N_738,N_775);
and U847 (N_847,N_770,N_733);
nor U848 (N_848,N_779,N_709);
or U849 (N_849,N_740,N_781);
or U850 (N_850,N_785,N_753);
nor U851 (N_851,N_746,N_762);
xor U852 (N_852,N_769,N_754);
xor U853 (N_853,N_755,N_741);
and U854 (N_854,N_748,N_764);
and U855 (N_855,N_774,N_744);
nand U856 (N_856,N_734,N_705);
or U857 (N_857,N_749,N_775);
nand U858 (N_858,N_785,N_722);
nor U859 (N_859,N_723,N_779);
and U860 (N_860,N_732,N_746);
xnor U861 (N_861,N_742,N_790);
or U862 (N_862,N_701,N_709);
or U863 (N_863,N_720,N_734);
and U864 (N_864,N_728,N_783);
and U865 (N_865,N_708,N_701);
nand U866 (N_866,N_707,N_745);
or U867 (N_867,N_751,N_710);
xor U868 (N_868,N_712,N_760);
or U869 (N_869,N_740,N_744);
nor U870 (N_870,N_771,N_797);
nand U871 (N_871,N_761,N_754);
or U872 (N_872,N_739,N_708);
or U873 (N_873,N_767,N_788);
or U874 (N_874,N_724,N_701);
or U875 (N_875,N_724,N_745);
or U876 (N_876,N_728,N_765);
xnor U877 (N_877,N_760,N_705);
and U878 (N_878,N_711,N_770);
nor U879 (N_879,N_713,N_712);
xnor U880 (N_880,N_772,N_765);
xor U881 (N_881,N_713,N_724);
and U882 (N_882,N_732,N_786);
or U883 (N_883,N_788,N_716);
nor U884 (N_884,N_724,N_740);
nand U885 (N_885,N_750,N_798);
nor U886 (N_886,N_767,N_774);
and U887 (N_887,N_765,N_700);
nand U888 (N_888,N_743,N_729);
nor U889 (N_889,N_709,N_771);
nand U890 (N_890,N_715,N_703);
xnor U891 (N_891,N_728,N_768);
nand U892 (N_892,N_729,N_759);
nor U893 (N_893,N_747,N_789);
and U894 (N_894,N_733,N_791);
or U895 (N_895,N_784,N_738);
or U896 (N_896,N_744,N_749);
nand U897 (N_897,N_737,N_787);
nor U898 (N_898,N_761,N_783);
and U899 (N_899,N_790,N_740);
and U900 (N_900,N_809,N_873);
or U901 (N_901,N_870,N_813);
and U902 (N_902,N_899,N_865);
nor U903 (N_903,N_867,N_863);
nand U904 (N_904,N_830,N_857);
and U905 (N_905,N_835,N_883);
nand U906 (N_906,N_890,N_898);
nor U907 (N_907,N_892,N_810);
nor U908 (N_908,N_874,N_849);
nand U909 (N_909,N_827,N_822);
and U910 (N_910,N_882,N_819);
nand U911 (N_911,N_864,N_846);
nor U912 (N_912,N_842,N_887);
nand U913 (N_913,N_801,N_877);
or U914 (N_914,N_820,N_866);
and U915 (N_915,N_812,N_802);
nand U916 (N_916,N_800,N_847);
nand U917 (N_917,N_868,N_843);
nand U918 (N_918,N_897,N_854);
nor U919 (N_919,N_829,N_845);
and U920 (N_920,N_886,N_816);
and U921 (N_921,N_851,N_824);
nand U922 (N_922,N_831,N_855);
nand U923 (N_923,N_885,N_838);
and U924 (N_924,N_862,N_841);
or U925 (N_925,N_858,N_875);
nand U926 (N_926,N_837,N_821);
and U927 (N_927,N_869,N_814);
nor U928 (N_928,N_806,N_893);
and U929 (N_929,N_884,N_828);
or U930 (N_930,N_815,N_811);
nand U931 (N_931,N_894,N_836);
nand U932 (N_932,N_859,N_804);
and U933 (N_933,N_833,N_803);
nand U934 (N_934,N_844,N_876);
nor U935 (N_935,N_881,N_888);
nor U936 (N_936,N_861,N_896);
nor U937 (N_937,N_839,N_823);
nand U938 (N_938,N_860,N_808);
nor U939 (N_939,N_832,N_834);
nand U940 (N_940,N_856,N_878);
nor U941 (N_941,N_871,N_872);
and U942 (N_942,N_817,N_826);
xnor U943 (N_943,N_891,N_880);
and U944 (N_944,N_879,N_889);
nor U945 (N_945,N_807,N_818);
or U946 (N_946,N_852,N_850);
nor U947 (N_947,N_805,N_853);
or U948 (N_948,N_848,N_825);
or U949 (N_949,N_895,N_840);
nor U950 (N_950,N_829,N_855);
xor U951 (N_951,N_817,N_860);
or U952 (N_952,N_858,N_831);
or U953 (N_953,N_856,N_860);
and U954 (N_954,N_863,N_824);
xor U955 (N_955,N_815,N_861);
nor U956 (N_956,N_820,N_835);
and U957 (N_957,N_859,N_824);
and U958 (N_958,N_837,N_891);
xnor U959 (N_959,N_879,N_869);
nor U960 (N_960,N_892,N_814);
nand U961 (N_961,N_819,N_817);
or U962 (N_962,N_813,N_848);
xnor U963 (N_963,N_830,N_862);
nor U964 (N_964,N_882,N_875);
xor U965 (N_965,N_809,N_857);
nand U966 (N_966,N_869,N_873);
xor U967 (N_967,N_825,N_837);
and U968 (N_968,N_865,N_869);
xnor U969 (N_969,N_800,N_843);
xnor U970 (N_970,N_883,N_890);
and U971 (N_971,N_818,N_828);
and U972 (N_972,N_814,N_842);
nor U973 (N_973,N_803,N_862);
xor U974 (N_974,N_826,N_849);
and U975 (N_975,N_804,N_847);
and U976 (N_976,N_805,N_882);
nand U977 (N_977,N_839,N_859);
or U978 (N_978,N_851,N_822);
or U979 (N_979,N_884,N_800);
nand U980 (N_980,N_885,N_876);
nor U981 (N_981,N_885,N_877);
or U982 (N_982,N_893,N_890);
nand U983 (N_983,N_815,N_804);
nand U984 (N_984,N_874,N_801);
nand U985 (N_985,N_879,N_837);
nand U986 (N_986,N_880,N_801);
nand U987 (N_987,N_805,N_844);
and U988 (N_988,N_870,N_837);
nor U989 (N_989,N_827,N_844);
nor U990 (N_990,N_880,N_832);
nand U991 (N_991,N_897,N_894);
nand U992 (N_992,N_879,N_867);
nor U993 (N_993,N_803,N_876);
nor U994 (N_994,N_899,N_846);
and U995 (N_995,N_820,N_852);
nand U996 (N_996,N_882,N_845);
or U997 (N_997,N_854,N_805);
nor U998 (N_998,N_843,N_815);
nor U999 (N_999,N_876,N_802);
and U1000 (N_1000,N_959,N_979);
xor U1001 (N_1001,N_996,N_961);
and U1002 (N_1002,N_922,N_945);
nor U1003 (N_1003,N_918,N_925);
and U1004 (N_1004,N_970,N_929);
and U1005 (N_1005,N_964,N_900);
nor U1006 (N_1006,N_946,N_921);
nor U1007 (N_1007,N_980,N_937);
and U1008 (N_1008,N_948,N_906);
nand U1009 (N_1009,N_956,N_974);
nand U1010 (N_1010,N_963,N_997);
and U1011 (N_1011,N_966,N_901);
nor U1012 (N_1012,N_954,N_969);
and U1013 (N_1013,N_942,N_923);
nand U1014 (N_1014,N_953,N_935);
nor U1015 (N_1015,N_911,N_902);
and U1016 (N_1016,N_934,N_932);
nor U1017 (N_1017,N_943,N_951);
nand U1018 (N_1018,N_917,N_949);
and U1019 (N_1019,N_947,N_968);
nand U1020 (N_1020,N_965,N_988);
nand U1021 (N_1021,N_987,N_958);
nand U1022 (N_1022,N_940,N_989);
nand U1023 (N_1023,N_983,N_905);
xnor U1024 (N_1024,N_972,N_978);
and U1025 (N_1025,N_975,N_916);
nor U1026 (N_1026,N_971,N_941);
nand U1027 (N_1027,N_903,N_981);
or U1028 (N_1028,N_967,N_982);
or U1029 (N_1029,N_992,N_952);
nor U1030 (N_1030,N_994,N_936);
or U1031 (N_1031,N_924,N_912);
nand U1032 (N_1032,N_990,N_920);
nor U1033 (N_1033,N_909,N_985);
nor U1034 (N_1034,N_919,N_986);
or U1035 (N_1035,N_991,N_938);
or U1036 (N_1036,N_976,N_950);
and U1037 (N_1037,N_973,N_993);
or U1038 (N_1038,N_977,N_962);
and U1039 (N_1039,N_930,N_995);
nand U1040 (N_1040,N_914,N_944);
nor U1041 (N_1041,N_926,N_928);
or U1042 (N_1042,N_915,N_904);
nand U1043 (N_1043,N_931,N_955);
nand U1044 (N_1044,N_999,N_927);
nand U1045 (N_1045,N_910,N_933);
nand U1046 (N_1046,N_998,N_907);
nor U1047 (N_1047,N_957,N_984);
xor U1048 (N_1048,N_913,N_908);
and U1049 (N_1049,N_939,N_960);
xnor U1050 (N_1050,N_939,N_929);
or U1051 (N_1051,N_996,N_901);
or U1052 (N_1052,N_957,N_944);
nor U1053 (N_1053,N_926,N_999);
nor U1054 (N_1054,N_934,N_939);
or U1055 (N_1055,N_980,N_908);
or U1056 (N_1056,N_951,N_962);
nor U1057 (N_1057,N_996,N_999);
and U1058 (N_1058,N_945,N_912);
xnor U1059 (N_1059,N_992,N_953);
and U1060 (N_1060,N_985,N_943);
and U1061 (N_1061,N_905,N_993);
nor U1062 (N_1062,N_909,N_956);
xor U1063 (N_1063,N_946,N_933);
nor U1064 (N_1064,N_977,N_950);
and U1065 (N_1065,N_944,N_989);
xnor U1066 (N_1066,N_915,N_939);
and U1067 (N_1067,N_977,N_914);
nand U1068 (N_1068,N_934,N_970);
nand U1069 (N_1069,N_979,N_947);
nand U1070 (N_1070,N_901,N_964);
and U1071 (N_1071,N_974,N_975);
nor U1072 (N_1072,N_987,N_977);
and U1073 (N_1073,N_984,N_949);
and U1074 (N_1074,N_990,N_989);
nor U1075 (N_1075,N_907,N_914);
nand U1076 (N_1076,N_919,N_963);
and U1077 (N_1077,N_927,N_982);
xor U1078 (N_1078,N_930,N_924);
and U1079 (N_1079,N_932,N_992);
nand U1080 (N_1080,N_909,N_936);
and U1081 (N_1081,N_961,N_934);
or U1082 (N_1082,N_975,N_965);
xnor U1083 (N_1083,N_947,N_966);
and U1084 (N_1084,N_929,N_917);
nor U1085 (N_1085,N_926,N_948);
or U1086 (N_1086,N_988,N_968);
nand U1087 (N_1087,N_944,N_984);
or U1088 (N_1088,N_941,N_901);
nand U1089 (N_1089,N_951,N_965);
or U1090 (N_1090,N_926,N_914);
or U1091 (N_1091,N_910,N_913);
nand U1092 (N_1092,N_996,N_976);
or U1093 (N_1093,N_908,N_987);
and U1094 (N_1094,N_909,N_915);
and U1095 (N_1095,N_951,N_970);
nand U1096 (N_1096,N_968,N_964);
nor U1097 (N_1097,N_900,N_943);
nor U1098 (N_1098,N_987,N_952);
nor U1099 (N_1099,N_936,N_954);
or U1100 (N_1100,N_1008,N_1044);
and U1101 (N_1101,N_1069,N_1045);
nand U1102 (N_1102,N_1047,N_1026);
or U1103 (N_1103,N_1057,N_1094);
and U1104 (N_1104,N_1021,N_1049);
and U1105 (N_1105,N_1041,N_1017);
xor U1106 (N_1106,N_1046,N_1007);
or U1107 (N_1107,N_1059,N_1071);
nor U1108 (N_1108,N_1089,N_1043);
nor U1109 (N_1109,N_1067,N_1006);
nand U1110 (N_1110,N_1083,N_1033);
and U1111 (N_1111,N_1036,N_1015);
or U1112 (N_1112,N_1072,N_1056);
nand U1113 (N_1113,N_1080,N_1086);
or U1114 (N_1114,N_1020,N_1016);
nor U1115 (N_1115,N_1031,N_1004);
or U1116 (N_1116,N_1097,N_1084);
or U1117 (N_1117,N_1060,N_1035);
or U1118 (N_1118,N_1091,N_1019);
nor U1119 (N_1119,N_1062,N_1048);
and U1120 (N_1120,N_1024,N_1055);
nand U1121 (N_1121,N_1018,N_1088);
or U1122 (N_1122,N_1030,N_1013);
nand U1123 (N_1123,N_1025,N_1065);
nor U1124 (N_1124,N_1087,N_1038);
or U1125 (N_1125,N_1077,N_1098);
nand U1126 (N_1126,N_1092,N_1011);
nand U1127 (N_1127,N_1029,N_1078);
and U1128 (N_1128,N_1028,N_1034);
nand U1129 (N_1129,N_1051,N_1023);
or U1130 (N_1130,N_1027,N_1093);
nor U1131 (N_1131,N_1002,N_1068);
and U1132 (N_1132,N_1037,N_1096);
nor U1133 (N_1133,N_1042,N_1085);
xor U1134 (N_1134,N_1099,N_1054);
nor U1135 (N_1135,N_1064,N_1074);
xnor U1136 (N_1136,N_1076,N_1040);
or U1137 (N_1137,N_1009,N_1095);
xor U1138 (N_1138,N_1050,N_1005);
nor U1139 (N_1139,N_1082,N_1014);
xnor U1140 (N_1140,N_1058,N_1032);
nand U1141 (N_1141,N_1073,N_1075);
nor U1142 (N_1142,N_1070,N_1079);
nand U1143 (N_1143,N_1022,N_1066);
xor U1144 (N_1144,N_1010,N_1039);
nand U1145 (N_1145,N_1000,N_1001);
nand U1146 (N_1146,N_1063,N_1061);
and U1147 (N_1147,N_1012,N_1052);
or U1148 (N_1148,N_1090,N_1081);
nor U1149 (N_1149,N_1053,N_1003);
and U1150 (N_1150,N_1091,N_1021);
or U1151 (N_1151,N_1088,N_1004);
nand U1152 (N_1152,N_1006,N_1052);
or U1153 (N_1153,N_1007,N_1050);
or U1154 (N_1154,N_1097,N_1035);
or U1155 (N_1155,N_1017,N_1056);
and U1156 (N_1156,N_1005,N_1035);
xor U1157 (N_1157,N_1040,N_1025);
nand U1158 (N_1158,N_1096,N_1033);
and U1159 (N_1159,N_1030,N_1048);
xor U1160 (N_1160,N_1058,N_1013);
nand U1161 (N_1161,N_1043,N_1039);
and U1162 (N_1162,N_1005,N_1073);
or U1163 (N_1163,N_1064,N_1022);
nand U1164 (N_1164,N_1018,N_1022);
nand U1165 (N_1165,N_1001,N_1091);
nand U1166 (N_1166,N_1010,N_1055);
and U1167 (N_1167,N_1074,N_1078);
nand U1168 (N_1168,N_1007,N_1098);
nand U1169 (N_1169,N_1036,N_1071);
and U1170 (N_1170,N_1031,N_1073);
nand U1171 (N_1171,N_1031,N_1090);
and U1172 (N_1172,N_1024,N_1045);
or U1173 (N_1173,N_1025,N_1056);
and U1174 (N_1174,N_1074,N_1057);
and U1175 (N_1175,N_1068,N_1048);
nand U1176 (N_1176,N_1023,N_1036);
and U1177 (N_1177,N_1043,N_1061);
and U1178 (N_1178,N_1065,N_1070);
xor U1179 (N_1179,N_1016,N_1012);
nor U1180 (N_1180,N_1032,N_1055);
nor U1181 (N_1181,N_1069,N_1094);
and U1182 (N_1182,N_1049,N_1050);
and U1183 (N_1183,N_1056,N_1086);
and U1184 (N_1184,N_1064,N_1045);
nor U1185 (N_1185,N_1049,N_1080);
or U1186 (N_1186,N_1062,N_1076);
or U1187 (N_1187,N_1070,N_1091);
nand U1188 (N_1188,N_1026,N_1055);
nor U1189 (N_1189,N_1082,N_1044);
or U1190 (N_1190,N_1015,N_1098);
nor U1191 (N_1191,N_1039,N_1008);
or U1192 (N_1192,N_1093,N_1065);
and U1193 (N_1193,N_1020,N_1014);
nand U1194 (N_1194,N_1014,N_1073);
xor U1195 (N_1195,N_1023,N_1000);
xnor U1196 (N_1196,N_1099,N_1064);
or U1197 (N_1197,N_1061,N_1098);
nor U1198 (N_1198,N_1012,N_1029);
or U1199 (N_1199,N_1014,N_1021);
xnor U1200 (N_1200,N_1169,N_1186);
nand U1201 (N_1201,N_1179,N_1133);
or U1202 (N_1202,N_1191,N_1193);
nor U1203 (N_1203,N_1182,N_1102);
xor U1204 (N_1204,N_1123,N_1175);
nor U1205 (N_1205,N_1177,N_1103);
nand U1206 (N_1206,N_1163,N_1138);
or U1207 (N_1207,N_1160,N_1106);
xor U1208 (N_1208,N_1170,N_1114);
nor U1209 (N_1209,N_1146,N_1121);
nor U1210 (N_1210,N_1132,N_1116);
nand U1211 (N_1211,N_1101,N_1111);
and U1212 (N_1212,N_1153,N_1126);
and U1213 (N_1213,N_1198,N_1155);
or U1214 (N_1214,N_1176,N_1105);
nand U1215 (N_1215,N_1168,N_1144);
and U1216 (N_1216,N_1174,N_1154);
nand U1217 (N_1217,N_1189,N_1173);
nand U1218 (N_1218,N_1143,N_1115);
nand U1219 (N_1219,N_1108,N_1166);
or U1220 (N_1220,N_1159,N_1180);
and U1221 (N_1221,N_1199,N_1149);
nor U1222 (N_1222,N_1158,N_1122);
nor U1223 (N_1223,N_1140,N_1184);
xnor U1224 (N_1224,N_1145,N_1142);
nor U1225 (N_1225,N_1104,N_1109);
or U1226 (N_1226,N_1152,N_1110);
xor U1227 (N_1227,N_1190,N_1181);
or U1228 (N_1228,N_1119,N_1137);
nor U1229 (N_1229,N_1125,N_1100);
nand U1230 (N_1230,N_1130,N_1187);
nor U1231 (N_1231,N_1150,N_1120);
xnor U1232 (N_1232,N_1194,N_1129);
nand U1233 (N_1233,N_1197,N_1127);
nand U1234 (N_1234,N_1117,N_1156);
nor U1235 (N_1235,N_1136,N_1183);
and U1236 (N_1236,N_1185,N_1131);
nand U1237 (N_1237,N_1128,N_1192);
and U1238 (N_1238,N_1139,N_1178);
and U1239 (N_1239,N_1157,N_1118);
nor U1240 (N_1240,N_1107,N_1161);
or U1241 (N_1241,N_1195,N_1124);
or U1242 (N_1242,N_1135,N_1148);
or U1243 (N_1243,N_1196,N_1162);
and U1244 (N_1244,N_1172,N_1164);
nand U1245 (N_1245,N_1147,N_1151);
nand U1246 (N_1246,N_1188,N_1134);
nand U1247 (N_1247,N_1167,N_1112);
nand U1248 (N_1248,N_1141,N_1171);
nor U1249 (N_1249,N_1113,N_1165);
or U1250 (N_1250,N_1181,N_1150);
nor U1251 (N_1251,N_1124,N_1106);
nand U1252 (N_1252,N_1159,N_1188);
nand U1253 (N_1253,N_1124,N_1191);
nor U1254 (N_1254,N_1186,N_1131);
nand U1255 (N_1255,N_1117,N_1151);
or U1256 (N_1256,N_1111,N_1173);
and U1257 (N_1257,N_1192,N_1108);
nor U1258 (N_1258,N_1143,N_1144);
nor U1259 (N_1259,N_1112,N_1149);
nor U1260 (N_1260,N_1152,N_1130);
nand U1261 (N_1261,N_1183,N_1174);
xor U1262 (N_1262,N_1146,N_1190);
and U1263 (N_1263,N_1122,N_1172);
xor U1264 (N_1264,N_1103,N_1194);
and U1265 (N_1265,N_1175,N_1198);
and U1266 (N_1266,N_1115,N_1128);
nor U1267 (N_1267,N_1164,N_1194);
nand U1268 (N_1268,N_1135,N_1166);
nand U1269 (N_1269,N_1180,N_1162);
nand U1270 (N_1270,N_1198,N_1133);
xor U1271 (N_1271,N_1185,N_1190);
nor U1272 (N_1272,N_1132,N_1184);
and U1273 (N_1273,N_1127,N_1145);
and U1274 (N_1274,N_1189,N_1186);
or U1275 (N_1275,N_1150,N_1190);
nand U1276 (N_1276,N_1137,N_1187);
nor U1277 (N_1277,N_1163,N_1136);
nand U1278 (N_1278,N_1161,N_1160);
xnor U1279 (N_1279,N_1167,N_1178);
nand U1280 (N_1280,N_1178,N_1156);
and U1281 (N_1281,N_1148,N_1171);
xnor U1282 (N_1282,N_1132,N_1194);
nand U1283 (N_1283,N_1127,N_1164);
and U1284 (N_1284,N_1196,N_1113);
nand U1285 (N_1285,N_1110,N_1190);
and U1286 (N_1286,N_1106,N_1147);
and U1287 (N_1287,N_1179,N_1180);
nand U1288 (N_1288,N_1158,N_1147);
nor U1289 (N_1289,N_1188,N_1131);
or U1290 (N_1290,N_1174,N_1108);
nor U1291 (N_1291,N_1132,N_1130);
nor U1292 (N_1292,N_1149,N_1117);
and U1293 (N_1293,N_1198,N_1139);
and U1294 (N_1294,N_1158,N_1127);
nor U1295 (N_1295,N_1129,N_1121);
nand U1296 (N_1296,N_1152,N_1195);
nand U1297 (N_1297,N_1163,N_1173);
nor U1298 (N_1298,N_1138,N_1116);
nand U1299 (N_1299,N_1165,N_1156);
nor U1300 (N_1300,N_1278,N_1200);
nor U1301 (N_1301,N_1248,N_1281);
nand U1302 (N_1302,N_1298,N_1211);
and U1303 (N_1303,N_1240,N_1273);
xor U1304 (N_1304,N_1229,N_1255);
and U1305 (N_1305,N_1236,N_1241);
and U1306 (N_1306,N_1271,N_1239);
nand U1307 (N_1307,N_1272,N_1270);
nor U1308 (N_1308,N_1256,N_1243);
and U1309 (N_1309,N_1296,N_1290);
xnor U1310 (N_1310,N_1208,N_1263);
nor U1311 (N_1311,N_1247,N_1244);
and U1312 (N_1312,N_1284,N_1253);
and U1313 (N_1313,N_1213,N_1238);
nand U1314 (N_1314,N_1232,N_1210);
and U1315 (N_1315,N_1203,N_1280);
and U1316 (N_1316,N_1275,N_1258);
nor U1317 (N_1317,N_1282,N_1265);
or U1318 (N_1318,N_1286,N_1214);
nor U1319 (N_1319,N_1204,N_1259);
or U1320 (N_1320,N_1212,N_1264);
or U1321 (N_1321,N_1268,N_1225);
or U1322 (N_1322,N_1215,N_1262);
nor U1323 (N_1323,N_1227,N_1218);
nor U1324 (N_1324,N_1234,N_1267);
and U1325 (N_1325,N_1260,N_1216);
or U1326 (N_1326,N_1249,N_1285);
nor U1327 (N_1327,N_1261,N_1231);
xor U1328 (N_1328,N_1201,N_1230);
nand U1329 (N_1329,N_1276,N_1217);
or U1330 (N_1330,N_1219,N_1233);
nand U1331 (N_1331,N_1279,N_1205);
or U1332 (N_1332,N_1254,N_1207);
or U1333 (N_1333,N_1289,N_1224);
and U1334 (N_1334,N_1293,N_1297);
and U1335 (N_1335,N_1283,N_1257);
nor U1336 (N_1336,N_1250,N_1252);
and U1337 (N_1337,N_1292,N_1299);
or U1338 (N_1338,N_1245,N_1223);
and U1339 (N_1339,N_1202,N_1206);
and U1340 (N_1340,N_1269,N_1266);
or U1341 (N_1341,N_1226,N_1220);
nor U1342 (N_1342,N_1221,N_1228);
nand U1343 (N_1343,N_1288,N_1251);
xnor U1344 (N_1344,N_1209,N_1291);
xnor U1345 (N_1345,N_1287,N_1235);
and U1346 (N_1346,N_1277,N_1222);
and U1347 (N_1347,N_1242,N_1237);
or U1348 (N_1348,N_1295,N_1246);
and U1349 (N_1349,N_1274,N_1294);
nor U1350 (N_1350,N_1252,N_1273);
or U1351 (N_1351,N_1222,N_1287);
or U1352 (N_1352,N_1214,N_1212);
nand U1353 (N_1353,N_1245,N_1213);
nor U1354 (N_1354,N_1267,N_1255);
nor U1355 (N_1355,N_1283,N_1275);
or U1356 (N_1356,N_1252,N_1262);
nand U1357 (N_1357,N_1295,N_1230);
nor U1358 (N_1358,N_1266,N_1256);
or U1359 (N_1359,N_1253,N_1275);
nand U1360 (N_1360,N_1234,N_1228);
and U1361 (N_1361,N_1246,N_1229);
and U1362 (N_1362,N_1256,N_1292);
or U1363 (N_1363,N_1233,N_1258);
and U1364 (N_1364,N_1239,N_1264);
nand U1365 (N_1365,N_1252,N_1214);
or U1366 (N_1366,N_1240,N_1243);
nand U1367 (N_1367,N_1284,N_1256);
xor U1368 (N_1368,N_1259,N_1208);
nor U1369 (N_1369,N_1269,N_1243);
or U1370 (N_1370,N_1239,N_1275);
or U1371 (N_1371,N_1207,N_1231);
and U1372 (N_1372,N_1289,N_1259);
and U1373 (N_1373,N_1287,N_1219);
and U1374 (N_1374,N_1236,N_1245);
and U1375 (N_1375,N_1230,N_1242);
nand U1376 (N_1376,N_1278,N_1276);
nor U1377 (N_1377,N_1275,N_1291);
nor U1378 (N_1378,N_1201,N_1239);
nor U1379 (N_1379,N_1293,N_1261);
nor U1380 (N_1380,N_1257,N_1236);
or U1381 (N_1381,N_1269,N_1231);
nand U1382 (N_1382,N_1215,N_1204);
nand U1383 (N_1383,N_1228,N_1237);
xor U1384 (N_1384,N_1282,N_1202);
and U1385 (N_1385,N_1211,N_1239);
nand U1386 (N_1386,N_1269,N_1284);
nor U1387 (N_1387,N_1231,N_1295);
xor U1388 (N_1388,N_1209,N_1207);
xor U1389 (N_1389,N_1215,N_1201);
and U1390 (N_1390,N_1206,N_1228);
or U1391 (N_1391,N_1266,N_1299);
nand U1392 (N_1392,N_1266,N_1273);
or U1393 (N_1393,N_1235,N_1238);
nand U1394 (N_1394,N_1279,N_1216);
nor U1395 (N_1395,N_1217,N_1233);
and U1396 (N_1396,N_1253,N_1296);
and U1397 (N_1397,N_1269,N_1251);
and U1398 (N_1398,N_1283,N_1201);
or U1399 (N_1399,N_1213,N_1230);
or U1400 (N_1400,N_1328,N_1377);
nand U1401 (N_1401,N_1378,N_1387);
nand U1402 (N_1402,N_1363,N_1366);
or U1403 (N_1403,N_1367,N_1354);
nor U1404 (N_1404,N_1340,N_1358);
nor U1405 (N_1405,N_1344,N_1309);
nor U1406 (N_1406,N_1323,N_1395);
or U1407 (N_1407,N_1389,N_1332);
nor U1408 (N_1408,N_1311,N_1372);
nand U1409 (N_1409,N_1368,N_1350);
nor U1410 (N_1410,N_1370,N_1351);
or U1411 (N_1411,N_1374,N_1365);
or U1412 (N_1412,N_1385,N_1315);
nand U1413 (N_1413,N_1313,N_1347);
nor U1414 (N_1414,N_1357,N_1304);
or U1415 (N_1415,N_1337,N_1376);
nor U1416 (N_1416,N_1348,N_1383);
and U1417 (N_1417,N_1303,N_1391);
nor U1418 (N_1418,N_1375,N_1335);
or U1419 (N_1419,N_1359,N_1382);
or U1420 (N_1420,N_1356,N_1331);
nand U1421 (N_1421,N_1314,N_1310);
nor U1422 (N_1422,N_1381,N_1343);
and U1423 (N_1423,N_1353,N_1321);
or U1424 (N_1424,N_1362,N_1393);
or U1425 (N_1425,N_1326,N_1327);
and U1426 (N_1426,N_1301,N_1345);
or U1427 (N_1427,N_1352,N_1364);
nand U1428 (N_1428,N_1338,N_1324);
nand U1429 (N_1429,N_1336,N_1341);
or U1430 (N_1430,N_1388,N_1380);
nand U1431 (N_1431,N_1342,N_1334);
nand U1432 (N_1432,N_1318,N_1394);
or U1433 (N_1433,N_1308,N_1302);
nand U1434 (N_1434,N_1325,N_1346);
or U1435 (N_1435,N_1317,N_1390);
nor U1436 (N_1436,N_1319,N_1386);
and U1437 (N_1437,N_1316,N_1312);
or U1438 (N_1438,N_1355,N_1320);
and U1439 (N_1439,N_1307,N_1306);
or U1440 (N_1440,N_1329,N_1330);
or U1441 (N_1441,N_1300,N_1361);
xor U1442 (N_1442,N_1396,N_1392);
or U1443 (N_1443,N_1360,N_1369);
nor U1444 (N_1444,N_1322,N_1399);
nor U1445 (N_1445,N_1305,N_1333);
or U1446 (N_1446,N_1371,N_1339);
xor U1447 (N_1447,N_1349,N_1384);
nand U1448 (N_1448,N_1398,N_1379);
and U1449 (N_1449,N_1373,N_1397);
and U1450 (N_1450,N_1314,N_1322);
or U1451 (N_1451,N_1362,N_1334);
and U1452 (N_1452,N_1376,N_1317);
nor U1453 (N_1453,N_1335,N_1322);
or U1454 (N_1454,N_1381,N_1368);
and U1455 (N_1455,N_1348,N_1303);
nor U1456 (N_1456,N_1382,N_1328);
or U1457 (N_1457,N_1360,N_1375);
or U1458 (N_1458,N_1329,N_1335);
or U1459 (N_1459,N_1346,N_1386);
nand U1460 (N_1460,N_1398,N_1342);
or U1461 (N_1461,N_1352,N_1357);
or U1462 (N_1462,N_1314,N_1300);
nand U1463 (N_1463,N_1380,N_1309);
and U1464 (N_1464,N_1341,N_1319);
nand U1465 (N_1465,N_1319,N_1312);
and U1466 (N_1466,N_1313,N_1364);
and U1467 (N_1467,N_1354,N_1327);
and U1468 (N_1468,N_1374,N_1307);
and U1469 (N_1469,N_1329,N_1337);
or U1470 (N_1470,N_1376,N_1346);
or U1471 (N_1471,N_1376,N_1340);
nor U1472 (N_1472,N_1339,N_1359);
or U1473 (N_1473,N_1349,N_1370);
and U1474 (N_1474,N_1363,N_1330);
and U1475 (N_1475,N_1312,N_1322);
and U1476 (N_1476,N_1318,N_1392);
nor U1477 (N_1477,N_1316,N_1317);
and U1478 (N_1478,N_1371,N_1354);
nor U1479 (N_1479,N_1336,N_1378);
or U1480 (N_1480,N_1381,N_1388);
nor U1481 (N_1481,N_1397,N_1387);
or U1482 (N_1482,N_1346,N_1355);
or U1483 (N_1483,N_1366,N_1390);
and U1484 (N_1484,N_1369,N_1346);
or U1485 (N_1485,N_1309,N_1304);
nand U1486 (N_1486,N_1366,N_1339);
nor U1487 (N_1487,N_1311,N_1347);
nor U1488 (N_1488,N_1385,N_1367);
nor U1489 (N_1489,N_1374,N_1340);
and U1490 (N_1490,N_1371,N_1383);
nor U1491 (N_1491,N_1340,N_1347);
nand U1492 (N_1492,N_1330,N_1391);
nor U1493 (N_1493,N_1378,N_1392);
or U1494 (N_1494,N_1387,N_1368);
nand U1495 (N_1495,N_1363,N_1329);
and U1496 (N_1496,N_1376,N_1339);
xnor U1497 (N_1497,N_1355,N_1383);
nand U1498 (N_1498,N_1333,N_1321);
xnor U1499 (N_1499,N_1321,N_1351);
nand U1500 (N_1500,N_1478,N_1431);
xor U1501 (N_1501,N_1453,N_1495);
or U1502 (N_1502,N_1406,N_1451);
or U1503 (N_1503,N_1487,N_1475);
and U1504 (N_1504,N_1452,N_1417);
nor U1505 (N_1505,N_1428,N_1419);
nor U1506 (N_1506,N_1454,N_1456);
and U1507 (N_1507,N_1459,N_1421);
nor U1508 (N_1508,N_1492,N_1461);
nor U1509 (N_1509,N_1489,N_1462);
nand U1510 (N_1510,N_1436,N_1424);
or U1511 (N_1511,N_1444,N_1483);
xnor U1512 (N_1512,N_1496,N_1407);
or U1513 (N_1513,N_1411,N_1498);
or U1514 (N_1514,N_1423,N_1410);
or U1515 (N_1515,N_1439,N_1438);
nor U1516 (N_1516,N_1445,N_1484);
or U1517 (N_1517,N_1471,N_1480);
and U1518 (N_1518,N_1460,N_1450);
nor U1519 (N_1519,N_1499,N_1441);
nor U1520 (N_1520,N_1432,N_1415);
and U1521 (N_1521,N_1486,N_1490);
or U1522 (N_1522,N_1402,N_1469);
and U1523 (N_1523,N_1408,N_1440);
and U1524 (N_1524,N_1463,N_1425);
nand U1525 (N_1525,N_1429,N_1443);
nand U1526 (N_1526,N_1482,N_1473);
nand U1527 (N_1527,N_1400,N_1422);
nor U1528 (N_1528,N_1457,N_1493);
nand U1529 (N_1529,N_1464,N_1420);
and U1530 (N_1530,N_1404,N_1474);
and U1531 (N_1531,N_1466,N_1435);
xor U1532 (N_1532,N_1485,N_1477);
and U1533 (N_1533,N_1458,N_1403);
or U1534 (N_1534,N_1430,N_1413);
nor U1535 (N_1535,N_1470,N_1412);
or U1536 (N_1536,N_1447,N_1416);
nor U1537 (N_1537,N_1427,N_1405);
xor U1538 (N_1538,N_1448,N_1434);
or U1539 (N_1539,N_1497,N_1426);
and U1540 (N_1540,N_1437,N_1488);
nand U1541 (N_1541,N_1442,N_1418);
nor U1542 (N_1542,N_1467,N_1409);
nor U1543 (N_1543,N_1494,N_1491);
and U1544 (N_1544,N_1433,N_1449);
nand U1545 (N_1545,N_1472,N_1455);
or U1546 (N_1546,N_1468,N_1446);
nand U1547 (N_1547,N_1481,N_1401);
and U1548 (N_1548,N_1414,N_1465);
and U1549 (N_1549,N_1476,N_1479);
and U1550 (N_1550,N_1447,N_1415);
or U1551 (N_1551,N_1411,N_1415);
nor U1552 (N_1552,N_1418,N_1459);
and U1553 (N_1553,N_1453,N_1443);
or U1554 (N_1554,N_1452,N_1428);
nor U1555 (N_1555,N_1463,N_1470);
and U1556 (N_1556,N_1482,N_1446);
nand U1557 (N_1557,N_1444,N_1485);
nor U1558 (N_1558,N_1473,N_1447);
nor U1559 (N_1559,N_1414,N_1482);
or U1560 (N_1560,N_1464,N_1430);
and U1561 (N_1561,N_1479,N_1425);
xor U1562 (N_1562,N_1432,N_1417);
nor U1563 (N_1563,N_1412,N_1469);
nand U1564 (N_1564,N_1401,N_1473);
nor U1565 (N_1565,N_1470,N_1486);
or U1566 (N_1566,N_1436,N_1484);
nor U1567 (N_1567,N_1493,N_1492);
nand U1568 (N_1568,N_1489,N_1491);
nor U1569 (N_1569,N_1475,N_1441);
nand U1570 (N_1570,N_1407,N_1452);
and U1571 (N_1571,N_1411,N_1486);
nand U1572 (N_1572,N_1450,N_1482);
and U1573 (N_1573,N_1449,N_1482);
and U1574 (N_1574,N_1404,N_1417);
nor U1575 (N_1575,N_1480,N_1427);
and U1576 (N_1576,N_1450,N_1474);
nor U1577 (N_1577,N_1442,N_1438);
or U1578 (N_1578,N_1471,N_1453);
nor U1579 (N_1579,N_1445,N_1467);
or U1580 (N_1580,N_1491,N_1462);
nand U1581 (N_1581,N_1457,N_1459);
or U1582 (N_1582,N_1492,N_1495);
and U1583 (N_1583,N_1469,N_1462);
and U1584 (N_1584,N_1456,N_1483);
nand U1585 (N_1585,N_1490,N_1477);
and U1586 (N_1586,N_1435,N_1428);
or U1587 (N_1587,N_1431,N_1402);
or U1588 (N_1588,N_1498,N_1453);
and U1589 (N_1589,N_1412,N_1419);
nand U1590 (N_1590,N_1487,N_1481);
and U1591 (N_1591,N_1484,N_1467);
nor U1592 (N_1592,N_1438,N_1467);
nand U1593 (N_1593,N_1411,N_1424);
and U1594 (N_1594,N_1486,N_1446);
nor U1595 (N_1595,N_1429,N_1424);
nor U1596 (N_1596,N_1403,N_1421);
nor U1597 (N_1597,N_1481,N_1424);
or U1598 (N_1598,N_1424,N_1423);
and U1599 (N_1599,N_1491,N_1414);
or U1600 (N_1600,N_1553,N_1592);
nand U1601 (N_1601,N_1557,N_1582);
and U1602 (N_1602,N_1533,N_1549);
or U1603 (N_1603,N_1556,N_1558);
or U1604 (N_1604,N_1522,N_1586);
and U1605 (N_1605,N_1551,N_1535);
or U1606 (N_1606,N_1594,N_1525);
and U1607 (N_1607,N_1544,N_1580);
and U1608 (N_1608,N_1517,N_1502);
or U1609 (N_1609,N_1588,N_1572);
and U1610 (N_1610,N_1577,N_1538);
and U1611 (N_1611,N_1585,N_1515);
nor U1612 (N_1612,N_1598,N_1575);
nand U1613 (N_1613,N_1560,N_1569);
nor U1614 (N_1614,N_1563,N_1532);
nand U1615 (N_1615,N_1584,N_1540);
nand U1616 (N_1616,N_1587,N_1506);
nor U1617 (N_1617,N_1518,N_1581);
or U1618 (N_1618,N_1593,N_1512);
nor U1619 (N_1619,N_1537,N_1564);
nor U1620 (N_1620,N_1519,N_1555);
and U1621 (N_1621,N_1526,N_1591);
and U1622 (N_1622,N_1552,N_1507);
nor U1623 (N_1623,N_1562,N_1501);
nand U1624 (N_1624,N_1559,N_1528);
nor U1625 (N_1625,N_1510,N_1570);
and U1626 (N_1626,N_1503,N_1520);
nor U1627 (N_1627,N_1567,N_1590);
nor U1628 (N_1628,N_1524,N_1541);
xnor U1629 (N_1629,N_1542,N_1546);
or U1630 (N_1630,N_1523,N_1534);
or U1631 (N_1631,N_1548,N_1565);
or U1632 (N_1632,N_1583,N_1539);
or U1633 (N_1633,N_1596,N_1573);
or U1634 (N_1634,N_1529,N_1514);
nor U1635 (N_1635,N_1513,N_1561);
and U1636 (N_1636,N_1500,N_1571);
nand U1637 (N_1637,N_1574,N_1599);
or U1638 (N_1638,N_1554,N_1509);
or U1639 (N_1639,N_1543,N_1516);
and U1640 (N_1640,N_1531,N_1504);
xnor U1641 (N_1641,N_1536,N_1527);
or U1642 (N_1642,N_1505,N_1589);
xnor U1643 (N_1643,N_1568,N_1508);
and U1644 (N_1644,N_1511,N_1530);
or U1645 (N_1645,N_1597,N_1550);
and U1646 (N_1646,N_1521,N_1576);
nor U1647 (N_1647,N_1579,N_1547);
and U1648 (N_1648,N_1545,N_1595);
nor U1649 (N_1649,N_1578,N_1566);
nand U1650 (N_1650,N_1547,N_1506);
and U1651 (N_1651,N_1582,N_1522);
nand U1652 (N_1652,N_1510,N_1577);
nand U1653 (N_1653,N_1561,N_1571);
nor U1654 (N_1654,N_1585,N_1540);
nor U1655 (N_1655,N_1556,N_1513);
nor U1656 (N_1656,N_1563,N_1579);
or U1657 (N_1657,N_1511,N_1542);
or U1658 (N_1658,N_1544,N_1555);
nor U1659 (N_1659,N_1544,N_1502);
or U1660 (N_1660,N_1596,N_1535);
and U1661 (N_1661,N_1543,N_1587);
nand U1662 (N_1662,N_1572,N_1544);
nand U1663 (N_1663,N_1594,N_1592);
and U1664 (N_1664,N_1509,N_1511);
or U1665 (N_1665,N_1590,N_1501);
nand U1666 (N_1666,N_1588,N_1568);
xnor U1667 (N_1667,N_1550,N_1506);
nand U1668 (N_1668,N_1520,N_1594);
xor U1669 (N_1669,N_1590,N_1552);
nand U1670 (N_1670,N_1578,N_1519);
xnor U1671 (N_1671,N_1534,N_1591);
and U1672 (N_1672,N_1512,N_1598);
or U1673 (N_1673,N_1562,N_1572);
and U1674 (N_1674,N_1577,N_1554);
nand U1675 (N_1675,N_1542,N_1599);
and U1676 (N_1676,N_1582,N_1586);
and U1677 (N_1677,N_1505,N_1528);
xor U1678 (N_1678,N_1582,N_1592);
and U1679 (N_1679,N_1526,N_1573);
nor U1680 (N_1680,N_1543,N_1531);
nor U1681 (N_1681,N_1515,N_1503);
or U1682 (N_1682,N_1595,N_1526);
and U1683 (N_1683,N_1533,N_1582);
nor U1684 (N_1684,N_1512,N_1581);
and U1685 (N_1685,N_1552,N_1574);
and U1686 (N_1686,N_1536,N_1534);
nor U1687 (N_1687,N_1510,N_1592);
or U1688 (N_1688,N_1541,N_1517);
and U1689 (N_1689,N_1512,N_1597);
and U1690 (N_1690,N_1515,N_1525);
or U1691 (N_1691,N_1588,N_1511);
or U1692 (N_1692,N_1502,N_1573);
or U1693 (N_1693,N_1544,N_1573);
nor U1694 (N_1694,N_1596,N_1500);
or U1695 (N_1695,N_1576,N_1591);
or U1696 (N_1696,N_1510,N_1514);
xnor U1697 (N_1697,N_1572,N_1545);
or U1698 (N_1698,N_1589,N_1559);
and U1699 (N_1699,N_1521,N_1503);
or U1700 (N_1700,N_1651,N_1654);
nand U1701 (N_1701,N_1615,N_1663);
or U1702 (N_1702,N_1632,N_1688);
and U1703 (N_1703,N_1686,N_1687);
nor U1704 (N_1704,N_1690,N_1635);
xnor U1705 (N_1705,N_1618,N_1648);
nor U1706 (N_1706,N_1626,N_1667);
or U1707 (N_1707,N_1657,N_1645);
xnor U1708 (N_1708,N_1697,N_1656);
nor U1709 (N_1709,N_1676,N_1605);
or U1710 (N_1710,N_1642,N_1658);
xor U1711 (N_1711,N_1679,N_1602);
nor U1712 (N_1712,N_1673,N_1601);
and U1713 (N_1713,N_1627,N_1681);
nand U1714 (N_1714,N_1649,N_1613);
nor U1715 (N_1715,N_1680,N_1699);
nor U1716 (N_1716,N_1664,N_1689);
nand U1717 (N_1717,N_1671,N_1606);
nor U1718 (N_1718,N_1684,N_1604);
xor U1719 (N_1719,N_1625,N_1647);
or U1720 (N_1720,N_1655,N_1662);
or U1721 (N_1721,N_1638,N_1614);
and U1722 (N_1722,N_1650,N_1616);
or U1723 (N_1723,N_1659,N_1675);
or U1724 (N_1724,N_1660,N_1674);
nor U1725 (N_1725,N_1661,N_1668);
and U1726 (N_1726,N_1646,N_1665);
nor U1727 (N_1727,N_1682,N_1610);
and U1728 (N_1728,N_1644,N_1677);
xor U1729 (N_1729,N_1693,N_1640);
or U1730 (N_1730,N_1622,N_1685);
xnor U1731 (N_1731,N_1666,N_1696);
xnor U1732 (N_1732,N_1608,N_1636);
and U1733 (N_1733,N_1619,N_1670);
and U1734 (N_1734,N_1600,N_1611);
or U1735 (N_1735,N_1695,N_1698);
or U1736 (N_1736,N_1683,N_1628);
nor U1737 (N_1737,N_1653,N_1634);
nor U1738 (N_1738,N_1652,N_1617);
and U1739 (N_1739,N_1630,N_1621);
nor U1740 (N_1740,N_1633,N_1641);
nor U1741 (N_1741,N_1607,N_1637);
nand U1742 (N_1742,N_1603,N_1694);
and U1743 (N_1743,N_1612,N_1692);
or U1744 (N_1744,N_1620,N_1678);
or U1745 (N_1745,N_1691,N_1623);
or U1746 (N_1746,N_1672,N_1609);
nand U1747 (N_1747,N_1629,N_1643);
nand U1748 (N_1748,N_1631,N_1639);
nand U1749 (N_1749,N_1624,N_1669);
xnor U1750 (N_1750,N_1645,N_1613);
nor U1751 (N_1751,N_1671,N_1611);
or U1752 (N_1752,N_1656,N_1640);
or U1753 (N_1753,N_1653,N_1626);
and U1754 (N_1754,N_1658,N_1650);
and U1755 (N_1755,N_1607,N_1614);
or U1756 (N_1756,N_1618,N_1631);
nor U1757 (N_1757,N_1626,N_1627);
or U1758 (N_1758,N_1611,N_1652);
nor U1759 (N_1759,N_1697,N_1669);
nor U1760 (N_1760,N_1637,N_1695);
and U1761 (N_1761,N_1609,N_1662);
or U1762 (N_1762,N_1650,N_1671);
and U1763 (N_1763,N_1631,N_1671);
and U1764 (N_1764,N_1628,N_1637);
nor U1765 (N_1765,N_1651,N_1640);
nand U1766 (N_1766,N_1621,N_1625);
and U1767 (N_1767,N_1645,N_1614);
nand U1768 (N_1768,N_1677,N_1625);
and U1769 (N_1769,N_1670,N_1691);
or U1770 (N_1770,N_1601,N_1604);
and U1771 (N_1771,N_1696,N_1691);
and U1772 (N_1772,N_1695,N_1679);
and U1773 (N_1773,N_1627,N_1613);
xor U1774 (N_1774,N_1630,N_1624);
xnor U1775 (N_1775,N_1629,N_1612);
nand U1776 (N_1776,N_1653,N_1615);
nand U1777 (N_1777,N_1683,N_1666);
nor U1778 (N_1778,N_1663,N_1609);
xnor U1779 (N_1779,N_1661,N_1616);
and U1780 (N_1780,N_1616,N_1645);
or U1781 (N_1781,N_1663,N_1693);
and U1782 (N_1782,N_1603,N_1655);
or U1783 (N_1783,N_1655,N_1619);
nor U1784 (N_1784,N_1671,N_1601);
nor U1785 (N_1785,N_1639,N_1642);
nand U1786 (N_1786,N_1698,N_1613);
xor U1787 (N_1787,N_1653,N_1655);
nand U1788 (N_1788,N_1600,N_1622);
and U1789 (N_1789,N_1609,N_1654);
nor U1790 (N_1790,N_1668,N_1664);
and U1791 (N_1791,N_1671,N_1656);
and U1792 (N_1792,N_1677,N_1607);
nor U1793 (N_1793,N_1619,N_1645);
or U1794 (N_1794,N_1607,N_1666);
xnor U1795 (N_1795,N_1680,N_1611);
nand U1796 (N_1796,N_1690,N_1681);
and U1797 (N_1797,N_1645,N_1639);
xnor U1798 (N_1798,N_1606,N_1616);
xor U1799 (N_1799,N_1630,N_1642);
nand U1800 (N_1800,N_1787,N_1741);
nand U1801 (N_1801,N_1759,N_1776);
and U1802 (N_1802,N_1785,N_1798);
xnor U1803 (N_1803,N_1714,N_1723);
nand U1804 (N_1804,N_1764,N_1724);
and U1805 (N_1805,N_1718,N_1726);
or U1806 (N_1806,N_1789,N_1751);
xor U1807 (N_1807,N_1781,N_1775);
and U1808 (N_1808,N_1797,N_1712);
nand U1809 (N_1809,N_1732,N_1734);
nor U1810 (N_1810,N_1760,N_1778);
xnor U1811 (N_1811,N_1709,N_1737);
nor U1812 (N_1812,N_1743,N_1738);
nand U1813 (N_1813,N_1720,N_1711);
xor U1814 (N_1814,N_1773,N_1755);
or U1815 (N_1815,N_1747,N_1766);
nor U1816 (N_1816,N_1728,N_1742);
nor U1817 (N_1817,N_1750,N_1730);
nor U1818 (N_1818,N_1795,N_1727);
or U1819 (N_1819,N_1716,N_1763);
or U1820 (N_1820,N_1706,N_1792);
nor U1821 (N_1821,N_1765,N_1768);
or U1822 (N_1822,N_1774,N_1736);
nor U1823 (N_1823,N_1782,N_1721);
or U1824 (N_1824,N_1703,N_1746);
nand U1825 (N_1825,N_1796,N_1758);
and U1826 (N_1826,N_1739,N_1704);
or U1827 (N_1827,N_1702,N_1710);
nor U1828 (N_1828,N_1794,N_1744);
or U1829 (N_1829,N_1770,N_1757);
and U1830 (N_1830,N_1753,N_1707);
nand U1831 (N_1831,N_1779,N_1767);
nor U1832 (N_1832,N_1783,N_1788);
nand U1833 (N_1833,N_1748,N_1769);
or U1834 (N_1834,N_1756,N_1719);
nor U1835 (N_1835,N_1791,N_1749);
or U1836 (N_1836,N_1772,N_1780);
xor U1837 (N_1837,N_1722,N_1708);
nor U1838 (N_1838,N_1752,N_1777);
nand U1839 (N_1839,N_1735,N_1793);
or U1840 (N_1840,N_1784,N_1717);
nor U1841 (N_1841,N_1715,N_1725);
and U1842 (N_1842,N_1713,N_1786);
nand U1843 (N_1843,N_1754,N_1790);
or U1844 (N_1844,N_1740,N_1700);
nor U1845 (N_1845,N_1745,N_1771);
or U1846 (N_1846,N_1705,N_1761);
or U1847 (N_1847,N_1799,N_1729);
nor U1848 (N_1848,N_1733,N_1762);
or U1849 (N_1849,N_1701,N_1731);
nor U1850 (N_1850,N_1720,N_1779);
nor U1851 (N_1851,N_1781,N_1754);
nand U1852 (N_1852,N_1738,N_1714);
nor U1853 (N_1853,N_1702,N_1709);
or U1854 (N_1854,N_1728,N_1798);
and U1855 (N_1855,N_1736,N_1782);
nor U1856 (N_1856,N_1796,N_1713);
or U1857 (N_1857,N_1754,N_1788);
nand U1858 (N_1858,N_1785,N_1790);
or U1859 (N_1859,N_1798,N_1788);
or U1860 (N_1860,N_1776,N_1755);
nand U1861 (N_1861,N_1797,N_1705);
or U1862 (N_1862,N_1772,N_1732);
or U1863 (N_1863,N_1748,N_1786);
or U1864 (N_1864,N_1766,N_1786);
xor U1865 (N_1865,N_1799,N_1716);
nor U1866 (N_1866,N_1791,N_1736);
xor U1867 (N_1867,N_1723,N_1793);
or U1868 (N_1868,N_1741,N_1772);
or U1869 (N_1869,N_1799,N_1782);
or U1870 (N_1870,N_1710,N_1760);
nand U1871 (N_1871,N_1736,N_1784);
nor U1872 (N_1872,N_1723,N_1768);
or U1873 (N_1873,N_1750,N_1718);
nor U1874 (N_1874,N_1710,N_1787);
or U1875 (N_1875,N_1706,N_1766);
nand U1876 (N_1876,N_1733,N_1721);
or U1877 (N_1877,N_1757,N_1794);
nor U1878 (N_1878,N_1719,N_1772);
or U1879 (N_1879,N_1799,N_1791);
and U1880 (N_1880,N_1791,N_1768);
xor U1881 (N_1881,N_1789,N_1703);
or U1882 (N_1882,N_1752,N_1721);
and U1883 (N_1883,N_1726,N_1702);
nor U1884 (N_1884,N_1718,N_1759);
nor U1885 (N_1885,N_1723,N_1746);
or U1886 (N_1886,N_1702,N_1799);
nand U1887 (N_1887,N_1710,N_1743);
or U1888 (N_1888,N_1738,N_1747);
and U1889 (N_1889,N_1738,N_1774);
nor U1890 (N_1890,N_1797,N_1720);
or U1891 (N_1891,N_1758,N_1786);
nor U1892 (N_1892,N_1744,N_1714);
nand U1893 (N_1893,N_1737,N_1795);
or U1894 (N_1894,N_1755,N_1779);
xor U1895 (N_1895,N_1722,N_1707);
or U1896 (N_1896,N_1775,N_1702);
or U1897 (N_1897,N_1728,N_1715);
nor U1898 (N_1898,N_1799,N_1794);
or U1899 (N_1899,N_1735,N_1762);
xor U1900 (N_1900,N_1841,N_1889);
and U1901 (N_1901,N_1877,N_1830);
or U1902 (N_1902,N_1856,N_1848);
nand U1903 (N_1903,N_1855,N_1898);
nand U1904 (N_1904,N_1815,N_1891);
nor U1905 (N_1905,N_1821,N_1828);
nand U1906 (N_1906,N_1868,N_1819);
and U1907 (N_1907,N_1814,N_1862);
xnor U1908 (N_1908,N_1849,N_1853);
nor U1909 (N_1909,N_1852,N_1879);
nand U1910 (N_1910,N_1832,N_1854);
nand U1911 (N_1911,N_1873,N_1834);
xor U1912 (N_1912,N_1831,N_1803);
nor U1913 (N_1913,N_1822,N_1897);
nand U1914 (N_1914,N_1847,N_1837);
or U1915 (N_1915,N_1888,N_1857);
and U1916 (N_1916,N_1885,N_1836);
and U1917 (N_1917,N_1835,N_1818);
nor U1918 (N_1918,N_1858,N_1874);
nand U1919 (N_1919,N_1878,N_1866);
nor U1920 (N_1920,N_1850,N_1809);
and U1921 (N_1921,N_1802,N_1861);
and U1922 (N_1922,N_1880,N_1865);
or U1923 (N_1923,N_1844,N_1846);
nor U1924 (N_1924,N_1826,N_1833);
or U1925 (N_1925,N_1827,N_1838);
or U1926 (N_1926,N_1867,N_1871);
nand U1927 (N_1927,N_1881,N_1842);
or U1928 (N_1928,N_1816,N_1895);
or U1929 (N_1929,N_1869,N_1876);
and U1930 (N_1930,N_1886,N_1829);
nor U1931 (N_1931,N_1825,N_1807);
nor U1932 (N_1932,N_1804,N_1812);
or U1933 (N_1933,N_1882,N_1813);
nand U1934 (N_1934,N_1896,N_1859);
nor U1935 (N_1935,N_1890,N_1800);
or U1936 (N_1936,N_1845,N_1840);
and U1937 (N_1937,N_1805,N_1824);
nor U1938 (N_1938,N_1875,N_1860);
nor U1939 (N_1939,N_1864,N_1893);
nor U1940 (N_1940,N_1883,N_1839);
and U1941 (N_1941,N_1811,N_1872);
or U1942 (N_1942,N_1806,N_1810);
or U1943 (N_1943,N_1851,N_1801);
xnor U1944 (N_1944,N_1887,N_1808);
or U1945 (N_1945,N_1863,N_1843);
xor U1946 (N_1946,N_1823,N_1870);
nor U1947 (N_1947,N_1817,N_1820);
xor U1948 (N_1948,N_1894,N_1892);
or U1949 (N_1949,N_1884,N_1899);
nor U1950 (N_1950,N_1834,N_1856);
nand U1951 (N_1951,N_1864,N_1853);
xnor U1952 (N_1952,N_1881,N_1848);
nand U1953 (N_1953,N_1876,N_1841);
and U1954 (N_1954,N_1821,N_1868);
nor U1955 (N_1955,N_1841,N_1883);
or U1956 (N_1956,N_1832,N_1807);
and U1957 (N_1957,N_1857,N_1823);
xor U1958 (N_1958,N_1896,N_1868);
xnor U1959 (N_1959,N_1868,N_1839);
nand U1960 (N_1960,N_1894,N_1847);
nor U1961 (N_1961,N_1805,N_1814);
or U1962 (N_1962,N_1886,N_1863);
or U1963 (N_1963,N_1878,N_1813);
and U1964 (N_1964,N_1880,N_1838);
and U1965 (N_1965,N_1891,N_1862);
or U1966 (N_1966,N_1850,N_1821);
nor U1967 (N_1967,N_1896,N_1810);
or U1968 (N_1968,N_1884,N_1808);
nor U1969 (N_1969,N_1891,N_1879);
and U1970 (N_1970,N_1843,N_1813);
nor U1971 (N_1971,N_1881,N_1808);
or U1972 (N_1972,N_1849,N_1824);
nor U1973 (N_1973,N_1818,N_1841);
and U1974 (N_1974,N_1881,N_1868);
nor U1975 (N_1975,N_1893,N_1879);
and U1976 (N_1976,N_1889,N_1829);
and U1977 (N_1977,N_1884,N_1817);
and U1978 (N_1978,N_1820,N_1807);
and U1979 (N_1979,N_1864,N_1879);
and U1980 (N_1980,N_1858,N_1822);
or U1981 (N_1981,N_1846,N_1820);
or U1982 (N_1982,N_1894,N_1831);
or U1983 (N_1983,N_1894,N_1828);
xor U1984 (N_1984,N_1889,N_1880);
and U1985 (N_1985,N_1838,N_1894);
or U1986 (N_1986,N_1815,N_1801);
nand U1987 (N_1987,N_1837,N_1865);
xor U1988 (N_1988,N_1801,N_1859);
and U1989 (N_1989,N_1860,N_1829);
or U1990 (N_1990,N_1879,N_1884);
or U1991 (N_1991,N_1819,N_1847);
or U1992 (N_1992,N_1839,N_1865);
or U1993 (N_1993,N_1897,N_1896);
xnor U1994 (N_1994,N_1821,N_1808);
xor U1995 (N_1995,N_1891,N_1800);
nand U1996 (N_1996,N_1852,N_1869);
or U1997 (N_1997,N_1832,N_1833);
or U1998 (N_1998,N_1813,N_1855);
nand U1999 (N_1999,N_1834,N_1882);
nor U2000 (N_2000,N_1912,N_1991);
nand U2001 (N_2001,N_1947,N_1922);
nand U2002 (N_2002,N_1910,N_1934);
and U2003 (N_2003,N_1990,N_1917);
or U2004 (N_2004,N_1982,N_1953);
nand U2005 (N_2005,N_1913,N_1948);
or U2006 (N_2006,N_1929,N_1911);
and U2007 (N_2007,N_1995,N_1945);
nor U2008 (N_2008,N_1985,N_1957);
or U2009 (N_2009,N_1996,N_1942);
nand U2010 (N_2010,N_1973,N_1966);
and U2011 (N_2011,N_1908,N_1987);
and U2012 (N_2012,N_1964,N_1979);
and U2013 (N_2013,N_1943,N_1926);
or U2014 (N_2014,N_1967,N_1937);
nand U2015 (N_2015,N_1930,N_1921);
or U2016 (N_2016,N_1915,N_1909);
nand U2017 (N_2017,N_1997,N_1970);
nor U2018 (N_2018,N_1977,N_1932);
nor U2019 (N_2019,N_1975,N_1992);
or U2020 (N_2020,N_1935,N_1994);
nor U2021 (N_2021,N_1952,N_1924);
and U2022 (N_2022,N_1965,N_1931);
or U2023 (N_2023,N_1904,N_1989);
nand U2024 (N_2024,N_1981,N_1984);
and U2025 (N_2025,N_1958,N_1928);
nor U2026 (N_2026,N_1933,N_1941);
or U2027 (N_2027,N_1901,N_1902);
and U2028 (N_2028,N_1919,N_1914);
nor U2029 (N_2029,N_1944,N_1925);
and U2030 (N_2030,N_1905,N_1951);
and U2031 (N_2031,N_1923,N_1903);
and U2032 (N_2032,N_1972,N_1974);
nand U2033 (N_2033,N_1939,N_1988);
nor U2034 (N_2034,N_1916,N_1962);
or U2035 (N_2035,N_1968,N_1938);
xor U2036 (N_2036,N_1927,N_1976);
nand U2037 (N_2037,N_1971,N_1999);
nor U2038 (N_2038,N_1963,N_1900);
or U2039 (N_2039,N_1980,N_1959);
or U2040 (N_2040,N_1986,N_1906);
nor U2041 (N_2041,N_1998,N_1978);
nor U2042 (N_2042,N_1940,N_1936);
xnor U2043 (N_2043,N_1920,N_1961);
or U2044 (N_2044,N_1946,N_1907);
and U2045 (N_2045,N_1983,N_1993);
nand U2046 (N_2046,N_1950,N_1956);
nor U2047 (N_2047,N_1954,N_1949);
nor U2048 (N_2048,N_1918,N_1960);
or U2049 (N_2049,N_1969,N_1955);
nor U2050 (N_2050,N_1907,N_1977);
and U2051 (N_2051,N_1926,N_1918);
or U2052 (N_2052,N_1999,N_1923);
nor U2053 (N_2053,N_1924,N_1993);
and U2054 (N_2054,N_1929,N_1945);
nand U2055 (N_2055,N_1995,N_1917);
and U2056 (N_2056,N_1992,N_1999);
or U2057 (N_2057,N_1904,N_1974);
or U2058 (N_2058,N_1948,N_1904);
xnor U2059 (N_2059,N_1992,N_1905);
or U2060 (N_2060,N_1938,N_1926);
and U2061 (N_2061,N_1995,N_1932);
xnor U2062 (N_2062,N_1984,N_1965);
nand U2063 (N_2063,N_1969,N_1968);
nand U2064 (N_2064,N_1953,N_1936);
nand U2065 (N_2065,N_1997,N_1943);
or U2066 (N_2066,N_1993,N_1973);
or U2067 (N_2067,N_1939,N_1979);
nand U2068 (N_2068,N_1994,N_1902);
nor U2069 (N_2069,N_1994,N_1933);
nor U2070 (N_2070,N_1915,N_1918);
nor U2071 (N_2071,N_1931,N_1987);
nor U2072 (N_2072,N_1900,N_1927);
nand U2073 (N_2073,N_1987,N_1922);
or U2074 (N_2074,N_1911,N_1917);
nand U2075 (N_2075,N_1986,N_1995);
or U2076 (N_2076,N_1926,N_1960);
nand U2077 (N_2077,N_1972,N_1908);
or U2078 (N_2078,N_1925,N_1924);
or U2079 (N_2079,N_1901,N_1982);
and U2080 (N_2080,N_1906,N_1940);
or U2081 (N_2081,N_1935,N_1939);
nor U2082 (N_2082,N_1914,N_1991);
nor U2083 (N_2083,N_1968,N_1932);
and U2084 (N_2084,N_1916,N_1905);
nand U2085 (N_2085,N_1939,N_1914);
and U2086 (N_2086,N_1925,N_1993);
nor U2087 (N_2087,N_1916,N_1939);
xnor U2088 (N_2088,N_1963,N_1950);
or U2089 (N_2089,N_1994,N_1999);
nor U2090 (N_2090,N_1918,N_1941);
nand U2091 (N_2091,N_1924,N_1999);
nor U2092 (N_2092,N_1966,N_1961);
nor U2093 (N_2093,N_1991,N_1986);
nor U2094 (N_2094,N_1900,N_1933);
nand U2095 (N_2095,N_1901,N_1920);
and U2096 (N_2096,N_1998,N_1921);
nor U2097 (N_2097,N_1983,N_1925);
nand U2098 (N_2098,N_1991,N_1968);
nor U2099 (N_2099,N_1974,N_1926);
nor U2100 (N_2100,N_2001,N_2069);
nand U2101 (N_2101,N_2088,N_2018);
nor U2102 (N_2102,N_2079,N_2058);
and U2103 (N_2103,N_2024,N_2054);
and U2104 (N_2104,N_2081,N_2065);
or U2105 (N_2105,N_2023,N_2060);
nand U2106 (N_2106,N_2020,N_2002);
nand U2107 (N_2107,N_2011,N_2091);
and U2108 (N_2108,N_2074,N_2008);
or U2109 (N_2109,N_2010,N_2046);
and U2110 (N_2110,N_2077,N_2005);
or U2111 (N_2111,N_2044,N_2071);
nor U2112 (N_2112,N_2038,N_2098);
or U2113 (N_2113,N_2035,N_2097);
nor U2114 (N_2114,N_2029,N_2087);
or U2115 (N_2115,N_2043,N_2063);
or U2116 (N_2116,N_2013,N_2022);
xnor U2117 (N_2117,N_2070,N_2033);
nor U2118 (N_2118,N_2007,N_2084);
nand U2119 (N_2119,N_2004,N_2086);
or U2120 (N_2120,N_2080,N_2051);
and U2121 (N_2121,N_2036,N_2014);
and U2122 (N_2122,N_2021,N_2061);
xnor U2123 (N_2123,N_2093,N_2045);
nor U2124 (N_2124,N_2027,N_2025);
nor U2125 (N_2125,N_2019,N_2050);
or U2126 (N_2126,N_2083,N_2053);
nor U2127 (N_2127,N_2003,N_2030);
or U2128 (N_2128,N_2057,N_2040);
nand U2129 (N_2129,N_2016,N_2082);
and U2130 (N_2130,N_2078,N_2076);
or U2131 (N_2131,N_2094,N_2096);
nand U2132 (N_2132,N_2042,N_2055);
nand U2133 (N_2133,N_2099,N_2012);
and U2134 (N_2134,N_2015,N_2006);
or U2135 (N_2135,N_2041,N_2034);
and U2136 (N_2136,N_2047,N_2056);
nand U2137 (N_2137,N_2017,N_2048);
nor U2138 (N_2138,N_2037,N_2095);
nand U2139 (N_2139,N_2026,N_2090);
or U2140 (N_2140,N_2085,N_2028);
xor U2141 (N_2141,N_2072,N_2049);
xnor U2142 (N_2142,N_2067,N_2092);
nand U2143 (N_2143,N_2000,N_2031);
nor U2144 (N_2144,N_2068,N_2059);
nand U2145 (N_2145,N_2052,N_2073);
and U2146 (N_2146,N_2089,N_2064);
nor U2147 (N_2147,N_2062,N_2009);
nor U2148 (N_2148,N_2032,N_2066);
and U2149 (N_2149,N_2039,N_2075);
or U2150 (N_2150,N_2059,N_2061);
or U2151 (N_2151,N_2085,N_2076);
nand U2152 (N_2152,N_2035,N_2056);
and U2153 (N_2153,N_2084,N_2053);
or U2154 (N_2154,N_2087,N_2018);
nand U2155 (N_2155,N_2094,N_2044);
xor U2156 (N_2156,N_2087,N_2084);
nor U2157 (N_2157,N_2031,N_2007);
nand U2158 (N_2158,N_2002,N_2003);
and U2159 (N_2159,N_2015,N_2029);
nand U2160 (N_2160,N_2047,N_2060);
and U2161 (N_2161,N_2072,N_2073);
or U2162 (N_2162,N_2026,N_2064);
nor U2163 (N_2163,N_2079,N_2033);
nand U2164 (N_2164,N_2021,N_2012);
nor U2165 (N_2165,N_2041,N_2077);
or U2166 (N_2166,N_2067,N_2058);
nor U2167 (N_2167,N_2078,N_2037);
nor U2168 (N_2168,N_2061,N_2013);
and U2169 (N_2169,N_2034,N_2000);
nor U2170 (N_2170,N_2026,N_2021);
and U2171 (N_2171,N_2085,N_2052);
and U2172 (N_2172,N_2031,N_2099);
nand U2173 (N_2173,N_2014,N_2010);
nor U2174 (N_2174,N_2059,N_2082);
or U2175 (N_2175,N_2053,N_2058);
nor U2176 (N_2176,N_2053,N_2016);
and U2177 (N_2177,N_2045,N_2053);
or U2178 (N_2178,N_2050,N_2068);
nand U2179 (N_2179,N_2087,N_2085);
or U2180 (N_2180,N_2072,N_2024);
nand U2181 (N_2181,N_2082,N_2017);
xnor U2182 (N_2182,N_2084,N_2068);
or U2183 (N_2183,N_2090,N_2014);
xor U2184 (N_2184,N_2071,N_2078);
nor U2185 (N_2185,N_2044,N_2000);
xor U2186 (N_2186,N_2086,N_2027);
nand U2187 (N_2187,N_2066,N_2081);
xnor U2188 (N_2188,N_2091,N_2077);
nand U2189 (N_2189,N_2017,N_2094);
and U2190 (N_2190,N_2018,N_2016);
or U2191 (N_2191,N_2068,N_2002);
or U2192 (N_2192,N_2097,N_2064);
and U2193 (N_2193,N_2062,N_2090);
and U2194 (N_2194,N_2049,N_2017);
or U2195 (N_2195,N_2035,N_2028);
or U2196 (N_2196,N_2067,N_2076);
and U2197 (N_2197,N_2097,N_2006);
and U2198 (N_2198,N_2067,N_2066);
nor U2199 (N_2199,N_2005,N_2021);
and U2200 (N_2200,N_2116,N_2139);
or U2201 (N_2201,N_2138,N_2182);
nor U2202 (N_2202,N_2159,N_2176);
nor U2203 (N_2203,N_2170,N_2149);
nor U2204 (N_2204,N_2109,N_2106);
and U2205 (N_2205,N_2115,N_2123);
or U2206 (N_2206,N_2187,N_2144);
nor U2207 (N_2207,N_2146,N_2185);
nor U2208 (N_2208,N_2184,N_2136);
or U2209 (N_2209,N_2131,N_2105);
or U2210 (N_2210,N_2178,N_2108);
and U2211 (N_2211,N_2104,N_2151);
and U2212 (N_2212,N_2177,N_2143);
and U2213 (N_2213,N_2197,N_2158);
and U2214 (N_2214,N_2118,N_2125);
and U2215 (N_2215,N_2145,N_2169);
and U2216 (N_2216,N_2186,N_2100);
nor U2217 (N_2217,N_2124,N_2107);
or U2218 (N_2218,N_2193,N_2127);
nand U2219 (N_2219,N_2183,N_2128);
nor U2220 (N_2220,N_2126,N_2110);
nor U2221 (N_2221,N_2171,N_2164);
nand U2222 (N_2222,N_2167,N_2165);
and U2223 (N_2223,N_2163,N_2117);
and U2224 (N_2224,N_2111,N_2150);
nor U2225 (N_2225,N_2132,N_2134);
or U2226 (N_2226,N_2156,N_2129);
nand U2227 (N_2227,N_2162,N_2174);
nand U2228 (N_2228,N_2113,N_2173);
nor U2229 (N_2229,N_2192,N_2191);
and U2230 (N_2230,N_2168,N_2140);
xnor U2231 (N_2231,N_2101,N_2142);
nor U2232 (N_2232,N_2122,N_2160);
nand U2233 (N_2233,N_2119,N_2133);
nand U2234 (N_2234,N_2172,N_2152);
and U2235 (N_2235,N_2180,N_2154);
nand U2236 (N_2236,N_2135,N_2166);
or U2237 (N_2237,N_2188,N_2137);
and U2238 (N_2238,N_2161,N_2196);
or U2239 (N_2239,N_2194,N_2181);
or U2240 (N_2240,N_2190,N_2155);
or U2241 (N_2241,N_2148,N_2147);
and U2242 (N_2242,N_2130,N_2141);
nand U2243 (N_2243,N_2175,N_2199);
xor U2244 (N_2244,N_2121,N_2103);
or U2245 (N_2245,N_2120,N_2153);
xor U2246 (N_2246,N_2102,N_2195);
or U2247 (N_2247,N_2112,N_2114);
xnor U2248 (N_2248,N_2189,N_2179);
or U2249 (N_2249,N_2157,N_2198);
nor U2250 (N_2250,N_2197,N_2169);
nor U2251 (N_2251,N_2140,N_2146);
nand U2252 (N_2252,N_2160,N_2157);
and U2253 (N_2253,N_2180,N_2156);
xor U2254 (N_2254,N_2100,N_2153);
and U2255 (N_2255,N_2189,N_2184);
nand U2256 (N_2256,N_2174,N_2185);
or U2257 (N_2257,N_2148,N_2162);
or U2258 (N_2258,N_2127,N_2105);
nor U2259 (N_2259,N_2185,N_2134);
nand U2260 (N_2260,N_2169,N_2199);
or U2261 (N_2261,N_2104,N_2129);
nand U2262 (N_2262,N_2127,N_2115);
and U2263 (N_2263,N_2158,N_2152);
nand U2264 (N_2264,N_2135,N_2155);
nor U2265 (N_2265,N_2180,N_2142);
nor U2266 (N_2266,N_2117,N_2199);
xor U2267 (N_2267,N_2144,N_2123);
and U2268 (N_2268,N_2129,N_2161);
nand U2269 (N_2269,N_2166,N_2152);
and U2270 (N_2270,N_2161,N_2173);
and U2271 (N_2271,N_2187,N_2148);
or U2272 (N_2272,N_2126,N_2163);
nand U2273 (N_2273,N_2195,N_2161);
or U2274 (N_2274,N_2126,N_2156);
xnor U2275 (N_2275,N_2141,N_2109);
nand U2276 (N_2276,N_2176,N_2107);
nand U2277 (N_2277,N_2109,N_2140);
xor U2278 (N_2278,N_2157,N_2196);
nor U2279 (N_2279,N_2133,N_2124);
or U2280 (N_2280,N_2180,N_2175);
nand U2281 (N_2281,N_2121,N_2132);
nand U2282 (N_2282,N_2162,N_2135);
nand U2283 (N_2283,N_2132,N_2188);
nand U2284 (N_2284,N_2141,N_2145);
and U2285 (N_2285,N_2114,N_2128);
or U2286 (N_2286,N_2186,N_2173);
nand U2287 (N_2287,N_2142,N_2155);
and U2288 (N_2288,N_2178,N_2184);
and U2289 (N_2289,N_2184,N_2182);
or U2290 (N_2290,N_2102,N_2118);
or U2291 (N_2291,N_2147,N_2133);
and U2292 (N_2292,N_2142,N_2130);
or U2293 (N_2293,N_2125,N_2128);
nand U2294 (N_2294,N_2164,N_2184);
or U2295 (N_2295,N_2183,N_2173);
or U2296 (N_2296,N_2145,N_2146);
nand U2297 (N_2297,N_2161,N_2184);
nor U2298 (N_2298,N_2153,N_2132);
or U2299 (N_2299,N_2108,N_2186);
xnor U2300 (N_2300,N_2249,N_2201);
or U2301 (N_2301,N_2250,N_2219);
or U2302 (N_2302,N_2266,N_2211);
xor U2303 (N_2303,N_2267,N_2223);
nand U2304 (N_2304,N_2263,N_2280);
nor U2305 (N_2305,N_2256,N_2246);
nand U2306 (N_2306,N_2271,N_2216);
and U2307 (N_2307,N_2214,N_2231);
nor U2308 (N_2308,N_2285,N_2205);
nand U2309 (N_2309,N_2209,N_2255);
or U2310 (N_2310,N_2259,N_2227);
nor U2311 (N_2311,N_2228,N_2282);
nor U2312 (N_2312,N_2253,N_2274);
or U2313 (N_2313,N_2276,N_2208);
nand U2314 (N_2314,N_2203,N_2245);
nor U2315 (N_2315,N_2238,N_2236);
nor U2316 (N_2316,N_2269,N_2233);
or U2317 (N_2317,N_2287,N_2277);
xnor U2318 (N_2318,N_2217,N_2222);
xnor U2319 (N_2319,N_2232,N_2265);
nor U2320 (N_2320,N_2204,N_2237);
or U2321 (N_2321,N_2212,N_2252);
xor U2322 (N_2322,N_2234,N_2299);
and U2323 (N_2323,N_2218,N_2283);
nand U2324 (N_2324,N_2226,N_2296);
and U2325 (N_2325,N_2275,N_2221);
nor U2326 (N_2326,N_2284,N_2294);
nand U2327 (N_2327,N_2220,N_2290);
nor U2328 (N_2328,N_2281,N_2258);
nand U2329 (N_2329,N_2215,N_2210);
nand U2330 (N_2330,N_2279,N_2207);
and U2331 (N_2331,N_2240,N_2261);
and U2332 (N_2332,N_2242,N_2248);
or U2333 (N_2333,N_2298,N_2295);
nor U2334 (N_2334,N_2293,N_2257);
or U2335 (N_2335,N_2254,N_2213);
nor U2336 (N_2336,N_2272,N_2288);
or U2337 (N_2337,N_2264,N_2206);
nand U2338 (N_2338,N_2268,N_2292);
xor U2339 (N_2339,N_2291,N_2260);
nand U2340 (N_2340,N_2244,N_2286);
nand U2341 (N_2341,N_2247,N_2297);
nor U2342 (N_2342,N_2251,N_2202);
nor U2343 (N_2343,N_2235,N_2243);
and U2344 (N_2344,N_2289,N_2225);
and U2345 (N_2345,N_2273,N_2229);
or U2346 (N_2346,N_2200,N_2262);
nand U2347 (N_2347,N_2230,N_2224);
nor U2348 (N_2348,N_2239,N_2270);
nor U2349 (N_2349,N_2278,N_2241);
and U2350 (N_2350,N_2298,N_2203);
and U2351 (N_2351,N_2243,N_2232);
and U2352 (N_2352,N_2276,N_2284);
nand U2353 (N_2353,N_2217,N_2278);
nand U2354 (N_2354,N_2235,N_2223);
xor U2355 (N_2355,N_2281,N_2269);
or U2356 (N_2356,N_2292,N_2234);
nand U2357 (N_2357,N_2203,N_2219);
nand U2358 (N_2358,N_2201,N_2214);
or U2359 (N_2359,N_2219,N_2225);
or U2360 (N_2360,N_2298,N_2270);
and U2361 (N_2361,N_2257,N_2296);
nor U2362 (N_2362,N_2275,N_2220);
and U2363 (N_2363,N_2226,N_2212);
or U2364 (N_2364,N_2294,N_2286);
and U2365 (N_2365,N_2200,N_2261);
and U2366 (N_2366,N_2228,N_2276);
xnor U2367 (N_2367,N_2241,N_2225);
nand U2368 (N_2368,N_2297,N_2268);
nand U2369 (N_2369,N_2226,N_2208);
and U2370 (N_2370,N_2209,N_2298);
nand U2371 (N_2371,N_2238,N_2273);
nand U2372 (N_2372,N_2265,N_2240);
nand U2373 (N_2373,N_2256,N_2213);
and U2374 (N_2374,N_2204,N_2241);
nand U2375 (N_2375,N_2230,N_2264);
or U2376 (N_2376,N_2238,N_2217);
and U2377 (N_2377,N_2274,N_2294);
or U2378 (N_2378,N_2220,N_2297);
nor U2379 (N_2379,N_2280,N_2214);
nor U2380 (N_2380,N_2237,N_2241);
nand U2381 (N_2381,N_2283,N_2254);
nor U2382 (N_2382,N_2283,N_2214);
nand U2383 (N_2383,N_2237,N_2278);
nand U2384 (N_2384,N_2256,N_2250);
and U2385 (N_2385,N_2288,N_2279);
nor U2386 (N_2386,N_2230,N_2227);
or U2387 (N_2387,N_2298,N_2223);
nor U2388 (N_2388,N_2217,N_2205);
nor U2389 (N_2389,N_2221,N_2243);
and U2390 (N_2390,N_2240,N_2248);
or U2391 (N_2391,N_2264,N_2284);
nor U2392 (N_2392,N_2293,N_2279);
or U2393 (N_2393,N_2283,N_2266);
nand U2394 (N_2394,N_2223,N_2276);
and U2395 (N_2395,N_2213,N_2253);
or U2396 (N_2396,N_2252,N_2220);
nand U2397 (N_2397,N_2274,N_2273);
nand U2398 (N_2398,N_2265,N_2201);
or U2399 (N_2399,N_2287,N_2283);
and U2400 (N_2400,N_2305,N_2376);
and U2401 (N_2401,N_2380,N_2360);
nor U2402 (N_2402,N_2377,N_2372);
nand U2403 (N_2403,N_2317,N_2398);
nand U2404 (N_2404,N_2321,N_2378);
xnor U2405 (N_2405,N_2311,N_2396);
nand U2406 (N_2406,N_2339,N_2327);
and U2407 (N_2407,N_2385,N_2322);
nand U2408 (N_2408,N_2307,N_2346);
nor U2409 (N_2409,N_2375,N_2309);
and U2410 (N_2410,N_2394,N_2314);
and U2411 (N_2411,N_2369,N_2325);
and U2412 (N_2412,N_2323,N_2333);
or U2413 (N_2413,N_2379,N_2355);
or U2414 (N_2414,N_2395,N_2340);
nor U2415 (N_2415,N_2342,N_2338);
nand U2416 (N_2416,N_2310,N_2370);
nor U2417 (N_2417,N_2303,N_2374);
xnor U2418 (N_2418,N_2387,N_2391);
nor U2419 (N_2419,N_2330,N_2332);
or U2420 (N_2420,N_2383,N_2359);
nand U2421 (N_2421,N_2337,N_2357);
nand U2422 (N_2422,N_2354,N_2329);
nand U2423 (N_2423,N_2366,N_2368);
xnor U2424 (N_2424,N_2353,N_2304);
and U2425 (N_2425,N_2324,N_2386);
or U2426 (N_2426,N_2356,N_2318);
or U2427 (N_2427,N_2364,N_2300);
or U2428 (N_2428,N_2336,N_2328);
and U2429 (N_2429,N_2381,N_2331);
nand U2430 (N_2430,N_2313,N_2393);
nand U2431 (N_2431,N_2345,N_2341);
or U2432 (N_2432,N_2349,N_2358);
nor U2433 (N_2433,N_2308,N_2388);
nand U2434 (N_2434,N_2367,N_2389);
and U2435 (N_2435,N_2326,N_2397);
nand U2436 (N_2436,N_2363,N_2352);
nand U2437 (N_2437,N_2351,N_2350);
nor U2438 (N_2438,N_2392,N_2371);
nor U2439 (N_2439,N_2348,N_2320);
or U2440 (N_2440,N_2302,N_2312);
nand U2441 (N_2441,N_2315,N_2343);
or U2442 (N_2442,N_2390,N_2334);
or U2443 (N_2443,N_2382,N_2365);
and U2444 (N_2444,N_2373,N_2306);
and U2445 (N_2445,N_2384,N_2347);
and U2446 (N_2446,N_2344,N_2362);
and U2447 (N_2447,N_2361,N_2316);
and U2448 (N_2448,N_2335,N_2399);
xor U2449 (N_2449,N_2301,N_2319);
or U2450 (N_2450,N_2308,N_2319);
nor U2451 (N_2451,N_2334,N_2358);
and U2452 (N_2452,N_2337,N_2323);
or U2453 (N_2453,N_2380,N_2344);
and U2454 (N_2454,N_2333,N_2388);
nand U2455 (N_2455,N_2320,N_2398);
nand U2456 (N_2456,N_2395,N_2386);
nand U2457 (N_2457,N_2373,N_2391);
or U2458 (N_2458,N_2341,N_2336);
and U2459 (N_2459,N_2305,N_2390);
and U2460 (N_2460,N_2372,N_2341);
nand U2461 (N_2461,N_2314,N_2365);
and U2462 (N_2462,N_2313,N_2349);
xor U2463 (N_2463,N_2376,N_2383);
nand U2464 (N_2464,N_2335,N_2322);
nor U2465 (N_2465,N_2371,N_2304);
or U2466 (N_2466,N_2367,N_2388);
or U2467 (N_2467,N_2365,N_2388);
nand U2468 (N_2468,N_2326,N_2340);
or U2469 (N_2469,N_2309,N_2306);
or U2470 (N_2470,N_2302,N_2387);
and U2471 (N_2471,N_2396,N_2368);
xnor U2472 (N_2472,N_2314,N_2334);
nor U2473 (N_2473,N_2358,N_2361);
nand U2474 (N_2474,N_2309,N_2397);
or U2475 (N_2475,N_2336,N_2392);
xnor U2476 (N_2476,N_2311,N_2383);
nor U2477 (N_2477,N_2354,N_2361);
nor U2478 (N_2478,N_2310,N_2356);
or U2479 (N_2479,N_2377,N_2368);
nand U2480 (N_2480,N_2309,N_2390);
nor U2481 (N_2481,N_2333,N_2391);
and U2482 (N_2482,N_2356,N_2312);
nand U2483 (N_2483,N_2310,N_2364);
nor U2484 (N_2484,N_2397,N_2360);
xnor U2485 (N_2485,N_2334,N_2348);
nand U2486 (N_2486,N_2355,N_2301);
and U2487 (N_2487,N_2312,N_2392);
or U2488 (N_2488,N_2393,N_2330);
or U2489 (N_2489,N_2375,N_2359);
nand U2490 (N_2490,N_2302,N_2360);
nand U2491 (N_2491,N_2328,N_2357);
nor U2492 (N_2492,N_2371,N_2322);
nor U2493 (N_2493,N_2314,N_2333);
nor U2494 (N_2494,N_2349,N_2363);
and U2495 (N_2495,N_2323,N_2365);
nand U2496 (N_2496,N_2357,N_2386);
nand U2497 (N_2497,N_2384,N_2353);
nor U2498 (N_2498,N_2376,N_2382);
and U2499 (N_2499,N_2331,N_2306);
xor U2500 (N_2500,N_2482,N_2432);
or U2501 (N_2501,N_2444,N_2448);
or U2502 (N_2502,N_2400,N_2468);
and U2503 (N_2503,N_2481,N_2409);
and U2504 (N_2504,N_2424,N_2405);
nor U2505 (N_2505,N_2423,N_2492);
nand U2506 (N_2506,N_2494,N_2415);
nor U2507 (N_2507,N_2490,N_2437);
or U2508 (N_2508,N_2493,N_2410);
nor U2509 (N_2509,N_2429,N_2473);
nor U2510 (N_2510,N_2412,N_2440);
nand U2511 (N_2511,N_2485,N_2469);
nand U2512 (N_2512,N_2497,N_2445);
nand U2513 (N_2513,N_2470,N_2438);
and U2514 (N_2514,N_2406,N_2430);
xor U2515 (N_2515,N_2403,N_2461);
nor U2516 (N_2516,N_2465,N_2498);
or U2517 (N_2517,N_2407,N_2420);
nor U2518 (N_2518,N_2427,N_2466);
xor U2519 (N_2519,N_2446,N_2483);
or U2520 (N_2520,N_2433,N_2480);
or U2521 (N_2521,N_2453,N_2435);
and U2522 (N_2522,N_2431,N_2477);
or U2523 (N_2523,N_2411,N_2404);
nor U2524 (N_2524,N_2428,N_2458);
xnor U2525 (N_2525,N_2455,N_2489);
or U2526 (N_2526,N_2499,N_2422);
or U2527 (N_2527,N_2441,N_2421);
or U2528 (N_2528,N_2476,N_2450);
nand U2529 (N_2529,N_2449,N_2439);
or U2530 (N_2530,N_2401,N_2462);
nand U2531 (N_2531,N_2426,N_2447);
or U2532 (N_2532,N_2459,N_2484);
and U2533 (N_2533,N_2475,N_2495);
xnor U2534 (N_2534,N_2425,N_2436);
xor U2535 (N_2535,N_2467,N_2402);
nor U2536 (N_2536,N_2488,N_2418);
nor U2537 (N_2537,N_2454,N_2434);
nand U2538 (N_2538,N_2416,N_2442);
xor U2539 (N_2539,N_2463,N_2471);
nand U2540 (N_2540,N_2472,N_2478);
or U2541 (N_2541,N_2419,N_2487);
nand U2542 (N_2542,N_2460,N_2486);
nor U2543 (N_2543,N_2413,N_2417);
and U2544 (N_2544,N_2479,N_2496);
xnor U2545 (N_2545,N_2451,N_2491);
nand U2546 (N_2546,N_2457,N_2414);
and U2547 (N_2547,N_2452,N_2456);
xnor U2548 (N_2548,N_2443,N_2464);
nand U2549 (N_2549,N_2408,N_2474);
nand U2550 (N_2550,N_2489,N_2457);
and U2551 (N_2551,N_2448,N_2426);
xor U2552 (N_2552,N_2403,N_2453);
and U2553 (N_2553,N_2472,N_2480);
or U2554 (N_2554,N_2479,N_2494);
xor U2555 (N_2555,N_2407,N_2411);
nor U2556 (N_2556,N_2427,N_2407);
or U2557 (N_2557,N_2483,N_2485);
and U2558 (N_2558,N_2495,N_2419);
nor U2559 (N_2559,N_2409,N_2485);
nand U2560 (N_2560,N_2499,N_2431);
and U2561 (N_2561,N_2494,N_2463);
and U2562 (N_2562,N_2443,N_2441);
nor U2563 (N_2563,N_2411,N_2425);
xor U2564 (N_2564,N_2445,N_2488);
and U2565 (N_2565,N_2499,N_2434);
and U2566 (N_2566,N_2480,N_2481);
or U2567 (N_2567,N_2451,N_2422);
and U2568 (N_2568,N_2499,N_2426);
and U2569 (N_2569,N_2482,N_2483);
nand U2570 (N_2570,N_2440,N_2490);
nand U2571 (N_2571,N_2451,N_2445);
nand U2572 (N_2572,N_2440,N_2472);
and U2573 (N_2573,N_2424,N_2403);
xnor U2574 (N_2574,N_2459,N_2469);
nor U2575 (N_2575,N_2467,N_2406);
nand U2576 (N_2576,N_2486,N_2421);
nor U2577 (N_2577,N_2405,N_2414);
nor U2578 (N_2578,N_2466,N_2425);
nand U2579 (N_2579,N_2452,N_2454);
nor U2580 (N_2580,N_2421,N_2419);
and U2581 (N_2581,N_2484,N_2431);
nand U2582 (N_2582,N_2419,N_2452);
xor U2583 (N_2583,N_2414,N_2402);
and U2584 (N_2584,N_2428,N_2465);
nor U2585 (N_2585,N_2461,N_2428);
nand U2586 (N_2586,N_2439,N_2452);
and U2587 (N_2587,N_2480,N_2462);
nand U2588 (N_2588,N_2441,N_2492);
and U2589 (N_2589,N_2402,N_2421);
or U2590 (N_2590,N_2449,N_2414);
nor U2591 (N_2591,N_2430,N_2464);
nor U2592 (N_2592,N_2403,N_2428);
nand U2593 (N_2593,N_2491,N_2408);
and U2594 (N_2594,N_2474,N_2424);
or U2595 (N_2595,N_2487,N_2499);
nor U2596 (N_2596,N_2483,N_2408);
and U2597 (N_2597,N_2481,N_2442);
nand U2598 (N_2598,N_2474,N_2496);
and U2599 (N_2599,N_2471,N_2435);
nor U2600 (N_2600,N_2552,N_2503);
xor U2601 (N_2601,N_2570,N_2587);
nand U2602 (N_2602,N_2546,N_2512);
xor U2603 (N_2603,N_2586,N_2539);
xnor U2604 (N_2604,N_2514,N_2515);
nand U2605 (N_2605,N_2519,N_2589);
or U2606 (N_2606,N_2553,N_2581);
and U2607 (N_2607,N_2534,N_2579);
or U2608 (N_2608,N_2599,N_2598);
nor U2609 (N_2609,N_2595,N_2524);
and U2610 (N_2610,N_2569,N_2506);
or U2611 (N_2611,N_2535,N_2572);
nand U2612 (N_2612,N_2583,N_2510);
nor U2613 (N_2613,N_2543,N_2558);
nand U2614 (N_2614,N_2555,N_2544);
nor U2615 (N_2615,N_2550,N_2588);
and U2616 (N_2616,N_2575,N_2525);
nor U2617 (N_2617,N_2590,N_2574);
nor U2618 (N_2618,N_2585,N_2560);
nand U2619 (N_2619,N_2541,N_2573);
nand U2620 (N_2620,N_2542,N_2520);
and U2621 (N_2621,N_2549,N_2532);
or U2622 (N_2622,N_2538,N_2571);
nand U2623 (N_2623,N_2566,N_2513);
nand U2624 (N_2624,N_2511,N_2540);
nor U2625 (N_2625,N_2531,N_2580);
nor U2626 (N_2626,N_2527,N_2518);
and U2627 (N_2627,N_2530,N_2556);
and U2628 (N_2628,N_2576,N_2567);
nand U2629 (N_2629,N_2536,N_2521);
xnor U2630 (N_2630,N_2596,N_2529);
nor U2631 (N_2631,N_2562,N_2507);
and U2632 (N_2632,N_2509,N_2578);
nand U2633 (N_2633,N_2508,N_2548);
nand U2634 (N_2634,N_2577,N_2593);
nand U2635 (N_2635,N_2504,N_2505);
nor U2636 (N_2636,N_2528,N_2582);
nand U2637 (N_2637,N_2537,N_2554);
or U2638 (N_2638,N_2522,N_2559);
nor U2639 (N_2639,N_2551,N_2533);
or U2640 (N_2640,N_2502,N_2501);
and U2641 (N_2641,N_2547,N_2584);
nor U2642 (N_2642,N_2517,N_2516);
and U2643 (N_2643,N_2545,N_2597);
nand U2644 (N_2644,N_2568,N_2565);
nand U2645 (N_2645,N_2526,N_2557);
or U2646 (N_2646,N_2564,N_2563);
nand U2647 (N_2647,N_2594,N_2523);
nor U2648 (N_2648,N_2500,N_2561);
or U2649 (N_2649,N_2592,N_2591);
xnor U2650 (N_2650,N_2531,N_2570);
or U2651 (N_2651,N_2526,N_2511);
and U2652 (N_2652,N_2500,N_2521);
or U2653 (N_2653,N_2578,N_2530);
and U2654 (N_2654,N_2567,N_2538);
nor U2655 (N_2655,N_2507,N_2567);
or U2656 (N_2656,N_2588,N_2558);
nor U2657 (N_2657,N_2515,N_2569);
nand U2658 (N_2658,N_2584,N_2538);
nor U2659 (N_2659,N_2501,N_2520);
and U2660 (N_2660,N_2533,N_2528);
nor U2661 (N_2661,N_2548,N_2507);
nor U2662 (N_2662,N_2571,N_2566);
xnor U2663 (N_2663,N_2529,N_2579);
nand U2664 (N_2664,N_2509,N_2534);
nand U2665 (N_2665,N_2544,N_2573);
nand U2666 (N_2666,N_2565,N_2578);
or U2667 (N_2667,N_2546,N_2538);
nor U2668 (N_2668,N_2584,N_2589);
nand U2669 (N_2669,N_2579,N_2524);
or U2670 (N_2670,N_2568,N_2552);
and U2671 (N_2671,N_2535,N_2532);
or U2672 (N_2672,N_2529,N_2587);
xor U2673 (N_2673,N_2555,N_2511);
nor U2674 (N_2674,N_2587,N_2537);
nor U2675 (N_2675,N_2543,N_2539);
or U2676 (N_2676,N_2545,N_2574);
or U2677 (N_2677,N_2562,N_2599);
nand U2678 (N_2678,N_2555,N_2599);
nor U2679 (N_2679,N_2503,N_2580);
xnor U2680 (N_2680,N_2519,N_2590);
or U2681 (N_2681,N_2567,N_2591);
or U2682 (N_2682,N_2558,N_2538);
or U2683 (N_2683,N_2569,N_2535);
and U2684 (N_2684,N_2556,N_2594);
nand U2685 (N_2685,N_2528,N_2566);
nand U2686 (N_2686,N_2536,N_2538);
nand U2687 (N_2687,N_2531,N_2525);
nand U2688 (N_2688,N_2597,N_2523);
and U2689 (N_2689,N_2562,N_2559);
or U2690 (N_2690,N_2506,N_2560);
nand U2691 (N_2691,N_2556,N_2558);
and U2692 (N_2692,N_2570,N_2542);
xor U2693 (N_2693,N_2573,N_2566);
or U2694 (N_2694,N_2588,N_2522);
nor U2695 (N_2695,N_2548,N_2523);
nor U2696 (N_2696,N_2516,N_2572);
and U2697 (N_2697,N_2589,N_2570);
and U2698 (N_2698,N_2545,N_2520);
nand U2699 (N_2699,N_2534,N_2561);
nor U2700 (N_2700,N_2679,N_2696);
or U2701 (N_2701,N_2693,N_2653);
nand U2702 (N_2702,N_2612,N_2688);
nor U2703 (N_2703,N_2623,N_2644);
or U2704 (N_2704,N_2607,N_2656);
or U2705 (N_2705,N_2637,N_2662);
nor U2706 (N_2706,N_2604,N_2677);
nor U2707 (N_2707,N_2647,N_2622);
nand U2708 (N_2708,N_2699,N_2632);
and U2709 (N_2709,N_2617,N_2620);
nor U2710 (N_2710,N_2673,N_2659);
nand U2711 (N_2711,N_2651,N_2621);
or U2712 (N_2712,N_2675,N_2639);
nand U2713 (N_2713,N_2667,N_2600);
and U2714 (N_2714,N_2697,N_2650);
nand U2715 (N_2715,N_2661,N_2618);
and U2716 (N_2716,N_2641,N_2692);
nand U2717 (N_2717,N_2642,N_2648);
nand U2718 (N_2718,N_2646,N_2689);
or U2719 (N_2719,N_2624,N_2601);
nand U2720 (N_2720,N_2672,N_2665);
xor U2721 (N_2721,N_2669,N_2640);
and U2722 (N_2722,N_2671,N_2678);
and U2723 (N_2723,N_2652,N_2603);
and U2724 (N_2724,N_2638,N_2691);
nand U2725 (N_2725,N_2683,N_2660);
nor U2726 (N_2726,N_2611,N_2694);
nor U2727 (N_2727,N_2626,N_2666);
or U2728 (N_2728,N_2664,N_2629);
and U2729 (N_2729,N_2663,N_2627);
nor U2730 (N_2730,N_2645,N_2610);
nor U2731 (N_2731,N_2606,N_2628);
nand U2732 (N_2732,N_2630,N_2636);
nor U2733 (N_2733,N_2658,N_2643);
or U2734 (N_2734,N_2605,N_2619);
nand U2735 (N_2735,N_2614,N_2690);
or U2736 (N_2736,N_2657,N_2686);
xnor U2737 (N_2737,N_2616,N_2634);
and U2738 (N_2738,N_2615,N_2684);
and U2739 (N_2739,N_2698,N_2635);
or U2740 (N_2740,N_2654,N_2674);
nand U2741 (N_2741,N_2633,N_2682);
nand U2742 (N_2742,N_2655,N_2608);
nand U2743 (N_2743,N_2609,N_2685);
nand U2744 (N_2744,N_2625,N_2602);
nor U2745 (N_2745,N_2631,N_2687);
and U2746 (N_2746,N_2681,N_2649);
xnor U2747 (N_2747,N_2676,N_2680);
and U2748 (N_2748,N_2695,N_2670);
nor U2749 (N_2749,N_2613,N_2668);
or U2750 (N_2750,N_2619,N_2674);
or U2751 (N_2751,N_2660,N_2666);
or U2752 (N_2752,N_2605,N_2667);
xor U2753 (N_2753,N_2680,N_2696);
nand U2754 (N_2754,N_2636,N_2606);
and U2755 (N_2755,N_2668,N_2626);
and U2756 (N_2756,N_2621,N_2682);
nor U2757 (N_2757,N_2669,N_2663);
xnor U2758 (N_2758,N_2652,N_2606);
nand U2759 (N_2759,N_2617,N_2649);
and U2760 (N_2760,N_2631,N_2645);
and U2761 (N_2761,N_2630,N_2692);
nand U2762 (N_2762,N_2695,N_2646);
nor U2763 (N_2763,N_2677,N_2643);
nand U2764 (N_2764,N_2690,N_2624);
nor U2765 (N_2765,N_2669,N_2642);
or U2766 (N_2766,N_2626,N_2607);
and U2767 (N_2767,N_2645,N_2650);
and U2768 (N_2768,N_2680,N_2671);
nor U2769 (N_2769,N_2666,N_2608);
or U2770 (N_2770,N_2647,N_2600);
or U2771 (N_2771,N_2644,N_2613);
or U2772 (N_2772,N_2652,N_2620);
and U2773 (N_2773,N_2673,N_2625);
and U2774 (N_2774,N_2614,N_2605);
or U2775 (N_2775,N_2628,N_2685);
nor U2776 (N_2776,N_2680,N_2689);
and U2777 (N_2777,N_2630,N_2656);
or U2778 (N_2778,N_2620,N_2690);
and U2779 (N_2779,N_2663,N_2633);
or U2780 (N_2780,N_2612,N_2686);
nor U2781 (N_2781,N_2635,N_2634);
nand U2782 (N_2782,N_2670,N_2667);
or U2783 (N_2783,N_2602,N_2636);
nand U2784 (N_2784,N_2699,N_2609);
xor U2785 (N_2785,N_2613,N_2647);
or U2786 (N_2786,N_2689,N_2634);
nand U2787 (N_2787,N_2677,N_2629);
nor U2788 (N_2788,N_2602,N_2656);
and U2789 (N_2789,N_2624,N_2609);
nor U2790 (N_2790,N_2685,N_2637);
nor U2791 (N_2791,N_2600,N_2648);
nor U2792 (N_2792,N_2623,N_2630);
and U2793 (N_2793,N_2652,N_2650);
xnor U2794 (N_2794,N_2670,N_2637);
and U2795 (N_2795,N_2646,N_2606);
nand U2796 (N_2796,N_2698,N_2659);
xnor U2797 (N_2797,N_2675,N_2600);
and U2798 (N_2798,N_2610,N_2666);
or U2799 (N_2799,N_2664,N_2602);
and U2800 (N_2800,N_2760,N_2762);
and U2801 (N_2801,N_2758,N_2785);
nand U2802 (N_2802,N_2753,N_2712);
nor U2803 (N_2803,N_2771,N_2797);
nand U2804 (N_2804,N_2734,N_2798);
and U2805 (N_2805,N_2763,N_2786);
nor U2806 (N_2806,N_2755,N_2759);
nor U2807 (N_2807,N_2701,N_2775);
nand U2808 (N_2808,N_2793,N_2714);
and U2809 (N_2809,N_2750,N_2710);
or U2810 (N_2810,N_2732,N_2756);
nand U2811 (N_2811,N_2757,N_2720);
and U2812 (N_2812,N_2707,N_2725);
or U2813 (N_2813,N_2799,N_2796);
nand U2814 (N_2814,N_2746,N_2767);
and U2815 (N_2815,N_2773,N_2719);
xnor U2816 (N_2816,N_2791,N_2702);
nand U2817 (N_2817,N_2741,N_2718);
nor U2818 (N_2818,N_2735,N_2772);
or U2819 (N_2819,N_2788,N_2742);
nor U2820 (N_2820,N_2781,N_2715);
or U2821 (N_2821,N_2787,N_2790);
and U2822 (N_2822,N_2784,N_2739);
nor U2823 (N_2823,N_2737,N_2754);
nand U2824 (N_2824,N_2726,N_2795);
nand U2825 (N_2825,N_2709,N_2708);
and U2826 (N_2826,N_2764,N_2700);
nand U2827 (N_2827,N_2776,N_2778);
nand U2828 (N_2828,N_2711,N_2722);
or U2829 (N_2829,N_2706,N_2769);
xnor U2830 (N_2830,N_2723,N_2713);
nor U2831 (N_2831,N_2752,N_2724);
and U2832 (N_2832,N_2727,N_2731);
nand U2833 (N_2833,N_2703,N_2738);
and U2834 (N_2834,N_2749,N_2733);
and U2835 (N_2835,N_2751,N_2747);
nand U2836 (N_2836,N_2770,N_2744);
xnor U2837 (N_2837,N_2716,N_2774);
nor U2838 (N_2838,N_2782,N_2777);
or U2839 (N_2839,N_2704,N_2766);
nand U2840 (N_2840,N_2765,N_2780);
or U2841 (N_2841,N_2768,N_2728);
nor U2842 (N_2842,N_2736,N_2705);
xor U2843 (N_2843,N_2783,N_2748);
nand U2844 (N_2844,N_2717,N_2779);
or U2845 (N_2845,N_2745,N_2761);
nor U2846 (N_2846,N_2740,N_2730);
and U2847 (N_2847,N_2794,N_2789);
or U2848 (N_2848,N_2729,N_2743);
and U2849 (N_2849,N_2792,N_2721);
nand U2850 (N_2850,N_2749,N_2751);
nor U2851 (N_2851,N_2748,N_2746);
nor U2852 (N_2852,N_2783,N_2752);
nor U2853 (N_2853,N_2785,N_2782);
nand U2854 (N_2854,N_2731,N_2763);
nand U2855 (N_2855,N_2701,N_2768);
or U2856 (N_2856,N_2723,N_2792);
or U2857 (N_2857,N_2752,N_2743);
or U2858 (N_2858,N_2746,N_2765);
nor U2859 (N_2859,N_2774,N_2749);
and U2860 (N_2860,N_2720,N_2790);
nand U2861 (N_2861,N_2731,N_2783);
or U2862 (N_2862,N_2730,N_2710);
and U2863 (N_2863,N_2798,N_2711);
or U2864 (N_2864,N_2793,N_2775);
xnor U2865 (N_2865,N_2785,N_2733);
and U2866 (N_2866,N_2774,N_2768);
and U2867 (N_2867,N_2783,N_2779);
nand U2868 (N_2868,N_2790,N_2736);
and U2869 (N_2869,N_2797,N_2796);
nand U2870 (N_2870,N_2729,N_2711);
nor U2871 (N_2871,N_2753,N_2720);
xor U2872 (N_2872,N_2767,N_2723);
or U2873 (N_2873,N_2791,N_2778);
nor U2874 (N_2874,N_2743,N_2757);
nand U2875 (N_2875,N_2746,N_2783);
nand U2876 (N_2876,N_2773,N_2748);
or U2877 (N_2877,N_2761,N_2752);
or U2878 (N_2878,N_2775,N_2758);
or U2879 (N_2879,N_2783,N_2736);
or U2880 (N_2880,N_2790,N_2746);
and U2881 (N_2881,N_2708,N_2726);
nor U2882 (N_2882,N_2768,N_2789);
xor U2883 (N_2883,N_2737,N_2783);
nor U2884 (N_2884,N_2708,N_2735);
nor U2885 (N_2885,N_2710,N_2772);
nand U2886 (N_2886,N_2756,N_2785);
or U2887 (N_2887,N_2776,N_2713);
nor U2888 (N_2888,N_2745,N_2768);
nor U2889 (N_2889,N_2750,N_2759);
and U2890 (N_2890,N_2782,N_2704);
nand U2891 (N_2891,N_2765,N_2723);
and U2892 (N_2892,N_2707,N_2743);
and U2893 (N_2893,N_2765,N_2700);
or U2894 (N_2894,N_2761,N_2764);
xor U2895 (N_2895,N_2738,N_2736);
nor U2896 (N_2896,N_2705,N_2762);
nor U2897 (N_2897,N_2749,N_2760);
nand U2898 (N_2898,N_2755,N_2763);
and U2899 (N_2899,N_2714,N_2792);
nor U2900 (N_2900,N_2891,N_2850);
nand U2901 (N_2901,N_2807,N_2826);
or U2902 (N_2902,N_2866,N_2842);
or U2903 (N_2903,N_2887,N_2893);
nor U2904 (N_2904,N_2867,N_2897);
xnor U2905 (N_2905,N_2881,N_2809);
nor U2906 (N_2906,N_2864,N_2834);
xor U2907 (N_2907,N_2831,N_2824);
nor U2908 (N_2908,N_2840,N_2833);
nor U2909 (N_2909,N_2859,N_2822);
and U2910 (N_2910,N_2878,N_2839);
xor U2911 (N_2911,N_2821,N_2841);
nor U2912 (N_2912,N_2877,N_2800);
and U2913 (N_2913,N_2894,N_2813);
xnor U2914 (N_2914,N_2882,N_2848);
or U2915 (N_2915,N_2883,N_2898);
nand U2916 (N_2916,N_2836,N_2804);
xor U2917 (N_2917,N_2846,N_2817);
or U2918 (N_2918,N_2869,N_2827);
and U2919 (N_2919,N_2829,N_2858);
or U2920 (N_2920,N_2851,N_2828);
xnor U2921 (N_2921,N_2844,N_2899);
nor U2922 (N_2922,N_2888,N_2847);
nand U2923 (N_2923,N_2884,N_2806);
and U2924 (N_2924,N_2820,N_2870);
nand U2925 (N_2925,N_2805,N_2879);
or U2926 (N_2926,N_2819,N_2808);
nor U2927 (N_2927,N_2886,N_2815);
or U2928 (N_2928,N_2873,N_2801);
nor U2929 (N_2929,N_2843,N_2861);
or U2930 (N_2930,N_2832,N_2863);
nand U2931 (N_2931,N_2852,N_2890);
or U2932 (N_2932,N_2857,N_2854);
xor U2933 (N_2933,N_2811,N_2835);
or U2934 (N_2934,N_2872,N_2868);
or U2935 (N_2935,N_2856,N_2849);
nor U2936 (N_2936,N_2892,N_2895);
or U2937 (N_2937,N_2896,N_2860);
nor U2938 (N_2938,N_2889,N_2802);
nor U2939 (N_2939,N_2838,N_2830);
or U2940 (N_2940,N_2816,N_2825);
xor U2941 (N_2941,N_2874,N_2810);
or U2942 (N_2942,N_2814,N_2812);
and U2943 (N_2943,N_2855,N_2885);
or U2944 (N_2944,N_2862,N_2880);
nand U2945 (N_2945,N_2853,N_2845);
nand U2946 (N_2946,N_2871,N_2818);
nand U2947 (N_2947,N_2876,N_2803);
nor U2948 (N_2948,N_2865,N_2823);
and U2949 (N_2949,N_2837,N_2875);
nor U2950 (N_2950,N_2828,N_2872);
and U2951 (N_2951,N_2873,N_2847);
nor U2952 (N_2952,N_2826,N_2853);
or U2953 (N_2953,N_2849,N_2853);
or U2954 (N_2954,N_2801,N_2881);
and U2955 (N_2955,N_2876,N_2811);
and U2956 (N_2956,N_2870,N_2882);
nor U2957 (N_2957,N_2819,N_2890);
nand U2958 (N_2958,N_2809,N_2898);
or U2959 (N_2959,N_2893,N_2820);
nand U2960 (N_2960,N_2832,N_2883);
or U2961 (N_2961,N_2806,N_2858);
xnor U2962 (N_2962,N_2863,N_2888);
nand U2963 (N_2963,N_2861,N_2850);
or U2964 (N_2964,N_2816,N_2801);
or U2965 (N_2965,N_2885,N_2816);
and U2966 (N_2966,N_2828,N_2827);
and U2967 (N_2967,N_2826,N_2837);
xor U2968 (N_2968,N_2836,N_2824);
nand U2969 (N_2969,N_2869,N_2862);
nand U2970 (N_2970,N_2815,N_2892);
nand U2971 (N_2971,N_2839,N_2805);
xor U2972 (N_2972,N_2899,N_2891);
or U2973 (N_2973,N_2820,N_2832);
nand U2974 (N_2974,N_2880,N_2871);
or U2975 (N_2975,N_2838,N_2858);
nor U2976 (N_2976,N_2817,N_2855);
nor U2977 (N_2977,N_2800,N_2899);
or U2978 (N_2978,N_2853,N_2883);
nor U2979 (N_2979,N_2852,N_2889);
nand U2980 (N_2980,N_2805,N_2847);
nand U2981 (N_2981,N_2846,N_2894);
xor U2982 (N_2982,N_2810,N_2853);
and U2983 (N_2983,N_2890,N_2822);
and U2984 (N_2984,N_2854,N_2851);
or U2985 (N_2985,N_2870,N_2874);
nand U2986 (N_2986,N_2866,N_2863);
nor U2987 (N_2987,N_2868,N_2809);
xor U2988 (N_2988,N_2863,N_2891);
nand U2989 (N_2989,N_2868,N_2834);
or U2990 (N_2990,N_2839,N_2802);
or U2991 (N_2991,N_2833,N_2881);
and U2992 (N_2992,N_2883,N_2819);
nand U2993 (N_2993,N_2846,N_2857);
and U2994 (N_2994,N_2813,N_2805);
nand U2995 (N_2995,N_2803,N_2810);
and U2996 (N_2996,N_2872,N_2852);
xnor U2997 (N_2997,N_2881,N_2880);
xor U2998 (N_2998,N_2882,N_2825);
nand U2999 (N_2999,N_2896,N_2861);
nor UO_0 (O_0,N_2924,N_2963);
or UO_1 (O_1,N_2900,N_2960);
xor UO_2 (O_2,N_2983,N_2946);
nor UO_3 (O_3,N_2987,N_2942);
and UO_4 (O_4,N_2955,N_2927);
nand UO_5 (O_5,N_2976,N_2947);
nand UO_6 (O_6,N_2902,N_2934);
nor UO_7 (O_7,N_2998,N_2923);
nor UO_8 (O_8,N_2919,N_2977);
nor UO_9 (O_9,N_2995,N_2954);
nor UO_10 (O_10,N_2958,N_2997);
nand UO_11 (O_11,N_2922,N_2916);
or UO_12 (O_12,N_2933,N_2961);
nor UO_13 (O_13,N_2968,N_2910);
nor UO_14 (O_14,N_2921,N_2966);
and UO_15 (O_15,N_2974,N_2912);
nor UO_16 (O_16,N_2932,N_2979);
nand UO_17 (O_17,N_2957,N_2937);
xnor UO_18 (O_18,N_2973,N_2986);
nand UO_19 (O_19,N_2980,N_2972);
or UO_20 (O_20,N_2956,N_2920);
xnor UO_21 (O_21,N_2925,N_2944);
nor UO_22 (O_22,N_2943,N_2905);
or UO_23 (O_23,N_2938,N_2996);
xor UO_24 (O_24,N_2988,N_2964);
or UO_25 (O_25,N_2930,N_2978);
and UO_26 (O_26,N_2911,N_2941);
nand UO_27 (O_27,N_2909,N_2953);
or UO_28 (O_28,N_2904,N_2940);
nor UO_29 (O_29,N_2949,N_2907);
or UO_30 (O_30,N_2906,N_2982);
and UO_31 (O_31,N_2929,N_2975);
xor UO_32 (O_32,N_2948,N_2994);
or UO_33 (O_33,N_2962,N_2965);
nand UO_34 (O_34,N_2926,N_2991);
nor UO_35 (O_35,N_2928,N_2989);
or UO_36 (O_36,N_2993,N_2914);
nand UO_37 (O_37,N_2945,N_2915);
or UO_38 (O_38,N_2903,N_2918);
and UO_39 (O_39,N_2913,N_2939);
nor UO_40 (O_40,N_2952,N_2985);
or UO_41 (O_41,N_2931,N_2967);
and UO_42 (O_42,N_2969,N_2970);
or UO_43 (O_43,N_2959,N_2951);
and UO_44 (O_44,N_2917,N_2936);
nand UO_45 (O_45,N_2950,N_2971);
nand UO_46 (O_46,N_2935,N_2901);
nand UO_47 (O_47,N_2999,N_2992);
or UO_48 (O_48,N_2984,N_2990);
nor UO_49 (O_49,N_2908,N_2981);
or UO_50 (O_50,N_2966,N_2999);
nand UO_51 (O_51,N_2903,N_2905);
nor UO_52 (O_52,N_2973,N_2958);
or UO_53 (O_53,N_2936,N_2979);
nor UO_54 (O_54,N_2942,N_2903);
or UO_55 (O_55,N_2932,N_2947);
nor UO_56 (O_56,N_2980,N_2910);
and UO_57 (O_57,N_2971,N_2996);
or UO_58 (O_58,N_2943,N_2935);
nor UO_59 (O_59,N_2953,N_2958);
nand UO_60 (O_60,N_2978,N_2958);
nand UO_61 (O_61,N_2930,N_2922);
nor UO_62 (O_62,N_2967,N_2932);
and UO_63 (O_63,N_2996,N_2942);
and UO_64 (O_64,N_2943,N_2972);
nor UO_65 (O_65,N_2925,N_2938);
nor UO_66 (O_66,N_2917,N_2945);
nand UO_67 (O_67,N_2922,N_2959);
nor UO_68 (O_68,N_2983,N_2964);
nand UO_69 (O_69,N_2991,N_2976);
nor UO_70 (O_70,N_2968,N_2962);
nand UO_71 (O_71,N_2950,N_2980);
nor UO_72 (O_72,N_2914,N_2964);
xnor UO_73 (O_73,N_2941,N_2973);
nand UO_74 (O_74,N_2994,N_2996);
or UO_75 (O_75,N_2908,N_2989);
or UO_76 (O_76,N_2941,N_2948);
or UO_77 (O_77,N_2942,N_2954);
and UO_78 (O_78,N_2998,N_2986);
or UO_79 (O_79,N_2933,N_2951);
and UO_80 (O_80,N_2944,N_2986);
nor UO_81 (O_81,N_2974,N_2950);
nor UO_82 (O_82,N_2913,N_2996);
or UO_83 (O_83,N_2990,N_2941);
and UO_84 (O_84,N_2979,N_2940);
or UO_85 (O_85,N_2986,N_2902);
nor UO_86 (O_86,N_2914,N_2971);
nor UO_87 (O_87,N_2993,N_2984);
xnor UO_88 (O_88,N_2913,N_2976);
nor UO_89 (O_89,N_2956,N_2974);
nor UO_90 (O_90,N_2948,N_2932);
nor UO_91 (O_91,N_2956,N_2985);
nand UO_92 (O_92,N_2989,N_2939);
nor UO_93 (O_93,N_2917,N_2907);
and UO_94 (O_94,N_2931,N_2988);
xor UO_95 (O_95,N_2988,N_2951);
nor UO_96 (O_96,N_2951,N_2937);
and UO_97 (O_97,N_2928,N_2961);
and UO_98 (O_98,N_2927,N_2947);
and UO_99 (O_99,N_2987,N_2903);
nor UO_100 (O_100,N_2966,N_2950);
nand UO_101 (O_101,N_2953,N_2965);
or UO_102 (O_102,N_2913,N_2942);
nand UO_103 (O_103,N_2984,N_2928);
nand UO_104 (O_104,N_2929,N_2978);
and UO_105 (O_105,N_2994,N_2905);
and UO_106 (O_106,N_2910,N_2936);
xor UO_107 (O_107,N_2934,N_2982);
xnor UO_108 (O_108,N_2986,N_2975);
nor UO_109 (O_109,N_2928,N_2910);
nand UO_110 (O_110,N_2977,N_2988);
and UO_111 (O_111,N_2971,N_2930);
nor UO_112 (O_112,N_2952,N_2918);
and UO_113 (O_113,N_2993,N_2909);
and UO_114 (O_114,N_2960,N_2939);
nor UO_115 (O_115,N_2909,N_2985);
nand UO_116 (O_116,N_2992,N_2997);
nor UO_117 (O_117,N_2977,N_2936);
or UO_118 (O_118,N_2952,N_2987);
or UO_119 (O_119,N_2907,N_2920);
nand UO_120 (O_120,N_2941,N_2987);
nand UO_121 (O_121,N_2984,N_2903);
and UO_122 (O_122,N_2924,N_2984);
and UO_123 (O_123,N_2958,N_2970);
nand UO_124 (O_124,N_2913,N_2963);
or UO_125 (O_125,N_2914,N_2978);
or UO_126 (O_126,N_2943,N_2928);
and UO_127 (O_127,N_2985,N_2974);
nor UO_128 (O_128,N_2938,N_2977);
nand UO_129 (O_129,N_2915,N_2905);
nor UO_130 (O_130,N_2943,N_2993);
nand UO_131 (O_131,N_2976,N_2903);
and UO_132 (O_132,N_2911,N_2967);
nor UO_133 (O_133,N_2933,N_2921);
xor UO_134 (O_134,N_2920,N_2996);
or UO_135 (O_135,N_2903,N_2962);
xor UO_136 (O_136,N_2900,N_2978);
or UO_137 (O_137,N_2948,N_2960);
xor UO_138 (O_138,N_2926,N_2950);
and UO_139 (O_139,N_2911,N_2994);
nand UO_140 (O_140,N_2945,N_2998);
nor UO_141 (O_141,N_2991,N_2946);
nand UO_142 (O_142,N_2966,N_2940);
nand UO_143 (O_143,N_2990,N_2929);
xor UO_144 (O_144,N_2990,N_2919);
nor UO_145 (O_145,N_2971,N_2918);
or UO_146 (O_146,N_2994,N_2915);
or UO_147 (O_147,N_2955,N_2923);
or UO_148 (O_148,N_2979,N_2957);
xnor UO_149 (O_149,N_2905,N_2978);
and UO_150 (O_150,N_2970,N_2906);
and UO_151 (O_151,N_2927,N_2963);
nor UO_152 (O_152,N_2943,N_2966);
and UO_153 (O_153,N_2983,N_2971);
xor UO_154 (O_154,N_2929,N_2902);
nor UO_155 (O_155,N_2954,N_2920);
nor UO_156 (O_156,N_2953,N_2922);
and UO_157 (O_157,N_2973,N_2966);
nand UO_158 (O_158,N_2906,N_2987);
or UO_159 (O_159,N_2960,N_2989);
nand UO_160 (O_160,N_2909,N_2963);
or UO_161 (O_161,N_2989,N_2912);
nor UO_162 (O_162,N_2989,N_2900);
and UO_163 (O_163,N_2989,N_2927);
xor UO_164 (O_164,N_2947,N_2914);
nand UO_165 (O_165,N_2949,N_2928);
or UO_166 (O_166,N_2991,N_2900);
xor UO_167 (O_167,N_2945,N_2900);
nand UO_168 (O_168,N_2930,N_2942);
and UO_169 (O_169,N_2935,N_2903);
or UO_170 (O_170,N_2997,N_2946);
or UO_171 (O_171,N_2908,N_2946);
and UO_172 (O_172,N_2903,N_2926);
nand UO_173 (O_173,N_2993,N_2999);
and UO_174 (O_174,N_2920,N_2965);
nand UO_175 (O_175,N_2972,N_2934);
nand UO_176 (O_176,N_2979,N_2921);
nor UO_177 (O_177,N_2974,N_2988);
and UO_178 (O_178,N_2973,N_2939);
nor UO_179 (O_179,N_2967,N_2960);
nand UO_180 (O_180,N_2920,N_2962);
and UO_181 (O_181,N_2915,N_2953);
and UO_182 (O_182,N_2972,N_2962);
nand UO_183 (O_183,N_2931,N_2980);
nor UO_184 (O_184,N_2916,N_2915);
and UO_185 (O_185,N_2913,N_2971);
nand UO_186 (O_186,N_2983,N_2951);
nand UO_187 (O_187,N_2976,N_2926);
and UO_188 (O_188,N_2938,N_2992);
or UO_189 (O_189,N_2912,N_2935);
and UO_190 (O_190,N_2923,N_2902);
nand UO_191 (O_191,N_2990,N_2986);
or UO_192 (O_192,N_2934,N_2931);
nand UO_193 (O_193,N_2972,N_2910);
nand UO_194 (O_194,N_2930,N_2936);
or UO_195 (O_195,N_2971,N_2989);
xor UO_196 (O_196,N_2951,N_2999);
nand UO_197 (O_197,N_2998,N_2921);
or UO_198 (O_198,N_2965,N_2910);
nand UO_199 (O_199,N_2952,N_2983);
nand UO_200 (O_200,N_2938,N_2998);
and UO_201 (O_201,N_2934,N_2918);
nand UO_202 (O_202,N_2926,N_2998);
or UO_203 (O_203,N_2981,N_2950);
nor UO_204 (O_204,N_2926,N_2904);
xor UO_205 (O_205,N_2968,N_2966);
nand UO_206 (O_206,N_2990,N_2972);
nand UO_207 (O_207,N_2955,N_2946);
nor UO_208 (O_208,N_2929,N_2972);
and UO_209 (O_209,N_2929,N_2914);
and UO_210 (O_210,N_2940,N_2915);
nand UO_211 (O_211,N_2993,N_2960);
and UO_212 (O_212,N_2946,N_2970);
and UO_213 (O_213,N_2969,N_2947);
and UO_214 (O_214,N_2977,N_2963);
nand UO_215 (O_215,N_2970,N_2949);
or UO_216 (O_216,N_2929,N_2948);
nor UO_217 (O_217,N_2907,N_2937);
or UO_218 (O_218,N_2950,N_2935);
or UO_219 (O_219,N_2949,N_2940);
nand UO_220 (O_220,N_2914,N_2977);
and UO_221 (O_221,N_2970,N_2920);
or UO_222 (O_222,N_2957,N_2913);
or UO_223 (O_223,N_2960,N_2927);
nand UO_224 (O_224,N_2928,N_2946);
and UO_225 (O_225,N_2955,N_2993);
nor UO_226 (O_226,N_2953,N_2946);
nor UO_227 (O_227,N_2992,N_2906);
nor UO_228 (O_228,N_2961,N_2934);
or UO_229 (O_229,N_2958,N_2915);
nand UO_230 (O_230,N_2966,N_2942);
and UO_231 (O_231,N_2923,N_2961);
and UO_232 (O_232,N_2962,N_2989);
or UO_233 (O_233,N_2925,N_2983);
nor UO_234 (O_234,N_2992,N_2958);
and UO_235 (O_235,N_2900,N_2979);
or UO_236 (O_236,N_2917,N_2994);
nor UO_237 (O_237,N_2988,N_2991);
and UO_238 (O_238,N_2942,N_2961);
nor UO_239 (O_239,N_2995,N_2977);
nand UO_240 (O_240,N_2967,N_2991);
or UO_241 (O_241,N_2978,N_2992);
nand UO_242 (O_242,N_2966,N_2963);
nand UO_243 (O_243,N_2972,N_2978);
or UO_244 (O_244,N_2974,N_2979);
nor UO_245 (O_245,N_2940,N_2999);
nand UO_246 (O_246,N_2984,N_2922);
or UO_247 (O_247,N_2965,N_2983);
nor UO_248 (O_248,N_2952,N_2925);
or UO_249 (O_249,N_2943,N_2910);
nor UO_250 (O_250,N_2928,N_2906);
and UO_251 (O_251,N_2947,N_2963);
and UO_252 (O_252,N_2978,N_2935);
and UO_253 (O_253,N_2994,N_2957);
and UO_254 (O_254,N_2931,N_2928);
nor UO_255 (O_255,N_2954,N_2966);
nor UO_256 (O_256,N_2964,N_2939);
or UO_257 (O_257,N_2959,N_2976);
and UO_258 (O_258,N_2992,N_2935);
and UO_259 (O_259,N_2977,N_2935);
or UO_260 (O_260,N_2935,N_2983);
nand UO_261 (O_261,N_2927,N_2930);
xnor UO_262 (O_262,N_2993,N_2997);
and UO_263 (O_263,N_2913,N_2927);
nor UO_264 (O_264,N_2986,N_2921);
nor UO_265 (O_265,N_2917,N_2915);
nand UO_266 (O_266,N_2985,N_2947);
nor UO_267 (O_267,N_2965,N_2921);
xnor UO_268 (O_268,N_2920,N_2979);
nor UO_269 (O_269,N_2969,N_2946);
and UO_270 (O_270,N_2987,N_2968);
or UO_271 (O_271,N_2950,N_2925);
nor UO_272 (O_272,N_2988,N_2975);
nor UO_273 (O_273,N_2981,N_2924);
or UO_274 (O_274,N_2972,N_2915);
nand UO_275 (O_275,N_2954,N_2984);
or UO_276 (O_276,N_2908,N_2983);
or UO_277 (O_277,N_2967,N_2902);
xnor UO_278 (O_278,N_2931,N_2905);
nand UO_279 (O_279,N_2902,N_2952);
nor UO_280 (O_280,N_2937,N_2946);
and UO_281 (O_281,N_2956,N_2976);
xnor UO_282 (O_282,N_2971,N_2958);
or UO_283 (O_283,N_2903,N_2951);
and UO_284 (O_284,N_2905,N_2904);
or UO_285 (O_285,N_2949,N_2990);
and UO_286 (O_286,N_2955,N_2919);
or UO_287 (O_287,N_2963,N_2984);
or UO_288 (O_288,N_2973,N_2998);
xor UO_289 (O_289,N_2911,N_2945);
and UO_290 (O_290,N_2930,N_2921);
nor UO_291 (O_291,N_2976,N_2943);
and UO_292 (O_292,N_2956,N_2910);
and UO_293 (O_293,N_2908,N_2978);
and UO_294 (O_294,N_2960,N_2975);
nand UO_295 (O_295,N_2991,N_2929);
and UO_296 (O_296,N_2945,N_2930);
or UO_297 (O_297,N_2941,N_2947);
nor UO_298 (O_298,N_2989,N_2974);
or UO_299 (O_299,N_2977,N_2987);
and UO_300 (O_300,N_2992,N_2964);
or UO_301 (O_301,N_2941,N_2931);
nand UO_302 (O_302,N_2930,N_2917);
or UO_303 (O_303,N_2956,N_2980);
nor UO_304 (O_304,N_2906,N_2947);
xor UO_305 (O_305,N_2952,N_2910);
xor UO_306 (O_306,N_2950,N_2942);
or UO_307 (O_307,N_2905,N_2930);
xor UO_308 (O_308,N_2959,N_2980);
and UO_309 (O_309,N_2962,N_2982);
nor UO_310 (O_310,N_2989,N_2938);
or UO_311 (O_311,N_2973,N_2922);
nor UO_312 (O_312,N_2908,N_2960);
nand UO_313 (O_313,N_2994,N_2998);
nand UO_314 (O_314,N_2903,N_2963);
or UO_315 (O_315,N_2981,N_2938);
and UO_316 (O_316,N_2931,N_2919);
and UO_317 (O_317,N_2996,N_2933);
xnor UO_318 (O_318,N_2903,N_2991);
or UO_319 (O_319,N_2973,N_2982);
nor UO_320 (O_320,N_2986,N_2918);
nand UO_321 (O_321,N_2975,N_2983);
nor UO_322 (O_322,N_2975,N_2992);
and UO_323 (O_323,N_2915,N_2911);
and UO_324 (O_324,N_2953,N_2972);
nand UO_325 (O_325,N_2923,N_2945);
xor UO_326 (O_326,N_2980,N_2979);
or UO_327 (O_327,N_2947,N_2966);
nand UO_328 (O_328,N_2954,N_2922);
or UO_329 (O_329,N_2992,N_2947);
nand UO_330 (O_330,N_2937,N_2924);
or UO_331 (O_331,N_2904,N_2944);
or UO_332 (O_332,N_2942,N_2927);
or UO_333 (O_333,N_2905,N_2983);
nor UO_334 (O_334,N_2902,N_2949);
or UO_335 (O_335,N_2926,N_2933);
or UO_336 (O_336,N_2924,N_2985);
or UO_337 (O_337,N_2977,N_2956);
nand UO_338 (O_338,N_2903,N_2944);
nor UO_339 (O_339,N_2967,N_2985);
xnor UO_340 (O_340,N_2929,N_2973);
nand UO_341 (O_341,N_2979,N_2937);
xor UO_342 (O_342,N_2900,N_2902);
nand UO_343 (O_343,N_2991,N_2949);
or UO_344 (O_344,N_2955,N_2922);
xnor UO_345 (O_345,N_2952,N_2961);
xnor UO_346 (O_346,N_2935,N_2906);
and UO_347 (O_347,N_2965,N_2993);
or UO_348 (O_348,N_2935,N_2909);
or UO_349 (O_349,N_2934,N_2939);
and UO_350 (O_350,N_2990,N_2962);
or UO_351 (O_351,N_2903,N_2910);
nor UO_352 (O_352,N_2907,N_2947);
nor UO_353 (O_353,N_2981,N_2995);
xnor UO_354 (O_354,N_2937,N_2983);
and UO_355 (O_355,N_2930,N_2947);
and UO_356 (O_356,N_2901,N_2910);
nand UO_357 (O_357,N_2917,N_2998);
nand UO_358 (O_358,N_2958,N_2931);
xnor UO_359 (O_359,N_2953,N_2944);
nand UO_360 (O_360,N_2932,N_2958);
nor UO_361 (O_361,N_2924,N_2907);
nor UO_362 (O_362,N_2927,N_2932);
nand UO_363 (O_363,N_2990,N_2982);
xnor UO_364 (O_364,N_2993,N_2925);
nor UO_365 (O_365,N_2953,N_2933);
nand UO_366 (O_366,N_2901,N_2987);
and UO_367 (O_367,N_2959,N_2967);
nand UO_368 (O_368,N_2904,N_2985);
or UO_369 (O_369,N_2904,N_2987);
nand UO_370 (O_370,N_2965,N_2963);
or UO_371 (O_371,N_2902,N_2954);
nor UO_372 (O_372,N_2901,N_2970);
or UO_373 (O_373,N_2972,N_2981);
or UO_374 (O_374,N_2972,N_2940);
nor UO_375 (O_375,N_2984,N_2937);
xor UO_376 (O_376,N_2921,N_2918);
nand UO_377 (O_377,N_2996,N_2987);
or UO_378 (O_378,N_2976,N_2955);
nor UO_379 (O_379,N_2932,N_2943);
and UO_380 (O_380,N_2915,N_2926);
or UO_381 (O_381,N_2911,N_2969);
nand UO_382 (O_382,N_2960,N_2996);
or UO_383 (O_383,N_2945,N_2968);
or UO_384 (O_384,N_2901,N_2958);
nor UO_385 (O_385,N_2959,N_2906);
or UO_386 (O_386,N_2936,N_2944);
and UO_387 (O_387,N_2989,N_2965);
xor UO_388 (O_388,N_2916,N_2925);
xnor UO_389 (O_389,N_2901,N_2974);
nor UO_390 (O_390,N_2955,N_2930);
nor UO_391 (O_391,N_2943,N_2908);
nand UO_392 (O_392,N_2923,N_2905);
or UO_393 (O_393,N_2923,N_2927);
nand UO_394 (O_394,N_2991,N_2980);
and UO_395 (O_395,N_2955,N_2944);
nand UO_396 (O_396,N_2979,N_2969);
and UO_397 (O_397,N_2909,N_2962);
nand UO_398 (O_398,N_2957,N_2919);
or UO_399 (O_399,N_2977,N_2964);
or UO_400 (O_400,N_2932,N_2996);
xnor UO_401 (O_401,N_2995,N_2933);
or UO_402 (O_402,N_2951,N_2911);
or UO_403 (O_403,N_2936,N_2937);
nor UO_404 (O_404,N_2989,N_2907);
nand UO_405 (O_405,N_2912,N_2921);
and UO_406 (O_406,N_2914,N_2996);
nand UO_407 (O_407,N_2901,N_2975);
nand UO_408 (O_408,N_2901,N_2918);
nor UO_409 (O_409,N_2997,N_2920);
nor UO_410 (O_410,N_2984,N_2952);
nor UO_411 (O_411,N_2947,N_2903);
xor UO_412 (O_412,N_2973,N_2953);
or UO_413 (O_413,N_2917,N_2920);
nand UO_414 (O_414,N_2948,N_2955);
nor UO_415 (O_415,N_2985,N_2973);
nand UO_416 (O_416,N_2924,N_2962);
nand UO_417 (O_417,N_2950,N_2970);
nand UO_418 (O_418,N_2977,N_2969);
or UO_419 (O_419,N_2910,N_2961);
or UO_420 (O_420,N_2971,N_2909);
and UO_421 (O_421,N_2967,N_2954);
and UO_422 (O_422,N_2994,N_2916);
nor UO_423 (O_423,N_2914,N_2987);
xnor UO_424 (O_424,N_2974,N_2900);
nor UO_425 (O_425,N_2973,N_2990);
and UO_426 (O_426,N_2943,N_2989);
and UO_427 (O_427,N_2944,N_2997);
or UO_428 (O_428,N_2977,N_2999);
xnor UO_429 (O_429,N_2921,N_2970);
or UO_430 (O_430,N_2989,N_2926);
and UO_431 (O_431,N_2973,N_2925);
and UO_432 (O_432,N_2944,N_2926);
or UO_433 (O_433,N_2900,N_2924);
and UO_434 (O_434,N_2972,N_2966);
or UO_435 (O_435,N_2952,N_2951);
or UO_436 (O_436,N_2938,N_2922);
or UO_437 (O_437,N_2947,N_2925);
and UO_438 (O_438,N_2912,N_2964);
or UO_439 (O_439,N_2937,N_2975);
nand UO_440 (O_440,N_2901,N_2952);
or UO_441 (O_441,N_2949,N_2997);
or UO_442 (O_442,N_2919,N_2986);
nor UO_443 (O_443,N_2963,N_2904);
and UO_444 (O_444,N_2923,N_2971);
and UO_445 (O_445,N_2993,N_2917);
xor UO_446 (O_446,N_2917,N_2906);
nor UO_447 (O_447,N_2945,N_2970);
xnor UO_448 (O_448,N_2929,N_2928);
nor UO_449 (O_449,N_2916,N_2921);
nand UO_450 (O_450,N_2930,N_2992);
xnor UO_451 (O_451,N_2997,N_2939);
and UO_452 (O_452,N_2984,N_2970);
nor UO_453 (O_453,N_2918,N_2920);
and UO_454 (O_454,N_2907,N_2914);
nor UO_455 (O_455,N_2922,N_2931);
nor UO_456 (O_456,N_2917,N_2973);
or UO_457 (O_457,N_2934,N_2984);
or UO_458 (O_458,N_2937,N_2919);
nor UO_459 (O_459,N_2997,N_2922);
nor UO_460 (O_460,N_2959,N_2990);
or UO_461 (O_461,N_2914,N_2917);
xor UO_462 (O_462,N_2933,N_2917);
nand UO_463 (O_463,N_2973,N_2993);
and UO_464 (O_464,N_2936,N_2932);
or UO_465 (O_465,N_2907,N_2913);
nor UO_466 (O_466,N_2972,N_2948);
or UO_467 (O_467,N_2909,N_2970);
nand UO_468 (O_468,N_2941,N_2933);
nor UO_469 (O_469,N_2996,N_2901);
or UO_470 (O_470,N_2976,N_2936);
nor UO_471 (O_471,N_2913,N_2919);
and UO_472 (O_472,N_2931,N_2952);
nor UO_473 (O_473,N_2943,N_2923);
nand UO_474 (O_474,N_2909,N_2918);
xnor UO_475 (O_475,N_2971,N_2900);
xnor UO_476 (O_476,N_2993,N_2902);
and UO_477 (O_477,N_2987,N_2918);
and UO_478 (O_478,N_2912,N_2979);
and UO_479 (O_479,N_2976,N_2968);
nor UO_480 (O_480,N_2925,N_2956);
and UO_481 (O_481,N_2987,N_2928);
and UO_482 (O_482,N_2940,N_2996);
nand UO_483 (O_483,N_2979,N_2915);
or UO_484 (O_484,N_2936,N_2973);
nor UO_485 (O_485,N_2977,N_2900);
and UO_486 (O_486,N_2921,N_2984);
nand UO_487 (O_487,N_2971,N_2951);
and UO_488 (O_488,N_2971,N_2959);
or UO_489 (O_489,N_2926,N_2977);
nand UO_490 (O_490,N_2943,N_2939);
nand UO_491 (O_491,N_2976,N_2938);
and UO_492 (O_492,N_2921,N_2943);
and UO_493 (O_493,N_2969,N_2960);
nor UO_494 (O_494,N_2993,N_2963);
nor UO_495 (O_495,N_2951,N_2984);
or UO_496 (O_496,N_2906,N_2937);
nor UO_497 (O_497,N_2975,N_2944);
or UO_498 (O_498,N_2932,N_2912);
and UO_499 (O_499,N_2978,N_2989);
endmodule