module basic_500_3000_500_50_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_185,In_219);
or U1 (N_1,In_173,In_424);
and U2 (N_2,In_81,In_130);
or U3 (N_3,In_101,In_100);
or U4 (N_4,In_153,In_467);
nor U5 (N_5,In_107,In_393);
or U6 (N_6,In_160,In_19);
nor U7 (N_7,In_76,In_403);
nor U8 (N_8,In_225,In_460);
nand U9 (N_9,In_109,In_289);
and U10 (N_10,In_99,In_486);
nor U11 (N_11,In_406,In_151);
and U12 (N_12,In_417,In_230);
or U13 (N_13,In_194,In_4);
or U14 (N_14,In_431,In_146);
nand U15 (N_15,In_473,In_170);
nand U16 (N_16,In_368,In_58);
nand U17 (N_17,In_351,In_339);
nor U18 (N_18,In_1,In_484);
and U19 (N_19,In_17,In_377);
nor U20 (N_20,In_364,In_48);
nand U21 (N_21,In_399,In_366);
or U22 (N_22,In_45,In_189);
nor U23 (N_23,In_382,In_300);
nor U24 (N_24,In_443,In_348);
nor U25 (N_25,In_157,In_441);
nor U26 (N_26,In_329,In_416);
nand U27 (N_27,In_288,In_301);
nand U28 (N_28,In_217,In_131);
nor U29 (N_29,In_497,In_87);
nor U30 (N_30,In_453,In_421);
nor U31 (N_31,In_353,In_231);
and U32 (N_32,In_326,In_213);
nand U33 (N_33,In_498,In_226);
and U34 (N_34,In_178,In_165);
and U35 (N_35,In_51,In_295);
or U36 (N_36,In_207,In_40);
and U37 (N_37,In_396,In_73);
nand U38 (N_38,In_481,In_218);
nor U39 (N_39,In_80,In_162);
nor U40 (N_40,In_310,In_139);
and U41 (N_41,In_234,In_150);
or U42 (N_42,In_359,In_26);
or U43 (N_43,In_251,In_297);
and U44 (N_44,In_272,In_205);
nand U45 (N_45,In_240,In_463);
nand U46 (N_46,In_214,In_363);
nand U47 (N_47,In_129,In_132);
and U48 (N_48,In_23,In_450);
and U49 (N_49,In_346,In_337);
and U50 (N_50,In_57,In_287);
and U51 (N_51,In_321,In_386);
and U52 (N_52,In_456,In_415);
nor U53 (N_53,In_8,In_405);
nor U54 (N_54,In_422,In_10);
nor U55 (N_55,In_152,In_269);
nand U56 (N_56,In_490,In_53);
nor U57 (N_57,In_468,In_229);
and U58 (N_58,In_35,In_198);
or U59 (N_59,In_252,In_465);
nor U60 (N_60,In_277,In_340);
nor U61 (N_61,In_31,In_92);
and U62 (N_62,In_158,In_263);
or U63 (N_63,In_104,N_23);
nand U64 (N_64,In_330,In_85);
or U65 (N_65,In_286,In_390);
or U66 (N_66,In_246,N_43);
and U67 (N_67,In_476,In_262);
nand U68 (N_68,In_180,In_3);
nor U69 (N_69,In_241,N_0);
or U70 (N_70,In_454,In_462);
nand U71 (N_71,In_119,N_4);
nor U72 (N_72,In_404,In_313);
and U73 (N_73,In_163,N_47);
nor U74 (N_74,N_58,In_372);
and U75 (N_75,In_172,In_335);
or U76 (N_76,In_64,N_14);
nand U77 (N_77,In_125,In_376);
nor U78 (N_78,In_455,In_428);
nand U79 (N_79,In_39,In_44);
nand U80 (N_80,In_411,In_168);
and U81 (N_81,In_304,In_159);
and U82 (N_82,In_79,In_154);
nor U83 (N_83,In_400,In_319);
nand U84 (N_84,In_281,In_223);
or U85 (N_85,In_333,In_7);
nor U86 (N_86,In_265,In_466);
nor U87 (N_87,In_419,In_305);
and U88 (N_88,In_68,In_211);
nor U89 (N_89,In_120,In_429);
nand U90 (N_90,In_34,In_276);
nand U91 (N_91,In_121,N_2);
or U92 (N_92,In_56,In_117);
or U93 (N_93,In_140,In_361);
and U94 (N_94,In_123,N_10);
nor U95 (N_95,In_238,In_228);
or U96 (N_96,In_93,In_54);
nor U97 (N_97,In_282,In_259);
and U98 (N_98,In_334,In_290);
or U99 (N_99,In_439,In_271);
nor U100 (N_100,N_25,In_127);
nand U101 (N_101,In_284,In_145);
or U102 (N_102,In_25,In_134);
and U103 (N_103,In_86,In_447);
or U104 (N_104,In_95,In_414);
nor U105 (N_105,In_47,In_365);
and U106 (N_106,N_9,In_347);
nand U107 (N_107,In_360,In_378);
nor U108 (N_108,In_492,In_434);
or U109 (N_109,In_496,In_352);
nor U110 (N_110,In_320,In_397);
and U111 (N_111,N_29,In_187);
and U112 (N_112,In_115,In_314);
or U113 (N_113,In_206,In_482);
nor U114 (N_114,In_63,In_373);
nor U115 (N_115,In_208,In_477);
and U116 (N_116,In_294,N_42);
nand U117 (N_117,In_480,In_243);
nand U118 (N_118,In_489,In_283);
nor U119 (N_119,N_33,N_59);
nor U120 (N_120,In_487,N_94);
nand U121 (N_121,N_7,In_312);
nor U122 (N_122,N_86,In_28);
or U123 (N_123,In_128,In_98);
and U124 (N_124,In_438,In_379);
nor U125 (N_125,N_35,In_227);
nand U126 (N_126,In_324,N_107);
nand U127 (N_127,In_471,In_258);
nand U128 (N_128,In_82,In_188);
and U129 (N_129,In_495,N_18);
and U130 (N_130,In_237,N_38);
nand U131 (N_131,In_166,In_311);
and U132 (N_132,N_61,N_68);
nand U133 (N_133,N_84,In_70);
or U134 (N_134,In_285,In_202);
nor U135 (N_135,N_93,N_115);
nand U136 (N_136,In_317,In_142);
and U137 (N_137,N_81,In_137);
and U138 (N_138,N_63,N_15);
or U139 (N_139,In_449,In_233);
nand U140 (N_140,N_65,In_407);
nor U141 (N_141,In_33,In_112);
nand U142 (N_142,In_268,In_293);
nor U143 (N_143,In_327,In_303);
or U144 (N_144,N_26,In_362);
nor U145 (N_145,In_84,In_461);
or U146 (N_146,In_459,In_440);
nand U147 (N_147,In_74,In_418);
nand U148 (N_148,In_275,In_254);
or U149 (N_149,In_182,In_394);
or U150 (N_150,In_278,In_102);
and U151 (N_151,In_402,In_30);
nor U152 (N_152,In_91,In_469);
nor U153 (N_153,N_44,N_85);
nor U154 (N_154,In_156,In_221);
xnor U155 (N_155,In_385,N_3);
or U156 (N_156,In_302,In_343);
nand U157 (N_157,N_40,In_430);
xor U158 (N_158,In_369,In_413);
and U159 (N_159,In_485,In_446);
nand U160 (N_160,In_60,In_494);
and U161 (N_161,In_37,In_410);
and U162 (N_162,In_354,In_478);
nor U163 (N_163,In_14,In_260);
nand U164 (N_164,In_13,In_279);
nand U165 (N_165,N_83,In_204);
or U166 (N_166,In_200,In_280);
nand U167 (N_167,In_253,In_55);
and U168 (N_168,N_113,N_53);
nor U169 (N_169,In_437,N_56);
nor U170 (N_170,N_36,N_106);
nor U171 (N_171,N_60,In_38);
nand U172 (N_172,In_274,In_244);
nand U173 (N_173,N_31,In_59);
nand U174 (N_174,In_408,N_91);
or U175 (N_175,N_1,In_344);
nand U176 (N_176,In_9,In_291);
and U177 (N_177,In_436,In_349);
or U178 (N_178,N_116,N_52);
nand U179 (N_179,N_100,In_220);
or U180 (N_180,In_72,In_474);
and U181 (N_181,N_76,N_149);
or U182 (N_182,In_94,N_179);
or U183 (N_183,N_170,In_196);
nor U184 (N_184,In_398,In_245);
nand U185 (N_185,N_167,In_409);
nand U186 (N_186,In_83,In_21);
and U187 (N_187,N_134,In_432);
nor U188 (N_188,In_388,In_167);
and U189 (N_189,In_66,In_22);
nand U190 (N_190,In_342,In_266);
nor U191 (N_191,In_149,N_50);
or U192 (N_192,N_158,In_216);
and U193 (N_193,N_177,N_74);
nand U194 (N_194,In_5,N_136);
nor U195 (N_195,In_75,In_464);
nor U196 (N_196,In_380,In_209);
xor U197 (N_197,In_483,N_133);
nand U198 (N_198,In_78,In_247);
nand U199 (N_199,N_17,In_2);
nor U200 (N_200,In_164,In_36);
nor U201 (N_201,In_114,In_69);
or U202 (N_202,In_451,N_73);
and U203 (N_203,In_65,In_328);
nor U204 (N_204,In_118,In_97);
nor U205 (N_205,In_358,In_357);
nand U206 (N_206,N_130,N_57);
or U207 (N_207,N_168,N_64);
nand U208 (N_208,N_172,In_367);
or U209 (N_209,In_96,In_124);
nor U210 (N_210,In_331,In_106);
or U211 (N_211,N_62,N_151);
or U212 (N_212,In_249,N_110);
and U213 (N_213,N_54,N_166);
nand U214 (N_214,N_5,N_78);
or U215 (N_215,N_67,In_387);
and U216 (N_216,In_488,In_77);
or U217 (N_217,In_122,In_264);
nor U218 (N_218,N_46,N_111);
nor U219 (N_219,N_80,N_72);
nand U220 (N_220,N_16,N_164);
and U221 (N_221,In_235,N_105);
nor U222 (N_222,N_69,In_457);
nand U223 (N_223,In_49,N_154);
nand U224 (N_224,In_186,In_425);
or U225 (N_225,In_356,In_50);
nor U226 (N_226,In_318,N_127);
and U227 (N_227,N_48,N_126);
nor U228 (N_228,N_163,N_142);
nand U229 (N_229,N_144,N_77);
xnor U230 (N_230,In_191,N_176);
or U231 (N_231,In_236,In_267);
nor U232 (N_232,In_176,In_136);
nand U233 (N_233,In_133,N_92);
or U234 (N_234,N_41,N_139);
nand U235 (N_235,In_261,In_24);
and U236 (N_236,N_70,N_157);
nor U237 (N_237,N_143,In_203);
nor U238 (N_238,N_125,N_34);
and U239 (N_239,In_0,N_37);
nand U240 (N_240,In_105,In_61);
nand U241 (N_241,N_178,N_22);
and U242 (N_242,In_270,In_67);
nor U243 (N_243,In_381,N_227);
and U244 (N_244,In_442,N_88);
nor U245 (N_245,In_316,In_250);
nor U246 (N_246,In_52,In_423);
nand U247 (N_247,N_165,N_79);
nor U248 (N_248,In_309,N_104);
nor U249 (N_249,In_332,In_315);
nor U250 (N_250,N_108,N_228);
or U251 (N_251,In_384,N_90);
or U252 (N_252,In_201,N_184);
or U253 (N_253,In_448,N_233);
nor U254 (N_254,In_255,N_232);
nor U255 (N_255,N_236,N_82);
and U256 (N_256,N_103,N_152);
nor U257 (N_257,In_307,In_248);
nand U258 (N_258,N_204,N_206);
or U259 (N_259,N_49,In_296);
and U260 (N_260,In_126,In_42);
and U261 (N_261,N_218,In_401);
and U262 (N_262,N_128,N_20);
or U263 (N_263,In_323,N_219);
or U264 (N_264,In_155,N_195);
nor U265 (N_265,In_29,In_475);
nand U266 (N_266,In_370,N_141);
nand U267 (N_267,N_123,N_185);
nand U268 (N_268,In_41,N_239);
and U269 (N_269,In_239,N_124);
nand U270 (N_270,N_229,N_87);
or U271 (N_271,N_212,N_194);
nor U272 (N_272,In_103,N_45);
and U273 (N_273,In_43,In_371);
or U274 (N_274,N_122,N_193);
or U275 (N_275,In_46,N_117);
or U276 (N_276,N_155,N_171);
or U277 (N_277,In_147,In_111);
and U278 (N_278,N_137,N_148);
nor U279 (N_279,N_102,N_131);
nand U280 (N_280,In_89,N_169);
nor U281 (N_281,N_28,In_435);
and U282 (N_282,In_20,In_257);
nand U283 (N_283,N_120,In_144);
or U284 (N_284,N_132,In_273);
and U285 (N_285,In_88,N_188);
and U286 (N_286,In_325,N_199);
or U287 (N_287,N_129,In_197);
nor U288 (N_288,N_180,In_499);
nand U289 (N_289,N_32,In_27);
nand U290 (N_290,N_186,In_192);
nand U291 (N_291,N_183,N_220);
nor U292 (N_292,N_147,In_175);
nor U293 (N_293,In_212,N_51);
and U294 (N_294,N_8,In_392);
nor U295 (N_295,N_189,N_24);
nand U296 (N_296,In_215,In_62);
and U297 (N_297,N_203,In_184);
and U298 (N_298,N_197,N_217);
nand U299 (N_299,N_71,In_452);
nand U300 (N_300,In_395,In_383);
nor U301 (N_301,In_135,N_30);
or U302 (N_302,In_12,In_350);
nor U303 (N_303,In_374,N_192);
nand U304 (N_304,N_235,In_195);
and U305 (N_305,N_291,In_298);
and U306 (N_306,N_118,N_198);
or U307 (N_307,N_230,In_458);
or U308 (N_308,N_259,In_472);
and U309 (N_309,N_109,In_138);
nand U310 (N_310,N_250,N_205);
nor U311 (N_311,In_292,N_262);
nor U312 (N_312,In_183,N_182);
nor U313 (N_313,N_145,In_341);
nor U314 (N_314,N_238,In_171);
or U315 (N_315,N_276,N_279);
nand U316 (N_316,N_244,N_150);
and U317 (N_317,N_258,In_18);
or U318 (N_318,N_226,In_116);
nor U319 (N_319,N_19,In_412);
nor U320 (N_320,N_286,N_97);
and U321 (N_321,In_110,In_433);
nand U322 (N_322,N_271,N_89);
nor U323 (N_323,N_175,In_179);
or U324 (N_324,In_242,N_221);
nand U325 (N_325,N_214,N_285);
and U326 (N_326,N_162,N_275);
nand U327 (N_327,In_190,N_156);
nand U328 (N_328,N_264,In_345);
and U329 (N_329,N_202,N_245);
or U330 (N_330,N_12,N_247);
nand U331 (N_331,In_161,In_177);
or U332 (N_332,In_193,N_55);
or U333 (N_333,N_251,N_268);
and U334 (N_334,In_445,In_141);
and U335 (N_335,N_255,In_148);
and U336 (N_336,N_260,N_201);
nand U337 (N_337,In_336,In_181);
nand U338 (N_338,N_215,N_278);
nor U339 (N_339,In_210,In_11);
or U340 (N_340,In_493,N_6);
nand U341 (N_341,N_39,N_160);
or U342 (N_342,N_101,In_299);
or U343 (N_343,N_270,N_114);
and U344 (N_344,N_223,N_246);
and U345 (N_345,N_96,N_266);
nor U346 (N_346,In_232,In_108);
nor U347 (N_347,N_211,In_15);
nor U348 (N_348,N_296,N_249);
nor U349 (N_349,In_426,In_71);
or U350 (N_350,In_322,N_254);
nand U351 (N_351,N_234,N_95);
nor U352 (N_352,N_138,N_173);
or U353 (N_353,In_470,N_290);
or U354 (N_354,In_427,In_174);
or U355 (N_355,N_196,N_287);
and U356 (N_356,N_241,N_256);
nor U357 (N_357,N_272,N_281);
nand U358 (N_358,N_263,N_21);
and U359 (N_359,N_253,In_491);
or U360 (N_360,In_479,N_346);
and U361 (N_361,N_146,N_343);
or U362 (N_362,In_256,N_248);
or U363 (N_363,In_391,N_311);
nand U364 (N_364,N_351,N_11);
and U365 (N_365,N_354,N_333);
nor U366 (N_366,N_200,N_242);
or U367 (N_367,N_337,N_300);
or U368 (N_368,N_310,N_353);
nor U369 (N_369,N_305,N_315);
nand U370 (N_370,In_222,N_216);
or U371 (N_371,N_261,N_213);
and U372 (N_372,N_328,N_280);
nand U373 (N_373,N_336,N_293);
and U374 (N_374,N_358,In_169);
nand U375 (N_375,N_301,N_340);
or U376 (N_376,N_352,N_208);
nand U377 (N_377,N_99,N_252);
and U378 (N_378,N_295,N_314);
nor U379 (N_379,In_199,N_119);
or U380 (N_380,N_121,N_334);
nor U381 (N_381,In_355,N_135);
or U382 (N_382,N_341,In_143);
xnor U383 (N_383,N_348,N_303);
and U384 (N_384,N_283,N_66);
or U385 (N_385,N_322,N_13);
nand U386 (N_386,In_338,N_292);
xor U387 (N_387,N_282,N_331);
and U388 (N_388,N_330,In_308);
nand U389 (N_389,N_327,N_357);
and U390 (N_390,N_317,N_312);
nand U391 (N_391,In_306,N_174);
nand U392 (N_392,N_289,N_237);
or U393 (N_393,N_140,N_240);
nor U394 (N_394,N_27,N_347);
nor U395 (N_395,N_288,N_277);
and U396 (N_396,N_225,N_243);
nand U397 (N_397,N_350,N_257);
and U398 (N_398,N_316,N_153);
nor U399 (N_399,N_284,N_159);
and U400 (N_400,In_444,N_231);
or U401 (N_401,N_307,N_338);
or U402 (N_402,N_306,N_210);
nand U403 (N_403,N_304,N_98);
nand U404 (N_404,N_313,N_161);
nand U405 (N_405,N_187,N_349);
and U406 (N_406,N_326,In_6);
nand U407 (N_407,N_302,N_112);
or U408 (N_408,In_90,N_356);
nand U409 (N_409,N_345,N_297);
and U410 (N_410,N_191,N_75);
nor U411 (N_411,N_181,N_209);
nand U412 (N_412,In_16,In_420);
or U413 (N_413,N_325,In_113);
or U414 (N_414,In_32,N_318);
or U415 (N_415,N_222,N_335);
and U416 (N_416,N_267,N_323);
nor U417 (N_417,N_273,N_190);
nor U418 (N_418,N_299,N_321);
and U419 (N_419,N_324,N_298);
nand U420 (N_420,N_415,N_397);
or U421 (N_421,N_417,N_359);
or U422 (N_422,N_369,N_385);
and U423 (N_423,N_384,N_411);
nand U424 (N_424,N_375,N_387);
or U425 (N_425,N_389,N_376);
nand U426 (N_426,N_412,N_377);
or U427 (N_427,N_419,N_416);
nor U428 (N_428,N_372,N_400);
and U429 (N_429,N_378,N_410);
or U430 (N_430,N_371,N_407);
nand U431 (N_431,N_294,N_329);
or U432 (N_432,N_383,N_392);
nand U433 (N_433,In_224,N_274);
nand U434 (N_434,N_414,N_401);
nand U435 (N_435,N_308,N_363);
or U436 (N_436,N_224,N_409);
nand U437 (N_437,N_265,N_404);
or U438 (N_438,N_391,N_393);
and U439 (N_439,N_408,N_379);
nand U440 (N_440,N_381,N_332);
nand U441 (N_441,N_380,N_418);
nand U442 (N_442,N_370,N_207);
nor U443 (N_443,N_395,N_398);
and U444 (N_444,N_269,N_373);
nand U445 (N_445,N_361,N_403);
nor U446 (N_446,N_386,N_368);
and U447 (N_447,N_339,N_413);
nand U448 (N_448,N_320,N_366);
and U449 (N_449,N_394,N_362);
or U450 (N_450,N_374,N_365);
nor U451 (N_451,N_402,N_355);
and U452 (N_452,N_319,N_367);
xnor U453 (N_453,N_390,N_309);
nand U454 (N_454,N_344,N_388);
nand U455 (N_455,In_375,N_399);
and U456 (N_456,N_364,N_396);
or U457 (N_457,N_382,N_342);
nor U458 (N_458,N_406,In_389);
nor U459 (N_459,N_405,N_360);
nor U460 (N_460,N_342,N_399);
nor U461 (N_461,N_367,In_375);
nand U462 (N_462,N_398,N_329);
nand U463 (N_463,N_402,N_274);
and U464 (N_464,N_409,N_395);
or U465 (N_465,N_294,In_375);
and U466 (N_466,N_412,N_381);
or U467 (N_467,N_408,N_359);
nor U468 (N_468,N_409,In_375);
or U469 (N_469,N_404,N_416);
or U470 (N_470,N_377,N_370);
or U471 (N_471,N_390,N_384);
and U472 (N_472,N_408,N_381);
or U473 (N_473,N_355,N_375);
and U474 (N_474,N_393,N_394);
nand U475 (N_475,N_265,N_408);
nor U476 (N_476,N_392,N_386);
nor U477 (N_477,N_385,N_339);
nor U478 (N_478,N_294,N_400);
nand U479 (N_479,N_407,N_402);
nor U480 (N_480,N_471,N_478);
or U481 (N_481,N_421,N_422);
and U482 (N_482,N_442,N_476);
nand U483 (N_483,N_463,N_459);
nand U484 (N_484,N_449,N_479);
nor U485 (N_485,N_420,N_434);
or U486 (N_486,N_433,N_461);
or U487 (N_487,N_438,N_429);
or U488 (N_488,N_445,N_423);
and U489 (N_489,N_444,N_439);
and U490 (N_490,N_460,N_435);
or U491 (N_491,N_456,N_452);
nor U492 (N_492,N_440,N_454);
or U493 (N_493,N_467,N_468);
nand U494 (N_494,N_441,N_472);
nand U495 (N_495,N_446,N_464);
and U496 (N_496,N_465,N_436);
nand U497 (N_497,N_432,N_425);
or U498 (N_498,N_437,N_457);
or U499 (N_499,N_475,N_469);
or U500 (N_500,N_426,N_443);
or U501 (N_501,N_424,N_428);
or U502 (N_502,N_448,N_427);
nand U503 (N_503,N_450,N_473);
or U504 (N_504,N_451,N_470);
nor U505 (N_505,N_430,N_453);
or U506 (N_506,N_462,N_431);
and U507 (N_507,N_477,N_455);
and U508 (N_508,N_466,N_474);
or U509 (N_509,N_458,N_447);
nand U510 (N_510,N_472,N_436);
nor U511 (N_511,N_430,N_460);
nand U512 (N_512,N_456,N_473);
or U513 (N_513,N_431,N_439);
nand U514 (N_514,N_435,N_438);
nand U515 (N_515,N_432,N_434);
or U516 (N_516,N_423,N_462);
nand U517 (N_517,N_450,N_479);
or U518 (N_518,N_446,N_448);
and U519 (N_519,N_475,N_454);
nor U520 (N_520,N_454,N_420);
and U521 (N_521,N_442,N_446);
and U522 (N_522,N_425,N_467);
nor U523 (N_523,N_432,N_423);
nand U524 (N_524,N_468,N_451);
and U525 (N_525,N_453,N_443);
nand U526 (N_526,N_437,N_478);
xor U527 (N_527,N_465,N_466);
and U528 (N_528,N_457,N_440);
and U529 (N_529,N_461,N_438);
or U530 (N_530,N_462,N_454);
nand U531 (N_531,N_427,N_445);
nor U532 (N_532,N_420,N_436);
or U533 (N_533,N_464,N_435);
nor U534 (N_534,N_425,N_470);
and U535 (N_535,N_453,N_474);
nand U536 (N_536,N_456,N_440);
nand U537 (N_537,N_448,N_456);
nor U538 (N_538,N_457,N_430);
and U539 (N_539,N_435,N_475);
or U540 (N_540,N_523,N_527);
or U541 (N_541,N_524,N_514);
or U542 (N_542,N_511,N_502);
nor U543 (N_543,N_533,N_530);
nand U544 (N_544,N_506,N_510);
nor U545 (N_545,N_499,N_495);
nor U546 (N_546,N_509,N_528);
and U547 (N_547,N_491,N_537);
and U548 (N_548,N_484,N_516);
nand U549 (N_549,N_515,N_517);
nor U550 (N_550,N_508,N_519);
and U551 (N_551,N_518,N_485);
nand U552 (N_552,N_481,N_494);
or U553 (N_553,N_513,N_534);
or U554 (N_554,N_525,N_531);
nand U555 (N_555,N_529,N_501);
or U556 (N_556,N_483,N_504);
or U557 (N_557,N_488,N_492);
or U558 (N_558,N_535,N_487);
and U559 (N_559,N_522,N_520);
or U560 (N_560,N_486,N_498);
or U561 (N_561,N_503,N_532);
or U562 (N_562,N_539,N_482);
nand U563 (N_563,N_496,N_521);
nand U564 (N_564,N_489,N_500);
and U565 (N_565,N_490,N_536);
nand U566 (N_566,N_507,N_497);
or U567 (N_567,N_526,N_538);
xnor U568 (N_568,N_512,N_505);
and U569 (N_569,N_480,N_493);
or U570 (N_570,N_484,N_525);
or U571 (N_571,N_498,N_494);
and U572 (N_572,N_513,N_527);
nand U573 (N_573,N_530,N_486);
and U574 (N_574,N_499,N_534);
nor U575 (N_575,N_512,N_533);
nand U576 (N_576,N_486,N_491);
nor U577 (N_577,N_493,N_498);
and U578 (N_578,N_522,N_489);
nand U579 (N_579,N_523,N_485);
or U580 (N_580,N_517,N_508);
nand U581 (N_581,N_518,N_496);
nor U582 (N_582,N_539,N_493);
or U583 (N_583,N_500,N_496);
nor U584 (N_584,N_531,N_530);
or U585 (N_585,N_503,N_523);
or U586 (N_586,N_515,N_490);
nor U587 (N_587,N_485,N_487);
or U588 (N_588,N_514,N_505);
or U589 (N_589,N_510,N_483);
or U590 (N_590,N_536,N_498);
nand U591 (N_591,N_483,N_497);
nand U592 (N_592,N_483,N_495);
or U593 (N_593,N_509,N_501);
or U594 (N_594,N_487,N_521);
nor U595 (N_595,N_480,N_483);
or U596 (N_596,N_516,N_487);
nor U597 (N_597,N_496,N_533);
or U598 (N_598,N_483,N_485);
and U599 (N_599,N_522,N_494);
nand U600 (N_600,N_583,N_582);
or U601 (N_601,N_590,N_555);
and U602 (N_602,N_553,N_549);
nand U603 (N_603,N_565,N_552);
nand U604 (N_604,N_543,N_569);
and U605 (N_605,N_542,N_566);
and U606 (N_606,N_570,N_563);
or U607 (N_607,N_598,N_581);
or U608 (N_608,N_548,N_562);
nor U609 (N_609,N_579,N_597);
nand U610 (N_610,N_574,N_587);
and U611 (N_611,N_547,N_594);
and U612 (N_612,N_558,N_573);
or U613 (N_613,N_545,N_564);
or U614 (N_614,N_592,N_585);
nand U615 (N_615,N_567,N_550);
or U616 (N_616,N_578,N_557);
nor U617 (N_617,N_540,N_560);
nand U618 (N_618,N_561,N_568);
nor U619 (N_619,N_577,N_589);
and U620 (N_620,N_596,N_595);
xnor U621 (N_621,N_593,N_580);
xor U622 (N_622,N_586,N_599);
nand U623 (N_623,N_571,N_559);
nand U624 (N_624,N_575,N_572);
xor U625 (N_625,N_546,N_554);
or U626 (N_626,N_551,N_591);
or U627 (N_627,N_541,N_584);
and U628 (N_628,N_544,N_556);
and U629 (N_629,N_576,N_588);
and U630 (N_630,N_558,N_549);
or U631 (N_631,N_565,N_591);
and U632 (N_632,N_599,N_591);
nor U633 (N_633,N_576,N_547);
or U634 (N_634,N_574,N_575);
or U635 (N_635,N_554,N_571);
nand U636 (N_636,N_546,N_541);
nand U637 (N_637,N_561,N_581);
nand U638 (N_638,N_587,N_589);
nor U639 (N_639,N_550,N_589);
and U640 (N_640,N_546,N_545);
or U641 (N_641,N_556,N_558);
nand U642 (N_642,N_571,N_573);
and U643 (N_643,N_586,N_593);
nor U644 (N_644,N_566,N_599);
nand U645 (N_645,N_556,N_563);
or U646 (N_646,N_576,N_585);
nor U647 (N_647,N_590,N_540);
nand U648 (N_648,N_588,N_578);
and U649 (N_649,N_596,N_574);
nor U650 (N_650,N_570,N_589);
xnor U651 (N_651,N_570,N_556);
and U652 (N_652,N_595,N_547);
nand U653 (N_653,N_564,N_586);
or U654 (N_654,N_552,N_582);
nand U655 (N_655,N_580,N_569);
nand U656 (N_656,N_546,N_562);
xnor U657 (N_657,N_553,N_589);
nor U658 (N_658,N_593,N_548);
and U659 (N_659,N_558,N_576);
or U660 (N_660,N_623,N_627);
nor U661 (N_661,N_644,N_653);
nor U662 (N_662,N_600,N_618);
nand U663 (N_663,N_659,N_621);
nand U664 (N_664,N_639,N_654);
and U665 (N_665,N_646,N_645);
nor U666 (N_666,N_640,N_652);
or U667 (N_667,N_603,N_614);
and U668 (N_668,N_615,N_636);
nand U669 (N_669,N_601,N_658);
nor U670 (N_670,N_657,N_610);
and U671 (N_671,N_642,N_602);
and U672 (N_672,N_638,N_648);
nor U673 (N_673,N_622,N_634);
or U674 (N_674,N_637,N_641);
nand U675 (N_675,N_606,N_650);
or U676 (N_676,N_605,N_629);
or U677 (N_677,N_647,N_649);
nand U678 (N_678,N_635,N_655);
and U679 (N_679,N_624,N_612);
nor U680 (N_680,N_643,N_651);
nand U681 (N_681,N_604,N_609);
and U682 (N_682,N_626,N_619);
nand U683 (N_683,N_625,N_608);
nor U684 (N_684,N_616,N_607);
and U685 (N_685,N_617,N_633);
nor U686 (N_686,N_611,N_631);
or U687 (N_687,N_632,N_628);
nor U688 (N_688,N_656,N_613);
nor U689 (N_689,N_630,N_620);
and U690 (N_690,N_616,N_634);
nand U691 (N_691,N_648,N_639);
nor U692 (N_692,N_622,N_638);
and U693 (N_693,N_604,N_641);
or U694 (N_694,N_611,N_658);
nand U695 (N_695,N_621,N_626);
nand U696 (N_696,N_603,N_606);
nor U697 (N_697,N_607,N_652);
or U698 (N_698,N_611,N_625);
or U699 (N_699,N_614,N_630);
nor U700 (N_700,N_644,N_641);
and U701 (N_701,N_620,N_638);
nor U702 (N_702,N_630,N_638);
nand U703 (N_703,N_627,N_642);
and U704 (N_704,N_631,N_601);
or U705 (N_705,N_629,N_606);
or U706 (N_706,N_649,N_602);
and U707 (N_707,N_618,N_628);
and U708 (N_708,N_612,N_602);
nand U709 (N_709,N_651,N_612);
nor U710 (N_710,N_640,N_641);
nor U711 (N_711,N_604,N_603);
and U712 (N_712,N_637,N_642);
nor U713 (N_713,N_645,N_607);
nor U714 (N_714,N_651,N_638);
or U715 (N_715,N_633,N_641);
nand U716 (N_716,N_637,N_640);
and U717 (N_717,N_615,N_641);
and U718 (N_718,N_600,N_648);
nand U719 (N_719,N_654,N_621);
nand U720 (N_720,N_711,N_705);
or U721 (N_721,N_685,N_674);
nand U722 (N_722,N_687,N_661);
nand U723 (N_723,N_664,N_701);
nand U724 (N_724,N_663,N_681);
or U725 (N_725,N_706,N_708);
nand U726 (N_726,N_678,N_700);
nor U727 (N_727,N_689,N_719);
nor U728 (N_728,N_703,N_688);
nand U729 (N_729,N_698,N_683);
nand U730 (N_730,N_668,N_699);
nand U731 (N_731,N_714,N_673);
nor U732 (N_732,N_695,N_670);
nor U733 (N_733,N_686,N_671);
nand U734 (N_734,N_694,N_680);
nand U735 (N_735,N_667,N_660);
nor U736 (N_736,N_677,N_690);
nand U737 (N_737,N_716,N_672);
xnor U738 (N_738,N_682,N_710);
or U739 (N_739,N_675,N_669);
nor U740 (N_740,N_709,N_665);
and U741 (N_741,N_707,N_704);
nor U742 (N_742,N_717,N_684);
nand U743 (N_743,N_712,N_715);
or U744 (N_744,N_702,N_662);
nor U745 (N_745,N_697,N_691);
nand U746 (N_746,N_713,N_666);
and U747 (N_747,N_692,N_676);
and U748 (N_748,N_718,N_679);
nor U749 (N_749,N_693,N_696);
or U750 (N_750,N_692,N_719);
nor U751 (N_751,N_712,N_664);
nor U752 (N_752,N_716,N_688);
or U753 (N_753,N_664,N_670);
nand U754 (N_754,N_717,N_695);
and U755 (N_755,N_673,N_694);
or U756 (N_756,N_690,N_707);
or U757 (N_757,N_665,N_688);
nand U758 (N_758,N_684,N_705);
nand U759 (N_759,N_687,N_710);
nand U760 (N_760,N_702,N_688);
and U761 (N_761,N_686,N_696);
xor U762 (N_762,N_678,N_688);
or U763 (N_763,N_707,N_709);
nor U764 (N_764,N_710,N_672);
nor U765 (N_765,N_661,N_678);
nand U766 (N_766,N_718,N_708);
and U767 (N_767,N_675,N_685);
nand U768 (N_768,N_685,N_673);
nand U769 (N_769,N_663,N_666);
or U770 (N_770,N_712,N_661);
nand U771 (N_771,N_681,N_719);
nor U772 (N_772,N_681,N_675);
or U773 (N_773,N_678,N_701);
nor U774 (N_774,N_677,N_667);
and U775 (N_775,N_684,N_710);
or U776 (N_776,N_662,N_663);
or U777 (N_777,N_703,N_697);
and U778 (N_778,N_715,N_664);
nor U779 (N_779,N_695,N_672);
nor U780 (N_780,N_763,N_731);
nor U781 (N_781,N_725,N_727);
and U782 (N_782,N_752,N_772);
xnor U783 (N_783,N_732,N_765);
or U784 (N_784,N_762,N_767);
or U785 (N_785,N_720,N_742);
nand U786 (N_786,N_743,N_773);
nand U787 (N_787,N_777,N_745);
nand U788 (N_788,N_747,N_761);
nor U789 (N_789,N_754,N_735);
nand U790 (N_790,N_751,N_755);
nand U791 (N_791,N_750,N_760);
nor U792 (N_792,N_723,N_768);
and U793 (N_793,N_729,N_771);
nand U794 (N_794,N_730,N_722);
nand U795 (N_795,N_733,N_721);
nor U796 (N_796,N_753,N_737);
nor U797 (N_797,N_728,N_756);
and U798 (N_798,N_758,N_770);
nand U799 (N_799,N_739,N_744);
or U800 (N_800,N_736,N_741);
and U801 (N_801,N_766,N_734);
nand U802 (N_802,N_778,N_749);
or U803 (N_803,N_779,N_748);
nand U804 (N_804,N_759,N_724);
or U805 (N_805,N_769,N_757);
nor U806 (N_806,N_776,N_746);
and U807 (N_807,N_738,N_764);
or U808 (N_808,N_726,N_774);
and U809 (N_809,N_775,N_740);
nor U810 (N_810,N_731,N_757);
or U811 (N_811,N_766,N_755);
nor U812 (N_812,N_726,N_739);
nand U813 (N_813,N_770,N_771);
or U814 (N_814,N_776,N_755);
or U815 (N_815,N_775,N_765);
and U816 (N_816,N_774,N_766);
and U817 (N_817,N_759,N_735);
nand U818 (N_818,N_726,N_737);
nor U819 (N_819,N_720,N_752);
and U820 (N_820,N_776,N_737);
nor U821 (N_821,N_740,N_732);
nor U822 (N_822,N_777,N_746);
and U823 (N_823,N_721,N_752);
nor U824 (N_824,N_740,N_769);
nand U825 (N_825,N_760,N_741);
nand U826 (N_826,N_764,N_756);
or U827 (N_827,N_722,N_741);
nand U828 (N_828,N_778,N_731);
nand U829 (N_829,N_745,N_778);
or U830 (N_830,N_772,N_773);
nor U831 (N_831,N_734,N_764);
and U832 (N_832,N_742,N_765);
nor U833 (N_833,N_728,N_748);
nor U834 (N_834,N_753,N_745);
and U835 (N_835,N_736,N_755);
nand U836 (N_836,N_743,N_728);
or U837 (N_837,N_734,N_721);
nand U838 (N_838,N_755,N_768);
nor U839 (N_839,N_726,N_779);
and U840 (N_840,N_830,N_828);
nand U841 (N_841,N_829,N_823);
or U842 (N_842,N_811,N_806);
nand U843 (N_843,N_785,N_827);
nand U844 (N_844,N_822,N_836);
nor U845 (N_845,N_839,N_789);
nor U846 (N_846,N_809,N_820);
nand U847 (N_847,N_804,N_791);
nand U848 (N_848,N_833,N_784);
and U849 (N_849,N_801,N_824);
and U850 (N_850,N_819,N_815);
nor U851 (N_851,N_788,N_810);
nor U852 (N_852,N_821,N_781);
nand U853 (N_853,N_816,N_818);
nand U854 (N_854,N_795,N_838);
nor U855 (N_855,N_790,N_796);
and U856 (N_856,N_800,N_812);
or U857 (N_857,N_783,N_805);
and U858 (N_858,N_834,N_835);
and U859 (N_859,N_782,N_794);
nand U860 (N_860,N_817,N_787);
and U861 (N_861,N_793,N_814);
and U862 (N_862,N_802,N_799);
and U863 (N_863,N_792,N_831);
nor U864 (N_864,N_807,N_797);
and U865 (N_865,N_826,N_798);
or U866 (N_866,N_808,N_825);
or U867 (N_867,N_780,N_832);
or U868 (N_868,N_803,N_837);
nor U869 (N_869,N_786,N_813);
nand U870 (N_870,N_813,N_816);
and U871 (N_871,N_786,N_826);
or U872 (N_872,N_812,N_838);
nand U873 (N_873,N_789,N_801);
nor U874 (N_874,N_794,N_809);
and U875 (N_875,N_793,N_819);
nor U876 (N_876,N_827,N_797);
and U877 (N_877,N_804,N_810);
or U878 (N_878,N_838,N_836);
nand U879 (N_879,N_817,N_819);
nand U880 (N_880,N_807,N_826);
nor U881 (N_881,N_805,N_797);
nand U882 (N_882,N_795,N_785);
and U883 (N_883,N_829,N_821);
or U884 (N_884,N_833,N_800);
and U885 (N_885,N_793,N_834);
nand U886 (N_886,N_820,N_832);
and U887 (N_887,N_835,N_829);
nand U888 (N_888,N_824,N_783);
nand U889 (N_889,N_817,N_831);
nand U890 (N_890,N_799,N_812);
nand U891 (N_891,N_801,N_799);
or U892 (N_892,N_832,N_788);
nand U893 (N_893,N_837,N_802);
and U894 (N_894,N_782,N_785);
nor U895 (N_895,N_829,N_813);
nor U896 (N_896,N_810,N_826);
nand U897 (N_897,N_823,N_787);
and U898 (N_898,N_823,N_800);
or U899 (N_899,N_836,N_796);
nor U900 (N_900,N_886,N_887);
or U901 (N_901,N_872,N_854);
and U902 (N_902,N_840,N_868);
and U903 (N_903,N_880,N_889);
or U904 (N_904,N_873,N_857);
nor U905 (N_905,N_848,N_897);
xor U906 (N_906,N_891,N_853);
nor U907 (N_907,N_885,N_883);
and U908 (N_908,N_850,N_879);
or U909 (N_909,N_866,N_855);
nor U910 (N_910,N_876,N_860);
and U911 (N_911,N_862,N_893);
nor U912 (N_912,N_843,N_852);
nand U913 (N_913,N_845,N_864);
and U914 (N_914,N_878,N_858);
nand U915 (N_915,N_898,N_875);
nor U916 (N_916,N_842,N_849);
nor U917 (N_917,N_881,N_884);
and U918 (N_918,N_890,N_859);
and U919 (N_919,N_882,N_899);
and U920 (N_920,N_844,N_869);
nor U921 (N_921,N_861,N_867);
nor U922 (N_922,N_895,N_874);
or U923 (N_923,N_888,N_863);
and U924 (N_924,N_896,N_877);
and U925 (N_925,N_851,N_871);
and U926 (N_926,N_894,N_865);
xnor U927 (N_927,N_841,N_892);
nand U928 (N_928,N_847,N_856);
nor U929 (N_929,N_870,N_846);
and U930 (N_930,N_870,N_856);
nand U931 (N_931,N_893,N_854);
nor U932 (N_932,N_877,N_887);
nand U933 (N_933,N_891,N_877);
or U934 (N_934,N_846,N_896);
nand U935 (N_935,N_844,N_861);
nor U936 (N_936,N_857,N_848);
nand U937 (N_937,N_865,N_890);
and U938 (N_938,N_841,N_854);
or U939 (N_939,N_855,N_882);
or U940 (N_940,N_878,N_862);
nor U941 (N_941,N_846,N_877);
xor U942 (N_942,N_873,N_854);
nand U943 (N_943,N_899,N_888);
or U944 (N_944,N_885,N_887);
nor U945 (N_945,N_853,N_884);
or U946 (N_946,N_857,N_884);
and U947 (N_947,N_850,N_887);
or U948 (N_948,N_850,N_888);
nor U949 (N_949,N_852,N_859);
and U950 (N_950,N_887,N_867);
or U951 (N_951,N_868,N_851);
or U952 (N_952,N_844,N_853);
and U953 (N_953,N_885,N_884);
and U954 (N_954,N_897,N_856);
nand U955 (N_955,N_884,N_887);
or U956 (N_956,N_857,N_892);
and U957 (N_957,N_859,N_848);
nand U958 (N_958,N_843,N_888);
or U959 (N_959,N_848,N_852);
nand U960 (N_960,N_934,N_956);
nand U961 (N_961,N_913,N_912);
and U962 (N_962,N_927,N_903);
and U963 (N_963,N_948,N_937);
nor U964 (N_964,N_944,N_914);
or U965 (N_965,N_920,N_946);
and U966 (N_966,N_929,N_923);
nor U967 (N_967,N_945,N_958);
nand U968 (N_968,N_917,N_959);
nand U969 (N_969,N_939,N_932);
and U970 (N_970,N_925,N_950);
or U971 (N_971,N_900,N_928);
or U972 (N_972,N_919,N_953);
nor U973 (N_973,N_915,N_911);
nor U974 (N_974,N_908,N_952);
and U975 (N_975,N_926,N_922);
nor U976 (N_976,N_940,N_951);
and U977 (N_977,N_954,N_942);
nand U978 (N_978,N_906,N_902);
nor U979 (N_979,N_957,N_930);
nor U980 (N_980,N_907,N_949);
or U981 (N_981,N_910,N_909);
nor U982 (N_982,N_943,N_941);
and U983 (N_983,N_933,N_901);
nand U984 (N_984,N_904,N_905);
or U985 (N_985,N_916,N_918);
or U986 (N_986,N_936,N_938);
and U987 (N_987,N_947,N_921);
and U988 (N_988,N_924,N_935);
and U989 (N_989,N_955,N_931);
and U990 (N_990,N_927,N_918);
and U991 (N_991,N_906,N_923);
nor U992 (N_992,N_959,N_912);
nand U993 (N_993,N_921,N_949);
or U994 (N_994,N_948,N_939);
nor U995 (N_995,N_917,N_924);
and U996 (N_996,N_912,N_924);
nand U997 (N_997,N_934,N_952);
or U998 (N_998,N_944,N_931);
xor U999 (N_999,N_940,N_932);
or U1000 (N_1000,N_938,N_952);
and U1001 (N_1001,N_916,N_912);
and U1002 (N_1002,N_947,N_952);
nor U1003 (N_1003,N_928,N_919);
nand U1004 (N_1004,N_927,N_921);
and U1005 (N_1005,N_941,N_909);
and U1006 (N_1006,N_952,N_953);
nor U1007 (N_1007,N_956,N_939);
nor U1008 (N_1008,N_920,N_901);
nor U1009 (N_1009,N_926,N_958);
nand U1010 (N_1010,N_918,N_923);
nand U1011 (N_1011,N_904,N_906);
nand U1012 (N_1012,N_907,N_939);
or U1013 (N_1013,N_959,N_945);
nor U1014 (N_1014,N_929,N_932);
nor U1015 (N_1015,N_929,N_928);
or U1016 (N_1016,N_951,N_948);
or U1017 (N_1017,N_955,N_922);
nor U1018 (N_1018,N_921,N_932);
and U1019 (N_1019,N_958,N_901);
and U1020 (N_1020,N_990,N_1004);
and U1021 (N_1021,N_992,N_997);
nor U1022 (N_1022,N_979,N_1015);
nand U1023 (N_1023,N_1006,N_1017);
nand U1024 (N_1024,N_1009,N_975);
or U1025 (N_1025,N_999,N_1012);
or U1026 (N_1026,N_989,N_1007);
nand U1027 (N_1027,N_985,N_967);
nand U1028 (N_1028,N_986,N_1010);
or U1029 (N_1029,N_974,N_973);
and U1030 (N_1030,N_1008,N_977);
nor U1031 (N_1031,N_981,N_1016);
nor U1032 (N_1032,N_1001,N_998);
and U1033 (N_1033,N_1000,N_980);
or U1034 (N_1034,N_963,N_961);
or U1035 (N_1035,N_972,N_994);
nand U1036 (N_1036,N_983,N_996);
nand U1037 (N_1037,N_1011,N_987);
nand U1038 (N_1038,N_995,N_984);
nand U1039 (N_1039,N_968,N_1005);
and U1040 (N_1040,N_993,N_991);
nand U1041 (N_1041,N_1018,N_964);
and U1042 (N_1042,N_965,N_969);
or U1043 (N_1043,N_966,N_1014);
and U1044 (N_1044,N_982,N_1019);
nand U1045 (N_1045,N_970,N_962);
nand U1046 (N_1046,N_1013,N_960);
and U1047 (N_1047,N_976,N_1003);
nand U1048 (N_1048,N_971,N_988);
and U1049 (N_1049,N_978,N_1002);
and U1050 (N_1050,N_996,N_986);
nand U1051 (N_1051,N_992,N_995);
and U1052 (N_1052,N_991,N_1013);
nand U1053 (N_1053,N_996,N_1011);
or U1054 (N_1054,N_1001,N_1003);
and U1055 (N_1055,N_970,N_1015);
or U1056 (N_1056,N_994,N_1017);
nor U1057 (N_1057,N_989,N_1014);
nand U1058 (N_1058,N_1012,N_1015);
nor U1059 (N_1059,N_968,N_1007);
nor U1060 (N_1060,N_1001,N_992);
or U1061 (N_1061,N_971,N_998);
or U1062 (N_1062,N_968,N_991);
nand U1063 (N_1063,N_978,N_1009);
and U1064 (N_1064,N_963,N_988);
nor U1065 (N_1065,N_989,N_988);
and U1066 (N_1066,N_976,N_974);
or U1067 (N_1067,N_1007,N_965);
and U1068 (N_1068,N_1000,N_978);
nand U1069 (N_1069,N_1014,N_974);
nor U1070 (N_1070,N_1001,N_1013);
nor U1071 (N_1071,N_983,N_978);
nor U1072 (N_1072,N_976,N_975);
nand U1073 (N_1073,N_1018,N_967);
and U1074 (N_1074,N_981,N_964);
or U1075 (N_1075,N_963,N_982);
and U1076 (N_1076,N_1011,N_976);
or U1077 (N_1077,N_971,N_1007);
and U1078 (N_1078,N_996,N_990);
nor U1079 (N_1079,N_1016,N_964);
nand U1080 (N_1080,N_1030,N_1038);
nor U1081 (N_1081,N_1071,N_1064);
or U1082 (N_1082,N_1058,N_1070);
nand U1083 (N_1083,N_1078,N_1039);
nand U1084 (N_1084,N_1066,N_1056);
or U1085 (N_1085,N_1057,N_1027);
nand U1086 (N_1086,N_1077,N_1046);
nand U1087 (N_1087,N_1052,N_1065);
nand U1088 (N_1088,N_1026,N_1075);
or U1089 (N_1089,N_1048,N_1049);
nand U1090 (N_1090,N_1069,N_1032);
nand U1091 (N_1091,N_1031,N_1061);
and U1092 (N_1092,N_1047,N_1053);
and U1093 (N_1093,N_1054,N_1040);
nand U1094 (N_1094,N_1074,N_1028);
and U1095 (N_1095,N_1036,N_1062);
and U1096 (N_1096,N_1073,N_1037);
nand U1097 (N_1097,N_1042,N_1024);
or U1098 (N_1098,N_1072,N_1033);
nand U1099 (N_1099,N_1079,N_1020);
nand U1100 (N_1100,N_1045,N_1067);
and U1101 (N_1101,N_1044,N_1055);
nand U1102 (N_1102,N_1050,N_1025);
nor U1103 (N_1103,N_1068,N_1043);
nand U1104 (N_1104,N_1041,N_1060);
and U1105 (N_1105,N_1022,N_1063);
nor U1106 (N_1106,N_1076,N_1021);
nand U1107 (N_1107,N_1035,N_1023);
or U1108 (N_1108,N_1059,N_1034);
nand U1109 (N_1109,N_1029,N_1051);
nand U1110 (N_1110,N_1030,N_1036);
or U1111 (N_1111,N_1076,N_1065);
and U1112 (N_1112,N_1066,N_1023);
and U1113 (N_1113,N_1021,N_1078);
or U1114 (N_1114,N_1078,N_1049);
nand U1115 (N_1115,N_1032,N_1049);
or U1116 (N_1116,N_1064,N_1054);
nor U1117 (N_1117,N_1066,N_1073);
nor U1118 (N_1118,N_1036,N_1041);
and U1119 (N_1119,N_1068,N_1031);
nor U1120 (N_1120,N_1043,N_1027);
nand U1121 (N_1121,N_1029,N_1042);
and U1122 (N_1122,N_1049,N_1046);
or U1123 (N_1123,N_1048,N_1075);
or U1124 (N_1124,N_1071,N_1079);
or U1125 (N_1125,N_1044,N_1027);
nand U1126 (N_1126,N_1035,N_1068);
nand U1127 (N_1127,N_1043,N_1040);
or U1128 (N_1128,N_1052,N_1071);
and U1129 (N_1129,N_1043,N_1030);
and U1130 (N_1130,N_1033,N_1077);
and U1131 (N_1131,N_1060,N_1067);
nand U1132 (N_1132,N_1065,N_1044);
nand U1133 (N_1133,N_1076,N_1070);
nand U1134 (N_1134,N_1024,N_1032);
and U1135 (N_1135,N_1059,N_1063);
and U1136 (N_1136,N_1023,N_1058);
and U1137 (N_1137,N_1066,N_1060);
nand U1138 (N_1138,N_1062,N_1067);
or U1139 (N_1139,N_1073,N_1033);
and U1140 (N_1140,N_1132,N_1115);
or U1141 (N_1141,N_1121,N_1105);
nand U1142 (N_1142,N_1107,N_1096);
and U1143 (N_1143,N_1125,N_1129);
and U1144 (N_1144,N_1093,N_1137);
nand U1145 (N_1145,N_1110,N_1084);
nand U1146 (N_1146,N_1123,N_1081);
nand U1147 (N_1147,N_1091,N_1131);
nor U1148 (N_1148,N_1130,N_1124);
or U1149 (N_1149,N_1101,N_1102);
and U1150 (N_1150,N_1111,N_1094);
or U1151 (N_1151,N_1117,N_1128);
or U1152 (N_1152,N_1126,N_1095);
nand U1153 (N_1153,N_1106,N_1089);
nor U1154 (N_1154,N_1138,N_1136);
or U1155 (N_1155,N_1112,N_1109);
and U1156 (N_1156,N_1139,N_1085);
or U1157 (N_1157,N_1099,N_1087);
and U1158 (N_1158,N_1113,N_1098);
nor U1159 (N_1159,N_1100,N_1083);
nand U1160 (N_1160,N_1103,N_1088);
nand U1161 (N_1161,N_1118,N_1090);
nand U1162 (N_1162,N_1120,N_1133);
nand U1163 (N_1163,N_1134,N_1114);
or U1164 (N_1164,N_1080,N_1116);
nor U1165 (N_1165,N_1082,N_1104);
nand U1166 (N_1166,N_1127,N_1135);
nor U1167 (N_1167,N_1119,N_1097);
and U1168 (N_1168,N_1092,N_1122);
nand U1169 (N_1169,N_1108,N_1086);
or U1170 (N_1170,N_1102,N_1115);
xnor U1171 (N_1171,N_1117,N_1093);
or U1172 (N_1172,N_1132,N_1139);
or U1173 (N_1173,N_1087,N_1115);
xnor U1174 (N_1174,N_1089,N_1135);
and U1175 (N_1175,N_1113,N_1136);
nand U1176 (N_1176,N_1096,N_1125);
or U1177 (N_1177,N_1106,N_1102);
nor U1178 (N_1178,N_1106,N_1095);
nor U1179 (N_1179,N_1134,N_1109);
nor U1180 (N_1180,N_1125,N_1091);
xnor U1181 (N_1181,N_1084,N_1112);
or U1182 (N_1182,N_1138,N_1117);
or U1183 (N_1183,N_1090,N_1128);
nor U1184 (N_1184,N_1137,N_1132);
and U1185 (N_1185,N_1094,N_1100);
nand U1186 (N_1186,N_1130,N_1118);
nor U1187 (N_1187,N_1112,N_1095);
nand U1188 (N_1188,N_1082,N_1095);
nor U1189 (N_1189,N_1101,N_1129);
nand U1190 (N_1190,N_1094,N_1139);
and U1191 (N_1191,N_1116,N_1119);
and U1192 (N_1192,N_1117,N_1134);
or U1193 (N_1193,N_1118,N_1120);
and U1194 (N_1194,N_1118,N_1083);
and U1195 (N_1195,N_1133,N_1137);
nor U1196 (N_1196,N_1090,N_1108);
or U1197 (N_1197,N_1106,N_1104);
and U1198 (N_1198,N_1121,N_1088);
or U1199 (N_1199,N_1116,N_1113);
nand U1200 (N_1200,N_1184,N_1169);
and U1201 (N_1201,N_1186,N_1148);
and U1202 (N_1202,N_1187,N_1146);
nor U1203 (N_1203,N_1178,N_1190);
and U1204 (N_1204,N_1156,N_1185);
nand U1205 (N_1205,N_1142,N_1155);
nor U1206 (N_1206,N_1168,N_1177);
nand U1207 (N_1207,N_1152,N_1188);
and U1208 (N_1208,N_1163,N_1164);
and U1209 (N_1209,N_1165,N_1183);
nor U1210 (N_1210,N_1189,N_1154);
or U1211 (N_1211,N_1167,N_1161);
nand U1212 (N_1212,N_1176,N_1196);
and U1213 (N_1213,N_1150,N_1174);
and U1214 (N_1214,N_1149,N_1172);
nor U1215 (N_1215,N_1140,N_1193);
nand U1216 (N_1216,N_1141,N_1143);
and U1217 (N_1217,N_1181,N_1173);
nand U1218 (N_1218,N_1157,N_1199);
nor U1219 (N_1219,N_1198,N_1194);
nor U1220 (N_1220,N_1151,N_1170);
nor U1221 (N_1221,N_1147,N_1144);
and U1222 (N_1222,N_1160,N_1179);
and U1223 (N_1223,N_1197,N_1153);
and U1224 (N_1224,N_1159,N_1192);
nor U1225 (N_1225,N_1182,N_1166);
nand U1226 (N_1226,N_1195,N_1180);
nor U1227 (N_1227,N_1162,N_1158);
nor U1228 (N_1228,N_1171,N_1191);
nor U1229 (N_1229,N_1175,N_1145);
nand U1230 (N_1230,N_1180,N_1185);
or U1231 (N_1231,N_1141,N_1183);
and U1232 (N_1232,N_1185,N_1175);
nand U1233 (N_1233,N_1182,N_1184);
nand U1234 (N_1234,N_1168,N_1186);
or U1235 (N_1235,N_1188,N_1161);
nand U1236 (N_1236,N_1184,N_1153);
and U1237 (N_1237,N_1142,N_1179);
nor U1238 (N_1238,N_1167,N_1190);
or U1239 (N_1239,N_1175,N_1163);
nor U1240 (N_1240,N_1171,N_1168);
nor U1241 (N_1241,N_1143,N_1169);
nand U1242 (N_1242,N_1191,N_1157);
and U1243 (N_1243,N_1190,N_1195);
and U1244 (N_1244,N_1176,N_1148);
nor U1245 (N_1245,N_1186,N_1167);
or U1246 (N_1246,N_1151,N_1149);
and U1247 (N_1247,N_1181,N_1179);
xnor U1248 (N_1248,N_1191,N_1178);
and U1249 (N_1249,N_1164,N_1160);
nor U1250 (N_1250,N_1163,N_1182);
or U1251 (N_1251,N_1179,N_1143);
nand U1252 (N_1252,N_1194,N_1149);
or U1253 (N_1253,N_1161,N_1171);
nor U1254 (N_1254,N_1162,N_1161);
nand U1255 (N_1255,N_1154,N_1147);
or U1256 (N_1256,N_1154,N_1142);
nor U1257 (N_1257,N_1142,N_1171);
nand U1258 (N_1258,N_1183,N_1163);
and U1259 (N_1259,N_1174,N_1166);
and U1260 (N_1260,N_1214,N_1243);
and U1261 (N_1261,N_1259,N_1210);
nor U1262 (N_1262,N_1247,N_1205);
nor U1263 (N_1263,N_1229,N_1213);
xor U1264 (N_1264,N_1246,N_1217);
nand U1265 (N_1265,N_1258,N_1234);
or U1266 (N_1266,N_1225,N_1254);
nor U1267 (N_1267,N_1204,N_1220);
nor U1268 (N_1268,N_1226,N_1222);
or U1269 (N_1269,N_1218,N_1251);
nand U1270 (N_1270,N_1212,N_1202);
nor U1271 (N_1271,N_1232,N_1245);
or U1272 (N_1272,N_1227,N_1242);
nor U1273 (N_1273,N_1241,N_1253);
nand U1274 (N_1274,N_1211,N_1244);
nor U1275 (N_1275,N_1200,N_1224);
nand U1276 (N_1276,N_1228,N_1206);
nor U1277 (N_1277,N_1256,N_1209);
or U1278 (N_1278,N_1221,N_1231);
nand U1279 (N_1279,N_1255,N_1257);
or U1280 (N_1280,N_1203,N_1207);
nand U1281 (N_1281,N_1238,N_1230);
nor U1282 (N_1282,N_1201,N_1250);
nand U1283 (N_1283,N_1233,N_1248);
nand U1284 (N_1284,N_1239,N_1216);
or U1285 (N_1285,N_1240,N_1208);
and U1286 (N_1286,N_1223,N_1215);
or U1287 (N_1287,N_1236,N_1219);
or U1288 (N_1288,N_1237,N_1252);
or U1289 (N_1289,N_1249,N_1235);
nor U1290 (N_1290,N_1247,N_1232);
nor U1291 (N_1291,N_1225,N_1235);
or U1292 (N_1292,N_1207,N_1257);
or U1293 (N_1293,N_1223,N_1234);
and U1294 (N_1294,N_1231,N_1254);
and U1295 (N_1295,N_1222,N_1238);
nor U1296 (N_1296,N_1255,N_1245);
or U1297 (N_1297,N_1251,N_1253);
or U1298 (N_1298,N_1230,N_1220);
nand U1299 (N_1299,N_1241,N_1213);
nand U1300 (N_1300,N_1255,N_1211);
and U1301 (N_1301,N_1207,N_1227);
nor U1302 (N_1302,N_1234,N_1218);
and U1303 (N_1303,N_1237,N_1226);
or U1304 (N_1304,N_1234,N_1237);
or U1305 (N_1305,N_1215,N_1256);
or U1306 (N_1306,N_1225,N_1237);
or U1307 (N_1307,N_1210,N_1221);
and U1308 (N_1308,N_1224,N_1245);
nor U1309 (N_1309,N_1232,N_1215);
nand U1310 (N_1310,N_1226,N_1245);
or U1311 (N_1311,N_1225,N_1221);
or U1312 (N_1312,N_1222,N_1241);
and U1313 (N_1313,N_1256,N_1228);
nand U1314 (N_1314,N_1204,N_1247);
and U1315 (N_1315,N_1228,N_1216);
and U1316 (N_1316,N_1239,N_1224);
nand U1317 (N_1317,N_1243,N_1236);
nand U1318 (N_1318,N_1222,N_1259);
nand U1319 (N_1319,N_1234,N_1246);
nand U1320 (N_1320,N_1274,N_1273);
and U1321 (N_1321,N_1264,N_1285);
nor U1322 (N_1322,N_1265,N_1302);
nand U1323 (N_1323,N_1315,N_1313);
or U1324 (N_1324,N_1299,N_1288);
or U1325 (N_1325,N_1270,N_1303);
and U1326 (N_1326,N_1287,N_1271);
nand U1327 (N_1327,N_1283,N_1298);
or U1328 (N_1328,N_1279,N_1275);
nand U1329 (N_1329,N_1304,N_1294);
nand U1330 (N_1330,N_1295,N_1289);
nor U1331 (N_1331,N_1291,N_1307);
nand U1332 (N_1332,N_1293,N_1286);
nand U1333 (N_1333,N_1319,N_1300);
nand U1334 (N_1334,N_1284,N_1260);
and U1335 (N_1335,N_1268,N_1308);
or U1336 (N_1336,N_1282,N_1301);
or U1337 (N_1337,N_1309,N_1276);
or U1338 (N_1338,N_1281,N_1312);
or U1339 (N_1339,N_1292,N_1261);
nor U1340 (N_1340,N_1266,N_1297);
nor U1341 (N_1341,N_1314,N_1263);
nand U1342 (N_1342,N_1311,N_1305);
or U1343 (N_1343,N_1318,N_1306);
and U1344 (N_1344,N_1267,N_1269);
nor U1345 (N_1345,N_1296,N_1316);
and U1346 (N_1346,N_1280,N_1290);
nand U1347 (N_1347,N_1317,N_1278);
nor U1348 (N_1348,N_1272,N_1310);
nor U1349 (N_1349,N_1277,N_1262);
xnor U1350 (N_1350,N_1263,N_1291);
or U1351 (N_1351,N_1287,N_1280);
nor U1352 (N_1352,N_1302,N_1262);
and U1353 (N_1353,N_1315,N_1317);
and U1354 (N_1354,N_1290,N_1312);
or U1355 (N_1355,N_1310,N_1262);
nand U1356 (N_1356,N_1263,N_1283);
or U1357 (N_1357,N_1310,N_1287);
nand U1358 (N_1358,N_1266,N_1309);
nor U1359 (N_1359,N_1270,N_1279);
nand U1360 (N_1360,N_1266,N_1265);
or U1361 (N_1361,N_1262,N_1279);
and U1362 (N_1362,N_1310,N_1280);
and U1363 (N_1363,N_1307,N_1295);
or U1364 (N_1364,N_1271,N_1284);
or U1365 (N_1365,N_1317,N_1281);
nor U1366 (N_1366,N_1311,N_1266);
and U1367 (N_1367,N_1311,N_1273);
nand U1368 (N_1368,N_1287,N_1297);
nor U1369 (N_1369,N_1286,N_1297);
nand U1370 (N_1370,N_1280,N_1302);
or U1371 (N_1371,N_1275,N_1267);
nor U1372 (N_1372,N_1308,N_1302);
and U1373 (N_1373,N_1268,N_1260);
nand U1374 (N_1374,N_1297,N_1313);
nand U1375 (N_1375,N_1308,N_1307);
or U1376 (N_1376,N_1296,N_1270);
nor U1377 (N_1377,N_1270,N_1289);
or U1378 (N_1378,N_1266,N_1260);
nor U1379 (N_1379,N_1261,N_1313);
and U1380 (N_1380,N_1366,N_1354);
nand U1381 (N_1381,N_1369,N_1359);
nor U1382 (N_1382,N_1353,N_1374);
nor U1383 (N_1383,N_1363,N_1378);
and U1384 (N_1384,N_1348,N_1325);
nand U1385 (N_1385,N_1330,N_1364);
nand U1386 (N_1386,N_1341,N_1371);
nand U1387 (N_1387,N_1332,N_1376);
nor U1388 (N_1388,N_1343,N_1338);
nor U1389 (N_1389,N_1362,N_1334);
and U1390 (N_1390,N_1361,N_1368);
nor U1391 (N_1391,N_1352,N_1367);
nor U1392 (N_1392,N_1351,N_1349);
nand U1393 (N_1393,N_1347,N_1339);
and U1394 (N_1394,N_1337,N_1356);
or U1395 (N_1395,N_1344,N_1370);
and U1396 (N_1396,N_1379,N_1346);
nand U1397 (N_1397,N_1342,N_1324);
or U1398 (N_1398,N_1357,N_1328);
nand U1399 (N_1399,N_1326,N_1336);
nor U1400 (N_1400,N_1323,N_1321);
or U1401 (N_1401,N_1320,N_1350);
and U1402 (N_1402,N_1329,N_1322);
or U1403 (N_1403,N_1373,N_1375);
nand U1404 (N_1404,N_1358,N_1335);
nand U1405 (N_1405,N_1340,N_1377);
nor U1406 (N_1406,N_1360,N_1355);
or U1407 (N_1407,N_1365,N_1327);
or U1408 (N_1408,N_1333,N_1331);
nand U1409 (N_1409,N_1345,N_1372);
nand U1410 (N_1410,N_1378,N_1333);
and U1411 (N_1411,N_1376,N_1333);
nand U1412 (N_1412,N_1345,N_1323);
and U1413 (N_1413,N_1370,N_1367);
or U1414 (N_1414,N_1368,N_1359);
or U1415 (N_1415,N_1371,N_1362);
or U1416 (N_1416,N_1371,N_1323);
and U1417 (N_1417,N_1323,N_1354);
and U1418 (N_1418,N_1372,N_1375);
and U1419 (N_1419,N_1374,N_1376);
and U1420 (N_1420,N_1375,N_1344);
or U1421 (N_1421,N_1338,N_1340);
or U1422 (N_1422,N_1358,N_1362);
and U1423 (N_1423,N_1342,N_1328);
nand U1424 (N_1424,N_1322,N_1366);
nor U1425 (N_1425,N_1334,N_1349);
or U1426 (N_1426,N_1371,N_1334);
nor U1427 (N_1427,N_1339,N_1333);
nand U1428 (N_1428,N_1335,N_1342);
and U1429 (N_1429,N_1342,N_1347);
nand U1430 (N_1430,N_1377,N_1336);
nor U1431 (N_1431,N_1340,N_1348);
and U1432 (N_1432,N_1367,N_1376);
nor U1433 (N_1433,N_1343,N_1349);
or U1434 (N_1434,N_1322,N_1365);
nand U1435 (N_1435,N_1363,N_1323);
nor U1436 (N_1436,N_1375,N_1334);
nor U1437 (N_1437,N_1364,N_1352);
nor U1438 (N_1438,N_1327,N_1368);
nand U1439 (N_1439,N_1363,N_1347);
and U1440 (N_1440,N_1417,N_1382);
nand U1441 (N_1441,N_1432,N_1409);
nor U1442 (N_1442,N_1391,N_1429);
or U1443 (N_1443,N_1410,N_1386);
and U1444 (N_1444,N_1396,N_1383);
and U1445 (N_1445,N_1423,N_1392);
or U1446 (N_1446,N_1404,N_1439);
nor U1447 (N_1447,N_1416,N_1435);
or U1448 (N_1448,N_1437,N_1394);
or U1449 (N_1449,N_1415,N_1414);
or U1450 (N_1450,N_1433,N_1436);
or U1451 (N_1451,N_1434,N_1395);
or U1452 (N_1452,N_1398,N_1400);
nor U1453 (N_1453,N_1390,N_1402);
and U1454 (N_1454,N_1389,N_1425);
nor U1455 (N_1455,N_1422,N_1418);
or U1456 (N_1456,N_1403,N_1399);
nand U1457 (N_1457,N_1424,N_1385);
nand U1458 (N_1458,N_1438,N_1420);
and U1459 (N_1459,N_1388,N_1407);
nor U1460 (N_1460,N_1405,N_1381);
or U1461 (N_1461,N_1397,N_1428);
nor U1462 (N_1462,N_1406,N_1408);
or U1463 (N_1463,N_1401,N_1380);
or U1464 (N_1464,N_1413,N_1412);
and U1465 (N_1465,N_1421,N_1387);
nand U1466 (N_1466,N_1419,N_1431);
nand U1467 (N_1467,N_1393,N_1430);
nor U1468 (N_1468,N_1427,N_1411);
and U1469 (N_1469,N_1426,N_1384);
nor U1470 (N_1470,N_1400,N_1411);
nor U1471 (N_1471,N_1388,N_1436);
nor U1472 (N_1472,N_1399,N_1392);
nand U1473 (N_1473,N_1430,N_1383);
nand U1474 (N_1474,N_1433,N_1413);
and U1475 (N_1475,N_1390,N_1407);
nand U1476 (N_1476,N_1408,N_1433);
and U1477 (N_1477,N_1387,N_1418);
and U1478 (N_1478,N_1428,N_1415);
and U1479 (N_1479,N_1395,N_1420);
nand U1480 (N_1480,N_1428,N_1416);
and U1481 (N_1481,N_1386,N_1427);
nor U1482 (N_1482,N_1389,N_1407);
nor U1483 (N_1483,N_1422,N_1430);
or U1484 (N_1484,N_1384,N_1437);
and U1485 (N_1485,N_1401,N_1404);
and U1486 (N_1486,N_1433,N_1400);
or U1487 (N_1487,N_1414,N_1409);
or U1488 (N_1488,N_1435,N_1422);
nor U1489 (N_1489,N_1390,N_1391);
nor U1490 (N_1490,N_1385,N_1429);
nor U1491 (N_1491,N_1427,N_1407);
nand U1492 (N_1492,N_1427,N_1387);
nand U1493 (N_1493,N_1408,N_1424);
nand U1494 (N_1494,N_1383,N_1421);
or U1495 (N_1495,N_1394,N_1424);
nor U1496 (N_1496,N_1399,N_1439);
or U1497 (N_1497,N_1437,N_1403);
and U1498 (N_1498,N_1415,N_1393);
and U1499 (N_1499,N_1427,N_1396);
or U1500 (N_1500,N_1451,N_1445);
nor U1501 (N_1501,N_1481,N_1479);
or U1502 (N_1502,N_1462,N_1467);
and U1503 (N_1503,N_1474,N_1449);
or U1504 (N_1504,N_1485,N_1484);
nor U1505 (N_1505,N_1483,N_1450);
nand U1506 (N_1506,N_1459,N_1453);
nor U1507 (N_1507,N_1468,N_1442);
or U1508 (N_1508,N_1480,N_1487);
nor U1509 (N_1509,N_1497,N_1454);
and U1510 (N_1510,N_1471,N_1495);
and U1511 (N_1511,N_1457,N_1444);
nand U1512 (N_1512,N_1490,N_1498);
or U1513 (N_1513,N_1461,N_1456);
nand U1514 (N_1514,N_1488,N_1469);
and U1515 (N_1515,N_1478,N_1470);
nor U1516 (N_1516,N_1472,N_1443);
or U1517 (N_1517,N_1473,N_1463);
or U1518 (N_1518,N_1460,N_1499);
and U1519 (N_1519,N_1477,N_1493);
and U1520 (N_1520,N_1446,N_1447);
and U1521 (N_1521,N_1441,N_1491);
nand U1522 (N_1522,N_1489,N_1466);
nor U1523 (N_1523,N_1475,N_1448);
nand U1524 (N_1524,N_1476,N_1494);
nand U1525 (N_1525,N_1464,N_1482);
nand U1526 (N_1526,N_1465,N_1496);
nor U1527 (N_1527,N_1486,N_1492);
or U1528 (N_1528,N_1440,N_1458);
and U1529 (N_1529,N_1455,N_1452);
nand U1530 (N_1530,N_1475,N_1479);
or U1531 (N_1531,N_1441,N_1472);
and U1532 (N_1532,N_1454,N_1467);
or U1533 (N_1533,N_1458,N_1454);
xnor U1534 (N_1534,N_1479,N_1461);
and U1535 (N_1535,N_1492,N_1484);
nor U1536 (N_1536,N_1442,N_1494);
nand U1537 (N_1537,N_1466,N_1497);
nand U1538 (N_1538,N_1471,N_1442);
nand U1539 (N_1539,N_1473,N_1487);
nor U1540 (N_1540,N_1466,N_1485);
nor U1541 (N_1541,N_1440,N_1442);
nor U1542 (N_1542,N_1494,N_1457);
and U1543 (N_1543,N_1447,N_1499);
nand U1544 (N_1544,N_1498,N_1467);
or U1545 (N_1545,N_1497,N_1493);
nor U1546 (N_1546,N_1489,N_1463);
or U1547 (N_1547,N_1480,N_1448);
nor U1548 (N_1548,N_1464,N_1489);
nand U1549 (N_1549,N_1498,N_1453);
nand U1550 (N_1550,N_1480,N_1457);
and U1551 (N_1551,N_1488,N_1475);
or U1552 (N_1552,N_1462,N_1441);
or U1553 (N_1553,N_1457,N_1487);
or U1554 (N_1554,N_1451,N_1489);
and U1555 (N_1555,N_1470,N_1451);
and U1556 (N_1556,N_1463,N_1498);
and U1557 (N_1557,N_1494,N_1498);
and U1558 (N_1558,N_1477,N_1495);
or U1559 (N_1559,N_1473,N_1482);
nand U1560 (N_1560,N_1515,N_1513);
nand U1561 (N_1561,N_1507,N_1528);
and U1562 (N_1562,N_1521,N_1558);
or U1563 (N_1563,N_1542,N_1520);
and U1564 (N_1564,N_1554,N_1559);
nor U1565 (N_1565,N_1533,N_1556);
and U1566 (N_1566,N_1534,N_1510);
or U1567 (N_1567,N_1553,N_1555);
and U1568 (N_1568,N_1536,N_1509);
nor U1569 (N_1569,N_1547,N_1522);
nor U1570 (N_1570,N_1504,N_1508);
and U1571 (N_1571,N_1530,N_1527);
nand U1572 (N_1572,N_1548,N_1514);
xnor U1573 (N_1573,N_1501,N_1538);
nor U1574 (N_1574,N_1525,N_1552);
nor U1575 (N_1575,N_1535,N_1531);
and U1576 (N_1576,N_1537,N_1506);
nor U1577 (N_1577,N_1546,N_1512);
or U1578 (N_1578,N_1526,N_1545);
nand U1579 (N_1579,N_1519,N_1540);
nand U1580 (N_1580,N_1539,N_1550);
nand U1581 (N_1581,N_1524,N_1523);
nor U1582 (N_1582,N_1505,N_1511);
nand U1583 (N_1583,N_1541,N_1557);
nand U1584 (N_1584,N_1551,N_1518);
nor U1585 (N_1585,N_1544,N_1529);
nand U1586 (N_1586,N_1532,N_1500);
or U1587 (N_1587,N_1516,N_1503);
and U1588 (N_1588,N_1543,N_1502);
nor U1589 (N_1589,N_1549,N_1517);
or U1590 (N_1590,N_1528,N_1529);
nand U1591 (N_1591,N_1543,N_1544);
or U1592 (N_1592,N_1557,N_1544);
nand U1593 (N_1593,N_1549,N_1542);
or U1594 (N_1594,N_1516,N_1542);
and U1595 (N_1595,N_1535,N_1504);
or U1596 (N_1596,N_1544,N_1552);
nor U1597 (N_1597,N_1556,N_1547);
or U1598 (N_1598,N_1511,N_1504);
nand U1599 (N_1599,N_1504,N_1555);
nor U1600 (N_1600,N_1543,N_1554);
nor U1601 (N_1601,N_1521,N_1537);
nor U1602 (N_1602,N_1543,N_1532);
nor U1603 (N_1603,N_1552,N_1507);
and U1604 (N_1604,N_1531,N_1505);
nor U1605 (N_1605,N_1528,N_1527);
nor U1606 (N_1606,N_1524,N_1510);
nor U1607 (N_1607,N_1558,N_1525);
and U1608 (N_1608,N_1521,N_1517);
and U1609 (N_1609,N_1525,N_1532);
and U1610 (N_1610,N_1530,N_1542);
or U1611 (N_1611,N_1521,N_1534);
and U1612 (N_1612,N_1532,N_1521);
nor U1613 (N_1613,N_1543,N_1551);
nor U1614 (N_1614,N_1500,N_1520);
nand U1615 (N_1615,N_1515,N_1557);
nand U1616 (N_1616,N_1533,N_1506);
or U1617 (N_1617,N_1529,N_1547);
and U1618 (N_1618,N_1557,N_1555);
nand U1619 (N_1619,N_1545,N_1512);
nor U1620 (N_1620,N_1613,N_1608);
and U1621 (N_1621,N_1609,N_1584);
and U1622 (N_1622,N_1617,N_1596);
or U1623 (N_1623,N_1567,N_1598);
nor U1624 (N_1624,N_1612,N_1605);
xor U1625 (N_1625,N_1597,N_1570);
nand U1626 (N_1626,N_1564,N_1578);
nor U1627 (N_1627,N_1569,N_1574);
nand U1628 (N_1628,N_1561,N_1615);
nor U1629 (N_1629,N_1601,N_1585);
nand U1630 (N_1630,N_1575,N_1587);
and U1631 (N_1631,N_1616,N_1592);
nand U1632 (N_1632,N_1595,N_1600);
nor U1633 (N_1633,N_1602,N_1568);
nand U1634 (N_1634,N_1572,N_1618);
nor U1635 (N_1635,N_1591,N_1562);
or U1636 (N_1636,N_1619,N_1604);
nor U1637 (N_1637,N_1583,N_1582);
nand U1638 (N_1638,N_1571,N_1599);
or U1639 (N_1639,N_1566,N_1560);
nor U1640 (N_1640,N_1577,N_1603);
nand U1641 (N_1641,N_1576,N_1581);
or U1642 (N_1642,N_1573,N_1614);
nor U1643 (N_1643,N_1563,N_1586);
nor U1644 (N_1644,N_1588,N_1606);
nand U1645 (N_1645,N_1593,N_1611);
nor U1646 (N_1646,N_1594,N_1589);
or U1647 (N_1647,N_1580,N_1610);
or U1648 (N_1648,N_1590,N_1607);
nand U1649 (N_1649,N_1579,N_1565);
nor U1650 (N_1650,N_1588,N_1599);
or U1651 (N_1651,N_1575,N_1597);
nand U1652 (N_1652,N_1580,N_1578);
or U1653 (N_1653,N_1618,N_1601);
and U1654 (N_1654,N_1597,N_1619);
and U1655 (N_1655,N_1574,N_1562);
xnor U1656 (N_1656,N_1610,N_1569);
nor U1657 (N_1657,N_1586,N_1589);
or U1658 (N_1658,N_1567,N_1585);
and U1659 (N_1659,N_1610,N_1616);
nor U1660 (N_1660,N_1567,N_1615);
nand U1661 (N_1661,N_1568,N_1604);
nor U1662 (N_1662,N_1567,N_1596);
and U1663 (N_1663,N_1602,N_1584);
and U1664 (N_1664,N_1573,N_1611);
or U1665 (N_1665,N_1598,N_1579);
and U1666 (N_1666,N_1588,N_1600);
or U1667 (N_1667,N_1579,N_1575);
or U1668 (N_1668,N_1612,N_1589);
nor U1669 (N_1669,N_1573,N_1619);
nor U1670 (N_1670,N_1605,N_1582);
nand U1671 (N_1671,N_1570,N_1571);
or U1672 (N_1672,N_1612,N_1573);
nand U1673 (N_1673,N_1580,N_1615);
and U1674 (N_1674,N_1603,N_1565);
nand U1675 (N_1675,N_1618,N_1605);
and U1676 (N_1676,N_1585,N_1599);
nor U1677 (N_1677,N_1575,N_1618);
or U1678 (N_1678,N_1579,N_1600);
nor U1679 (N_1679,N_1585,N_1603);
nor U1680 (N_1680,N_1675,N_1671);
and U1681 (N_1681,N_1669,N_1623);
nor U1682 (N_1682,N_1635,N_1660);
or U1683 (N_1683,N_1661,N_1655);
or U1684 (N_1684,N_1672,N_1645);
nor U1685 (N_1685,N_1632,N_1621);
xnor U1686 (N_1686,N_1649,N_1657);
and U1687 (N_1687,N_1650,N_1663);
or U1688 (N_1688,N_1648,N_1643);
nand U1689 (N_1689,N_1638,N_1640);
nand U1690 (N_1690,N_1637,N_1639);
nand U1691 (N_1691,N_1642,N_1678);
nor U1692 (N_1692,N_1654,N_1644);
or U1693 (N_1693,N_1664,N_1641);
or U1694 (N_1694,N_1674,N_1627);
or U1695 (N_1695,N_1668,N_1626);
nand U1696 (N_1696,N_1662,N_1673);
nor U1697 (N_1697,N_1636,N_1625);
and U1698 (N_1698,N_1630,N_1629);
nand U1699 (N_1699,N_1651,N_1665);
nor U1700 (N_1700,N_1658,N_1646);
or U1701 (N_1701,N_1647,N_1666);
nor U1702 (N_1702,N_1659,N_1670);
or U1703 (N_1703,N_1628,N_1653);
or U1704 (N_1704,N_1622,N_1679);
nand U1705 (N_1705,N_1620,N_1656);
or U1706 (N_1706,N_1667,N_1652);
nor U1707 (N_1707,N_1677,N_1634);
nand U1708 (N_1708,N_1633,N_1676);
or U1709 (N_1709,N_1631,N_1624);
or U1710 (N_1710,N_1631,N_1635);
and U1711 (N_1711,N_1631,N_1677);
nand U1712 (N_1712,N_1637,N_1673);
and U1713 (N_1713,N_1657,N_1676);
or U1714 (N_1714,N_1639,N_1660);
or U1715 (N_1715,N_1672,N_1667);
nor U1716 (N_1716,N_1656,N_1661);
nand U1717 (N_1717,N_1674,N_1625);
nand U1718 (N_1718,N_1622,N_1642);
or U1719 (N_1719,N_1674,N_1638);
or U1720 (N_1720,N_1638,N_1677);
nor U1721 (N_1721,N_1633,N_1643);
and U1722 (N_1722,N_1670,N_1644);
xnor U1723 (N_1723,N_1622,N_1629);
nand U1724 (N_1724,N_1664,N_1652);
or U1725 (N_1725,N_1652,N_1675);
and U1726 (N_1726,N_1670,N_1621);
nor U1727 (N_1727,N_1637,N_1652);
nor U1728 (N_1728,N_1624,N_1632);
nand U1729 (N_1729,N_1672,N_1669);
nand U1730 (N_1730,N_1635,N_1627);
and U1731 (N_1731,N_1679,N_1678);
nand U1732 (N_1732,N_1627,N_1624);
nand U1733 (N_1733,N_1667,N_1647);
and U1734 (N_1734,N_1640,N_1651);
or U1735 (N_1735,N_1635,N_1644);
or U1736 (N_1736,N_1673,N_1676);
or U1737 (N_1737,N_1670,N_1653);
nor U1738 (N_1738,N_1665,N_1636);
or U1739 (N_1739,N_1655,N_1648);
and U1740 (N_1740,N_1688,N_1723);
nand U1741 (N_1741,N_1718,N_1690);
nor U1742 (N_1742,N_1700,N_1710);
nand U1743 (N_1743,N_1714,N_1728);
or U1744 (N_1744,N_1685,N_1702);
and U1745 (N_1745,N_1691,N_1738);
or U1746 (N_1746,N_1733,N_1687);
nor U1747 (N_1747,N_1735,N_1716);
or U1748 (N_1748,N_1721,N_1682);
and U1749 (N_1749,N_1698,N_1701);
nor U1750 (N_1750,N_1694,N_1699);
nand U1751 (N_1751,N_1734,N_1732);
and U1752 (N_1752,N_1693,N_1705);
and U1753 (N_1753,N_1689,N_1727);
nand U1754 (N_1754,N_1709,N_1725);
or U1755 (N_1755,N_1692,N_1736);
or U1756 (N_1756,N_1722,N_1717);
or U1757 (N_1757,N_1681,N_1680);
or U1758 (N_1758,N_1708,N_1719);
and U1759 (N_1759,N_1696,N_1686);
nand U1760 (N_1760,N_1730,N_1724);
or U1761 (N_1761,N_1737,N_1683);
nand U1762 (N_1762,N_1720,N_1707);
nand U1763 (N_1763,N_1695,N_1739);
nor U1764 (N_1764,N_1715,N_1697);
or U1765 (N_1765,N_1704,N_1706);
and U1766 (N_1766,N_1729,N_1726);
nor U1767 (N_1767,N_1713,N_1711);
or U1768 (N_1768,N_1684,N_1712);
or U1769 (N_1769,N_1731,N_1703);
or U1770 (N_1770,N_1733,N_1699);
nor U1771 (N_1771,N_1710,N_1697);
nor U1772 (N_1772,N_1711,N_1706);
nor U1773 (N_1773,N_1707,N_1702);
or U1774 (N_1774,N_1714,N_1725);
or U1775 (N_1775,N_1691,N_1680);
nor U1776 (N_1776,N_1716,N_1713);
nand U1777 (N_1777,N_1732,N_1726);
and U1778 (N_1778,N_1720,N_1698);
nand U1779 (N_1779,N_1707,N_1730);
nand U1780 (N_1780,N_1694,N_1695);
and U1781 (N_1781,N_1716,N_1722);
and U1782 (N_1782,N_1709,N_1692);
nor U1783 (N_1783,N_1730,N_1709);
nor U1784 (N_1784,N_1736,N_1682);
nand U1785 (N_1785,N_1704,N_1730);
xnor U1786 (N_1786,N_1729,N_1680);
nand U1787 (N_1787,N_1700,N_1695);
nor U1788 (N_1788,N_1722,N_1738);
or U1789 (N_1789,N_1725,N_1730);
nand U1790 (N_1790,N_1700,N_1696);
or U1791 (N_1791,N_1734,N_1721);
or U1792 (N_1792,N_1727,N_1733);
or U1793 (N_1793,N_1713,N_1724);
nor U1794 (N_1794,N_1701,N_1712);
and U1795 (N_1795,N_1705,N_1698);
nand U1796 (N_1796,N_1709,N_1699);
and U1797 (N_1797,N_1736,N_1713);
nand U1798 (N_1798,N_1681,N_1690);
or U1799 (N_1799,N_1719,N_1714);
or U1800 (N_1800,N_1754,N_1792);
or U1801 (N_1801,N_1760,N_1785);
nor U1802 (N_1802,N_1796,N_1741);
or U1803 (N_1803,N_1782,N_1790);
or U1804 (N_1804,N_1761,N_1799);
nor U1805 (N_1805,N_1765,N_1793);
or U1806 (N_1806,N_1773,N_1783);
or U1807 (N_1807,N_1768,N_1767);
and U1808 (N_1808,N_1750,N_1779);
nand U1809 (N_1809,N_1762,N_1746);
or U1810 (N_1810,N_1763,N_1791);
or U1811 (N_1811,N_1753,N_1780);
nor U1812 (N_1812,N_1742,N_1777);
nand U1813 (N_1813,N_1795,N_1744);
nor U1814 (N_1814,N_1764,N_1751);
or U1815 (N_1815,N_1743,N_1756);
nand U1816 (N_1816,N_1788,N_1787);
xnor U1817 (N_1817,N_1752,N_1786);
or U1818 (N_1818,N_1770,N_1766);
nor U1819 (N_1819,N_1758,N_1784);
and U1820 (N_1820,N_1769,N_1798);
or U1821 (N_1821,N_1781,N_1778);
or U1822 (N_1822,N_1745,N_1748);
nand U1823 (N_1823,N_1749,N_1771);
nand U1824 (N_1824,N_1789,N_1757);
and U1825 (N_1825,N_1776,N_1759);
nor U1826 (N_1826,N_1774,N_1775);
nand U1827 (N_1827,N_1747,N_1794);
or U1828 (N_1828,N_1772,N_1740);
and U1829 (N_1829,N_1755,N_1797);
nor U1830 (N_1830,N_1765,N_1790);
and U1831 (N_1831,N_1783,N_1744);
nand U1832 (N_1832,N_1758,N_1740);
nor U1833 (N_1833,N_1756,N_1753);
nor U1834 (N_1834,N_1761,N_1766);
nor U1835 (N_1835,N_1753,N_1748);
or U1836 (N_1836,N_1786,N_1784);
and U1837 (N_1837,N_1743,N_1765);
nor U1838 (N_1838,N_1775,N_1784);
or U1839 (N_1839,N_1788,N_1773);
nand U1840 (N_1840,N_1755,N_1746);
and U1841 (N_1841,N_1779,N_1771);
nor U1842 (N_1842,N_1786,N_1777);
nand U1843 (N_1843,N_1784,N_1795);
nor U1844 (N_1844,N_1766,N_1781);
and U1845 (N_1845,N_1765,N_1770);
or U1846 (N_1846,N_1795,N_1772);
nor U1847 (N_1847,N_1796,N_1787);
nand U1848 (N_1848,N_1746,N_1741);
and U1849 (N_1849,N_1774,N_1766);
nor U1850 (N_1850,N_1773,N_1758);
and U1851 (N_1851,N_1767,N_1793);
and U1852 (N_1852,N_1774,N_1782);
or U1853 (N_1853,N_1784,N_1773);
nand U1854 (N_1854,N_1749,N_1766);
nor U1855 (N_1855,N_1740,N_1779);
nand U1856 (N_1856,N_1787,N_1794);
nand U1857 (N_1857,N_1745,N_1755);
nand U1858 (N_1858,N_1789,N_1784);
nand U1859 (N_1859,N_1750,N_1751);
and U1860 (N_1860,N_1801,N_1822);
or U1861 (N_1861,N_1836,N_1855);
or U1862 (N_1862,N_1818,N_1849);
or U1863 (N_1863,N_1852,N_1803);
and U1864 (N_1864,N_1857,N_1827);
and U1865 (N_1865,N_1845,N_1839);
nor U1866 (N_1866,N_1829,N_1802);
or U1867 (N_1867,N_1812,N_1821);
or U1868 (N_1868,N_1811,N_1814);
or U1869 (N_1869,N_1858,N_1847);
or U1870 (N_1870,N_1832,N_1807);
nor U1871 (N_1871,N_1850,N_1842);
or U1872 (N_1872,N_1805,N_1813);
nand U1873 (N_1873,N_1837,N_1841);
or U1874 (N_1874,N_1834,N_1833);
and U1875 (N_1875,N_1819,N_1800);
and U1876 (N_1876,N_1816,N_1830);
nand U1877 (N_1877,N_1848,N_1835);
nor U1878 (N_1878,N_1825,N_1838);
nand U1879 (N_1879,N_1859,N_1815);
and U1880 (N_1880,N_1820,N_1817);
and U1881 (N_1881,N_1854,N_1843);
and U1882 (N_1882,N_1831,N_1810);
nor U1883 (N_1883,N_1804,N_1828);
nand U1884 (N_1884,N_1853,N_1851);
nand U1885 (N_1885,N_1826,N_1856);
nor U1886 (N_1886,N_1846,N_1844);
nor U1887 (N_1887,N_1824,N_1823);
nand U1888 (N_1888,N_1840,N_1809);
or U1889 (N_1889,N_1808,N_1806);
or U1890 (N_1890,N_1844,N_1858);
nand U1891 (N_1891,N_1850,N_1847);
and U1892 (N_1892,N_1846,N_1858);
nand U1893 (N_1893,N_1859,N_1810);
and U1894 (N_1894,N_1813,N_1808);
and U1895 (N_1895,N_1842,N_1831);
or U1896 (N_1896,N_1823,N_1821);
nor U1897 (N_1897,N_1857,N_1829);
nor U1898 (N_1898,N_1805,N_1855);
nor U1899 (N_1899,N_1809,N_1828);
or U1900 (N_1900,N_1800,N_1839);
nand U1901 (N_1901,N_1852,N_1843);
nand U1902 (N_1902,N_1809,N_1841);
or U1903 (N_1903,N_1821,N_1829);
nand U1904 (N_1904,N_1846,N_1819);
or U1905 (N_1905,N_1805,N_1808);
or U1906 (N_1906,N_1837,N_1816);
nor U1907 (N_1907,N_1815,N_1817);
and U1908 (N_1908,N_1827,N_1850);
and U1909 (N_1909,N_1853,N_1806);
or U1910 (N_1910,N_1831,N_1858);
nand U1911 (N_1911,N_1808,N_1838);
or U1912 (N_1912,N_1811,N_1822);
nor U1913 (N_1913,N_1848,N_1815);
nand U1914 (N_1914,N_1842,N_1856);
and U1915 (N_1915,N_1833,N_1850);
and U1916 (N_1916,N_1832,N_1854);
or U1917 (N_1917,N_1854,N_1801);
or U1918 (N_1918,N_1822,N_1800);
nor U1919 (N_1919,N_1815,N_1802);
nand U1920 (N_1920,N_1868,N_1909);
nor U1921 (N_1921,N_1895,N_1878);
nor U1922 (N_1922,N_1885,N_1892);
or U1923 (N_1923,N_1865,N_1884);
or U1924 (N_1924,N_1882,N_1873);
nand U1925 (N_1925,N_1880,N_1910);
and U1926 (N_1926,N_1901,N_1889);
nor U1927 (N_1927,N_1903,N_1870);
nand U1928 (N_1928,N_1916,N_1898);
nand U1929 (N_1929,N_1886,N_1861);
and U1930 (N_1930,N_1888,N_1912);
nand U1931 (N_1931,N_1871,N_1906);
nand U1932 (N_1932,N_1866,N_1917);
and U1933 (N_1933,N_1897,N_1876);
or U1934 (N_1934,N_1899,N_1890);
and U1935 (N_1935,N_1911,N_1918);
and U1936 (N_1936,N_1891,N_1908);
xor U1937 (N_1937,N_1863,N_1900);
or U1938 (N_1938,N_1874,N_1902);
or U1939 (N_1939,N_1919,N_1907);
nand U1940 (N_1940,N_1913,N_1881);
or U1941 (N_1941,N_1860,N_1864);
or U1942 (N_1942,N_1875,N_1893);
nand U1943 (N_1943,N_1915,N_1883);
or U1944 (N_1944,N_1877,N_1905);
xor U1945 (N_1945,N_1887,N_1867);
nand U1946 (N_1946,N_1904,N_1894);
or U1947 (N_1947,N_1869,N_1872);
nand U1948 (N_1948,N_1862,N_1914);
and U1949 (N_1949,N_1879,N_1896);
and U1950 (N_1950,N_1867,N_1862);
nand U1951 (N_1951,N_1874,N_1879);
or U1952 (N_1952,N_1864,N_1887);
nand U1953 (N_1953,N_1860,N_1884);
nand U1954 (N_1954,N_1872,N_1884);
or U1955 (N_1955,N_1913,N_1888);
nand U1956 (N_1956,N_1910,N_1919);
or U1957 (N_1957,N_1902,N_1900);
nor U1958 (N_1958,N_1861,N_1901);
nand U1959 (N_1959,N_1911,N_1915);
or U1960 (N_1960,N_1910,N_1890);
nand U1961 (N_1961,N_1860,N_1902);
nand U1962 (N_1962,N_1886,N_1897);
nand U1963 (N_1963,N_1887,N_1905);
nor U1964 (N_1964,N_1908,N_1872);
nor U1965 (N_1965,N_1869,N_1888);
or U1966 (N_1966,N_1886,N_1893);
nand U1967 (N_1967,N_1872,N_1910);
nor U1968 (N_1968,N_1904,N_1870);
and U1969 (N_1969,N_1870,N_1876);
nand U1970 (N_1970,N_1905,N_1915);
and U1971 (N_1971,N_1888,N_1908);
and U1972 (N_1972,N_1886,N_1909);
or U1973 (N_1973,N_1907,N_1900);
nor U1974 (N_1974,N_1906,N_1886);
and U1975 (N_1975,N_1907,N_1887);
nand U1976 (N_1976,N_1886,N_1918);
nor U1977 (N_1977,N_1892,N_1864);
nand U1978 (N_1978,N_1898,N_1860);
or U1979 (N_1979,N_1871,N_1862);
nor U1980 (N_1980,N_1955,N_1957);
or U1981 (N_1981,N_1973,N_1960);
xor U1982 (N_1982,N_1939,N_1943);
xor U1983 (N_1983,N_1938,N_1963);
nand U1984 (N_1984,N_1935,N_1930);
and U1985 (N_1985,N_1978,N_1923);
nand U1986 (N_1986,N_1931,N_1944);
nor U1987 (N_1987,N_1959,N_1940);
and U1988 (N_1988,N_1964,N_1946);
or U1989 (N_1989,N_1945,N_1937);
and U1990 (N_1990,N_1974,N_1962);
nor U1991 (N_1991,N_1950,N_1947);
and U1992 (N_1992,N_1941,N_1954);
nand U1993 (N_1993,N_1969,N_1965);
and U1994 (N_1994,N_1929,N_1920);
nand U1995 (N_1995,N_1951,N_1926);
and U1996 (N_1996,N_1948,N_1979);
nor U1997 (N_1997,N_1922,N_1968);
and U1998 (N_1998,N_1966,N_1952);
nor U1999 (N_1999,N_1932,N_1961);
or U2000 (N_2000,N_1977,N_1958);
nor U2001 (N_2001,N_1928,N_1976);
or U2002 (N_2002,N_1927,N_1956);
and U2003 (N_2003,N_1971,N_1933);
or U2004 (N_2004,N_1925,N_1970);
and U2005 (N_2005,N_1921,N_1975);
nor U2006 (N_2006,N_1967,N_1934);
nand U2007 (N_2007,N_1924,N_1949);
nand U2008 (N_2008,N_1936,N_1942);
nand U2009 (N_2009,N_1972,N_1953);
nand U2010 (N_2010,N_1963,N_1942);
nor U2011 (N_2011,N_1956,N_1944);
nand U2012 (N_2012,N_1923,N_1976);
nand U2013 (N_2013,N_1955,N_1927);
nor U2014 (N_2014,N_1974,N_1951);
or U2015 (N_2015,N_1957,N_1951);
or U2016 (N_2016,N_1946,N_1924);
nand U2017 (N_2017,N_1934,N_1923);
and U2018 (N_2018,N_1957,N_1943);
or U2019 (N_2019,N_1962,N_1935);
nand U2020 (N_2020,N_1952,N_1976);
nor U2021 (N_2021,N_1923,N_1964);
and U2022 (N_2022,N_1931,N_1977);
nand U2023 (N_2023,N_1971,N_1936);
nand U2024 (N_2024,N_1959,N_1929);
and U2025 (N_2025,N_1959,N_1942);
and U2026 (N_2026,N_1969,N_1958);
nand U2027 (N_2027,N_1957,N_1946);
and U2028 (N_2028,N_1960,N_1932);
nand U2029 (N_2029,N_1948,N_1968);
nor U2030 (N_2030,N_1936,N_1931);
and U2031 (N_2031,N_1952,N_1924);
or U2032 (N_2032,N_1955,N_1968);
nand U2033 (N_2033,N_1942,N_1965);
and U2034 (N_2034,N_1961,N_1928);
and U2035 (N_2035,N_1932,N_1921);
nor U2036 (N_2036,N_1941,N_1927);
and U2037 (N_2037,N_1930,N_1958);
nand U2038 (N_2038,N_1937,N_1940);
and U2039 (N_2039,N_1944,N_1941);
and U2040 (N_2040,N_2032,N_2006);
or U2041 (N_2041,N_1980,N_1989);
or U2042 (N_2042,N_2000,N_2010);
nor U2043 (N_2043,N_2031,N_1983);
and U2044 (N_2044,N_1993,N_2018);
and U2045 (N_2045,N_2008,N_1985);
nor U2046 (N_2046,N_2012,N_2014);
and U2047 (N_2047,N_1987,N_1995);
nor U2048 (N_2048,N_2009,N_1992);
nor U2049 (N_2049,N_1990,N_1991);
or U2050 (N_2050,N_2029,N_2016);
or U2051 (N_2051,N_1994,N_2005);
and U2052 (N_2052,N_2015,N_2027);
nand U2053 (N_2053,N_1997,N_1996);
or U2054 (N_2054,N_2023,N_2002);
nand U2055 (N_2055,N_1982,N_1999);
nand U2056 (N_2056,N_1986,N_2028);
nand U2057 (N_2057,N_2011,N_2007);
nand U2058 (N_2058,N_2001,N_2022);
or U2059 (N_2059,N_1981,N_2039);
nor U2060 (N_2060,N_2038,N_2017);
and U2061 (N_2061,N_2003,N_1984);
xnor U2062 (N_2062,N_2019,N_2034);
or U2063 (N_2063,N_2026,N_2037);
or U2064 (N_2064,N_1998,N_2004);
and U2065 (N_2065,N_2030,N_2036);
nand U2066 (N_2066,N_2020,N_2021);
nor U2067 (N_2067,N_2033,N_1988);
or U2068 (N_2068,N_2025,N_2024);
nand U2069 (N_2069,N_2035,N_2013);
nand U2070 (N_2070,N_2032,N_2007);
and U2071 (N_2071,N_2002,N_1996);
nor U2072 (N_2072,N_1990,N_1983);
or U2073 (N_2073,N_1984,N_2021);
nor U2074 (N_2074,N_1980,N_1995);
nand U2075 (N_2075,N_2037,N_2009);
and U2076 (N_2076,N_2000,N_2018);
nand U2077 (N_2077,N_1982,N_1993);
nand U2078 (N_2078,N_2025,N_2020);
and U2079 (N_2079,N_1980,N_2034);
nand U2080 (N_2080,N_2011,N_1995);
nand U2081 (N_2081,N_2030,N_1986);
or U2082 (N_2082,N_2033,N_1990);
nand U2083 (N_2083,N_1983,N_2005);
or U2084 (N_2084,N_1999,N_2026);
nor U2085 (N_2085,N_1990,N_2012);
nand U2086 (N_2086,N_2038,N_2012);
nand U2087 (N_2087,N_2033,N_2024);
nand U2088 (N_2088,N_1984,N_2015);
nor U2089 (N_2089,N_2010,N_2022);
nor U2090 (N_2090,N_1981,N_2009);
nand U2091 (N_2091,N_2016,N_2033);
nand U2092 (N_2092,N_1996,N_1988);
nand U2093 (N_2093,N_1987,N_2027);
nand U2094 (N_2094,N_2035,N_1988);
nand U2095 (N_2095,N_2034,N_1999);
or U2096 (N_2096,N_2022,N_2038);
or U2097 (N_2097,N_2027,N_2028);
and U2098 (N_2098,N_1995,N_2001);
and U2099 (N_2099,N_2032,N_2018);
and U2100 (N_2100,N_2076,N_2089);
and U2101 (N_2101,N_2044,N_2062);
and U2102 (N_2102,N_2086,N_2061);
and U2103 (N_2103,N_2058,N_2093);
and U2104 (N_2104,N_2048,N_2055);
nor U2105 (N_2105,N_2084,N_2082);
and U2106 (N_2106,N_2049,N_2081);
nand U2107 (N_2107,N_2090,N_2063);
nor U2108 (N_2108,N_2094,N_2050);
and U2109 (N_2109,N_2059,N_2045);
or U2110 (N_2110,N_2056,N_2091);
and U2111 (N_2111,N_2064,N_2053);
and U2112 (N_2112,N_2060,N_2042);
and U2113 (N_2113,N_2047,N_2079);
nor U2114 (N_2114,N_2052,N_2080);
and U2115 (N_2115,N_2073,N_2099);
and U2116 (N_2116,N_2054,N_2078);
nor U2117 (N_2117,N_2085,N_2041);
or U2118 (N_2118,N_2072,N_2065);
or U2119 (N_2119,N_2069,N_2083);
or U2120 (N_2120,N_2074,N_2077);
and U2121 (N_2121,N_2071,N_2075);
nor U2122 (N_2122,N_2098,N_2057);
nor U2123 (N_2123,N_2092,N_2066);
nor U2124 (N_2124,N_2051,N_2095);
nor U2125 (N_2125,N_2096,N_2070);
or U2126 (N_2126,N_2046,N_2088);
nand U2127 (N_2127,N_2068,N_2097);
and U2128 (N_2128,N_2040,N_2067);
nand U2129 (N_2129,N_2043,N_2087);
nor U2130 (N_2130,N_2078,N_2085);
and U2131 (N_2131,N_2060,N_2094);
nand U2132 (N_2132,N_2098,N_2068);
xor U2133 (N_2133,N_2040,N_2063);
and U2134 (N_2134,N_2067,N_2043);
nand U2135 (N_2135,N_2049,N_2099);
or U2136 (N_2136,N_2042,N_2073);
nand U2137 (N_2137,N_2052,N_2097);
nand U2138 (N_2138,N_2074,N_2069);
nand U2139 (N_2139,N_2080,N_2095);
and U2140 (N_2140,N_2083,N_2042);
nor U2141 (N_2141,N_2070,N_2060);
nor U2142 (N_2142,N_2081,N_2068);
or U2143 (N_2143,N_2092,N_2096);
nor U2144 (N_2144,N_2068,N_2087);
and U2145 (N_2145,N_2047,N_2086);
and U2146 (N_2146,N_2062,N_2053);
and U2147 (N_2147,N_2085,N_2069);
and U2148 (N_2148,N_2080,N_2082);
and U2149 (N_2149,N_2085,N_2059);
nor U2150 (N_2150,N_2096,N_2055);
and U2151 (N_2151,N_2048,N_2080);
nor U2152 (N_2152,N_2076,N_2074);
or U2153 (N_2153,N_2081,N_2080);
nand U2154 (N_2154,N_2077,N_2079);
and U2155 (N_2155,N_2063,N_2057);
and U2156 (N_2156,N_2081,N_2053);
and U2157 (N_2157,N_2093,N_2091);
or U2158 (N_2158,N_2079,N_2056);
nor U2159 (N_2159,N_2055,N_2064);
and U2160 (N_2160,N_2106,N_2124);
or U2161 (N_2161,N_2145,N_2105);
nor U2162 (N_2162,N_2111,N_2156);
or U2163 (N_2163,N_2130,N_2157);
and U2164 (N_2164,N_2159,N_2122);
and U2165 (N_2165,N_2151,N_2150);
nor U2166 (N_2166,N_2103,N_2131);
or U2167 (N_2167,N_2137,N_2109);
nor U2168 (N_2168,N_2135,N_2117);
or U2169 (N_2169,N_2154,N_2114);
nand U2170 (N_2170,N_2100,N_2107);
and U2171 (N_2171,N_2138,N_2118);
nor U2172 (N_2172,N_2128,N_2139);
nor U2173 (N_2173,N_2113,N_2125);
nand U2174 (N_2174,N_2116,N_2152);
nand U2175 (N_2175,N_2127,N_2149);
and U2176 (N_2176,N_2134,N_2123);
and U2177 (N_2177,N_2115,N_2148);
nor U2178 (N_2178,N_2104,N_2144);
or U2179 (N_2179,N_2110,N_2155);
and U2180 (N_2180,N_2140,N_2101);
nand U2181 (N_2181,N_2147,N_2120);
nor U2182 (N_2182,N_2132,N_2112);
nor U2183 (N_2183,N_2141,N_2153);
xnor U2184 (N_2184,N_2143,N_2121);
nand U2185 (N_2185,N_2146,N_2133);
and U2186 (N_2186,N_2129,N_2119);
or U2187 (N_2187,N_2142,N_2126);
or U2188 (N_2188,N_2136,N_2102);
nand U2189 (N_2189,N_2158,N_2108);
and U2190 (N_2190,N_2107,N_2106);
nand U2191 (N_2191,N_2135,N_2105);
nand U2192 (N_2192,N_2154,N_2111);
nand U2193 (N_2193,N_2156,N_2159);
nor U2194 (N_2194,N_2127,N_2107);
or U2195 (N_2195,N_2115,N_2128);
nand U2196 (N_2196,N_2115,N_2140);
and U2197 (N_2197,N_2131,N_2106);
and U2198 (N_2198,N_2149,N_2152);
nand U2199 (N_2199,N_2147,N_2121);
or U2200 (N_2200,N_2106,N_2156);
and U2201 (N_2201,N_2125,N_2104);
nand U2202 (N_2202,N_2104,N_2136);
nand U2203 (N_2203,N_2114,N_2134);
nand U2204 (N_2204,N_2108,N_2154);
nor U2205 (N_2205,N_2147,N_2151);
nor U2206 (N_2206,N_2157,N_2115);
or U2207 (N_2207,N_2110,N_2104);
nand U2208 (N_2208,N_2108,N_2136);
or U2209 (N_2209,N_2133,N_2142);
nand U2210 (N_2210,N_2150,N_2127);
nor U2211 (N_2211,N_2120,N_2101);
nand U2212 (N_2212,N_2122,N_2154);
or U2213 (N_2213,N_2136,N_2116);
nand U2214 (N_2214,N_2114,N_2131);
and U2215 (N_2215,N_2144,N_2134);
nand U2216 (N_2216,N_2146,N_2126);
or U2217 (N_2217,N_2123,N_2141);
nor U2218 (N_2218,N_2109,N_2134);
nand U2219 (N_2219,N_2131,N_2104);
or U2220 (N_2220,N_2187,N_2201);
nand U2221 (N_2221,N_2188,N_2192);
nor U2222 (N_2222,N_2183,N_2177);
or U2223 (N_2223,N_2169,N_2171);
and U2224 (N_2224,N_2213,N_2160);
or U2225 (N_2225,N_2173,N_2198);
nand U2226 (N_2226,N_2214,N_2191);
or U2227 (N_2227,N_2215,N_2202);
and U2228 (N_2228,N_2203,N_2168);
or U2229 (N_2229,N_2207,N_2167);
and U2230 (N_2230,N_2209,N_2217);
nor U2231 (N_2231,N_2208,N_2193);
nor U2232 (N_2232,N_2210,N_2205);
nor U2233 (N_2233,N_2181,N_2182);
or U2234 (N_2234,N_2219,N_2190);
and U2235 (N_2235,N_2206,N_2218);
xor U2236 (N_2236,N_2174,N_2189);
nor U2237 (N_2237,N_2186,N_2164);
nor U2238 (N_2238,N_2162,N_2175);
nand U2239 (N_2239,N_2216,N_2161);
and U2240 (N_2240,N_2180,N_2176);
nor U2241 (N_2241,N_2163,N_2172);
or U2242 (N_2242,N_2200,N_2212);
nand U2243 (N_2243,N_2195,N_2197);
nor U2244 (N_2244,N_2179,N_2170);
nand U2245 (N_2245,N_2211,N_2165);
and U2246 (N_2246,N_2185,N_2194);
or U2247 (N_2247,N_2199,N_2196);
nor U2248 (N_2248,N_2184,N_2166);
or U2249 (N_2249,N_2178,N_2204);
nand U2250 (N_2250,N_2208,N_2218);
or U2251 (N_2251,N_2199,N_2214);
nor U2252 (N_2252,N_2176,N_2169);
nand U2253 (N_2253,N_2208,N_2195);
nor U2254 (N_2254,N_2179,N_2164);
or U2255 (N_2255,N_2177,N_2160);
nor U2256 (N_2256,N_2202,N_2209);
nand U2257 (N_2257,N_2161,N_2217);
and U2258 (N_2258,N_2185,N_2164);
or U2259 (N_2259,N_2201,N_2174);
nand U2260 (N_2260,N_2192,N_2190);
nand U2261 (N_2261,N_2210,N_2181);
nor U2262 (N_2262,N_2197,N_2217);
nor U2263 (N_2263,N_2180,N_2174);
nand U2264 (N_2264,N_2167,N_2185);
and U2265 (N_2265,N_2172,N_2195);
and U2266 (N_2266,N_2191,N_2167);
nand U2267 (N_2267,N_2182,N_2193);
nand U2268 (N_2268,N_2164,N_2189);
nor U2269 (N_2269,N_2211,N_2192);
or U2270 (N_2270,N_2206,N_2171);
nand U2271 (N_2271,N_2179,N_2177);
nor U2272 (N_2272,N_2194,N_2166);
and U2273 (N_2273,N_2174,N_2214);
nor U2274 (N_2274,N_2182,N_2168);
nand U2275 (N_2275,N_2195,N_2218);
or U2276 (N_2276,N_2211,N_2169);
nor U2277 (N_2277,N_2175,N_2170);
nor U2278 (N_2278,N_2189,N_2161);
nand U2279 (N_2279,N_2181,N_2203);
and U2280 (N_2280,N_2231,N_2248);
nor U2281 (N_2281,N_2259,N_2275);
or U2282 (N_2282,N_2279,N_2262);
nor U2283 (N_2283,N_2274,N_2268);
nor U2284 (N_2284,N_2227,N_2255);
and U2285 (N_2285,N_2232,N_2272);
nand U2286 (N_2286,N_2253,N_2266);
and U2287 (N_2287,N_2247,N_2221);
nor U2288 (N_2288,N_2273,N_2225);
nand U2289 (N_2289,N_2270,N_2246);
nand U2290 (N_2290,N_2276,N_2250);
and U2291 (N_2291,N_2241,N_2226);
and U2292 (N_2292,N_2265,N_2244);
or U2293 (N_2293,N_2256,N_2243);
nor U2294 (N_2294,N_2257,N_2261);
or U2295 (N_2295,N_2229,N_2223);
and U2296 (N_2296,N_2235,N_2263);
nand U2297 (N_2297,N_2233,N_2267);
nor U2298 (N_2298,N_2240,N_2220);
nor U2299 (N_2299,N_2228,N_2254);
nand U2300 (N_2300,N_2239,N_2245);
and U2301 (N_2301,N_2242,N_2238);
and U2302 (N_2302,N_2249,N_2269);
or U2303 (N_2303,N_2258,N_2230);
and U2304 (N_2304,N_2236,N_2264);
nor U2305 (N_2305,N_2237,N_2277);
nand U2306 (N_2306,N_2251,N_2271);
nand U2307 (N_2307,N_2234,N_2224);
or U2308 (N_2308,N_2252,N_2278);
or U2309 (N_2309,N_2222,N_2260);
and U2310 (N_2310,N_2275,N_2231);
or U2311 (N_2311,N_2241,N_2261);
nand U2312 (N_2312,N_2221,N_2244);
or U2313 (N_2313,N_2263,N_2227);
nand U2314 (N_2314,N_2262,N_2223);
and U2315 (N_2315,N_2276,N_2264);
nand U2316 (N_2316,N_2237,N_2233);
and U2317 (N_2317,N_2247,N_2264);
or U2318 (N_2318,N_2266,N_2232);
and U2319 (N_2319,N_2271,N_2237);
and U2320 (N_2320,N_2246,N_2273);
nand U2321 (N_2321,N_2275,N_2249);
nor U2322 (N_2322,N_2244,N_2246);
and U2323 (N_2323,N_2220,N_2254);
and U2324 (N_2324,N_2253,N_2265);
nand U2325 (N_2325,N_2278,N_2233);
and U2326 (N_2326,N_2275,N_2224);
nand U2327 (N_2327,N_2242,N_2248);
or U2328 (N_2328,N_2276,N_2234);
nand U2329 (N_2329,N_2263,N_2256);
or U2330 (N_2330,N_2257,N_2270);
and U2331 (N_2331,N_2229,N_2270);
nand U2332 (N_2332,N_2235,N_2225);
or U2333 (N_2333,N_2237,N_2231);
nor U2334 (N_2334,N_2225,N_2237);
nand U2335 (N_2335,N_2225,N_2230);
or U2336 (N_2336,N_2269,N_2232);
nor U2337 (N_2337,N_2248,N_2250);
nor U2338 (N_2338,N_2255,N_2275);
nor U2339 (N_2339,N_2259,N_2257);
or U2340 (N_2340,N_2315,N_2319);
and U2341 (N_2341,N_2304,N_2303);
nand U2342 (N_2342,N_2323,N_2297);
or U2343 (N_2343,N_2318,N_2296);
or U2344 (N_2344,N_2295,N_2313);
nor U2345 (N_2345,N_2286,N_2330);
nor U2346 (N_2346,N_2335,N_2308);
nand U2347 (N_2347,N_2331,N_2293);
and U2348 (N_2348,N_2312,N_2284);
nor U2349 (N_2349,N_2291,N_2307);
or U2350 (N_2350,N_2326,N_2325);
nand U2351 (N_2351,N_2287,N_2328);
nor U2352 (N_2352,N_2339,N_2314);
and U2353 (N_2353,N_2310,N_2332);
and U2354 (N_2354,N_2336,N_2280);
or U2355 (N_2355,N_2299,N_2300);
or U2356 (N_2356,N_2288,N_2337);
nand U2357 (N_2357,N_2338,N_2306);
and U2358 (N_2358,N_2298,N_2301);
xor U2359 (N_2359,N_2333,N_2302);
nor U2360 (N_2360,N_2309,N_2329);
nand U2361 (N_2361,N_2283,N_2320);
and U2362 (N_2362,N_2311,N_2324);
and U2363 (N_2363,N_2321,N_2282);
nor U2364 (N_2364,N_2316,N_2290);
nor U2365 (N_2365,N_2294,N_2327);
or U2366 (N_2366,N_2281,N_2305);
and U2367 (N_2367,N_2334,N_2317);
nor U2368 (N_2368,N_2289,N_2322);
nand U2369 (N_2369,N_2285,N_2292);
or U2370 (N_2370,N_2302,N_2309);
nand U2371 (N_2371,N_2307,N_2286);
nor U2372 (N_2372,N_2300,N_2310);
nand U2373 (N_2373,N_2284,N_2294);
nand U2374 (N_2374,N_2290,N_2291);
or U2375 (N_2375,N_2320,N_2327);
nor U2376 (N_2376,N_2301,N_2317);
nand U2377 (N_2377,N_2304,N_2332);
and U2378 (N_2378,N_2303,N_2293);
nand U2379 (N_2379,N_2338,N_2307);
nand U2380 (N_2380,N_2330,N_2309);
nand U2381 (N_2381,N_2333,N_2309);
and U2382 (N_2382,N_2334,N_2293);
nand U2383 (N_2383,N_2325,N_2336);
nor U2384 (N_2384,N_2313,N_2288);
nand U2385 (N_2385,N_2285,N_2331);
xor U2386 (N_2386,N_2315,N_2322);
nand U2387 (N_2387,N_2318,N_2288);
nor U2388 (N_2388,N_2305,N_2283);
or U2389 (N_2389,N_2316,N_2281);
nor U2390 (N_2390,N_2319,N_2286);
xnor U2391 (N_2391,N_2332,N_2305);
and U2392 (N_2392,N_2309,N_2311);
and U2393 (N_2393,N_2334,N_2332);
nand U2394 (N_2394,N_2311,N_2285);
nand U2395 (N_2395,N_2282,N_2337);
nand U2396 (N_2396,N_2298,N_2313);
or U2397 (N_2397,N_2304,N_2294);
nand U2398 (N_2398,N_2314,N_2289);
and U2399 (N_2399,N_2308,N_2303);
or U2400 (N_2400,N_2376,N_2371);
and U2401 (N_2401,N_2341,N_2356);
nor U2402 (N_2402,N_2347,N_2361);
and U2403 (N_2403,N_2398,N_2354);
nor U2404 (N_2404,N_2379,N_2358);
and U2405 (N_2405,N_2399,N_2381);
nor U2406 (N_2406,N_2368,N_2388);
nor U2407 (N_2407,N_2340,N_2382);
nand U2408 (N_2408,N_2390,N_2349);
xor U2409 (N_2409,N_2396,N_2350);
or U2410 (N_2410,N_2352,N_2366);
nor U2411 (N_2411,N_2370,N_2360);
nor U2412 (N_2412,N_2357,N_2345);
nand U2413 (N_2413,N_2355,N_2359);
and U2414 (N_2414,N_2351,N_2392);
nor U2415 (N_2415,N_2362,N_2373);
nor U2416 (N_2416,N_2389,N_2363);
or U2417 (N_2417,N_2353,N_2391);
or U2418 (N_2418,N_2397,N_2385);
nor U2419 (N_2419,N_2393,N_2378);
or U2420 (N_2420,N_2383,N_2364);
or U2421 (N_2421,N_2374,N_2375);
and U2422 (N_2422,N_2369,N_2365);
or U2423 (N_2423,N_2384,N_2377);
or U2424 (N_2424,N_2346,N_2387);
nand U2425 (N_2425,N_2380,N_2343);
or U2426 (N_2426,N_2395,N_2372);
or U2427 (N_2427,N_2344,N_2348);
nand U2428 (N_2428,N_2394,N_2342);
nand U2429 (N_2429,N_2367,N_2386);
and U2430 (N_2430,N_2388,N_2377);
nand U2431 (N_2431,N_2378,N_2381);
nor U2432 (N_2432,N_2371,N_2399);
or U2433 (N_2433,N_2379,N_2374);
or U2434 (N_2434,N_2341,N_2378);
nor U2435 (N_2435,N_2368,N_2366);
and U2436 (N_2436,N_2399,N_2383);
nand U2437 (N_2437,N_2373,N_2389);
nand U2438 (N_2438,N_2367,N_2389);
or U2439 (N_2439,N_2388,N_2375);
nor U2440 (N_2440,N_2375,N_2360);
nand U2441 (N_2441,N_2385,N_2345);
and U2442 (N_2442,N_2352,N_2364);
and U2443 (N_2443,N_2370,N_2376);
and U2444 (N_2444,N_2383,N_2356);
and U2445 (N_2445,N_2359,N_2373);
and U2446 (N_2446,N_2341,N_2352);
and U2447 (N_2447,N_2358,N_2375);
nand U2448 (N_2448,N_2360,N_2342);
nor U2449 (N_2449,N_2359,N_2363);
nand U2450 (N_2450,N_2354,N_2362);
nand U2451 (N_2451,N_2372,N_2380);
or U2452 (N_2452,N_2346,N_2360);
nor U2453 (N_2453,N_2342,N_2386);
and U2454 (N_2454,N_2345,N_2340);
nor U2455 (N_2455,N_2365,N_2347);
nor U2456 (N_2456,N_2391,N_2344);
nand U2457 (N_2457,N_2388,N_2341);
or U2458 (N_2458,N_2365,N_2380);
nor U2459 (N_2459,N_2376,N_2394);
and U2460 (N_2460,N_2415,N_2431);
nand U2461 (N_2461,N_2402,N_2434);
nor U2462 (N_2462,N_2443,N_2406);
and U2463 (N_2463,N_2416,N_2439);
nor U2464 (N_2464,N_2449,N_2401);
and U2465 (N_2465,N_2448,N_2451);
or U2466 (N_2466,N_2408,N_2435);
nand U2467 (N_2467,N_2407,N_2457);
or U2468 (N_2468,N_2445,N_2420);
or U2469 (N_2469,N_2453,N_2436);
nor U2470 (N_2470,N_2452,N_2413);
or U2471 (N_2471,N_2440,N_2428);
xor U2472 (N_2472,N_2446,N_2410);
nor U2473 (N_2473,N_2455,N_2404);
nor U2474 (N_2474,N_2441,N_2429);
or U2475 (N_2475,N_2454,N_2403);
or U2476 (N_2476,N_2423,N_2409);
nor U2477 (N_2477,N_2433,N_2425);
or U2478 (N_2478,N_2456,N_2400);
or U2479 (N_2479,N_2421,N_2427);
or U2480 (N_2480,N_2422,N_2438);
and U2481 (N_2481,N_2432,N_2450);
or U2482 (N_2482,N_2424,N_2418);
nand U2483 (N_2483,N_2419,N_2444);
nand U2484 (N_2484,N_2459,N_2412);
or U2485 (N_2485,N_2447,N_2417);
or U2486 (N_2486,N_2437,N_2411);
and U2487 (N_2487,N_2430,N_2458);
or U2488 (N_2488,N_2414,N_2405);
nand U2489 (N_2489,N_2442,N_2426);
nand U2490 (N_2490,N_2414,N_2424);
nor U2491 (N_2491,N_2452,N_2449);
nor U2492 (N_2492,N_2430,N_2434);
or U2493 (N_2493,N_2412,N_2457);
nand U2494 (N_2494,N_2448,N_2408);
and U2495 (N_2495,N_2421,N_2448);
and U2496 (N_2496,N_2444,N_2452);
nor U2497 (N_2497,N_2421,N_2458);
and U2498 (N_2498,N_2410,N_2447);
or U2499 (N_2499,N_2424,N_2439);
nand U2500 (N_2500,N_2405,N_2416);
or U2501 (N_2501,N_2450,N_2417);
nor U2502 (N_2502,N_2433,N_2426);
or U2503 (N_2503,N_2432,N_2455);
and U2504 (N_2504,N_2432,N_2418);
nor U2505 (N_2505,N_2417,N_2440);
nor U2506 (N_2506,N_2404,N_2414);
or U2507 (N_2507,N_2438,N_2421);
nand U2508 (N_2508,N_2419,N_2418);
nand U2509 (N_2509,N_2422,N_2402);
nand U2510 (N_2510,N_2407,N_2422);
nor U2511 (N_2511,N_2448,N_2404);
or U2512 (N_2512,N_2405,N_2444);
or U2513 (N_2513,N_2426,N_2446);
and U2514 (N_2514,N_2418,N_2430);
or U2515 (N_2515,N_2424,N_2427);
nand U2516 (N_2516,N_2451,N_2439);
and U2517 (N_2517,N_2440,N_2407);
or U2518 (N_2518,N_2446,N_2428);
and U2519 (N_2519,N_2425,N_2428);
nand U2520 (N_2520,N_2476,N_2474);
or U2521 (N_2521,N_2516,N_2509);
and U2522 (N_2522,N_2479,N_2470);
and U2523 (N_2523,N_2464,N_2488);
or U2524 (N_2524,N_2510,N_2481);
nand U2525 (N_2525,N_2478,N_2466);
nor U2526 (N_2526,N_2512,N_2501);
or U2527 (N_2527,N_2504,N_2500);
and U2528 (N_2528,N_2495,N_2503);
nand U2529 (N_2529,N_2505,N_2484);
and U2530 (N_2530,N_2465,N_2507);
nand U2531 (N_2531,N_2511,N_2477);
or U2532 (N_2532,N_2469,N_2498);
and U2533 (N_2533,N_2462,N_2508);
nor U2534 (N_2534,N_2460,N_2513);
nor U2535 (N_2535,N_2482,N_2497);
or U2536 (N_2536,N_2514,N_2473);
nor U2537 (N_2537,N_2485,N_2467);
nor U2538 (N_2538,N_2471,N_2494);
and U2539 (N_2539,N_2491,N_2461);
or U2540 (N_2540,N_2506,N_2492);
or U2541 (N_2541,N_2518,N_2499);
nand U2542 (N_2542,N_2468,N_2489);
and U2543 (N_2543,N_2487,N_2480);
and U2544 (N_2544,N_2493,N_2502);
and U2545 (N_2545,N_2472,N_2486);
nand U2546 (N_2546,N_2483,N_2517);
nand U2547 (N_2547,N_2496,N_2519);
nor U2548 (N_2548,N_2490,N_2475);
and U2549 (N_2549,N_2515,N_2463);
or U2550 (N_2550,N_2514,N_2487);
nor U2551 (N_2551,N_2511,N_2478);
nor U2552 (N_2552,N_2509,N_2468);
or U2553 (N_2553,N_2511,N_2513);
nand U2554 (N_2554,N_2473,N_2489);
nand U2555 (N_2555,N_2500,N_2511);
or U2556 (N_2556,N_2473,N_2483);
and U2557 (N_2557,N_2480,N_2468);
nor U2558 (N_2558,N_2509,N_2503);
nand U2559 (N_2559,N_2465,N_2463);
nand U2560 (N_2560,N_2476,N_2478);
nand U2561 (N_2561,N_2466,N_2482);
and U2562 (N_2562,N_2465,N_2477);
nor U2563 (N_2563,N_2473,N_2509);
nand U2564 (N_2564,N_2496,N_2495);
or U2565 (N_2565,N_2480,N_2509);
nor U2566 (N_2566,N_2501,N_2507);
or U2567 (N_2567,N_2498,N_2460);
or U2568 (N_2568,N_2515,N_2516);
and U2569 (N_2569,N_2481,N_2460);
nand U2570 (N_2570,N_2470,N_2503);
or U2571 (N_2571,N_2497,N_2495);
or U2572 (N_2572,N_2463,N_2496);
or U2573 (N_2573,N_2504,N_2473);
and U2574 (N_2574,N_2479,N_2500);
or U2575 (N_2575,N_2465,N_2495);
nor U2576 (N_2576,N_2504,N_2494);
and U2577 (N_2577,N_2499,N_2516);
and U2578 (N_2578,N_2463,N_2489);
nor U2579 (N_2579,N_2462,N_2484);
or U2580 (N_2580,N_2571,N_2556);
nand U2581 (N_2581,N_2560,N_2563);
nand U2582 (N_2582,N_2541,N_2565);
nor U2583 (N_2583,N_2579,N_2532);
and U2584 (N_2584,N_2543,N_2528);
nand U2585 (N_2585,N_2566,N_2536);
and U2586 (N_2586,N_2538,N_2534);
or U2587 (N_2587,N_2554,N_2570);
nand U2588 (N_2588,N_2520,N_2575);
nor U2589 (N_2589,N_2548,N_2555);
and U2590 (N_2590,N_2559,N_2527);
nand U2591 (N_2591,N_2525,N_2549);
and U2592 (N_2592,N_2562,N_2533);
nor U2593 (N_2593,N_2531,N_2546);
nor U2594 (N_2594,N_2568,N_2567);
or U2595 (N_2595,N_2522,N_2553);
nand U2596 (N_2596,N_2576,N_2574);
and U2597 (N_2597,N_2577,N_2564);
nand U2598 (N_2598,N_2537,N_2572);
or U2599 (N_2599,N_2547,N_2557);
nand U2600 (N_2600,N_2551,N_2578);
and U2601 (N_2601,N_2545,N_2526);
nor U2602 (N_2602,N_2529,N_2535);
nor U2603 (N_2603,N_2540,N_2550);
or U2604 (N_2604,N_2552,N_2523);
nand U2605 (N_2605,N_2539,N_2521);
or U2606 (N_2606,N_2542,N_2530);
nor U2607 (N_2607,N_2573,N_2558);
nand U2608 (N_2608,N_2544,N_2561);
or U2609 (N_2609,N_2569,N_2524);
nand U2610 (N_2610,N_2571,N_2574);
and U2611 (N_2611,N_2560,N_2574);
or U2612 (N_2612,N_2567,N_2572);
and U2613 (N_2613,N_2529,N_2555);
and U2614 (N_2614,N_2544,N_2552);
nor U2615 (N_2615,N_2540,N_2525);
and U2616 (N_2616,N_2528,N_2557);
nand U2617 (N_2617,N_2534,N_2562);
nor U2618 (N_2618,N_2563,N_2543);
nor U2619 (N_2619,N_2537,N_2527);
nand U2620 (N_2620,N_2533,N_2534);
or U2621 (N_2621,N_2536,N_2577);
or U2622 (N_2622,N_2576,N_2564);
nor U2623 (N_2623,N_2554,N_2541);
or U2624 (N_2624,N_2560,N_2523);
or U2625 (N_2625,N_2541,N_2562);
nand U2626 (N_2626,N_2565,N_2579);
nand U2627 (N_2627,N_2550,N_2529);
or U2628 (N_2628,N_2525,N_2537);
or U2629 (N_2629,N_2578,N_2548);
and U2630 (N_2630,N_2566,N_2542);
or U2631 (N_2631,N_2547,N_2548);
or U2632 (N_2632,N_2568,N_2563);
or U2633 (N_2633,N_2526,N_2557);
nand U2634 (N_2634,N_2541,N_2537);
or U2635 (N_2635,N_2523,N_2553);
nor U2636 (N_2636,N_2550,N_2573);
and U2637 (N_2637,N_2531,N_2541);
nand U2638 (N_2638,N_2561,N_2578);
or U2639 (N_2639,N_2566,N_2569);
nand U2640 (N_2640,N_2591,N_2618);
nand U2641 (N_2641,N_2624,N_2597);
and U2642 (N_2642,N_2613,N_2600);
or U2643 (N_2643,N_2610,N_2634);
nand U2644 (N_2644,N_2635,N_2617);
and U2645 (N_2645,N_2627,N_2585);
nor U2646 (N_2646,N_2636,N_2599);
or U2647 (N_2647,N_2598,N_2614);
nand U2648 (N_2648,N_2630,N_2590);
and U2649 (N_2649,N_2593,N_2601);
nand U2650 (N_2650,N_2638,N_2631);
nor U2651 (N_2651,N_2609,N_2639);
or U2652 (N_2652,N_2588,N_2594);
nand U2653 (N_2653,N_2604,N_2611);
or U2654 (N_2654,N_2616,N_2623);
and U2655 (N_2655,N_2592,N_2608);
nand U2656 (N_2656,N_2582,N_2615);
or U2657 (N_2657,N_2629,N_2602);
or U2658 (N_2658,N_2581,N_2619);
nor U2659 (N_2659,N_2626,N_2595);
or U2660 (N_2660,N_2637,N_2625);
nand U2661 (N_2661,N_2603,N_2633);
nand U2662 (N_2662,N_2580,N_2589);
nor U2663 (N_2663,N_2584,N_2606);
or U2664 (N_2664,N_2612,N_2622);
nor U2665 (N_2665,N_2621,N_2605);
or U2666 (N_2666,N_2586,N_2596);
nand U2667 (N_2667,N_2587,N_2583);
or U2668 (N_2668,N_2607,N_2628);
nand U2669 (N_2669,N_2620,N_2632);
or U2670 (N_2670,N_2604,N_2593);
or U2671 (N_2671,N_2623,N_2592);
and U2672 (N_2672,N_2614,N_2625);
and U2673 (N_2673,N_2596,N_2599);
and U2674 (N_2674,N_2620,N_2584);
or U2675 (N_2675,N_2616,N_2611);
and U2676 (N_2676,N_2631,N_2594);
or U2677 (N_2677,N_2615,N_2607);
nand U2678 (N_2678,N_2615,N_2627);
nand U2679 (N_2679,N_2613,N_2585);
nand U2680 (N_2680,N_2607,N_2593);
nor U2681 (N_2681,N_2618,N_2581);
or U2682 (N_2682,N_2612,N_2584);
or U2683 (N_2683,N_2598,N_2600);
and U2684 (N_2684,N_2607,N_2630);
nor U2685 (N_2685,N_2600,N_2617);
nand U2686 (N_2686,N_2634,N_2608);
and U2687 (N_2687,N_2590,N_2592);
nor U2688 (N_2688,N_2622,N_2617);
and U2689 (N_2689,N_2593,N_2629);
nor U2690 (N_2690,N_2593,N_2625);
or U2691 (N_2691,N_2623,N_2635);
nand U2692 (N_2692,N_2624,N_2614);
nor U2693 (N_2693,N_2635,N_2611);
nor U2694 (N_2694,N_2615,N_2585);
or U2695 (N_2695,N_2606,N_2591);
or U2696 (N_2696,N_2632,N_2584);
or U2697 (N_2697,N_2625,N_2616);
or U2698 (N_2698,N_2623,N_2599);
nand U2699 (N_2699,N_2618,N_2600);
or U2700 (N_2700,N_2680,N_2676);
or U2701 (N_2701,N_2651,N_2679);
and U2702 (N_2702,N_2656,N_2699);
nor U2703 (N_2703,N_2675,N_2668);
or U2704 (N_2704,N_2689,N_2684);
nand U2705 (N_2705,N_2694,N_2690);
or U2706 (N_2706,N_2678,N_2698);
nand U2707 (N_2707,N_2665,N_2677);
and U2708 (N_2708,N_2648,N_2673);
or U2709 (N_2709,N_2682,N_2666);
nor U2710 (N_2710,N_2697,N_2661);
or U2711 (N_2711,N_2658,N_2644);
nor U2712 (N_2712,N_2686,N_2667);
nor U2713 (N_2713,N_2659,N_2654);
or U2714 (N_2714,N_2693,N_2655);
nor U2715 (N_2715,N_2641,N_2649);
or U2716 (N_2716,N_2688,N_2653);
and U2717 (N_2717,N_2662,N_2660);
and U2718 (N_2718,N_2672,N_2691);
or U2719 (N_2719,N_2643,N_2685);
and U2720 (N_2720,N_2695,N_2692);
nor U2721 (N_2721,N_2674,N_2640);
and U2722 (N_2722,N_2670,N_2657);
and U2723 (N_2723,N_2664,N_2647);
nand U2724 (N_2724,N_2683,N_2687);
nand U2725 (N_2725,N_2642,N_2681);
or U2726 (N_2726,N_2646,N_2645);
nand U2727 (N_2727,N_2671,N_2663);
nand U2728 (N_2728,N_2669,N_2650);
nand U2729 (N_2729,N_2696,N_2652);
nor U2730 (N_2730,N_2696,N_2698);
and U2731 (N_2731,N_2665,N_2659);
and U2732 (N_2732,N_2661,N_2645);
nand U2733 (N_2733,N_2640,N_2683);
or U2734 (N_2734,N_2682,N_2684);
xnor U2735 (N_2735,N_2643,N_2675);
and U2736 (N_2736,N_2666,N_2684);
nand U2737 (N_2737,N_2669,N_2679);
nand U2738 (N_2738,N_2687,N_2674);
or U2739 (N_2739,N_2694,N_2657);
and U2740 (N_2740,N_2684,N_2672);
and U2741 (N_2741,N_2679,N_2647);
nand U2742 (N_2742,N_2669,N_2675);
nor U2743 (N_2743,N_2697,N_2649);
or U2744 (N_2744,N_2658,N_2656);
nand U2745 (N_2745,N_2691,N_2664);
and U2746 (N_2746,N_2662,N_2663);
or U2747 (N_2747,N_2694,N_2671);
nand U2748 (N_2748,N_2657,N_2684);
or U2749 (N_2749,N_2664,N_2662);
xor U2750 (N_2750,N_2647,N_2671);
and U2751 (N_2751,N_2664,N_2687);
nor U2752 (N_2752,N_2676,N_2663);
nand U2753 (N_2753,N_2661,N_2695);
and U2754 (N_2754,N_2683,N_2646);
or U2755 (N_2755,N_2697,N_2669);
and U2756 (N_2756,N_2646,N_2692);
nand U2757 (N_2757,N_2690,N_2689);
and U2758 (N_2758,N_2663,N_2670);
nor U2759 (N_2759,N_2664,N_2646);
and U2760 (N_2760,N_2741,N_2718);
nand U2761 (N_2761,N_2708,N_2727);
and U2762 (N_2762,N_2713,N_2705);
nand U2763 (N_2763,N_2715,N_2750);
nand U2764 (N_2764,N_2701,N_2721);
nand U2765 (N_2765,N_2726,N_2746);
or U2766 (N_2766,N_2755,N_2738);
and U2767 (N_2767,N_2757,N_2749);
or U2768 (N_2768,N_2744,N_2712);
nand U2769 (N_2769,N_2745,N_2722);
nor U2770 (N_2770,N_2711,N_2747);
nand U2771 (N_2771,N_2742,N_2736);
nor U2772 (N_2772,N_2717,N_2756);
nand U2773 (N_2773,N_2707,N_2728);
nor U2774 (N_2774,N_2734,N_2740);
nand U2775 (N_2775,N_2724,N_2743);
and U2776 (N_2776,N_2739,N_2759);
nand U2777 (N_2777,N_2748,N_2723);
nand U2778 (N_2778,N_2710,N_2733);
nand U2779 (N_2779,N_2719,N_2754);
nand U2780 (N_2780,N_2703,N_2735);
nand U2781 (N_2781,N_2720,N_2729);
and U2782 (N_2782,N_2731,N_2730);
and U2783 (N_2783,N_2753,N_2709);
nand U2784 (N_2784,N_2752,N_2706);
nand U2785 (N_2785,N_2732,N_2725);
nor U2786 (N_2786,N_2737,N_2704);
nor U2787 (N_2787,N_2714,N_2751);
or U2788 (N_2788,N_2700,N_2716);
and U2789 (N_2789,N_2702,N_2758);
nand U2790 (N_2790,N_2727,N_2744);
nor U2791 (N_2791,N_2746,N_2712);
and U2792 (N_2792,N_2704,N_2741);
or U2793 (N_2793,N_2717,N_2713);
and U2794 (N_2794,N_2722,N_2737);
nor U2795 (N_2795,N_2708,N_2703);
nor U2796 (N_2796,N_2725,N_2729);
nand U2797 (N_2797,N_2720,N_2747);
nor U2798 (N_2798,N_2758,N_2751);
or U2799 (N_2799,N_2726,N_2740);
nor U2800 (N_2800,N_2701,N_2729);
and U2801 (N_2801,N_2740,N_2750);
or U2802 (N_2802,N_2752,N_2721);
nand U2803 (N_2803,N_2709,N_2718);
and U2804 (N_2804,N_2711,N_2737);
and U2805 (N_2805,N_2751,N_2742);
and U2806 (N_2806,N_2754,N_2753);
and U2807 (N_2807,N_2724,N_2728);
and U2808 (N_2808,N_2756,N_2754);
and U2809 (N_2809,N_2750,N_2739);
or U2810 (N_2810,N_2701,N_2702);
nand U2811 (N_2811,N_2737,N_2703);
or U2812 (N_2812,N_2705,N_2706);
nor U2813 (N_2813,N_2749,N_2713);
nor U2814 (N_2814,N_2751,N_2748);
nor U2815 (N_2815,N_2703,N_2732);
nand U2816 (N_2816,N_2730,N_2712);
nand U2817 (N_2817,N_2728,N_2702);
nor U2818 (N_2818,N_2743,N_2728);
nor U2819 (N_2819,N_2719,N_2727);
and U2820 (N_2820,N_2772,N_2760);
nand U2821 (N_2821,N_2761,N_2801);
and U2822 (N_2822,N_2798,N_2768);
nor U2823 (N_2823,N_2762,N_2792);
or U2824 (N_2824,N_2769,N_2811);
or U2825 (N_2825,N_2806,N_2816);
or U2826 (N_2826,N_2786,N_2795);
nand U2827 (N_2827,N_2788,N_2810);
nand U2828 (N_2828,N_2799,N_2804);
and U2829 (N_2829,N_2815,N_2789);
or U2830 (N_2830,N_2809,N_2797);
and U2831 (N_2831,N_2767,N_2779);
or U2832 (N_2832,N_2800,N_2778);
or U2833 (N_2833,N_2817,N_2773);
or U2834 (N_2834,N_2814,N_2794);
or U2835 (N_2835,N_2781,N_2787);
or U2836 (N_2836,N_2785,N_2783);
and U2837 (N_2837,N_2802,N_2782);
and U2838 (N_2838,N_2819,N_2812);
and U2839 (N_2839,N_2793,N_2765);
and U2840 (N_2840,N_2803,N_2766);
nand U2841 (N_2841,N_2780,N_2807);
nor U2842 (N_2842,N_2818,N_2770);
nand U2843 (N_2843,N_2791,N_2771);
or U2844 (N_2844,N_2805,N_2764);
and U2845 (N_2845,N_2774,N_2776);
or U2846 (N_2846,N_2796,N_2784);
and U2847 (N_2847,N_2775,N_2763);
or U2848 (N_2848,N_2777,N_2808);
nand U2849 (N_2849,N_2813,N_2790);
or U2850 (N_2850,N_2781,N_2806);
nand U2851 (N_2851,N_2763,N_2788);
or U2852 (N_2852,N_2788,N_2796);
and U2853 (N_2853,N_2767,N_2789);
and U2854 (N_2854,N_2793,N_2798);
and U2855 (N_2855,N_2766,N_2794);
nor U2856 (N_2856,N_2778,N_2811);
xor U2857 (N_2857,N_2802,N_2796);
nand U2858 (N_2858,N_2801,N_2814);
nand U2859 (N_2859,N_2785,N_2819);
or U2860 (N_2860,N_2785,N_2811);
nor U2861 (N_2861,N_2788,N_2819);
nor U2862 (N_2862,N_2765,N_2790);
or U2863 (N_2863,N_2760,N_2778);
or U2864 (N_2864,N_2787,N_2804);
or U2865 (N_2865,N_2782,N_2765);
and U2866 (N_2866,N_2767,N_2787);
nor U2867 (N_2867,N_2775,N_2781);
and U2868 (N_2868,N_2784,N_2810);
and U2869 (N_2869,N_2763,N_2785);
and U2870 (N_2870,N_2809,N_2792);
nor U2871 (N_2871,N_2771,N_2768);
or U2872 (N_2872,N_2805,N_2763);
or U2873 (N_2873,N_2784,N_2806);
nand U2874 (N_2874,N_2765,N_2819);
or U2875 (N_2875,N_2819,N_2782);
and U2876 (N_2876,N_2816,N_2783);
nor U2877 (N_2877,N_2760,N_2813);
xor U2878 (N_2878,N_2778,N_2816);
and U2879 (N_2879,N_2805,N_2806);
and U2880 (N_2880,N_2855,N_2872);
and U2881 (N_2881,N_2821,N_2820);
and U2882 (N_2882,N_2824,N_2835);
nand U2883 (N_2883,N_2857,N_2871);
and U2884 (N_2884,N_2828,N_2830);
or U2885 (N_2885,N_2852,N_2825);
nand U2886 (N_2886,N_2849,N_2879);
and U2887 (N_2887,N_2860,N_2866);
nor U2888 (N_2888,N_2874,N_2838);
and U2889 (N_2889,N_2844,N_2826);
and U2890 (N_2890,N_2869,N_2878);
nor U2891 (N_2891,N_2827,N_2851);
nor U2892 (N_2892,N_2854,N_2867);
and U2893 (N_2893,N_2861,N_2846);
nand U2894 (N_2894,N_2842,N_2875);
and U2895 (N_2895,N_2843,N_2831);
or U2896 (N_2896,N_2876,N_2834);
nor U2897 (N_2897,N_2873,N_2836);
nand U2898 (N_2898,N_2823,N_2868);
or U2899 (N_2899,N_2864,N_2850);
nor U2900 (N_2900,N_2862,N_2841);
nor U2901 (N_2901,N_2847,N_2837);
and U2902 (N_2902,N_2853,N_2848);
or U2903 (N_2903,N_2822,N_2839);
xor U2904 (N_2904,N_2840,N_2870);
nand U2905 (N_2905,N_2865,N_2856);
nor U2906 (N_2906,N_2833,N_2829);
or U2907 (N_2907,N_2877,N_2859);
or U2908 (N_2908,N_2858,N_2845);
and U2909 (N_2909,N_2863,N_2832);
nor U2910 (N_2910,N_2844,N_2868);
or U2911 (N_2911,N_2867,N_2847);
and U2912 (N_2912,N_2830,N_2848);
or U2913 (N_2913,N_2857,N_2830);
nand U2914 (N_2914,N_2856,N_2877);
nor U2915 (N_2915,N_2834,N_2823);
nor U2916 (N_2916,N_2856,N_2879);
and U2917 (N_2917,N_2832,N_2852);
nor U2918 (N_2918,N_2842,N_2836);
nor U2919 (N_2919,N_2830,N_2840);
nor U2920 (N_2920,N_2848,N_2856);
nor U2921 (N_2921,N_2864,N_2855);
nor U2922 (N_2922,N_2837,N_2838);
and U2923 (N_2923,N_2846,N_2873);
and U2924 (N_2924,N_2865,N_2825);
nor U2925 (N_2925,N_2876,N_2854);
nand U2926 (N_2926,N_2825,N_2876);
nor U2927 (N_2927,N_2827,N_2873);
or U2928 (N_2928,N_2853,N_2863);
nor U2929 (N_2929,N_2833,N_2872);
nand U2930 (N_2930,N_2872,N_2830);
nand U2931 (N_2931,N_2849,N_2835);
nand U2932 (N_2932,N_2839,N_2857);
and U2933 (N_2933,N_2868,N_2878);
or U2934 (N_2934,N_2822,N_2821);
nand U2935 (N_2935,N_2857,N_2849);
and U2936 (N_2936,N_2867,N_2857);
or U2937 (N_2937,N_2839,N_2831);
nor U2938 (N_2938,N_2824,N_2828);
nand U2939 (N_2939,N_2833,N_2839);
or U2940 (N_2940,N_2930,N_2898);
or U2941 (N_2941,N_2890,N_2912);
nand U2942 (N_2942,N_2904,N_2886);
or U2943 (N_2943,N_2935,N_2915);
nor U2944 (N_2944,N_2919,N_2920);
nand U2945 (N_2945,N_2888,N_2916);
and U2946 (N_2946,N_2880,N_2899);
nand U2947 (N_2947,N_2936,N_2923);
and U2948 (N_2948,N_2938,N_2934);
nand U2949 (N_2949,N_2894,N_2910);
nand U2950 (N_2950,N_2933,N_2918);
or U2951 (N_2951,N_2911,N_2928);
and U2952 (N_2952,N_2893,N_2925);
nor U2953 (N_2953,N_2937,N_2885);
nand U2954 (N_2954,N_2907,N_2909);
nand U2955 (N_2955,N_2884,N_2902);
and U2956 (N_2956,N_2931,N_2905);
and U2957 (N_2957,N_2922,N_2887);
nand U2958 (N_2958,N_2921,N_2900);
and U2959 (N_2959,N_2883,N_2917);
or U2960 (N_2960,N_2881,N_2914);
nor U2961 (N_2961,N_2901,N_2908);
nand U2962 (N_2962,N_2932,N_2903);
nor U2963 (N_2963,N_2882,N_2891);
or U2964 (N_2964,N_2924,N_2892);
nor U2965 (N_2965,N_2895,N_2896);
nand U2966 (N_2966,N_2927,N_2939);
and U2967 (N_2967,N_2913,N_2926);
and U2968 (N_2968,N_2929,N_2897);
nor U2969 (N_2969,N_2889,N_2906);
or U2970 (N_2970,N_2937,N_2910);
xor U2971 (N_2971,N_2900,N_2919);
and U2972 (N_2972,N_2927,N_2883);
nor U2973 (N_2973,N_2882,N_2930);
nand U2974 (N_2974,N_2935,N_2913);
and U2975 (N_2975,N_2939,N_2923);
xnor U2976 (N_2976,N_2928,N_2915);
nand U2977 (N_2977,N_2931,N_2925);
nor U2978 (N_2978,N_2911,N_2880);
nand U2979 (N_2979,N_2928,N_2932);
nand U2980 (N_2980,N_2904,N_2897);
nor U2981 (N_2981,N_2893,N_2901);
or U2982 (N_2982,N_2932,N_2905);
nand U2983 (N_2983,N_2906,N_2898);
nor U2984 (N_2984,N_2901,N_2891);
and U2985 (N_2985,N_2901,N_2884);
and U2986 (N_2986,N_2923,N_2916);
nor U2987 (N_2987,N_2900,N_2883);
or U2988 (N_2988,N_2914,N_2902);
nor U2989 (N_2989,N_2893,N_2899);
nand U2990 (N_2990,N_2935,N_2920);
and U2991 (N_2991,N_2931,N_2911);
nand U2992 (N_2992,N_2888,N_2923);
or U2993 (N_2993,N_2885,N_2932);
or U2994 (N_2994,N_2893,N_2910);
and U2995 (N_2995,N_2885,N_2888);
and U2996 (N_2996,N_2886,N_2921);
nand U2997 (N_2997,N_2921,N_2930);
or U2998 (N_2998,N_2881,N_2892);
and U2999 (N_2999,N_2887,N_2885);
nor UO_0 (O_0,N_2972,N_2950);
nor UO_1 (O_1,N_2995,N_2986);
nor UO_2 (O_2,N_2994,N_2958);
or UO_3 (O_3,N_2945,N_2957);
nand UO_4 (O_4,N_2999,N_2956);
and UO_5 (O_5,N_2962,N_2946);
and UO_6 (O_6,N_2959,N_2961);
or UO_7 (O_7,N_2951,N_2940);
or UO_8 (O_8,N_2990,N_2979);
or UO_9 (O_9,N_2965,N_2977);
or UO_10 (O_10,N_2984,N_2996);
xor UO_11 (O_11,N_2941,N_2970);
nor UO_12 (O_12,N_2967,N_2983);
nand UO_13 (O_13,N_2942,N_2981);
nand UO_14 (O_14,N_2980,N_2964);
nand UO_15 (O_15,N_2943,N_2989);
and UO_16 (O_16,N_2949,N_2973);
and UO_17 (O_17,N_2954,N_2988);
nand UO_18 (O_18,N_2963,N_2971);
or UO_19 (O_19,N_2955,N_2944);
nand UO_20 (O_20,N_2978,N_2966);
nor UO_21 (O_21,N_2991,N_2948);
nor UO_22 (O_22,N_2976,N_2985);
nand UO_23 (O_23,N_2960,N_2975);
nand UO_24 (O_24,N_2982,N_2969);
nand UO_25 (O_25,N_2998,N_2992);
or UO_26 (O_26,N_2974,N_2968);
nor UO_27 (O_27,N_2997,N_2952);
xor UO_28 (O_28,N_2987,N_2993);
nand UO_29 (O_29,N_2947,N_2953);
or UO_30 (O_30,N_2985,N_2943);
nor UO_31 (O_31,N_2994,N_2948);
and UO_32 (O_32,N_2984,N_2944);
or UO_33 (O_33,N_2997,N_2959);
nor UO_34 (O_34,N_2974,N_2948);
and UO_35 (O_35,N_2948,N_2957);
nor UO_36 (O_36,N_2993,N_2983);
or UO_37 (O_37,N_2985,N_2959);
or UO_38 (O_38,N_2961,N_2993);
or UO_39 (O_39,N_2957,N_2988);
nand UO_40 (O_40,N_2953,N_2961);
xor UO_41 (O_41,N_2965,N_2994);
or UO_42 (O_42,N_2984,N_2994);
or UO_43 (O_43,N_2985,N_2996);
and UO_44 (O_44,N_2977,N_2940);
and UO_45 (O_45,N_2993,N_2964);
nand UO_46 (O_46,N_2971,N_2982);
nor UO_47 (O_47,N_2992,N_2982);
nor UO_48 (O_48,N_2986,N_2953);
nand UO_49 (O_49,N_2977,N_2991);
nand UO_50 (O_50,N_2951,N_2986);
and UO_51 (O_51,N_2978,N_2960);
nor UO_52 (O_52,N_2992,N_2974);
nand UO_53 (O_53,N_2966,N_2942);
or UO_54 (O_54,N_2962,N_2941);
nand UO_55 (O_55,N_2983,N_2958);
nand UO_56 (O_56,N_2974,N_2947);
and UO_57 (O_57,N_2991,N_2965);
nand UO_58 (O_58,N_2949,N_2989);
nand UO_59 (O_59,N_2943,N_2966);
nor UO_60 (O_60,N_2965,N_2988);
nand UO_61 (O_61,N_2979,N_2956);
and UO_62 (O_62,N_2973,N_2968);
or UO_63 (O_63,N_2940,N_2996);
and UO_64 (O_64,N_2941,N_2989);
or UO_65 (O_65,N_2994,N_2946);
and UO_66 (O_66,N_2943,N_2976);
and UO_67 (O_67,N_2944,N_2991);
or UO_68 (O_68,N_2975,N_2966);
or UO_69 (O_69,N_2965,N_2986);
and UO_70 (O_70,N_2949,N_2964);
nand UO_71 (O_71,N_2946,N_2977);
and UO_72 (O_72,N_2948,N_2940);
nor UO_73 (O_73,N_2960,N_2980);
or UO_74 (O_74,N_2970,N_2983);
nor UO_75 (O_75,N_2977,N_2949);
or UO_76 (O_76,N_2940,N_2966);
or UO_77 (O_77,N_2942,N_2960);
nand UO_78 (O_78,N_2977,N_2948);
and UO_79 (O_79,N_2979,N_2963);
nor UO_80 (O_80,N_2941,N_2978);
or UO_81 (O_81,N_2991,N_2956);
and UO_82 (O_82,N_2958,N_2949);
and UO_83 (O_83,N_2980,N_2975);
nand UO_84 (O_84,N_2978,N_2982);
or UO_85 (O_85,N_2942,N_2941);
or UO_86 (O_86,N_2976,N_2971);
and UO_87 (O_87,N_2981,N_2983);
and UO_88 (O_88,N_2982,N_2943);
nand UO_89 (O_89,N_2956,N_2971);
nor UO_90 (O_90,N_2947,N_2990);
or UO_91 (O_91,N_2971,N_2958);
nand UO_92 (O_92,N_2992,N_2961);
and UO_93 (O_93,N_2975,N_2998);
nor UO_94 (O_94,N_2996,N_2951);
nand UO_95 (O_95,N_2988,N_2995);
nand UO_96 (O_96,N_2946,N_2988);
or UO_97 (O_97,N_2978,N_2953);
and UO_98 (O_98,N_2952,N_2946);
and UO_99 (O_99,N_2942,N_2974);
or UO_100 (O_100,N_2958,N_2981);
or UO_101 (O_101,N_2961,N_2979);
or UO_102 (O_102,N_2949,N_2960);
nor UO_103 (O_103,N_2970,N_2980);
and UO_104 (O_104,N_2978,N_2956);
nor UO_105 (O_105,N_2979,N_2946);
and UO_106 (O_106,N_2951,N_2954);
nor UO_107 (O_107,N_2994,N_2950);
or UO_108 (O_108,N_2960,N_2940);
or UO_109 (O_109,N_2945,N_2940);
nor UO_110 (O_110,N_2985,N_2991);
nand UO_111 (O_111,N_2963,N_2950);
and UO_112 (O_112,N_2944,N_2983);
or UO_113 (O_113,N_2951,N_2965);
and UO_114 (O_114,N_2999,N_2984);
and UO_115 (O_115,N_2990,N_2957);
nand UO_116 (O_116,N_2984,N_2989);
and UO_117 (O_117,N_2951,N_2980);
nand UO_118 (O_118,N_2953,N_2989);
nor UO_119 (O_119,N_2941,N_2971);
nor UO_120 (O_120,N_2956,N_2984);
nor UO_121 (O_121,N_2977,N_2983);
or UO_122 (O_122,N_2964,N_2966);
and UO_123 (O_123,N_2941,N_2976);
nand UO_124 (O_124,N_2941,N_2958);
or UO_125 (O_125,N_2967,N_2954);
and UO_126 (O_126,N_2984,N_2952);
nand UO_127 (O_127,N_2994,N_2991);
nand UO_128 (O_128,N_2961,N_2998);
xnor UO_129 (O_129,N_2951,N_2981);
nand UO_130 (O_130,N_2943,N_2946);
and UO_131 (O_131,N_2980,N_2998);
nand UO_132 (O_132,N_2974,N_2989);
and UO_133 (O_133,N_2958,N_2972);
nand UO_134 (O_134,N_2950,N_2955);
nor UO_135 (O_135,N_2977,N_2945);
xnor UO_136 (O_136,N_2996,N_2955);
nand UO_137 (O_137,N_2982,N_2998);
nand UO_138 (O_138,N_2949,N_2997);
nor UO_139 (O_139,N_2954,N_2982);
and UO_140 (O_140,N_2953,N_2943);
and UO_141 (O_141,N_2985,N_2953);
and UO_142 (O_142,N_2941,N_2986);
nand UO_143 (O_143,N_2940,N_2952);
nand UO_144 (O_144,N_2966,N_2994);
nor UO_145 (O_145,N_2954,N_2985);
nand UO_146 (O_146,N_2946,N_2945);
or UO_147 (O_147,N_2983,N_2954);
and UO_148 (O_148,N_2991,N_2960);
nand UO_149 (O_149,N_2955,N_2978);
or UO_150 (O_150,N_2971,N_2944);
nand UO_151 (O_151,N_2957,N_2942);
and UO_152 (O_152,N_2976,N_2959);
or UO_153 (O_153,N_2989,N_2990);
nor UO_154 (O_154,N_2953,N_2944);
or UO_155 (O_155,N_2976,N_2998);
nand UO_156 (O_156,N_2999,N_2978);
nor UO_157 (O_157,N_2954,N_2997);
or UO_158 (O_158,N_2977,N_2990);
nor UO_159 (O_159,N_2952,N_2983);
nand UO_160 (O_160,N_2952,N_2971);
and UO_161 (O_161,N_2954,N_2974);
or UO_162 (O_162,N_2964,N_2969);
nand UO_163 (O_163,N_2948,N_2963);
nand UO_164 (O_164,N_2984,N_2997);
or UO_165 (O_165,N_2963,N_2986);
and UO_166 (O_166,N_2995,N_2960);
nand UO_167 (O_167,N_2990,N_2966);
or UO_168 (O_168,N_2998,N_2967);
or UO_169 (O_169,N_2981,N_2971);
nor UO_170 (O_170,N_2940,N_2941);
nor UO_171 (O_171,N_2947,N_2941);
nor UO_172 (O_172,N_2992,N_2981);
nor UO_173 (O_173,N_2968,N_2951);
and UO_174 (O_174,N_2965,N_2956);
nand UO_175 (O_175,N_2948,N_2966);
nor UO_176 (O_176,N_2970,N_2944);
or UO_177 (O_177,N_2982,N_2981);
nor UO_178 (O_178,N_2948,N_2995);
nor UO_179 (O_179,N_2961,N_2947);
and UO_180 (O_180,N_2969,N_2973);
nand UO_181 (O_181,N_2982,N_2987);
or UO_182 (O_182,N_2980,N_2949);
or UO_183 (O_183,N_2954,N_2987);
and UO_184 (O_184,N_2964,N_2977);
or UO_185 (O_185,N_2965,N_2941);
nor UO_186 (O_186,N_2991,N_2954);
nand UO_187 (O_187,N_2996,N_2982);
xnor UO_188 (O_188,N_2950,N_2996);
nor UO_189 (O_189,N_2965,N_2946);
nor UO_190 (O_190,N_2986,N_2961);
and UO_191 (O_191,N_2993,N_2958);
and UO_192 (O_192,N_2957,N_2959);
nor UO_193 (O_193,N_2946,N_2967);
nand UO_194 (O_194,N_2983,N_2942);
or UO_195 (O_195,N_2976,N_2997);
and UO_196 (O_196,N_2987,N_2984);
nor UO_197 (O_197,N_2972,N_2998);
nand UO_198 (O_198,N_2964,N_2983);
or UO_199 (O_199,N_2958,N_2957);
and UO_200 (O_200,N_2988,N_2952);
nor UO_201 (O_201,N_2988,N_2978);
and UO_202 (O_202,N_2980,N_2966);
nor UO_203 (O_203,N_2973,N_2943);
and UO_204 (O_204,N_2988,N_2993);
nand UO_205 (O_205,N_2994,N_2960);
or UO_206 (O_206,N_2964,N_2943);
and UO_207 (O_207,N_2960,N_2993);
nand UO_208 (O_208,N_2965,N_2998);
nand UO_209 (O_209,N_2991,N_2983);
or UO_210 (O_210,N_2946,N_2975);
and UO_211 (O_211,N_2954,N_2948);
nand UO_212 (O_212,N_2953,N_2972);
or UO_213 (O_213,N_2991,N_2959);
and UO_214 (O_214,N_2978,N_2983);
and UO_215 (O_215,N_2967,N_2993);
and UO_216 (O_216,N_2969,N_2986);
or UO_217 (O_217,N_2969,N_2988);
and UO_218 (O_218,N_2991,N_2970);
nand UO_219 (O_219,N_2956,N_2945);
nor UO_220 (O_220,N_2974,N_2969);
nor UO_221 (O_221,N_2945,N_2989);
or UO_222 (O_222,N_2944,N_2961);
nor UO_223 (O_223,N_2973,N_2954);
or UO_224 (O_224,N_2997,N_2969);
nor UO_225 (O_225,N_2986,N_2950);
nor UO_226 (O_226,N_2952,N_2989);
nand UO_227 (O_227,N_2967,N_2973);
nand UO_228 (O_228,N_2948,N_2962);
nand UO_229 (O_229,N_2954,N_2977);
or UO_230 (O_230,N_2966,N_2955);
and UO_231 (O_231,N_2996,N_2971);
or UO_232 (O_232,N_2990,N_2999);
and UO_233 (O_233,N_2951,N_2988);
nor UO_234 (O_234,N_2986,N_2968);
or UO_235 (O_235,N_2991,N_2978);
or UO_236 (O_236,N_2975,N_2969);
or UO_237 (O_237,N_2943,N_2987);
nor UO_238 (O_238,N_2948,N_2947);
or UO_239 (O_239,N_2966,N_2972);
and UO_240 (O_240,N_2956,N_2958);
or UO_241 (O_241,N_2998,N_2974);
and UO_242 (O_242,N_2951,N_2976);
or UO_243 (O_243,N_2966,N_2941);
nor UO_244 (O_244,N_2981,N_2953);
and UO_245 (O_245,N_2990,N_2974);
nor UO_246 (O_246,N_2997,N_2973);
and UO_247 (O_247,N_2971,N_2955);
or UO_248 (O_248,N_2999,N_2981);
nand UO_249 (O_249,N_2952,N_2948);
nor UO_250 (O_250,N_2962,N_2998);
and UO_251 (O_251,N_2994,N_2972);
nor UO_252 (O_252,N_2947,N_2951);
and UO_253 (O_253,N_2969,N_2999);
nand UO_254 (O_254,N_2991,N_2997);
nor UO_255 (O_255,N_2957,N_2941);
nor UO_256 (O_256,N_2997,N_2947);
and UO_257 (O_257,N_2962,N_2986);
or UO_258 (O_258,N_2960,N_2948);
nand UO_259 (O_259,N_2956,N_2996);
and UO_260 (O_260,N_2943,N_2940);
nand UO_261 (O_261,N_2966,N_2988);
and UO_262 (O_262,N_2973,N_2970);
nand UO_263 (O_263,N_2995,N_2943);
or UO_264 (O_264,N_2952,N_2955);
nor UO_265 (O_265,N_2989,N_2964);
nand UO_266 (O_266,N_2986,N_2960);
nand UO_267 (O_267,N_2985,N_2958);
and UO_268 (O_268,N_2981,N_2998);
nor UO_269 (O_269,N_2972,N_2943);
and UO_270 (O_270,N_2945,N_2976);
nand UO_271 (O_271,N_2956,N_2973);
and UO_272 (O_272,N_2966,N_2971);
and UO_273 (O_273,N_2943,N_2988);
nor UO_274 (O_274,N_2984,N_2988);
and UO_275 (O_275,N_2953,N_2964);
or UO_276 (O_276,N_2987,N_2977);
nand UO_277 (O_277,N_2982,N_2990);
and UO_278 (O_278,N_2989,N_2980);
or UO_279 (O_279,N_2949,N_2948);
nor UO_280 (O_280,N_2993,N_2990);
or UO_281 (O_281,N_2982,N_2946);
nand UO_282 (O_282,N_2957,N_2980);
or UO_283 (O_283,N_2985,N_2982);
and UO_284 (O_284,N_2975,N_2951);
and UO_285 (O_285,N_2969,N_2979);
or UO_286 (O_286,N_2979,N_2987);
and UO_287 (O_287,N_2946,N_2949);
and UO_288 (O_288,N_2970,N_2947);
and UO_289 (O_289,N_2997,N_2948);
or UO_290 (O_290,N_2985,N_2992);
or UO_291 (O_291,N_2983,N_2969);
nand UO_292 (O_292,N_2980,N_2997);
or UO_293 (O_293,N_2998,N_2949);
nor UO_294 (O_294,N_2959,N_2969);
or UO_295 (O_295,N_2965,N_2985);
nand UO_296 (O_296,N_2996,N_2957);
nor UO_297 (O_297,N_2948,N_2990);
or UO_298 (O_298,N_2965,N_2999);
or UO_299 (O_299,N_2955,N_2983);
or UO_300 (O_300,N_2966,N_2977);
and UO_301 (O_301,N_2989,N_2960);
or UO_302 (O_302,N_2963,N_2969);
nand UO_303 (O_303,N_2974,N_2984);
xor UO_304 (O_304,N_2945,N_2947);
nor UO_305 (O_305,N_2983,N_2960);
nand UO_306 (O_306,N_2962,N_2950);
and UO_307 (O_307,N_2955,N_2995);
nor UO_308 (O_308,N_2961,N_2997);
nand UO_309 (O_309,N_2977,N_2961);
nand UO_310 (O_310,N_2954,N_2959);
nor UO_311 (O_311,N_2985,N_2968);
or UO_312 (O_312,N_2962,N_2989);
nand UO_313 (O_313,N_2949,N_2944);
nand UO_314 (O_314,N_2972,N_2968);
nand UO_315 (O_315,N_2984,N_2943);
nor UO_316 (O_316,N_2965,N_2961);
and UO_317 (O_317,N_2958,N_2989);
or UO_318 (O_318,N_2978,N_2981);
nand UO_319 (O_319,N_2943,N_2970);
nor UO_320 (O_320,N_2952,N_2970);
nor UO_321 (O_321,N_2956,N_2957);
and UO_322 (O_322,N_2950,N_2945);
nand UO_323 (O_323,N_2960,N_2979);
and UO_324 (O_324,N_2976,N_2981);
nand UO_325 (O_325,N_2988,N_2945);
nor UO_326 (O_326,N_2974,N_2958);
or UO_327 (O_327,N_2971,N_2974);
nand UO_328 (O_328,N_2964,N_2942);
and UO_329 (O_329,N_2992,N_2971);
nand UO_330 (O_330,N_2971,N_2977);
nand UO_331 (O_331,N_2982,N_2963);
or UO_332 (O_332,N_2979,N_2940);
nor UO_333 (O_333,N_2997,N_2977);
or UO_334 (O_334,N_2943,N_2967);
and UO_335 (O_335,N_2954,N_2966);
or UO_336 (O_336,N_2964,N_2940);
nand UO_337 (O_337,N_2961,N_2971);
or UO_338 (O_338,N_2959,N_2964);
and UO_339 (O_339,N_2960,N_2953);
nor UO_340 (O_340,N_2973,N_2945);
or UO_341 (O_341,N_2991,N_2951);
nand UO_342 (O_342,N_2949,N_2951);
and UO_343 (O_343,N_2958,N_2945);
nor UO_344 (O_344,N_2941,N_2944);
and UO_345 (O_345,N_2995,N_2940);
nor UO_346 (O_346,N_2950,N_2940);
or UO_347 (O_347,N_2993,N_2998);
or UO_348 (O_348,N_2986,N_2993);
xor UO_349 (O_349,N_2989,N_2999);
nand UO_350 (O_350,N_2944,N_2996);
nor UO_351 (O_351,N_2971,N_2947);
nand UO_352 (O_352,N_2942,N_2961);
or UO_353 (O_353,N_2944,N_2958);
nor UO_354 (O_354,N_2956,N_2962);
nand UO_355 (O_355,N_2960,N_2999);
nor UO_356 (O_356,N_2953,N_2975);
nor UO_357 (O_357,N_2980,N_2983);
and UO_358 (O_358,N_2987,N_2941);
nor UO_359 (O_359,N_2999,N_2968);
or UO_360 (O_360,N_2989,N_2988);
nand UO_361 (O_361,N_2988,N_2975);
or UO_362 (O_362,N_2983,N_2943);
and UO_363 (O_363,N_2951,N_2989);
and UO_364 (O_364,N_2991,N_2947);
and UO_365 (O_365,N_2980,N_2973);
or UO_366 (O_366,N_2998,N_2969);
nor UO_367 (O_367,N_2990,N_2968);
nor UO_368 (O_368,N_2965,N_2974);
nor UO_369 (O_369,N_2972,N_2959);
nor UO_370 (O_370,N_2990,N_2956);
nand UO_371 (O_371,N_2969,N_2977);
or UO_372 (O_372,N_2997,N_2995);
nand UO_373 (O_373,N_2946,N_2997);
and UO_374 (O_374,N_2955,N_2993);
nand UO_375 (O_375,N_2973,N_2962);
nor UO_376 (O_376,N_2948,N_2968);
nand UO_377 (O_377,N_2980,N_2945);
nor UO_378 (O_378,N_2985,N_2966);
or UO_379 (O_379,N_2972,N_2963);
and UO_380 (O_380,N_2963,N_2964);
nand UO_381 (O_381,N_2944,N_2977);
nand UO_382 (O_382,N_2970,N_2966);
nand UO_383 (O_383,N_2960,N_2951);
nand UO_384 (O_384,N_2968,N_2978);
and UO_385 (O_385,N_2951,N_2944);
nand UO_386 (O_386,N_2993,N_2971);
nor UO_387 (O_387,N_2981,N_2943);
and UO_388 (O_388,N_2942,N_2955);
or UO_389 (O_389,N_2994,N_2945);
nand UO_390 (O_390,N_2951,N_2957);
nand UO_391 (O_391,N_2987,N_2964);
xor UO_392 (O_392,N_2968,N_2947);
and UO_393 (O_393,N_2999,N_2942);
nand UO_394 (O_394,N_2982,N_2959);
nor UO_395 (O_395,N_2988,N_2985);
or UO_396 (O_396,N_2981,N_2956);
or UO_397 (O_397,N_2953,N_2988);
nor UO_398 (O_398,N_2994,N_2959);
nor UO_399 (O_399,N_2998,N_2978);
and UO_400 (O_400,N_2946,N_2941);
or UO_401 (O_401,N_2988,N_2976);
or UO_402 (O_402,N_2943,N_2941);
or UO_403 (O_403,N_2966,N_2996);
nand UO_404 (O_404,N_2957,N_2995);
or UO_405 (O_405,N_2977,N_2941);
nor UO_406 (O_406,N_2973,N_2944);
nor UO_407 (O_407,N_2983,N_2990);
nor UO_408 (O_408,N_2943,N_2994);
nor UO_409 (O_409,N_2964,N_2955);
and UO_410 (O_410,N_2960,N_2972);
or UO_411 (O_411,N_2969,N_2992);
nand UO_412 (O_412,N_2977,N_2973);
or UO_413 (O_413,N_2958,N_2953);
or UO_414 (O_414,N_2983,N_2968);
or UO_415 (O_415,N_2946,N_2996);
and UO_416 (O_416,N_2940,N_2984);
and UO_417 (O_417,N_2951,N_2973);
nor UO_418 (O_418,N_2998,N_2956);
nand UO_419 (O_419,N_2987,N_2960);
and UO_420 (O_420,N_2989,N_2957);
nand UO_421 (O_421,N_2964,N_2974);
nand UO_422 (O_422,N_2969,N_2955);
and UO_423 (O_423,N_2981,N_2965);
or UO_424 (O_424,N_2954,N_2964);
nand UO_425 (O_425,N_2962,N_2958);
nand UO_426 (O_426,N_2973,N_2992);
and UO_427 (O_427,N_2950,N_2970);
nor UO_428 (O_428,N_2972,N_2999);
nor UO_429 (O_429,N_2987,N_2996);
or UO_430 (O_430,N_2957,N_2968);
and UO_431 (O_431,N_2957,N_2947);
nand UO_432 (O_432,N_2961,N_2954);
and UO_433 (O_433,N_2945,N_2952);
or UO_434 (O_434,N_2966,N_2981);
nand UO_435 (O_435,N_2951,N_2966);
and UO_436 (O_436,N_2994,N_2947);
or UO_437 (O_437,N_2958,N_2964);
nand UO_438 (O_438,N_2957,N_2974);
or UO_439 (O_439,N_2966,N_2974);
nand UO_440 (O_440,N_2983,N_2982);
nor UO_441 (O_441,N_2961,N_2960);
or UO_442 (O_442,N_2944,N_2948);
and UO_443 (O_443,N_2987,N_2959);
and UO_444 (O_444,N_2974,N_2975);
nor UO_445 (O_445,N_2981,N_2973);
nor UO_446 (O_446,N_2955,N_2987);
nor UO_447 (O_447,N_2995,N_2964);
nor UO_448 (O_448,N_2959,N_2956);
and UO_449 (O_449,N_2975,N_2978);
and UO_450 (O_450,N_2945,N_2993);
xor UO_451 (O_451,N_2963,N_2997);
or UO_452 (O_452,N_2992,N_2955);
or UO_453 (O_453,N_2972,N_2974);
nand UO_454 (O_454,N_2962,N_2944);
or UO_455 (O_455,N_2963,N_2999);
or UO_456 (O_456,N_2990,N_2950);
nand UO_457 (O_457,N_2958,N_2996);
and UO_458 (O_458,N_2979,N_2983);
nor UO_459 (O_459,N_2986,N_2982);
nor UO_460 (O_460,N_2989,N_2993);
nand UO_461 (O_461,N_2970,N_2946);
or UO_462 (O_462,N_2990,N_2945);
or UO_463 (O_463,N_2986,N_2996);
nand UO_464 (O_464,N_2958,N_2960);
nand UO_465 (O_465,N_2961,N_2948);
nor UO_466 (O_466,N_2999,N_2991);
nand UO_467 (O_467,N_2986,N_2955);
or UO_468 (O_468,N_2970,N_2975);
nand UO_469 (O_469,N_2951,N_2995);
nand UO_470 (O_470,N_2992,N_2944);
or UO_471 (O_471,N_2955,N_2972);
nand UO_472 (O_472,N_2974,N_2943);
or UO_473 (O_473,N_2953,N_2955);
nor UO_474 (O_474,N_2989,N_2977);
nand UO_475 (O_475,N_2946,N_2974);
nor UO_476 (O_476,N_2981,N_2985);
nand UO_477 (O_477,N_2972,N_2985);
nor UO_478 (O_478,N_2967,N_2987);
nor UO_479 (O_479,N_2949,N_2995);
nand UO_480 (O_480,N_2972,N_2992);
nor UO_481 (O_481,N_2980,N_2953);
and UO_482 (O_482,N_2996,N_2942);
or UO_483 (O_483,N_2964,N_2950);
and UO_484 (O_484,N_2973,N_2964);
nand UO_485 (O_485,N_2977,N_2974);
nand UO_486 (O_486,N_2991,N_2996);
nand UO_487 (O_487,N_2956,N_2966);
nand UO_488 (O_488,N_2997,N_2962);
and UO_489 (O_489,N_2966,N_2950);
or UO_490 (O_490,N_2965,N_2954);
nand UO_491 (O_491,N_2984,N_2961);
and UO_492 (O_492,N_2985,N_2989);
nand UO_493 (O_493,N_2992,N_2990);
and UO_494 (O_494,N_2945,N_2981);
xnor UO_495 (O_495,N_2980,N_2948);
nand UO_496 (O_496,N_2945,N_2969);
nand UO_497 (O_497,N_2970,N_2967);
and UO_498 (O_498,N_2976,N_2955);
nor UO_499 (O_499,N_2968,N_2998);
endmodule