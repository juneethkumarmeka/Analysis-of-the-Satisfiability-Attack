module basic_500_3000_500_15_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xor U0 (N_0,In_124,In_304);
xnor U1 (N_1,In_20,In_131);
nand U2 (N_2,In_177,In_192);
xor U3 (N_3,In_487,In_82);
and U4 (N_4,In_447,In_418);
nand U5 (N_5,In_452,In_331);
nor U6 (N_6,In_383,In_499);
nand U7 (N_7,In_8,In_135);
or U8 (N_8,In_88,In_468);
and U9 (N_9,In_337,In_220);
nand U10 (N_10,In_457,In_187);
or U11 (N_11,In_108,In_342);
or U12 (N_12,In_287,In_214);
nor U13 (N_13,In_444,In_264);
nand U14 (N_14,In_492,In_190);
xnor U15 (N_15,In_181,In_169);
nor U16 (N_16,In_285,In_228);
or U17 (N_17,In_47,In_308);
or U18 (N_18,In_407,In_204);
or U19 (N_19,In_385,In_146);
nand U20 (N_20,In_394,In_266);
nand U21 (N_21,In_224,In_134);
and U22 (N_22,In_55,In_436);
and U23 (N_23,In_262,In_327);
xor U24 (N_24,In_302,In_74);
nand U25 (N_25,In_199,In_207);
nor U26 (N_26,In_116,In_217);
nand U27 (N_27,In_363,In_222);
or U28 (N_28,In_281,In_320);
nand U29 (N_29,In_380,In_73);
nor U30 (N_30,In_6,In_361);
xnor U31 (N_31,In_58,In_85);
nor U32 (N_32,In_369,In_141);
and U33 (N_33,In_7,In_84);
nand U34 (N_34,In_432,In_422);
nor U35 (N_35,In_333,In_32);
or U36 (N_36,In_38,In_184);
nand U37 (N_37,In_392,In_283);
or U38 (N_38,In_317,In_196);
nand U39 (N_39,In_482,In_93);
nand U40 (N_40,In_273,In_276);
and U41 (N_41,In_99,In_185);
and U42 (N_42,In_257,In_12);
and U43 (N_43,In_296,In_90);
or U44 (N_44,In_386,In_255);
or U45 (N_45,In_293,In_51);
nand U46 (N_46,In_338,In_19);
xnor U47 (N_47,In_315,In_357);
nor U48 (N_48,In_230,In_106);
nand U49 (N_49,In_388,In_269);
and U50 (N_50,In_147,In_391);
or U51 (N_51,In_140,In_493);
and U52 (N_52,In_119,In_201);
and U53 (N_53,In_424,In_367);
or U54 (N_54,In_270,In_61);
nor U55 (N_55,In_408,In_200);
xor U56 (N_56,In_234,In_110);
xnor U57 (N_57,In_247,In_485);
or U58 (N_58,In_491,In_4);
nor U59 (N_59,In_25,In_133);
xnor U60 (N_60,In_87,In_384);
xnor U61 (N_61,In_465,In_243);
xnor U62 (N_62,In_488,In_414);
nor U63 (N_63,In_328,In_301);
nand U64 (N_64,In_368,In_105);
xor U65 (N_65,In_313,In_372);
nand U66 (N_66,In_80,In_377);
nand U67 (N_67,In_43,In_129);
nor U68 (N_68,In_14,In_341);
or U69 (N_69,In_433,In_59);
or U70 (N_70,In_23,In_280);
nor U71 (N_71,In_162,In_278);
and U72 (N_72,In_183,In_178);
nand U73 (N_73,In_197,In_261);
nand U74 (N_74,In_164,In_344);
nand U75 (N_75,In_481,In_490);
or U76 (N_76,In_21,In_467);
nor U77 (N_77,In_271,In_48);
nand U78 (N_78,In_168,In_477);
or U79 (N_79,In_448,In_390);
nor U80 (N_80,In_460,In_494);
nand U81 (N_81,In_473,In_451);
or U82 (N_82,In_314,In_104);
or U83 (N_83,In_226,In_152);
and U84 (N_84,In_321,In_299);
nand U85 (N_85,In_113,In_34);
nand U86 (N_86,In_239,In_286);
nand U87 (N_87,In_66,In_282);
and U88 (N_88,In_441,In_98);
xnor U89 (N_89,In_475,In_193);
nor U90 (N_90,In_236,In_160);
or U91 (N_91,In_289,In_91);
or U92 (N_92,In_428,In_86);
and U93 (N_93,In_415,In_175);
and U94 (N_94,In_150,In_248);
and U95 (N_95,In_225,In_348);
xnor U96 (N_96,In_268,In_145);
nor U97 (N_97,In_332,In_254);
or U98 (N_98,In_443,In_495);
nand U99 (N_99,In_366,In_202);
nor U100 (N_100,In_118,In_421);
nand U101 (N_101,In_470,In_362);
or U102 (N_102,In_159,In_126);
or U103 (N_103,In_65,In_155);
nor U104 (N_104,In_330,In_29);
and U105 (N_105,In_396,In_212);
and U106 (N_106,In_191,In_256);
and U107 (N_107,In_137,In_426);
and U108 (N_108,In_478,In_253);
and U109 (N_109,In_401,In_456);
or U110 (N_110,In_486,In_339);
and U111 (N_111,In_358,In_103);
and U112 (N_112,In_36,In_128);
or U113 (N_113,In_322,In_431);
or U114 (N_114,In_307,In_354);
or U115 (N_115,In_397,In_346);
and U116 (N_116,In_284,In_437);
nor U117 (N_117,In_345,In_132);
xor U118 (N_118,In_3,In_425);
xnor U119 (N_119,In_483,In_434);
xnor U120 (N_120,In_497,In_123);
or U121 (N_121,In_355,In_218);
nor U122 (N_122,In_259,In_381);
and U123 (N_123,In_420,In_265);
nor U124 (N_124,In_144,In_62);
nand U125 (N_125,In_423,In_455);
and U126 (N_126,In_79,In_233);
or U127 (N_127,In_379,In_306);
nand U128 (N_128,In_1,In_438);
or U129 (N_129,In_472,In_263);
xnor U130 (N_130,In_311,In_430);
or U131 (N_131,In_68,In_165);
nand U132 (N_132,In_2,In_359);
nand U133 (N_133,In_210,In_153);
or U134 (N_134,In_142,In_458);
and U135 (N_135,In_179,In_411);
nand U136 (N_136,In_112,In_274);
or U137 (N_137,In_292,In_462);
nor U138 (N_138,In_42,In_417);
nand U139 (N_139,In_52,In_101);
and U140 (N_140,In_72,In_245);
nand U141 (N_141,In_33,In_238);
or U142 (N_142,In_240,In_40);
and U143 (N_143,In_413,In_291);
nor U144 (N_144,In_387,In_406);
or U145 (N_145,In_77,In_275);
xor U146 (N_146,In_27,In_16);
nor U147 (N_147,In_241,In_139);
and U148 (N_148,In_167,In_251);
xor U149 (N_149,In_158,In_298);
and U150 (N_150,In_400,In_429);
or U151 (N_151,In_120,In_75);
nand U152 (N_152,In_449,In_35);
nand U153 (N_153,In_409,In_114);
nand U154 (N_154,In_17,In_67);
or U155 (N_155,In_136,In_10);
or U156 (N_156,In_297,In_189);
xnor U157 (N_157,In_439,In_166);
nor U158 (N_158,In_182,In_111);
nor U159 (N_159,In_360,In_252);
xor U160 (N_160,In_365,In_300);
nor U161 (N_161,In_350,In_326);
xnor U162 (N_162,In_419,In_30);
nand U163 (N_163,In_54,In_246);
or U164 (N_164,In_356,In_229);
nand U165 (N_165,In_352,In_279);
nor U166 (N_166,In_46,In_435);
or U167 (N_167,In_45,In_28);
and U168 (N_168,In_63,In_39);
xnor U169 (N_169,In_97,In_49);
xor U170 (N_170,In_410,In_31);
nor U171 (N_171,In_498,In_476);
nand U172 (N_172,In_375,In_156);
and U173 (N_173,In_471,In_316);
or U174 (N_174,In_170,In_53);
xnor U175 (N_175,In_267,In_26);
or U176 (N_176,In_107,In_41);
nand U177 (N_177,In_95,In_496);
or U178 (N_178,In_393,In_474);
or U179 (N_179,In_454,In_398);
nand U180 (N_180,In_399,In_353);
nand U181 (N_181,In_102,In_213);
nor U182 (N_182,In_195,In_89);
and U183 (N_183,In_389,In_60);
and U184 (N_184,In_446,In_157);
and U185 (N_185,In_24,In_403);
nand U186 (N_186,In_161,In_215);
or U187 (N_187,In_83,In_223);
nand U188 (N_188,In_76,In_219);
and U189 (N_189,In_249,In_371);
or U190 (N_190,In_5,In_427);
nor U191 (N_191,In_64,In_71);
xnor U192 (N_192,In_237,In_312);
nor U193 (N_193,In_69,In_370);
and U194 (N_194,In_347,In_176);
nor U195 (N_195,In_303,In_318);
and U196 (N_196,In_378,In_295);
xnor U197 (N_197,In_288,In_172);
nor U198 (N_198,In_412,In_149);
and U199 (N_199,In_489,In_13);
and U200 (N_200,In_211,N_130);
nand U201 (N_201,N_20,N_127);
and U202 (N_202,In_203,In_221);
or U203 (N_203,In_395,N_197);
nor U204 (N_204,N_104,N_164);
or U205 (N_205,N_150,In_469);
or U206 (N_206,N_165,In_463);
or U207 (N_207,In_81,N_152);
or U208 (N_208,N_80,N_196);
nor U209 (N_209,In_18,N_12);
nor U210 (N_210,N_180,In_480);
or U211 (N_211,In_9,N_6);
nor U212 (N_212,N_143,In_231);
and U213 (N_213,N_126,N_70);
xnor U214 (N_214,N_101,N_192);
and U215 (N_215,In_376,N_147);
nor U216 (N_216,In_484,N_75);
nor U217 (N_217,In_216,N_184);
nor U218 (N_218,N_145,N_117);
xnor U219 (N_219,N_4,N_124);
or U220 (N_220,N_106,N_29);
xor U221 (N_221,N_69,N_142);
xor U222 (N_222,N_44,N_33);
and U223 (N_223,In_242,N_7);
nor U224 (N_224,In_277,N_157);
or U225 (N_225,N_32,In_96);
nand U226 (N_226,N_84,N_108);
nor U227 (N_227,N_120,In_479);
nor U228 (N_228,N_53,N_25);
nand U229 (N_229,N_36,In_148);
nand U230 (N_230,N_11,N_131);
or U231 (N_231,In_272,N_110);
or U232 (N_232,N_85,N_139);
or U233 (N_233,N_95,In_171);
nor U234 (N_234,In_206,N_27);
or U235 (N_235,N_86,N_26);
and U236 (N_236,In_37,N_185);
nor U237 (N_237,N_96,In_15);
and U238 (N_238,In_22,N_138);
or U239 (N_239,In_244,N_156);
or U240 (N_240,N_30,N_47);
and U241 (N_241,In_374,N_10);
or U242 (N_242,N_188,N_22);
or U243 (N_243,In_174,In_349);
nor U244 (N_244,N_122,N_64);
xnor U245 (N_245,In_325,N_116);
nand U246 (N_246,N_15,N_191);
or U247 (N_247,N_48,N_55);
xnor U248 (N_248,In_416,N_58);
and U249 (N_249,N_92,N_163);
nor U250 (N_250,N_83,N_194);
nor U251 (N_251,In_115,N_19);
or U252 (N_252,In_336,In_94);
nor U253 (N_253,N_0,N_37);
nor U254 (N_254,N_1,N_113);
or U255 (N_255,N_59,N_24);
or U256 (N_256,In_208,N_62);
nor U257 (N_257,N_154,In_194);
nor U258 (N_258,In_323,N_119);
and U259 (N_259,In_334,In_186);
xor U260 (N_260,N_193,N_111);
nand U261 (N_261,N_88,N_146);
nand U262 (N_262,N_93,N_105);
and U263 (N_263,N_121,N_65);
or U264 (N_264,In_117,N_66);
nor U265 (N_265,N_129,In_57);
nand U266 (N_266,In_109,N_2);
and U267 (N_267,N_41,In_442);
xnor U268 (N_268,N_123,N_49);
or U269 (N_269,In_335,In_404);
or U270 (N_270,N_57,N_94);
nand U271 (N_271,N_161,N_195);
nand U272 (N_272,N_102,N_177);
and U273 (N_273,N_174,N_109);
nand U274 (N_274,N_40,N_90);
xor U275 (N_275,N_9,In_143);
nor U276 (N_276,N_133,N_35);
xnor U277 (N_277,N_103,N_81);
nand U278 (N_278,N_67,In_402);
and U279 (N_279,N_182,In_154);
and U280 (N_280,N_141,In_151);
nor U281 (N_281,In_440,N_8);
nor U282 (N_282,N_149,In_44);
xnor U283 (N_283,N_43,In_324);
or U284 (N_284,N_134,In_198);
xor U285 (N_285,N_140,N_176);
and U286 (N_286,In_205,N_42);
and U287 (N_287,In_163,N_14);
nand U288 (N_288,In_459,N_76);
nor U289 (N_289,N_87,N_190);
and U290 (N_290,N_68,In_138);
nand U291 (N_291,N_31,In_340);
and U292 (N_292,N_148,N_173);
nand U293 (N_293,N_160,N_186);
or U294 (N_294,N_162,N_136);
xor U295 (N_295,N_155,N_74);
and U296 (N_296,N_50,In_309);
and U297 (N_297,N_51,N_151);
nand U298 (N_298,N_79,N_17);
and U299 (N_299,N_166,N_89);
nor U300 (N_300,N_91,N_112);
nand U301 (N_301,N_82,N_71);
nand U302 (N_302,In_364,In_180);
nor U303 (N_303,In_209,N_18);
nor U304 (N_304,N_16,N_34);
nand U305 (N_305,N_125,N_115);
nand U306 (N_306,N_183,N_99);
or U307 (N_307,N_5,In_382);
or U308 (N_308,N_135,In_258);
nor U309 (N_309,In_260,N_189);
and U310 (N_310,N_77,In_405);
xor U311 (N_311,N_169,N_128);
or U312 (N_312,N_171,N_23);
and U313 (N_313,In_319,In_122);
and U314 (N_314,In_127,In_450);
xor U315 (N_315,N_132,In_188);
nand U316 (N_316,N_54,In_173);
or U317 (N_317,In_329,N_61);
nor U318 (N_318,N_198,In_130);
or U319 (N_319,N_45,N_118);
nand U320 (N_320,N_97,N_73);
nor U321 (N_321,N_178,N_137);
or U322 (N_322,In_250,N_13);
or U323 (N_323,N_72,N_167);
nor U324 (N_324,In_373,N_60);
or U325 (N_325,N_172,N_179);
nand U326 (N_326,N_39,In_125);
or U327 (N_327,In_305,N_153);
and U328 (N_328,N_187,In_466);
nand U329 (N_329,In_92,In_56);
and U330 (N_330,In_461,N_181);
or U331 (N_331,In_11,In_232);
xor U332 (N_332,N_144,N_46);
and U333 (N_333,N_175,N_98);
and U334 (N_334,N_199,N_114);
and U335 (N_335,In_100,N_158);
nand U336 (N_336,In_453,N_52);
nor U337 (N_337,In_290,In_235);
and U338 (N_338,N_21,N_63);
and U339 (N_339,In_445,In_50);
or U340 (N_340,N_3,In_294);
nor U341 (N_341,N_38,N_28);
nand U342 (N_342,In_70,In_464);
nor U343 (N_343,N_107,N_170);
nor U344 (N_344,N_78,N_56);
and U345 (N_345,In_78,In_343);
nand U346 (N_346,In_0,In_310);
nand U347 (N_347,In_121,N_168);
xnor U348 (N_348,In_227,N_100);
and U349 (N_349,In_351,N_159);
or U350 (N_350,N_117,N_130);
nand U351 (N_351,N_178,In_56);
and U352 (N_352,N_184,N_7);
and U353 (N_353,N_86,In_143);
nand U354 (N_354,N_152,N_74);
or U355 (N_355,N_73,N_57);
or U356 (N_356,In_340,N_71);
nor U357 (N_357,In_151,N_43);
or U358 (N_358,N_173,N_0);
xnor U359 (N_359,N_87,In_440);
nor U360 (N_360,N_71,N_180);
or U361 (N_361,In_232,N_104);
xnor U362 (N_362,N_133,N_150);
and U363 (N_363,In_109,N_60);
nand U364 (N_364,In_203,N_106);
or U365 (N_365,N_85,N_181);
and U366 (N_366,N_76,In_290);
nor U367 (N_367,N_135,N_32);
or U368 (N_368,N_135,In_416);
nor U369 (N_369,N_46,In_364);
and U370 (N_370,In_450,N_145);
nor U371 (N_371,N_178,N_150);
nor U372 (N_372,N_47,In_290);
and U373 (N_373,N_186,N_83);
and U374 (N_374,N_176,N_187);
nor U375 (N_375,In_329,In_127);
and U376 (N_376,N_142,N_138);
nand U377 (N_377,N_38,N_113);
and U378 (N_378,In_205,In_171);
and U379 (N_379,In_334,In_188);
nand U380 (N_380,N_111,In_309);
or U381 (N_381,In_171,In_11);
xor U382 (N_382,In_15,N_47);
and U383 (N_383,N_156,In_121);
nand U384 (N_384,N_69,N_122);
nor U385 (N_385,N_144,N_88);
nand U386 (N_386,N_8,N_1);
nor U387 (N_387,In_335,N_173);
nand U388 (N_388,N_183,N_146);
nor U389 (N_389,In_232,N_123);
and U390 (N_390,In_209,N_42);
and U391 (N_391,In_94,In_57);
nor U392 (N_392,N_82,N_109);
nand U393 (N_393,In_186,N_180);
nor U394 (N_394,In_232,In_374);
nor U395 (N_395,N_122,N_116);
xor U396 (N_396,N_41,N_43);
nand U397 (N_397,In_15,N_194);
and U398 (N_398,N_165,In_173);
xnor U399 (N_399,In_221,N_128);
xnor U400 (N_400,N_296,N_204);
nor U401 (N_401,N_326,N_248);
and U402 (N_402,N_333,N_295);
and U403 (N_403,N_325,N_267);
and U404 (N_404,N_301,N_351);
or U405 (N_405,N_327,N_268);
xnor U406 (N_406,N_346,N_228);
and U407 (N_407,N_377,N_396);
nand U408 (N_408,N_320,N_354);
or U409 (N_409,N_348,N_332);
or U410 (N_410,N_321,N_276);
or U411 (N_411,N_271,N_318);
xor U412 (N_412,N_331,N_249);
nor U413 (N_413,N_219,N_270);
xor U414 (N_414,N_293,N_283);
xor U415 (N_415,N_306,N_334);
nand U416 (N_416,N_361,N_252);
nor U417 (N_417,N_399,N_227);
or U418 (N_418,N_277,N_207);
xnor U419 (N_419,N_387,N_261);
and U420 (N_420,N_221,N_230);
nor U421 (N_421,N_217,N_202);
or U422 (N_422,N_244,N_257);
nand U423 (N_423,N_305,N_250);
nor U424 (N_424,N_258,N_292);
and U425 (N_425,N_350,N_224);
nand U426 (N_426,N_315,N_393);
or U427 (N_427,N_253,N_307);
nor U428 (N_428,N_269,N_367);
and U429 (N_429,N_245,N_226);
nor U430 (N_430,N_213,N_200);
and U431 (N_431,N_355,N_254);
or U432 (N_432,N_343,N_237);
nand U433 (N_433,N_304,N_233);
or U434 (N_434,N_286,N_349);
xnor U435 (N_435,N_323,N_360);
or U436 (N_436,N_357,N_372);
nor U437 (N_437,N_395,N_239);
or U438 (N_438,N_266,N_235);
and U439 (N_439,N_282,N_225);
nand U440 (N_440,N_251,N_375);
or U441 (N_441,N_340,N_339);
and U442 (N_442,N_329,N_300);
and U443 (N_443,N_297,N_214);
xor U444 (N_444,N_309,N_308);
nand U445 (N_445,N_263,N_338);
and U446 (N_446,N_347,N_311);
and U447 (N_447,N_241,N_264);
nand U448 (N_448,N_246,N_390);
or U449 (N_449,N_287,N_206);
nor U450 (N_450,N_376,N_290);
nor U451 (N_451,N_201,N_280);
xor U452 (N_452,N_319,N_322);
and U453 (N_453,N_256,N_313);
nor U454 (N_454,N_312,N_366);
xnor U455 (N_455,N_341,N_299);
nand U456 (N_456,N_216,N_281);
nor U457 (N_457,N_310,N_223);
nor U458 (N_458,N_385,N_302);
and U459 (N_459,N_337,N_234);
and U460 (N_460,N_262,N_398);
nor U461 (N_461,N_232,N_284);
xnor U462 (N_462,N_345,N_324);
nand U463 (N_463,N_274,N_285);
and U464 (N_464,N_247,N_342);
and U465 (N_465,N_255,N_384);
nor U466 (N_466,N_383,N_211);
xor U467 (N_467,N_364,N_330);
nor U468 (N_468,N_231,N_272);
xor U469 (N_469,N_335,N_397);
nand U470 (N_470,N_381,N_278);
nand U471 (N_471,N_275,N_358);
or U472 (N_472,N_273,N_215);
nand U473 (N_473,N_208,N_218);
xnor U474 (N_474,N_289,N_298);
xor U475 (N_475,N_210,N_369);
or U476 (N_476,N_291,N_389);
or U477 (N_477,N_317,N_279);
or U478 (N_478,N_394,N_222);
nand U479 (N_479,N_382,N_242);
and U480 (N_480,N_379,N_386);
nor U481 (N_481,N_356,N_288);
nand U482 (N_482,N_363,N_388);
or U483 (N_483,N_353,N_365);
xor U484 (N_484,N_236,N_371);
nand U485 (N_485,N_370,N_240);
nand U486 (N_486,N_205,N_391);
or U487 (N_487,N_362,N_294);
and U488 (N_488,N_212,N_209);
or U489 (N_489,N_229,N_314);
and U490 (N_490,N_374,N_373);
nand U491 (N_491,N_316,N_344);
and U492 (N_492,N_352,N_303);
and U493 (N_493,N_368,N_336);
nor U494 (N_494,N_243,N_238);
nand U495 (N_495,N_378,N_359);
nor U496 (N_496,N_260,N_380);
or U497 (N_497,N_259,N_203);
nand U498 (N_498,N_392,N_265);
nor U499 (N_499,N_328,N_220);
or U500 (N_500,N_378,N_230);
nand U501 (N_501,N_392,N_373);
and U502 (N_502,N_291,N_335);
nand U503 (N_503,N_280,N_238);
and U504 (N_504,N_358,N_323);
and U505 (N_505,N_320,N_208);
nor U506 (N_506,N_239,N_342);
and U507 (N_507,N_253,N_385);
and U508 (N_508,N_295,N_275);
or U509 (N_509,N_277,N_340);
nor U510 (N_510,N_286,N_250);
or U511 (N_511,N_347,N_284);
or U512 (N_512,N_308,N_339);
or U513 (N_513,N_277,N_311);
xnor U514 (N_514,N_202,N_271);
and U515 (N_515,N_260,N_217);
nor U516 (N_516,N_357,N_342);
and U517 (N_517,N_255,N_241);
or U518 (N_518,N_268,N_301);
nor U519 (N_519,N_382,N_233);
or U520 (N_520,N_218,N_244);
nand U521 (N_521,N_294,N_219);
nand U522 (N_522,N_322,N_279);
or U523 (N_523,N_389,N_300);
nor U524 (N_524,N_210,N_394);
and U525 (N_525,N_376,N_365);
nor U526 (N_526,N_331,N_298);
xnor U527 (N_527,N_324,N_234);
or U528 (N_528,N_255,N_355);
nor U529 (N_529,N_324,N_292);
xnor U530 (N_530,N_212,N_218);
xnor U531 (N_531,N_331,N_361);
and U532 (N_532,N_251,N_308);
and U533 (N_533,N_305,N_357);
or U534 (N_534,N_385,N_369);
nand U535 (N_535,N_280,N_256);
nand U536 (N_536,N_215,N_396);
or U537 (N_537,N_341,N_257);
xor U538 (N_538,N_327,N_251);
nor U539 (N_539,N_251,N_380);
or U540 (N_540,N_275,N_329);
and U541 (N_541,N_364,N_352);
and U542 (N_542,N_375,N_262);
or U543 (N_543,N_276,N_366);
nor U544 (N_544,N_302,N_281);
nor U545 (N_545,N_200,N_284);
and U546 (N_546,N_235,N_268);
or U547 (N_547,N_277,N_309);
or U548 (N_548,N_359,N_350);
nor U549 (N_549,N_258,N_215);
nand U550 (N_550,N_261,N_279);
xor U551 (N_551,N_289,N_234);
or U552 (N_552,N_393,N_310);
nor U553 (N_553,N_223,N_262);
and U554 (N_554,N_258,N_399);
nand U555 (N_555,N_335,N_370);
nand U556 (N_556,N_289,N_373);
and U557 (N_557,N_281,N_279);
or U558 (N_558,N_283,N_248);
xnor U559 (N_559,N_335,N_376);
nor U560 (N_560,N_282,N_303);
and U561 (N_561,N_361,N_376);
nand U562 (N_562,N_258,N_389);
and U563 (N_563,N_279,N_394);
and U564 (N_564,N_386,N_256);
nand U565 (N_565,N_256,N_289);
or U566 (N_566,N_326,N_263);
nand U567 (N_567,N_223,N_385);
or U568 (N_568,N_337,N_381);
nor U569 (N_569,N_299,N_245);
and U570 (N_570,N_249,N_294);
xor U571 (N_571,N_292,N_280);
or U572 (N_572,N_328,N_306);
and U573 (N_573,N_274,N_215);
nor U574 (N_574,N_270,N_326);
nor U575 (N_575,N_395,N_319);
or U576 (N_576,N_207,N_331);
and U577 (N_577,N_266,N_245);
and U578 (N_578,N_275,N_379);
xor U579 (N_579,N_249,N_364);
and U580 (N_580,N_246,N_311);
or U581 (N_581,N_347,N_384);
nand U582 (N_582,N_356,N_240);
and U583 (N_583,N_242,N_398);
or U584 (N_584,N_227,N_209);
or U585 (N_585,N_357,N_363);
and U586 (N_586,N_372,N_335);
or U587 (N_587,N_328,N_280);
nand U588 (N_588,N_312,N_349);
or U589 (N_589,N_306,N_363);
nor U590 (N_590,N_305,N_274);
and U591 (N_591,N_314,N_294);
and U592 (N_592,N_361,N_234);
nor U593 (N_593,N_360,N_377);
nor U594 (N_594,N_278,N_303);
nand U595 (N_595,N_215,N_271);
nor U596 (N_596,N_392,N_290);
nand U597 (N_597,N_208,N_232);
or U598 (N_598,N_338,N_346);
nor U599 (N_599,N_315,N_246);
and U600 (N_600,N_590,N_598);
and U601 (N_601,N_473,N_531);
and U602 (N_602,N_566,N_567);
or U603 (N_603,N_532,N_546);
and U604 (N_604,N_413,N_434);
xor U605 (N_605,N_487,N_483);
nor U606 (N_606,N_520,N_594);
and U607 (N_607,N_445,N_444);
and U608 (N_608,N_543,N_454);
xor U609 (N_609,N_541,N_429);
nor U610 (N_610,N_408,N_556);
nand U611 (N_611,N_419,N_485);
or U612 (N_612,N_506,N_563);
and U613 (N_613,N_425,N_587);
nor U614 (N_614,N_493,N_466);
or U615 (N_615,N_544,N_458);
nand U616 (N_616,N_499,N_521);
or U617 (N_617,N_443,N_406);
and U618 (N_618,N_470,N_421);
nor U619 (N_619,N_568,N_488);
nand U620 (N_620,N_472,N_562);
and U621 (N_621,N_441,N_513);
nand U622 (N_622,N_599,N_480);
or U623 (N_623,N_518,N_498);
or U624 (N_624,N_420,N_536);
or U625 (N_625,N_423,N_401);
nor U626 (N_626,N_400,N_553);
nor U627 (N_627,N_517,N_565);
or U628 (N_628,N_502,N_433);
nor U629 (N_629,N_555,N_559);
nand U630 (N_630,N_507,N_503);
nor U631 (N_631,N_428,N_404);
and U632 (N_632,N_554,N_579);
nand U633 (N_633,N_582,N_596);
and U634 (N_634,N_560,N_448);
nor U635 (N_635,N_572,N_505);
or U636 (N_636,N_501,N_528);
nor U637 (N_637,N_508,N_535);
and U638 (N_638,N_539,N_500);
nand U639 (N_639,N_405,N_494);
and U640 (N_640,N_452,N_591);
or U641 (N_641,N_504,N_446);
nand U642 (N_642,N_489,N_426);
nand U643 (N_643,N_422,N_550);
or U644 (N_644,N_456,N_542);
xor U645 (N_645,N_496,N_573);
or U646 (N_646,N_585,N_457);
nor U647 (N_647,N_595,N_484);
nor U648 (N_648,N_436,N_529);
or U649 (N_649,N_537,N_577);
or U650 (N_650,N_450,N_525);
nor U651 (N_651,N_491,N_435);
nor U652 (N_652,N_575,N_411);
or U653 (N_653,N_402,N_409);
or U654 (N_654,N_515,N_407);
nand U655 (N_655,N_417,N_453);
xnor U656 (N_656,N_516,N_574);
or U657 (N_657,N_589,N_463);
nand U658 (N_658,N_469,N_476);
xnor U659 (N_659,N_460,N_490);
and U660 (N_660,N_526,N_569);
and U661 (N_661,N_486,N_547);
and U662 (N_662,N_468,N_509);
xnor U663 (N_663,N_530,N_475);
or U664 (N_664,N_449,N_586);
and U665 (N_665,N_471,N_557);
and U666 (N_666,N_512,N_578);
nand U667 (N_667,N_519,N_451);
nand U668 (N_668,N_558,N_534);
nor U669 (N_669,N_495,N_551);
nor U670 (N_670,N_479,N_482);
or U671 (N_671,N_455,N_548);
or U672 (N_672,N_415,N_510);
or U673 (N_673,N_410,N_474);
or U674 (N_674,N_465,N_431);
nand U675 (N_675,N_497,N_561);
or U676 (N_676,N_523,N_564);
or U677 (N_677,N_492,N_583);
or U678 (N_678,N_527,N_437);
or U679 (N_679,N_414,N_467);
xor U680 (N_680,N_412,N_432);
nand U681 (N_681,N_570,N_403);
or U682 (N_682,N_580,N_576);
nand U683 (N_683,N_592,N_427);
or U684 (N_684,N_552,N_424);
and U685 (N_685,N_538,N_522);
nor U686 (N_686,N_540,N_439);
nor U687 (N_687,N_478,N_581);
nor U688 (N_688,N_571,N_593);
nor U689 (N_689,N_511,N_464);
nor U690 (N_690,N_461,N_533);
nand U691 (N_691,N_430,N_549);
or U692 (N_692,N_416,N_584);
nor U693 (N_693,N_588,N_462);
and U694 (N_694,N_477,N_524);
xor U695 (N_695,N_514,N_418);
nor U696 (N_696,N_481,N_438);
xnor U697 (N_697,N_442,N_440);
and U698 (N_698,N_545,N_597);
and U699 (N_699,N_459,N_447);
xor U700 (N_700,N_537,N_430);
nor U701 (N_701,N_504,N_473);
nor U702 (N_702,N_585,N_498);
nor U703 (N_703,N_579,N_526);
or U704 (N_704,N_416,N_517);
nor U705 (N_705,N_429,N_580);
nand U706 (N_706,N_410,N_490);
or U707 (N_707,N_487,N_592);
and U708 (N_708,N_546,N_450);
or U709 (N_709,N_432,N_581);
or U710 (N_710,N_487,N_462);
or U711 (N_711,N_401,N_580);
and U712 (N_712,N_480,N_508);
nand U713 (N_713,N_448,N_504);
and U714 (N_714,N_534,N_400);
or U715 (N_715,N_527,N_451);
nand U716 (N_716,N_567,N_550);
nor U717 (N_717,N_538,N_419);
and U718 (N_718,N_563,N_458);
and U719 (N_719,N_418,N_572);
or U720 (N_720,N_561,N_513);
nor U721 (N_721,N_542,N_403);
xnor U722 (N_722,N_432,N_562);
nand U723 (N_723,N_460,N_484);
nor U724 (N_724,N_557,N_422);
and U725 (N_725,N_436,N_431);
and U726 (N_726,N_430,N_412);
and U727 (N_727,N_524,N_402);
and U728 (N_728,N_511,N_478);
nor U729 (N_729,N_507,N_473);
nor U730 (N_730,N_407,N_473);
or U731 (N_731,N_463,N_578);
nand U732 (N_732,N_555,N_535);
nor U733 (N_733,N_526,N_538);
or U734 (N_734,N_406,N_515);
nand U735 (N_735,N_570,N_482);
nand U736 (N_736,N_495,N_418);
or U737 (N_737,N_587,N_480);
nor U738 (N_738,N_597,N_528);
or U739 (N_739,N_552,N_504);
nor U740 (N_740,N_544,N_548);
nor U741 (N_741,N_588,N_567);
nor U742 (N_742,N_450,N_550);
nor U743 (N_743,N_492,N_509);
and U744 (N_744,N_533,N_555);
nor U745 (N_745,N_573,N_448);
or U746 (N_746,N_434,N_452);
nand U747 (N_747,N_541,N_554);
or U748 (N_748,N_477,N_537);
nor U749 (N_749,N_513,N_449);
or U750 (N_750,N_412,N_437);
and U751 (N_751,N_443,N_565);
nor U752 (N_752,N_512,N_594);
nor U753 (N_753,N_519,N_521);
or U754 (N_754,N_554,N_414);
or U755 (N_755,N_559,N_542);
nor U756 (N_756,N_503,N_475);
or U757 (N_757,N_536,N_566);
nand U758 (N_758,N_454,N_516);
xor U759 (N_759,N_506,N_405);
xor U760 (N_760,N_532,N_407);
nand U761 (N_761,N_580,N_574);
nand U762 (N_762,N_556,N_426);
and U763 (N_763,N_571,N_505);
and U764 (N_764,N_537,N_525);
nor U765 (N_765,N_562,N_496);
and U766 (N_766,N_546,N_504);
nand U767 (N_767,N_566,N_418);
nor U768 (N_768,N_568,N_513);
and U769 (N_769,N_510,N_490);
nor U770 (N_770,N_426,N_471);
or U771 (N_771,N_514,N_462);
nand U772 (N_772,N_557,N_496);
and U773 (N_773,N_592,N_448);
and U774 (N_774,N_431,N_502);
or U775 (N_775,N_432,N_592);
nor U776 (N_776,N_453,N_569);
nor U777 (N_777,N_565,N_550);
nor U778 (N_778,N_480,N_472);
xnor U779 (N_779,N_424,N_463);
or U780 (N_780,N_556,N_480);
nor U781 (N_781,N_457,N_487);
xnor U782 (N_782,N_455,N_462);
nand U783 (N_783,N_402,N_445);
and U784 (N_784,N_497,N_565);
xor U785 (N_785,N_597,N_425);
nor U786 (N_786,N_590,N_410);
xor U787 (N_787,N_412,N_444);
and U788 (N_788,N_413,N_579);
nor U789 (N_789,N_566,N_564);
and U790 (N_790,N_593,N_440);
and U791 (N_791,N_551,N_594);
or U792 (N_792,N_561,N_591);
nor U793 (N_793,N_523,N_596);
nand U794 (N_794,N_468,N_592);
and U795 (N_795,N_429,N_495);
nor U796 (N_796,N_593,N_434);
and U797 (N_797,N_595,N_416);
and U798 (N_798,N_420,N_558);
and U799 (N_799,N_524,N_466);
or U800 (N_800,N_753,N_729);
and U801 (N_801,N_600,N_654);
nand U802 (N_802,N_641,N_738);
and U803 (N_803,N_665,N_702);
nor U804 (N_804,N_652,N_675);
nor U805 (N_805,N_679,N_698);
nor U806 (N_806,N_662,N_636);
nand U807 (N_807,N_669,N_666);
xor U808 (N_808,N_667,N_746);
or U809 (N_809,N_605,N_703);
and U810 (N_810,N_619,N_755);
and U811 (N_811,N_677,N_762);
nor U812 (N_812,N_766,N_763);
or U813 (N_813,N_716,N_715);
and U814 (N_814,N_752,N_771);
nor U815 (N_815,N_642,N_777);
nand U816 (N_816,N_646,N_783);
and U817 (N_817,N_709,N_603);
nand U818 (N_818,N_734,N_781);
and U819 (N_819,N_782,N_727);
nand U820 (N_820,N_658,N_606);
nand U821 (N_821,N_712,N_701);
or U822 (N_822,N_651,N_699);
nand U823 (N_823,N_747,N_649);
and U824 (N_824,N_770,N_614);
nor U825 (N_825,N_750,N_639);
and U826 (N_826,N_791,N_625);
xnor U827 (N_827,N_706,N_618);
or U828 (N_828,N_722,N_756);
nand U829 (N_829,N_720,N_668);
nor U830 (N_830,N_688,N_789);
nand U831 (N_831,N_692,N_772);
nor U832 (N_832,N_723,N_615);
nor U833 (N_833,N_725,N_761);
nand U834 (N_834,N_681,N_683);
nand U835 (N_835,N_684,N_645);
xor U836 (N_836,N_638,N_784);
nor U837 (N_837,N_704,N_690);
xor U838 (N_838,N_656,N_631);
nor U839 (N_839,N_735,N_686);
xnor U840 (N_840,N_775,N_713);
and U841 (N_841,N_621,N_643);
and U842 (N_842,N_624,N_663);
or U843 (N_843,N_793,N_653);
or U844 (N_844,N_764,N_790);
nor U845 (N_845,N_673,N_691);
nand U846 (N_846,N_736,N_648);
nand U847 (N_847,N_717,N_796);
nor U848 (N_848,N_628,N_697);
nand U849 (N_849,N_602,N_767);
nand U850 (N_850,N_728,N_757);
and U851 (N_851,N_607,N_644);
or U852 (N_852,N_694,N_730);
nand U853 (N_853,N_732,N_740);
nand U854 (N_854,N_604,N_630);
and U855 (N_855,N_795,N_632);
nand U856 (N_856,N_612,N_733);
and U857 (N_857,N_637,N_758);
or U858 (N_858,N_797,N_659);
nor U859 (N_859,N_609,N_759);
nand U860 (N_860,N_792,N_798);
nor U861 (N_861,N_743,N_687);
nor U862 (N_862,N_776,N_640);
nor U863 (N_863,N_633,N_705);
and U864 (N_864,N_724,N_622);
nor U865 (N_865,N_616,N_708);
nor U866 (N_866,N_696,N_635);
or U867 (N_867,N_657,N_678);
or U868 (N_868,N_749,N_664);
and U869 (N_869,N_794,N_744);
nand U870 (N_870,N_780,N_661);
and U871 (N_871,N_751,N_670);
nor U872 (N_872,N_672,N_676);
nand U873 (N_873,N_647,N_745);
nor U874 (N_874,N_680,N_634);
xor U875 (N_875,N_693,N_748);
nand U876 (N_876,N_769,N_765);
or U877 (N_877,N_710,N_601);
nand U878 (N_878,N_718,N_695);
or U879 (N_879,N_650,N_627);
and U880 (N_880,N_685,N_760);
nor U881 (N_881,N_788,N_617);
nor U882 (N_882,N_700,N_608);
and U883 (N_883,N_741,N_786);
and U884 (N_884,N_689,N_768);
nor U885 (N_885,N_799,N_671);
nand U886 (N_886,N_739,N_623);
nor U887 (N_887,N_629,N_613);
or U888 (N_888,N_787,N_655);
nand U889 (N_889,N_674,N_778);
or U890 (N_890,N_754,N_611);
nand U891 (N_891,N_626,N_731);
and U892 (N_892,N_714,N_620);
or U893 (N_893,N_742,N_737);
or U894 (N_894,N_721,N_660);
nor U895 (N_895,N_707,N_774);
nand U896 (N_896,N_726,N_773);
and U897 (N_897,N_719,N_785);
nand U898 (N_898,N_610,N_682);
and U899 (N_899,N_779,N_711);
nand U900 (N_900,N_795,N_651);
nor U901 (N_901,N_618,N_665);
nor U902 (N_902,N_668,N_777);
nand U903 (N_903,N_673,N_642);
nand U904 (N_904,N_769,N_764);
nand U905 (N_905,N_785,N_761);
nand U906 (N_906,N_612,N_730);
nand U907 (N_907,N_631,N_782);
or U908 (N_908,N_659,N_740);
nand U909 (N_909,N_664,N_716);
nand U910 (N_910,N_785,N_769);
nand U911 (N_911,N_657,N_619);
nor U912 (N_912,N_638,N_769);
and U913 (N_913,N_665,N_781);
and U914 (N_914,N_692,N_754);
and U915 (N_915,N_684,N_652);
nor U916 (N_916,N_657,N_721);
nor U917 (N_917,N_721,N_600);
xor U918 (N_918,N_618,N_649);
nor U919 (N_919,N_607,N_616);
xor U920 (N_920,N_790,N_689);
and U921 (N_921,N_690,N_664);
or U922 (N_922,N_716,N_604);
nand U923 (N_923,N_654,N_787);
and U924 (N_924,N_742,N_653);
xor U925 (N_925,N_713,N_718);
xor U926 (N_926,N_603,N_609);
or U927 (N_927,N_676,N_651);
nand U928 (N_928,N_713,N_672);
and U929 (N_929,N_648,N_691);
and U930 (N_930,N_682,N_781);
or U931 (N_931,N_713,N_681);
or U932 (N_932,N_695,N_760);
and U933 (N_933,N_667,N_682);
and U934 (N_934,N_700,N_793);
nor U935 (N_935,N_674,N_763);
nand U936 (N_936,N_652,N_747);
and U937 (N_937,N_689,N_770);
or U938 (N_938,N_666,N_643);
or U939 (N_939,N_653,N_693);
and U940 (N_940,N_773,N_671);
and U941 (N_941,N_728,N_702);
or U942 (N_942,N_716,N_643);
nand U943 (N_943,N_622,N_781);
xor U944 (N_944,N_687,N_784);
nand U945 (N_945,N_662,N_698);
and U946 (N_946,N_783,N_636);
xor U947 (N_947,N_777,N_709);
or U948 (N_948,N_643,N_698);
and U949 (N_949,N_750,N_752);
nand U950 (N_950,N_643,N_623);
nor U951 (N_951,N_769,N_697);
and U952 (N_952,N_615,N_746);
nor U953 (N_953,N_785,N_657);
nor U954 (N_954,N_647,N_609);
or U955 (N_955,N_669,N_743);
or U956 (N_956,N_730,N_681);
nand U957 (N_957,N_612,N_703);
and U958 (N_958,N_654,N_709);
xor U959 (N_959,N_671,N_623);
and U960 (N_960,N_684,N_732);
nand U961 (N_961,N_691,N_634);
nand U962 (N_962,N_609,N_699);
and U963 (N_963,N_712,N_704);
nor U964 (N_964,N_762,N_687);
or U965 (N_965,N_730,N_699);
and U966 (N_966,N_690,N_717);
nor U967 (N_967,N_637,N_613);
nor U968 (N_968,N_650,N_632);
and U969 (N_969,N_605,N_718);
or U970 (N_970,N_749,N_746);
and U971 (N_971,N_647,N_744);
and U972 (N_972,N_616,N_733);
or U973 (N_973,N_764,N_732);
nand U974 (N_974,N_757,N_717);
and U975 (N_975,N_633,N_629);
xnor U976 (N_976,N_703,N_760);
nand U977 (N_977,N_751,N_657);
nand U978 (N_978,N_609,N_629);
and U979 (N_979,N_655,N_641);
or U980 (N_980,N_755,N_719);
nand U981 (N_981,N_649,N_619);
nor U982 (N_982,N_615,N_796);
nor U983 (N_983,N_779,N_767);
and U984 (N_984,N_624,N_620);
nor U985 (N_985,N_691,N_665);
nand U986 (N_986,N_665,N_782);
or U987 (N_987,N_684,N_751);
nor U988 (N_988,N_674,N_768);
and U989 (N_989,N_794,N_754);
or U990 (N_990,N_721,N_674);
and U991 (N_991,N_632,N_692);
or U992 (N_992,N_745,N_735);
or U993 (N_993,N_778,N_721);
and U994 (N_994,N_722,N_689);
nand U995 (N_995,N_788,N_663);
nor U996 (N_996,N_787,N_732);
or U997 (N_997,N_647,N_725);
and U998 (N_998,N_725,N_707);
nand U999 (N_999,N_770,N_619);
and U1000 (N_1000,N_837,N_957);
or U1001 (N_1001,N_836,N_946);
and U1002 (N_1002,N_930,N_903);
or U1003 (N_1003,N_962,N_810);
nand U1004 (N_1004,N_952,N_990);
and U1005 (N_1005,N_823,N_864);
and U1006 (N_1006,N_993,N_937);
or U1007 (N_1007,N_901,N_983);
nand U1008 (N_1008,N_817,N_908);
nand U1009 (N_1009,N_964,N_967);
xnor U1010 (N_1010,N_831,N_882);
nor U1011 (N_1011,N_911,N_899);
nand U1012 (N_1012,N_948,N_917);
or U1013 (N_1013,N_924,N_879);
nand U1014 (N_1014,N_803,N_805);
nand U1015 (N_1015,N_960,N_986);
or U1016 (N_1016,N_942,N_921);
nor U1017 (N_1017,N_828,N_873);
or U1018 (N_1018,N_996,N_900);
nand U1019 (N_1019,N_929,N_884);
xnor U1020 (N_1020,N_825,N_926);
nand U1021 (N_1021,N_856,N_992);
nor U1022 (N_1022,N_984,N_991);
or U1023 (N_1023,N_916,N_886);
nand U1024 (N_1024,N_940,N_982);
nand U1025 (N_1025,N_976,N_889);
nor U1026 (N_1026,N_941,N_872);
nand U1027 (N_1027,N_947,N_968);
xnor U1028 (N_1028,N_913,N_865);
nand U1029 (N_1029,N_909,N_860);
and U1030 (N_1030,N_905,N_923);
nand U1031 (N_1031,N_954,N_800);
xnor U1032 (N_1032,N_859,N_877);
nand U1033 (N_1033,N_822,N_896);
nand U1034 (N_1034,N_863,N_919);
and U1035 (N_1035,N_980,N_829);
and U1036 (N_1036,N_955,N_802);
nor U1037 (N_1037,N_981,N_806);
nand U1038 (N_1038,N_875,N_857);
and U1039 (N_1039,N_910,N_809);
and U1040 (N_1040,N_876,N_804);
and U1041 (N_1041,N_943,N_840);
nand U1042 (N_1042,N_850,N_973);
or U1043 (N_1043,N_848,N_961);
nand U1044 (N_1044,N_931,N_861);
xnor U1045 (N_1045,N_914,N_934);
xor U1046 (N_1046,N_912,N_813);
nor U1047 (N_1047,N_963,N_883);
nand U1048 (N_1048,N_834,N_922);
or U1049 (N_1049,N_958,N_826);
and U1050 (N_1050,N_999,N_808);
or U1051 (N_1051,N_972,N_956);
nor U1052 (N_1052,N_936,N_892);
or U1053 (N_1053,N_844,N_807);
nand U1054 (N_1054,N_869,N_938);
or U1055 (N_1055,N_979,N_812);
nor U1056 (N_1056,N_835,N_858);
nor U1057 (N_1057,N_855,N_814);
xnor U1058 (N_1058,N_945,N_902);
nand U1059 (N_1059,N_890,N_851);
xnor U1060 (N_1060,N_888,N_853);
nand U1061 (N_1061,N_951,N_885);
nand U1062 (N_1062,N_880,N_918);
nand U1063 (N_1063,N_927,N_995);
or U1064 (N_1064,N_849,N_878);
or U1065 (N_1065,N_868,N_985);
and U1066 (N_1066,N_891,N_895);
nor U1067 (N_1067,N_998,N_841);
nand U1068 (N_1068,N_871,N_907);
nor U1069 (N_1069,N_994,N_987);
nor U1070 (N_1070,N_854,N_839);
or U1071 (N_1071,N_824,N_953);
nand U1072 (N_1072,N_977,N_874);
nand U1073 (N_1073,N_820,N_971);
nand U1074 (N_1074,N_939,N_898);
nand U1075 (N_1075,N_978,N_897);
and U1076 (N_1076,N_969,N_950);
and U1077 (N_1077,N_887,N_842);
and U1078 (N_1078,N_833,N_997);
and U1079 (N_1079,N_838,N_989);
nand U1080 (N_1080,N_846,N_915);
or U1081 (N_1081,N_965,N_816);
or U1082 (N_1082,N_845,N_866);
nor U1083 (N_1083,N_815,N_811);
nand U1084 (N_1084,N_906,N_830);
nor U1085 (N_1085,N_975,N_949);
and U1086 (N_1086,N_894,N_852);
and U1087 (N_1087,N_818,N_867);
or U1088 (N_1088,N_801,N_843);
and U1089 (N_1089,N_827,N_819);
nand U1090 (N_1090,N_933,N_821);
nor U1091 (N_1091,N_870,N_904);
xnor U1092 (N_1092,N_928,N_944);
or U1093 (N_1093,N_932,N_966);
and U1094 (N_1094,N_925,N_881);
nand U1095 (N_1095,N_935,N_847);
or U1096 (N_1096,N_974,N_959);
and U1097 (N_1097,N_862,N_988);
and U1098 (N_1098,N_970,N_893);
and U1099 (N_1099,N_832,N_920);
or U1100 (N_1100,N_848,N_882);
nand U1101 (N_1101,N_908,N_993);
or U1102 (N_1102,N_936,N_820);
xor U1103 (N_1103,N_930,N_869);
nand U1104 (N_1104,N_834,N_921);
or U1105 (N_1105,N_884,N_904);
nand U1106 (N_1106,N_961,N_941);
nand U1107 (N_1107,N_956,N_950);
or U1108 (N_1108,N_810,N_816);
nand U1109 (N_1109,N_988,N_866);
or U1110 (N_1110,N_909,N_951);
or U1111 (N_1111,N_970,N_856);
or U1112 (N_1112,N_858,N_863);
and U1113 (N_1113,N_834,N_952);
nor U1114 (N_1114,N_994,N_984);
and U1115 (N_1115,N_954,N_904);
or U1116 (N_1116,N_977,N_958);
xor U1117 (N_1117,N_884,N_936);
nand U1118 (N_1118,N_872,N_980);
and U1119 (N_1119,N_957,N_862);
xor U1120 (N_1120,N_961,N_810);
or U1121 (N_1121,N_896,N_976);
and U1122 (N_1122,N_955,N_927);
xnor U1123 (N_1123,N_968,N_932);
or U1124 (N_1124,N_989,N_999);
xnor U1125 (N_1125,N_937,N_923);
or U1126 (N_1126,N_955,N_858);
nand U1127 (N_1127,N_854,N_943);
and U1128 (N_1128,N_863,N_949);
nor U1129 (N_1129,N_928,N_843);
nand U1130 (N_1130,N_953,N_935);
nor U1131 (N_1131,N_833,N_808);
nor U1132 (N_1132,N_883,N_937);
xnor U1133 (N_1133,N_896,N_901);
or U1134 (N_1134,N_808,N_802);
or U1135 (N_1135,N_954,N_920);
or U1136 (N_1136,N_881,N_852);
and U1137 (N_1137,N_846,N_813);
or U1138 (N_1138,N_905,N_865);
nand U1139 (N_1139,N_941,N_915);
and U1140 (N_1140,N_809,N_998);
nand U1141 (N_1141,N_868,N_953);
and U1142 (N_1142,N_835,N_822);
nand U1143 (N_1143,N_902,N_837);
nor U1144 (N_1144,N_920,N_899);
nand U1145 (N_1145,N_888,N_809);
or U1146 (N_1146,N_921,N_803);
nand U1147 (N_1147,N_840,N_869);
nor U1148 (N_1148,N_829,N_985);
or U1149 (N_1149,N_966,N_892);
and U1150 (N_1150,N_986,N_901);
nor U1151 (N_1151,N_840,N_882);
nand U1152 (N_1152,N_914,N_932);
or U1153 (N_1153,N_975,N_952);
nor U1154 (N_1154,N_836,N_835);
nor U1155 (N_1155,N_950,N_892);
nand U1156 (N_1156,N_812,N_900);
xor U1157 (N_1157,N_980,N_918);
xnor U1158 (N_1158,N_804,N_979);
or U1159 (N_1159,N_913,N_924);
nor U1160 (N_1160,N_825,N_929);
and U1161 (N_1161,N_855,N_991);
and U1162 (N_1162,N_947,N_840);
xnor U1163 (N_1163,N_893,N_855);
nand U1164 (N_1164,N_966,N_858);
and U1165 (N_1165,N_801,N_895);
nor U1166 (N_1166,N_805,N_838);
and U1167 (N_1167,N_882,N_917);
nand U1168 (N_1168,N_989,N_955);
nor U1169 (N_1169,N_897,N_957);
nor U1170 (N_1170,N_943,N_949);
nand U1171 (N_1171,N_939,N_833);
nand U1172 (N_1172,N_821,N_978);
xor U1173 (N_1173,N_810,N_951);
or U1174 (N_1174,N_976,N_834);
nand U1175 (N_1175,N_865,N_896);
xor U1176 (N_1176,N_992,N_819);
and U1177 (N_1177,N_944,N_882);
nand U1178 (N_1178,N_970,N_968);
nand U1179 (N_1179,N_859,N_983);
nor U1180 (N_1180,N_886,N_843);
xnor U1181 (N_1181,N_960,N_802);
nor U1182 (N_1182,N_841,N_874);
and U1183 (N_1183,N_879,N_931);
nor U1184 (N_1184,N_999,N_982);
nor U1185 (N_1185,N_800,N_992);
or U1186 (N_1186,N_849,N_934);
nor U1187 (N_1187,N_896,N_828);
and U1188 (N_1188,N_941,N_864);
nand U1189 (N_1189,N_997,N_976);
and U1190 (N_1190,N_997,N_887);
or U1191 (N_1191,N_976,N_965);
nand U1192 (N_1192,N_927,N_836);
or U1193 (N_1193,N_835,N_916);
nor U1194 (N_1194,N_951,N_958);
or U1195 (N_1195,N_824,N_882);
and U1196 (N_1196,N_803,N_947);
and U1197 (N_1197,N_803,N_834);
nor U1198 (N_1198,N_949,N_986);
nand U1199 (N_1199,N_966,N_815);
nor U1200 (N_1200,N_1145,N_1000);
or U1201 (N_1201,N_1012,N_1055);
xor U1202 (N_1202,N_1184,N_1177);
and U1203 (N_1203,N_1005,N_1147);
and U1204 (N_1204,N_1071,N_1130);
nor U1205 (N_1205,N_1070,N_1060);
or U1206 (N_1206,N_1132,N_1142);
nand U1207 (N_1207,N_1093,N_1042);
and U1208 (N_1208,N_1191,N_1043);
or U1209 (N_1209,N_1056,N_1054);
xnor U1210 (N_1210,N_1032,N_1098);
or U1211 (N_1211,N_1090,N_1065);
nor U1212 (N_1212,N_1140,N_1009);
and U1213 (N_1213,N_1161,N_1024);
xor U1214 (N_1214,N_1044,N_1175);
nor U1215 (N_1215,N_1006,N_1180);
nor U1216 (N_1216,N_1114,N_1007);
nor U1217 (N_1217,N_1035,N_1016);
xnor U1218 (N_1218,N_1089,N_1051);
nand U1219 (N_1219,N_1010,N_1077);
or U1220 (N_1220,N_1001,N_1127);
xnor U1221 (N_1221,N_1170,N_1030);
or U1222 (N_1222,N_1112,N_1198);
nor U1223 (N_1223,N_1072,N_1081);
nand U1224 (N_1224,N_1146,N_1154);
nor U1225 (N_1225,N_1156,N_1064);
and U1226 (N_1226,N_1078,N_1125);
xor U1227 (N_1227,N_1040,N_1068);
nand U1228 (N_1228,N_1015,N_1188);
and U1229 (N_1229,N_1088,N_1189);
and U1230 (N_1230,N_1166,N_1013);
or U1231 (N_1231,N_1002,N_1186);
nand U1232 (N_1232,N_1105,N_1158);
nand U1233 (N_1233,N_1058,N_1197);
nor U1234 (N_1234,N_1144,N_1107);
and U1235 (N_1235,N_1086,N_1092);
or U1236 (N_1236,N_1022,N_1136);
nand U1237 (N_1237,N_1118,N_1168);
xor U1238 (N_1238,N_1134,N_1187);
nand U1239 (N_1239,N_1033,N_1052);
and U1240 (N_1240,N_1159,N_1023);
xor U1241 (N_1241,N_1131,N_1063);
xor U1242 (N_1242,N_1047,N_1182);
and U1243 (N_1243,N_1190,N_1128);
nor U1244 (N_1244,N_1113,N_1094);
or U1245 (N_1245,N_1126,N_1179);
nor U1246 (N_1246,N_1139,N_1157);
nor U1247 (N_1247,N_1116,N_1103);
nor U1248 (N_1248,N_1048,N_1020);
or U1249 (N_1249,N_1162,N_1014);
and U1250 (N_1250,N_1028,N_1057);
and U1251 (N_1251,N_1026,N_1102);
nor U1252 (N_1252,N_1029,N_1031);
or U1253 (N_1253,N_1066,N_1120);
and U1254 (N_1254,N_1017,N_1101);
and U1255 (N_1255,N_1111,N_1165);
nor U1256 (N_1256,N_1059,N_1195);
and U1257 (N_1257,N_1019,N_1176);
nand U1258 (N_1258,N_1034,N_1172);
nor U1259 (N_1259,N_1192,N_1108);
or U1260 (N_1260,N_1149,N_1080);
and U1261 (N_1261,N_1074,N_1138);
and U1262 (N_1262,N_1129,N_1153);
nor U1263 (N_1263,N_1003,N_1046);
nand U1264 (N_1264,N_1109,N_1119);
and U1265 (N_1265,N_1163,N_1038);
nor U1266 (N_1266,N_1152,N_1025);
nand U1267 (N_1267,N_1141,N_1036);
nor U1268 (N_1268,N_1084,N_1027);
or U1269 (N_1269,N_1150,N_1050);
and U1270 (N_1270,N_1075,N_1039);
nor U1271 (N_1271,N_1167,N_1091);
and U1272 (N_1272,N_1011,N_1037);
nand U1273 (N_1273,N_1135,N_1067);
nand U1274 (N_1274,N_1160,N_1124);
xnor U1275 (N_1275,N_1004,N_1123);
or U1276 (N_1276,N_1121,N_1174);
and U1277 (N_1277,N_1008,N_1169);
nand U1278 (N_1278,N_1143,N_1181);
nor U1279 (N_1279,N_1095,N_1122);
nor U1280 (N_1280,N_1097,N_1106);
or U1281 (N_1281,N_1076,N_1041);
nor U1282 (N_1282,N_1148,N_1117);
and U1283 (N_1283,N_1069,N_1178);
or U1284 (N_1284,N_1099,N_1082);
and U1285 (N_1285,N_1045,N_1083);
and U1286 (N_1286,N_1073,N_1087);
or U1287 (N_1287,N_1110,N_1185);
nor U1288 (N_1288,N_1171,N_1053);
nor U1289 (N_1289,N_1183,N_1115);
nand U1290 (N_1290,N_1062,N_1155);
nor U1291 (N_1291,N_1194,N_1085);
nand U1292 (N_1292,N_1173,N_1196);
nand U1293 (N_1293,N_1021,N_1079);
nand U1294 (N_1294,N_1193,N_1096);
or U1295 (N_1295,N_1061,N_1049);
and U1296 (N_1296,N_1104,N_1199);
and U1297 (N_1297,N_1151,N_1100);
and U1298 (N_1298,N_1133,N_1018);
nand U1299 (N_1299,N_1137,N_1164);
nor U1300 (N_1300,N_1014,N_1118);
and U1301 (N_1301,N_1017,N_1150);
nor U1302 (N_1302,N_1039,N_1038);
and U1303 (N_1303,N_1199,N_1057);
nor U1304 (N_1304,N_1085,N_1053);
nor U1305 (N_1305,N_1196,N_1145);
and U1306 (N_1306,N_1051,N_1111);
or U1307 (N_1307,N_1195,N_1092);
and U1308 (N_1308,N_1030,N_1052);
and U1309 (N_1309,N_1071,N_1024);
or U1310 (N_1310,N_1095,N_1097);
nor U1311 (N_1311,N_1090,N_1186);
nand U1312 (N_1312,N_1187,N_1036);
nor U1313 (N_1313,N_1181,N_1008);
and U1314 (N_1314,N_1036,N_1035);
and U1315 (N_1315,N_1063,N_1087);
or U1316 (N_1316,N_1094,N_1035);
and U1317 (N_1317,N_1162,N_1081);
nor U1318 (N_1318,N_1174,N_1099);
xor U1319 (N_1319,N_1061,N_1189);
nor U1320 (N_1320,N_1093,N_1145);
nand U1321 (N_1321,N_1158,N_1037);
nand U1322 (N_1322,N_1057,N_1065);
nor U1323 (N_1323,N_1068,N_1192);
and U1324 (N_1324,N_1036,N_1140);
and U1325 (N_1325,N_1150,N_1076);
nand U1326 (N_1326,N_1182,N_1134);
and U1327 (N_1327,N_1062,N_1139);
and U1328 (N_1328,N_1181,N_1196);
nor U1329 (N_1329,N_1024,N_1195);
nor U1330 (N_1330,N_1184,N_1045);
nor U1331 (N_1331,N_1021,N_1139);
nor U1332 (N_1332,N_1173,N_1037);
xnor U1333 (N_1333,N_1012,N_1107);
or U1334 (N_1334,N_1115,N_1056);
nand U1335 (N_1335,N_1070,N_1160);
or U1336 (N_1336,N_1044,N_1139);
nand U1337 (N_1337,N_1126,N_1069);
or U1338 (N_1338,N_1114,N_1149);
and U1339 (N_1339,N_1105,N_1151);
nor U1340 (N_1340,N_1153,N_1127);
or U1341 (N_1341,N_1162,N_1019);
xnor U1342 (N_1342,N_1067,N_1045);
or U1343 (N_1343,N_1008,N_1129);
nor U1344 (N_1344,N_1112,N_1177);
nand U1345 (N_1345,N_1050,N_1022);
or U1346 (N_1346,N_1051,N_1086);
and U1347 (N_1347,N_1005,N_1143);
nand U1348 (N_1348,N_1057,N_1038);
nor U1349 (N_1349,N_1112,N_1099);
and U1350 (N_1350,N_1157,N_1003);
nor U1351 (N_1351,N_1137,N_1040);
or U1352 (N_1352,N_1065,N_1039);
nor U1353 (N_1353,N_1003,N_1074);
or U1354 (N_1354,N_1055,N_1169);
and U1355 (N_1355,N_1067,N_1109);
or U1356 (N_1356,N_1056,N_1001);
xnor U1357 (N_1357,N_1039,N_1052);
nor U1358 (N_1358,N_1129,N_1027);
xnor U1359 (N_1359,N_1085,N_1143);
nand U1360 (N_1360,N_1172,N_1058);
xor U1361 (N_1361,N_1024,N_1079);
xnor U1362 (N_1362,N_1143,N_1100);
nor U1363 (N_1363,N_1049,N_1193);
xor U1364 (N_1364,N_1101,N_1124);
and U1365 (N_1365,N_1161,N_1064);
and U1366 (N_1366,N_1191,N_1146);
and U1367 (N_1367,N_1148,N_1154);
nand U1368 (N_1368,N_1188,N_1057);
and U1369 (N_1369,N_1137,N_1067);
nor U1370 (N_1370,N_1121,N_1060);
and U1371 (N_1371,N_1192,N_1140);
and U1372 (N_1372,N_1021,N_1054);
or U1373 (N_1373,N_1063,N_1194);
or U1374 (N_1374,N_1053,N_1126);
and U1375 (N_1375,N_1199,N_1125);
or U1376 (N_1376,N_1167,N_1126);
nor U1377 (N_1377,N_1125,N_1080);
and U1378 (N_1378,N_1076,N_1138);
nand U1379 (N_1379,N_1028,N_1102);
nor U1380 (N_1380,N_1187,N_1054);
and U1381 (N_1381,N_1153,N_1198);
nor U1382 (N_1382,N_1155,N_1046);
or U1383 (N_1383,N_1152,N_1077);
or U1384 (N_1384,N_1144,N_1114);
nand U1385 (N_1385,N_1097,N_1137);
and U1386 (N_1386,N_1177,N_1183);
and U1387 (N_1387,N_1175,N_1164);
nand U1388 (N_1388,N_1064,N_1054);
or U1389 (N_1389,N_1194,N_1180);
xor U1390 (N_1390,N_1081,N_1157);
nand U1391 (N_1391,N_1044,N_1097);
nor U1392 (N_1392,N_1185,N_1028);
nor U1393 (N_1393,N_1135,N_1102);
or U1394 (N_1394,N_1038,N_1143);
and U1395 (N_1395,N_1088,N_1151);
xnor U1396 (N_1396,N_1069,N_1190);
and U1397 (N_1397,N_1105,N_1040);
and U1398 (N_1398,N_1034,N_1096);
and U1399 (N_1399,N_1059,N_1028);
nand U1400 (N_1400,N_1268,N_1252);
nand U1401 (N_1401,N_1250,N_1240);
xnor U1402 (N_1402,N_1342,N_1289);
nand U1403 (N_1403,N_1355,N_1200);
xor U1404 (N_1404,N_1388,N_1339);
and U1405 (N_1405,N_1318,N_1354);
or U1406 (N_1406,N_1255,N_1203);
nor U1407 (N_1407,N_1310,N_1211);
nor U1408 (N_1408,N_1273,N_1338);
nor U1409 (N_1409,N_1283,N_1396);
or U1410 (N_1410,N_1311,N_1257);
nand U1411 (N_1411,N_1208,N_1306);
or U1412 (N_1412,N_1393,N_1253);
nand U1413 (N_1413,N_1372,N_1321);
or U1414 (N_1414,N_1374,N_1242);
nand U1415 (N_1415,N_1266,N_1366);
or U1416 (N_1416,N_1316,N_1299);
or U1417 (N_1417,N_1336,N_1233);
nor U1418 (N_1418,N_1226,N_1352);
nor U1419 (N_1419,N_1219,N_1216);
nor U1420 (N_1420,N_1385,N_1389);
and U1421 (N_1421,N_1308,N_1262);
and U1422 (N_1422,N_1313,N_1247);
and U1423 (N_1423,N_1204,N_1300);
or U1424 (N_1424,N_1319,N_1391);
and U1425 (N_1425,N_1357,N_1291);
or U1426 (N_1426,N_1274,N_1373);
nor U1427 (N_1427,N_1224,N_1229);
nor U1428 (N_1428,N_1230,N_1205);
or U1429 (N_1429,N_1383,N_1235);
or U1430 (N_1430,N_1303,N_1239);
nor U1431 (N_1431,N_1202,N_1363);
or U1432 (N_1432,N_1260,N_1387);
and U1433 (N_1433,N_1277,N_1217);
nand U1434 (N_1434,N_1328,N_1290);
nor U1435 (N_1435,N_1375,N_1390);
or U1436 (N_1436,N_1309,N_1256);
nor U1437 (N_1437,N_1296,N_1399);
xnor U1438 (N_1438,N_1265,N_1331);
nor U1439 (N_1439,N_1218,N_1294);
or U1440 (N_1440,N_1379,N_1359);
nor U1441 (N_1441,N_1210,N_1370);
nand U1442 (N_1442,N_1329,N_1312);
nand U1443 (N_1443,N_1254,N_1243);
or U1444 (N_1444,N_1215,N_1271);
nand U1445 (N_1445,N_1330,N_1351);
nor U1446 (N_1446,N_1378,N_1276);
nand U1447 (N_1447,N_1275,N_1349);
xnor U1448 (N_1448,N_1207,N_1209);
or U1449 (N_1449,N_1384,N_1246);
or U1450 (N_1450,N_1244,N_1381);
xnor U1451 (N_1451,N_1327,N_1236);
nand U1452 (N_1452,N_1223,N_1371);
nor U1453 (N_1453,N_1392,N_1263);
or U1454 (N_1454,N_1295,N_1347);
xnor U1455 (N_1455,N_1343,N_1232);
and U1456 (N_1456,N_1241,N_1345);
xor U1457 (N_1457,N_1325,N_1293);
nor U1458 (N_1458,N_1358,N_1398);
nor U1459 (N_1459,N_1287,N_1285);
nand U1460 (N_1460,N_1228,N_1238);
and U1461 (N_1461,N_1245,N_1315);
nor U1462 (N_1462,N_1320,N_1380);
nand U1463 (N_1463,N_1333,N_1297);
nand U1464 (N_1464,N_1261,N_1346);
nand U1465 (N_1465,N_1341,N_1222);
xnor U1466 (N_1466,N_1348,N_1369);
or U1467 (N_1467,N_1284,N_1365);
nand U1468 (N_1468,N_1367,N_1377);
nand U1469 (N_1469,N_1227,N_1281);
nor U1470 (N_1470,N_1364,N_1258);
and U1471 (N_1471,N_1272,N_1350);
and U1472 (N_1472,N_1225,N_1324);
and U1473 (N_1473,N_1237,N_1301);
nand U1474 (N_1474,N_1322,N_1386);
and U1475 (N_1475,N_1353,N_1340);
nor U1476 (N_1476,N_1356,N_1314);
and U1477 (N_1477,N_1280,N_1360);
nand U1478 (N_1478,N_1326,N_1269);
nand U1479 (N_1479,N_1362,N_1361);
and U1480 (N_1480,N_1307,N_1335);
nor U1481 (N_1481,N_1288,N_1286);
nor U1482 (N_1482,N_1368,N_1395);
or U1483 (N_1483,N_1323,N_1337);
nand U1484 (N_1484,N_1332,N_1305);
and U1485 (N_1485,N_1201,N_1251);
nor U1486 (N_1486,N_1264,N_1206);
or U1487 (N_1487,N_1279,N_1317);
xor U1488 (N_1488,N_1397,N_1213);
and U1489 (N_1489,N_1376,N_1304);
nor U1490 (N_1490,N_1249,N_1270);
nand U1491 (N_1491,N_1221,N_1382);
nand U1492 (N_1492,N_1234,N_1220);
nand U1493 (N_1493,N_1248,N_1344);
nand U1494 (N_1494,N_1259,N_1278);
and U1495 (N_1495,N_1302,N_1334);
nand U1496 (N_1496,N_1282,N_1394);
or U1497 (N_1497,N_1298,N_1212);
nand U1498 (N_1498,N_1292,N_1231);
or U1499 (N_1499,N_1214,N_1267);
and U1500 (N_1500,N_1366,N_1276);
nand U1501 (N_1501,N_1380,N_1268);
xor U1502 (N_1502,N_1310,N_1220);
or U1503 (N_1503,N_1353,N_1218);
or U1504 (N_1504,N_1304,N_1295);
nand U1505 (N_1505,N_1323,N_1369);
xor U1506 (N_1506,N_1374,N_1273);
nor U1507 (N_1507,N_1211,N_1253);
nand U1508 (N_1508,N_1265,N_1268);
and U1509 (N_1509,N_1286,N_1287);
xor U1510 (N_1510,N_1389,N_1275);
and U1511 (N_1511,N_1368,N_1334);
nand U1512 (N_1512,N_1217,N_1339);
nand U1513 (N_1513,N_1276,N_1283);
and U1514 (N_1514,N_1267,N_1344);
and U1515 (N_1515,N_1247,N_1269);
nor U1516 (N_1516,N_1319,N_1263);
nand U1517 (N_1517,N_1257,N_1232);
or U1518 (N_1518,N_1321,N_1286);
and U1519 (N_1519,N_1275,N_1309);
nand U1520 (N_1520,N_1231,N_1280);
or U1521 (N_1521,N_1229,N_1364);
nand U1522 (N_1522,N_1366,N_1316);
nor U1523 (N_1523,N_1279,N_1386);
and U1524 (N_1524,N_1366,N_1337);
xnor U1525 (N_1525,N_1389,N_1355);
and U1526 (N_1526,N_1271,N_1261);
nand U1527 (N_1527,N_1353,N_1276);
and U1528 (N_1528,N_1267,N_1326);
nand U1529 (N_1529,N_1332,N_1395);
nand U1530 (N_1530,N_1330,N_1207);
xnor U1531 (N_1531,N_1272,N_1202);
and U1532 (N_1532,N_1226,N_1313);
or U1533 (N_1533,N_1213,N_1336);
nand U1534 (N_1534,N_1203,N_1345);
xnor U1535 (N_1535,N_1324,N_1346);
or U1536 (N_1536,N_1242,N_1325);
nor U1537 (N_1537,N_1291,N_1344);
or U1538 (N_1538,N_1381,N_1308);
and U1539 (N_1539,N_1373,N_1336);
nor U1540 (N_1540,N_1368,N_1303);
and U1541 (N_1541,N_1362,N_1298);
nand U1542 (N_1542,N_1298,N_1260);
and U1543 (N_1543,N_1392,N_1311);
or U1544 (N_1544,N_1397,N_1308);
nand U1545 (N_1545,N_1260,N_1245);
nor U1546 (N_1546,N_1209,N_1366);
nand U1547 (N_1547,N_1367,N_1242);
nand U1548 (N_1548,N_1233,N_1381);
nand U1549 (N_1549,N_1345,N_1217);
nor U1550 (N_1550,N_1383,N_1328);
or U1551 (N_1551,N_1243,N_1211);
or U1552 (N_1552,N_1279,N_1264);
and U1553 (N_1553,N_1287,N_1289);
or U1554 (N_1554,N_1308,N_1331);
nor U1555 (N_1555,N_1387,N_1320);
or U1556 (N_1556,N_1217,N_1355);
nor U1557 (N_1557,N_1307,N_1209);
and U1558 (N_1558,N_1359,N_1390);
and U1559 (N_1559,N_1388,N_1248);
nand U1560 (N_1560,N_1387,N_1361);
or U1561 (N_1561,N_1396,N_1342);
nand U1562 (N_1562,N_1220,N_1207);
nor U1563 (N_1563,N_1236,N_1365);
and U1564 (N_1564,N_1284,N_1384);
and U1565 (N_1565,N_1328,N_1365);
or U1566 (N_1566,N_1239,N_1357);
nor U1567 (N_1567,N_1255,N_1263);
and U1568 (N_1568,N_1289,N_1211);
or U1569 (N_1569,N_1286,N_1275);
and U1570 (N_1570,N_1315,N_1385);
nor U1571 (N_1571,N_1261,N_1307);
nand U1572 (N_1572,N_1334,N_1335);
nor U1573 (N_1573,N_1378,N_1353);
or U1574 (N_1574,N_1369,N_1271);
or U1575 (N_1575,N_1362,N_1331);
xor U1576 (N_1576,N_1230,N_1348);
and U1577 (N_1577,N_1332,N_1271);
or U1578 (N_1578,N_1343,N_1373);
and U1579 (N_1579,N_1219,N_1285);
nand U1580 (N_1580,N_1392,N_1266);
or U1581 (N_1581,N_1284,N_1234);
xor U1582 (N_1582,N_1263,N_1239);
nand U1583 (N_1583,N_1298,N_1328);
nand U1584 (N_1584,N_1387,N_1371);
and U1585 (N_1585,N_1358,N_1355);
or U1586 (N_1586,N_1329,N_1350);
or U1587 (N_1587,N_1310,N_1208);
or U1588 (N_1588,N_1290,N_1390);
nor U1589 (N_1589,N_1335,N_1218);
or U1590 (N_1590,N_1281,N_1315);
nand U1591 (N_1591,N_1363,N_1390);
nor U1592 (N_1592,N_1336,N_1396);
nor U1593 (N_1593,N_1254,N_1210);
nand U1594 (N_1594,N_1246,N_1219);
and U1595 (N_1595,N_1235,N_1326);
nand U1596 (N_1596,N_1353,N_1376);
nand U1597 (N_1597,N_1246,N_1279);
nand U1598 (N_1598,N_1223,N_1298);
nor U1599 (N_1599,N_1226,N_1228);
nand U1600 (N_1600,N_1527,N_1550);
nand U1601 (N_1601,N_1431,N_1595);
and U1602 (N_1602,N_1545,N_1581);
nor U1603 (N_1603,N_1566,N_1551);
nand U1604 (N_1604,N_1511,N_1484);
or U1605 (N_1605,N_1517,N_1478);
nand U1606 (N_1606,N_1435,N_1421);
nor U1607 (N_1607,N_1419,N_1403);
or U1608 (N_1608,N_1492,N_1575);
nand U1609 (N_1609,N_1573,N_1570);
nand U1610 (N_1610,N_1490,N_1475);
nand U1611 (N_1611,N_1474,N_1587);
nand U1612 (N_1612,N_1506,N_1548);
nand U1613 (N_1613,N_1466,N_1503);
or U1614 (N_1614,N_1430,N_1510);
nand U1615 (N_1615,N_1443,N_1469);
or U1616 (N_1616,N_1540,N_1442);
nor U1617 (N_1617,N_1557,N_1446);
nand U1618 (N_1618,N_1516,N_1565);
nor U1619 (N_1619,N_1468,N_1562);
nor U1620 (N_1620,N_1445,N_1571);
or U1621 (N_1621,N_1589,N_1505);
nor U1622 (N_1622,N_1494,N_1464);
or U1623 (N_1623,N_1546,N_1487);
nor U1624 (N_1624,N_1448,N_1463);
nor U1625 (N_1625,N_1454,N_1501);
nor U1626 (N_1626,N_1453,N_1499);
nand U1627 (N_1627,N_1572,N_1496);
and U1628 (N_1628,N_1576,N_1569);
or U1629 (N_1629,N_1436,N_1529);
nor U1630 (N_1630,N_1561,N_1476);
nor U1631 (N_1631,N_1567,N_1525);
or U1632 (N_1632,N_1486,N_1524);
or U1633 (N_1633,N_1542,N_1416);
nand U1634 (N_1634,N_1521,N_1405);
and U1635 (N_1635,N_1554,N_1444);
and U1636 (N_1636,N_1426,N_1509);
or U1637 (N_1637,N_1513,N_1401);
or U1638 (N_1638,N_1456,N_1584);
or U1639 (N_1639,N_1532,N_1479);
nand U1640 (N_1640,N_1408,N_1497);
or U1641 (N_1641,N_1585,N_1417);
and U1642 (N_1642,N_1438,N_1520);
or U1643 (N_1643,N_1472,N_1564);
nor U1644 (N_1644,N_1433,N_1493);
nor U1645 (N_1645,N_1526,N_1578);
nand U1646 (N_1646,N_1514,N_1413);
or U1647 (N_1647,N_1425,N_1579);
nand U1648 (N_1648,N_1414,N_1488);
nor U1649 (N_1649,N_1498,N_1535);
and U1650 (N_1650,N_1591,N_1491);
and U1651 (N_1651,N_1536,N_1537);
xor U1652 (N_1652,N_1541,N_1507);
and U1653 (N_1653,N_1553,N_1410);
xor U1654 (N_1654,N_1485,N_1512);
nand U1655 (N_1655,N_1409,N_1404);
nor U1656 (N_1656,N_1500,N_1559);
nor U1657 (N_1657,N_1422,N_1462);
and U1658 (N_1658,N_1577,N_1593);
xor U1659 (N_1659,N_1523,N_1495);
nor U1660 (N_1660,N_1598,N_1406);
nand U1661 (N_1661,N_1519,N_1539);
nor U1662 (N_1662,N_1465,N_1534);
or U1663 (N_1663,N_1411,N_1481);
or U1664 (N_1664,N_1504,N_1455);
or U1665 (N_1665,N_1480,N_1471);
and U1666 (N_1666,N_1580,N_1450);
xor U1667 (N_1667,N_1460,N_1508);
xor U1668 (N_1668,N_1522,N_1558);
nor U1669 (N_1669,N_1458,N_1586);
nor U1670 (N_1670,N_1418,N_1531);
and U1671 (N_1671,N_1467,N_1432);
xor U1672 (N_1672,N_1563,N_1449);
nor U1673 (N_1673,N_1515,N_1544);
nor U1674 (N_1674,N_1568,N_1549);
nor U1675 (N_1675,N_1447,N_1489);
and U1676 (N_1676,N_1574,N_1428);
nand U1677 (N_1677,N_1461,N_1583);
and U1678 (N_1678,N_1560,N_1594);
or U1679 (N_1679,N_1420,N_1439);
nand U1680 (N_1680,N_1470,N_1502);
or U1681 (N_1681,N_1407,N_1543);
or U1682 (N_1682,N_1423,N_1555);
xor U1683 (N_1683,N_1477,N_1412);
and U1684 (N_1684,N_1483,N_1588);
nand U1685 (N_1685,N_1528,N_1552);
nand U1686 (N_1686,N_1538,N_1518);
nand U1687 (N_1687,N_1437,N_1473);
nor U1688 (N_1688,N_1400,N_1556);
nor U1689 (N_1689,N_1590,N_1452);
and U1690 (N_1690,N_1451,N_1440);
nand U1691 (N_1691,N_1533,N_1597);
nor U1692 (N_1692,N_1429,N_1427);
nor U1693 (N_1693,N_1459,N_1530);
or U1694 (N_1694,N_1596,N_1434);
nand U1695 (N_1695,N_1482,N_1582);
xor U1696 (N_1696,N_1441,N_1599);
nor U1697 (N_1697,N_1592,N_1457);
nor U1698 (N_1698,N_1424,N_1415);
and U1699 (N_1699,N_1547,N_1402);
or U1700 (N_1700,N_1408,N_1480);
nand U1701 (N_1701,N_1479,N_1588);
xor U1702 (N_1702,N_1513,N_1593);
and U1703 (N_1703,N_1455,N_1424);
or U1704 (N_1704,N_1491,N_1574);
nor U1705 (N_1705,N_1590,N_1584);
xor U1706 (N_1706,N_1413,N_1460);
or U1707 (N_1707,N_1442,N_1511);
and U1708 (N_1708,N_1433,N_1594);
nor U1709 (N_1709,N_1574,N_1480);
or U1710 (N_1710,N_1454,N_1451);
xor U1711 (N_1711,N_1550,N_1412);
nand U1712 (N_1712,N_1517,N_1558);
and U1713 (N_1713,N_1444,N_1577);
xnor U1714 (N_1714,N_1408,N_1455);
or U1715 (N_1715,N_1597,N_1562);
or U1716 (N_1716,N_1434,N_1508);
or U1717 (N_1717,N_1436,N_1496);
xor U1718 (N_1718,N_1441,N_1423);
nand U1719 (N_1719,N_1532,N_1496);
nand U1720 (N_1720,N_1533,N_1441);
nand U1721 (N_1721,N_1586,N_1465);
and U1722 (N_1722,N_1402,N_1461);
or U1723 (N_1723,N_1557,N_1472);
nand U1724 (N_1724,N_1570,N_1413);
and U1725 (N_1725,N_1535,N_1430);
xnor U1726 (N_1726,N_1531,N_1483);
nand U1727 (N_1727,N_1574,N_1594);
and U1728 (N_1728,N_1420,N_1408);
xnor U1729 (N_1729,N_1466,N_1498);
or U1730 (N_1730,N_1516,N_1523);
xnor U1731 (N_1731,N_1458,N_1441);
xnor U1732 (N_1732,N_1578,N_1441);
nand U1733 (N_1733,N_1482,N_1519);
or U1734 (N_1734,N_1549,N_1496);
or U1735 (N_1735,N_1592,N_1453);
and U1736 (N_1736,N_1444,N_1586);
and U1737 (N_1737,N_1582,N_1580);
or U1738 (N_1738,N_1508,N_1592);
and U1739 (N_1739,N_1480,N_1550);
or U1740 (N_1740,N_1400,N_1583);
or U1741 (N_1741,N_1442,N_1422);
and U1742 (N_1742,N_1436,N_1587);
and U1743 (N_1743,N_1445,N_1521);
and U1744 (N_1744,N_1501,N_1588);
nand U1745 (N_1745,N_1493,N_1580);
xnor U1746 (N_1746,N_1537,N_1402);
and U1747 (N_1747,N_1504,N_1437);
nor U1748 (N_1748,N_1439,N_1410);
nand U1749 (N_1749,N_1546,N_1468);
or U1750 (N_1750,N_1498,N_1555);
nand U1751 (N_1751,N_1494,N_1572);
xor U1752 (N_1752,N_1531,N_1500);
and U1753 (N_1753,N_1545,N_1465);
and U1754 (N_1754,N_1555,N_1575);
nor U1755 (N_1755,N_1448,N_1460);
xnor U1756 (N_1756,N_1558,N_1496);
nor U1757 (N_1757,N_1572,N_1557);
or U1758 (N_1758,N_1444,N_1498);
xnor U1759 (N_1759,N_1422,N_1428);
and U1760 (N_1760,N_1464,N_1455);
and U1761 (N_1761,N_1420,N_1586);
and U1762 (N_1762,N_1568,N_1402);
nand U1763 (N_1763,N_1423,N_1557);
xnor U1764 (N_1764,N_1549,N_1595);
nand U1765 (N_1765,N_1586,N_1435);
nand U1766 (N_1766,N_1491,N_1542);
or U1767 (N_1767,N_1483,N_1490);
and U1768 (N_1768,N_1417,N_1504);
and U1769 (N_1769,N_1586,N_1493);
or U1770 (N_1770,N_1488,N_1498);
nor U1771 (N_1771,N_1474,N_1424);
or U1772 (N_1772,N_1483,N_1597);
nand U1773 (N_1773,N_1429,N_1430);
nor U1774 (N_1774,N_1414,N_1424);
nor U1775 (N_1775,N_1536,N_1474);
or U1776 (N_1776,N_1401,N_1413);
nor U1777 (N_1777,N_1487,N_1508);
and U1778 (N_1778,N_1597,N_1532);
or U1779 (N_1779,N_1522,N_1505);
nand U1780 (N_1780,N_1463,N_1432);
and U1781 (N_1781,N_1404,N_1492);
and U1782 (N_1782,N_1583,N_1438);
nand U1783 (N_1783,N_1535,N_1435);
nor U1784 (N_1784,N_1413,N_1506);
and U1785 (N_1785,N_1540,N_1451);
nand U1786 (N_1786,N_1505,N_1519);
xnor U1787 (N_1787,N_1579,N_1418);
and U1788 (N_1788,N_1525,N_1497);
or U1789 (N_1789,N_1579,N_1486);
nor U1790 (N_1790,N_1488,N_1553);
or U1791 (N_1791,N_1566,N_1530);
xnor U1792 (N_1792,N_1539,N_1592);
nor U1793 (N_1793,N_1447,N_1418);
nand U1794 (N_1794,N_1407,N_1405);
nor U1795 (N_1795,N_1582,N_1475);
nand U1796 (N_1796,N_1510,N_1477);
xnor U1797 (N_1797,N_1475,N_1515);
nand U1798 (N_1798,N_1477,N_1552);
and U1799 (N_1799,N_1586,N_1421);
and U1800 (N_1800,N_1717,N_1716);
or U1801 (N_1801,N_1738,N_1646);
and U1802 (N_1802,N_1644,N_1675);
and U1803 (N_1803,N_1712,N_1792);
nand U1804 (N_1804,N_1768,N_1650);
or U1805 (N_1805,N_1776,N_1631);
nor U1806 (N_1806,N_1658,N_1711);
nor U1807 (N_1807,N_1622,N_1672);
and U1808 (N_1808,N_1721,N_1726);
or U1809 (N_1809,N_1641,N_1742);
or U1810 (N_1810,N_1702,N_1795);
nor U1811 (N_1811,N_1627,N_1680);
nand U1812 (N_1812,N_1770,N_1777);
or U1813 (N_1813,N_1699,N_1784);
nand U1814 (N_1814,N_1608,N_1610);
nand U1815 (N_1815,N_1660,N_1730);
or U1816 (N_1816,N_1718,N_1625);
or U1817 (N_1817,N_1630,N_1665);
and U1818 (N_1818,N_1753,N_1612);
nand U1819 (N_1819,N_1760,N_1629);
nor U1820 (N_1820,N_1744,N_1766);
nor U1821 (N_1821,N_1727,N_1689);
nand U1822 (N_1822,N_1657,N_1663);
nand U1823 (N_1823,N_1750,N_1626);
nor U1824 (N_1824,N_1791,N_1743);
and U1825 (N_1825,N_1692,N_1648);
nor U1826 (N_1826,N_1705,N_1772);
nor U1827 (N_1827,N_1737,N_1676);
and U1828 (N_1828,N_1670,N_1634);
and U1829 (N_1829,N_1731,N_1653);
nor U1830 (N_1830,N_1624,N_1667);
nor U1831 (N_1831,N_1681,N_1707);
nor U1832 (N_1832,N_1618,N_1682);
nor U1833 (N_1833,N_1762,N_1715);
nor U1834 (N_1834,N_1633,N_1756);
and U1835 (N_1835,N_1602,N_1684);
and U1836 (N_1836,N_1723,N_1751);
nand U1837 (N_1837,N_1786,N_1790);
nand U1838 (N_1838,N_1655,N_1673);
and U1839 (N_1839,N_1773,N_1606);
xor U1840 (N_1840,N_1708,N_1788);
and U1841 (N_1841,N_1669,N_1604);
or U1842 (N_1842,N_1685,N_1799);
xor U1843 (N_1843,N_1628,N_1656);
xor U1844 (N_1844,N_1782,N_1700);
nand U1845 (N_1845,N_1758,N_1639);
or U1846 (N_1846,N_1763,N_1796);
or U1847 (N_1847,N_1746,N_1764);
nor U1848 (N_1848,N_1607,N_1703);
nand U1849 (N_1849,N_1601,N_1710);
or U1850 (N_1850,N_1704,N_1706);
nand U1851 (N_1851,N_1749,N_1739);
and U1852 (N_1852,N_1771,N_1611);
or U1853 (N_1853,N_1785,N_1761);
and U1854 (N_1854,N_1609,N_1613);
nor U1855 (N_1855,N_1798,N_1740);
xor U1856 (N_1856,N_1695,N_1637);
nor U1857 (N_1857,N_1623,N_1619);
or U1858 (N_1858,N_1769,N_1635);
and U1859 (N_1859,N_1620,N_1666);
nor U1860 (N_1860,N_1720,N_1678);
nand U1861 (N_1861,N_1779,N_1748);
nor U1862 (N_1862,N_1775,N_1719);
nand U1863 (N_1863,N_1645,N_1747);
and U1864 (N_1864,N_1668,N_1724);
nand U1865 (N_1865,N_1632,N_1725);
nand U1866 (N_1866,N_1643,N_1793);
nor U1867 (N_1867,N_1603,N_1651);
nor U1868 (N_1868,N_1652,N_1600);
nand U1869 (N_1869,N_1638,N_1781);
and U1870 (N_1870,N_1759,N_1696);
nor U1871 (N_1871,N_1778,N_1614);
nand U1872 (N_1872,N_1732,N_1755);
or U1873 (N_1873,N_1780,N_1621);
and U1874 (N_1874,N_1714,N_1642);
or U1875 (N_1875,N_1617,N_1736);
or U1876 (N_1876,N_1662,N_1679);
and U1877 (N_1877,N_1733,N_1664);
xnor U1878 (N_1878,N_1728,N_1783);
nor U1879 (N_1879,N_1734,N_1757);
and U1880 (N_1880,N_1729,N_1649);
nor U1881 (N_1881,N_1674,N_1654);
xnor U1882 (N_1882,N_1794,N_1741);
nor U1883 (N_1883,N_1774,N_1647);
nor U1884 (N_1884,N_1694,N_1690);
nor U1885 (N_1885,N_1735,N_1754);
nor U1886 (N_1886,N_1752,N_1686);
nor U1887 (N_1887,N_1698,N_1797);
nand U1888 (N_1888,N_1767,N_1787);
and U1889 (N_1889,N_1688,N_1683);
and U1890 (N_1890,N_1616,N_1709);
or U1891 (N_1891,N_1605,N_1691);
nand U1892 (N_1892,N_1615,N_1745);
or U1893 (N_1893,N_1661,N_1722);
nand U1894 (N_1894,N_1671,N_1697);
xor U1895 (N_1895,N_1687,N_1677);
nor U1896 (N_1896,N_1693,N_1713);
or U1897 (N_1897,N_1765,N_1789);
and U1898 (N_1898,N_1701,N_1640);
nor U1899 (N_1899,N_1659,N_1636);
nor U1900 (N_1900,N_1749,N_1679);
or U1901 (N_1901,N_1667,N_1683);
nor U1902 (N_1902,N_1664,N_1672);
and U1903 (N_1903,N_1657,N_1637);
and U1904 (N_1904,N_1778,N_1640);
and U1905 (N_1905,N_1621,N_1723);
or U1906 (N_1906,N_1735,N_1688);
xnor U1907 (N_1907,N_1777,N_1725);
and U1908 (N_1908,N_1655,N_1646);
nor U1909 (N_1909,N_1613,N_1725);
or U1910 (N_1910,N_1766,N_1710);
or U1911 (N_1911,N_1649,N_1601);
or U1912 (N_1912,N_1751,N_1712);
or U1913 (N_1913,N_1772,N_1693);
and U1914 (N_1914,N_1758,N_1779);
nor U1915 (N_1915,N_1685,N_1673);
or U1916 (N_1916,N_1779,N_1642);
or U1917 (N_1917,N_1794,N_1693);
or U1918 (N_1918,N_1775,N_1646);
nand U1919 (N_1919,N_1704,N_1754);
xor U1920 (N_1920,N_1763,N_1774);
nand U1921 (N_1921,N_1783,N_1770);
and U1922 (N_1922,N_1607,N_1619);
or U1923 (N_1923,N_1725,N_1653);
xnor U1924 (N_1924,N_1602,N_1790);
and U1925 (N_1925,N_1762,N_1770);
or U1926 (N_1926,N_1706,N_1720);
nor U1927 (N_1927,N_1741,N_1615);
nor U1928 (N_1928,N_1708,N_1711);
nand U1929 (N_1929,N_1788,N_1713);
nand U1930 (N_1930,N_1701,N_1747);
or U1931 (N_1931,N_1621,N_1671);
nand U1932 (N_1932,N_1665,N_1677);
nand U1933 (N_1933,N_1611,N_1765);
nor U1934 (N_1934,N_1734,N_1670);
nand U1935 (N_1935,N_1606,N_1648);
xor U1936 (N_1936,N_1732,N_1675);
and U1937 (N_1937,N_1725,N_1691);
nor U1938 (N_1938,N_1780,N_1735);
nand U1939 (N_1939,N_1767,N_1713);
nor U1940 (N_1940,N_1633,N_1676);
and U1941 (N_1941,N_1760,N_1729);
or U1942 (N_1942,N_1649,N_1783);
nor U1943 (N_1943,N_1603,N_1758);
nand U1944 (N_1944,N_1665,N_1709);
and U1945 (N_1945,N_1716,N_1749);
and U1946 (N_1946,N_1622,N_1662);
nor U1947 (N_1947,N_1625,N_1779);
or U1948 (N_1948,N_1740,N_1746);
xor U1949 (N_1949,N_1775,N_1636);
nor U1950 (N_1950,N_1637,N_1726);
or U1951 (N_1951,N_1613,N_1750);
xnor U1952 (N_1952,N_1625,N_1624);
nand U1953 (N_1953,N_1692,N_1611);
nand U1954 (N_1954,N_1748,N_1763);
or U1955 (N_1955,N_1658,N_1600);
nor U1956 (N_1956,N_1666,N_1661);
nor U1957 (N_1957,N_1664,N_1710);
and U1958 (N_1958,N_1661,N_1763);
xnor U1959 (N_1959,N_1674,N_1774);
and U1960 (N_1960,N_1625,N_1759);
nand U1961 (N_1961,N_1727,N_1736);
or U1962 (N_1962,N_1724,N_1798);
nor U1963 (N_1963,N_1677,N_1627);
nor U1964 (N_1964,N_1793,N_1626);
nand U1965 (N_1965,N_1675,N_1708);
nand U1966 (N_1966,N_1736,N_1639);
xnor U1967 (N_1967,N_1796,N_1749);
nor U1968 (N_1968,N_1748,N_1774);
or U1969 (N_1969,N_1624,N_1687);
and U1970 (N_1970,N_1620,N_1720);
nand U1971 (N_1971,N_1790,N_1776);
nand U1972 (N_1972,N_1731,N_1751);
or U1973 (N_1973,N_1768,N_1756);
and U1974 (N_1974,N_1671,N_1685);
nand U1975 (N_1975,N_1752,N_1668);
nor U1976 (N_1976,N_1795,N_1620);
and U1977 (N_1977,N_1641,N_1763);
nor U1978 (N_1978,N_1674,N_1667);
and U1979 (N_1979,N_1670,N_1665);
and U1980 (N_1980,N_1777,N_1650);
nand U1981 (N_1981,N_1768,N_1701);
nand U1982 (N_1982,N_1676,N_1630);
nor U1983 (N_1983,N_1687,N_1772);
nor U1984 (N_1984,N_1669,N_1793);
xor U1985 (N_1985,N_1616,N_1717);
or U1986 (N_1986,N_1792,N_1781);
nor U1987 (N_1987,N_1639,N_1770);
nor U1988 (N_1988,N_1762,N_1686);
or U1989 (N_1989,N_1686,N_1699);
nor U1990 (N_1990,N_1604,N_1795);
nand U1991 (N_1991,N_1722,N_1633);
nor U1992 (N_1992,N_1717,N_1738);
or U1993 (N_1993,N_1736,N_1657);
nand U1994 (N_1994,N_1619,N_1644);
or U1995 (N_1995,N_1719,N_1729);
nor U1996 (N_1996,N_1710,N_1780);
or U1997 (N_1997,N_1772,N_1697);
xnor U1998 (N_1998,N_1673,N_1710);
or U1999 (N_1999,N_1678,N_1793);
xnor U2000 (N_2000,N_1883,N_1818);
or U2001 (N_2001,N_1817,N_1992);
and U2002 (N_2002,N_1861,N_1850);
xnor U2003 (N_2003,N_1921,N_1840);
and U2004 (N_2004,N_1815,N_1887);
and U2005 (N_2005,N_1917,N_1969);
or U2006 (N_2006,N_1916,N_1837);
xnor U2007 (N_2007,N_1984,N_1985);
and U2008 (N_2008,N_1943,N_1871);
and U2009 (N_2009,N_1967,N_1972);
and U2010 (N_2010,N_1875,N_1841);
xnor U2011 (N_2011,N_1965,N_1877);
or U2012 (N_2012,N_1983,N_1940);
xor U2013 (N_2013,N_1987,N_1957);
nand U2014 (N_2014,N_1941,N_1829);
nor U2015 (N_2015,N_1931,N_1919);
or U2016 (N_2016,N_1801,N_1935);
or U2017 (N_2017,N_1933,N_1962);
nand U2018 (N_2018,N_1844,N_1907);
and U2019 (N_2019,N_1963,N_1993);
nand U2020 (N_2020,N_1975,N_1858);
or U2021 (N_2021,N_1839,N_1989);
nand U2022 (N_2022,N_1833,N_1869);
nor U2023 (N_2023,N_1816,N_1878);
and U2024 (N_2024,N_1947,N_1981);
and U2025 (N_2025,N_1823,N_1835);
or U2026 (N_2026,N_1929,N_1930);
or U2027 (N_2027,N_1942,N_1855);
or U2028 (N_2028,N_1843,N_1889);
and U2029 (N_2029,N_1954,N_1934);
xor U2030 (N_2030,N_1892,N_1831);
and U2031 (N_2031,N_1863,N_1970);
and U2032 (N_2032,N_1902,N_1828);
nand U2033 (N_2033,N_1853,N_1925);
or U2034 (N_2034,N_1979,N_1956);
nand U2035 (N_2035,N_1856,N_1959);
nand U2036 (N_2036,N_1882,N_1950);
nor U2037 (N_2037,N_1918,N_1923);
nand U2038 (N_2038,N_1982,N_1926);
nand U2039 (N_2039,N_1859,N_1913);
nand U2040 (N_2040,N_1802,N_1980);
xnor U2041 (N_2041,N_1958,N_1945);
nor U2042 (N_2042,N_1805,N_1881);
nand U2043 (N_2043,N_1827,N_1949);
and U2044 (N_2044,N_1819,N_1922);
xor U2045 (N_2045,N_1998,N_1909);
and U2046 (N_2046,N_1852,N_1914);
nor U2047 (N_2047,N_1910,N_1822);
and U2048 (N_2048,N_1834,N_1994);
nand U2049 (N_2049,N_1857,N_1860);
and U2050 (N_2050,N_1814,N_1873);
and U2051 (N_2051,N_1847,N_1865);
nand U2052 (N_2052,N_1904,N_1888);
nor U2053 (N_2053,N_1826,N_1920);
or U2054 (N_2054,N_1899,N_1948);
or U2055 (N_2055,N_1825,N_1915);
xor U2056 (N_2056,N_1867,N_1806);
nor U2057 (N_2057,N_1905,N_1986);
nand U2058 (N_2058,N_1848,N_1936);
nor U2059 (N_2059,N_1812,N_1976);
and U2060 (N_2060,N_1811,N_1820);
nor U2061 (N_2061,N_1866,N_1898);
nor U2062 (N_2062,N_1971,N_1932);
nor U2063 (N_2063,N_1809,N_1938);
or U2064 (N_2064,N_1912,N_1851);
xnor U2065 (N_2065,N_1842,N_1991);
or U2066 (N_2066,N_1995,N_1928);
nand U2067 (N_2067,N_1830,N_1953);
nor U2068 (N_2068,N_1832,N_1961);
nand U2069 (N_2069,N_1821,N_1804);
nor U2070 (N_2070,N_1813,N_1846);
or U2071 (N_2071,N_1974,N_1960);
and U2072 (N_2072,N_1990,N_1901);
and U2073 (N_2073,N_1824,N_1897);
xor U2074 (N_2074,N_1868,N_1885);
nor U2075 (N_2075,N_1911,N_1999);
and U2076 (N_2076,N_1803,N_1880);
nand U2077 (N_2077,N_1968,N_1951);
or U2078 (N_2078,N_1973,N_1876);
nand U2079 (N_2079,N_1808,N_1893);
or U2080 (N_2080,N_1838,N_1937);
or U2081 (N_2081,N_1807,N_1946);
or U2082 (N_2082,N_1886,N_1810);
nand U2083 (N_2083,N_1964,N_1864);
or U2084 (N_2084,N_1939,N_1908);
or U2085 (N_2085,N_1874,N_1800);
and U2086 (N_2086,N_1906,N_1894);
or U2087 (N_2087,N_1879,N_1978);
nand U2088 (N_2088,N_1996,N_1895);
nor U2089 (N_2089,N_1896,N_1872);
nor U2090 (N_2090,N_1845,N_1870);
or U2091 (N_2091,N_1988,N_1927);
nor U2092 (N_2092,N_1900,N_1952);
and U2093 (N_2093,N_1849,N_1903);
and U2094 (N_2094,N_1890,N_1862);
and U2095 (N_2095,N_1854,N_1884);
nor U2096 (N_2096,N_1944,N_1836);
and U2097 (N_2097,N_1924,N_1977);
nand U2098 (N_2098,N_1997,N_1955);
nor U2099 (N_2099,N_1966,N_1891);
and U2100 (N_2100,N_1923,N_1823);
or U2101 (N_2101,N_1861,N_1937);
and U2102 (N_2102,N_1959,N_1965);
or U2103 (N_2103,N_1936,N_1962);
and U2104 (N_2104,N_1902,N_1917);
and U2105 (N_2105,N_1859,N_1850);
or U2106 (N_2106,N_1912,N_1874);
nand U2107 (N_2107,N_1887,N_1934);
or U2108 (N_2108,N_1804,N_1963);
and U2109 (N_2109,N_1839,N_1849);
nand U2110 (N_2110,N_1830,N_1994);
nor U2111 (N_2111,N_1877,N_1819);
or U2112 (N_2112,N_1802,N_1990);
and U2113 (N_2113,N_1846,N_1983);
xor U2114 (N_2114,N_1941,N_1995);
xor U2115 (N_2115,N_1804,N_1984);
nand U2116 (N_2116,N_1802,N_1982);
nand U2117 (N_2117,N_1972,N_1847);
nor U2118 (N_2118,N_1887,N_1966);
or U2119 (N_2119,N_1971,N_1922);
and U2120 (N_2120,N_1929,N_1935);
nand U2121 (N_2121,N_1919,N_1832);
nor U2122 (N_2122,N_1950,N_1963);
and U2123 (N_2123,N_1939,N_1830);
nand U2124 (N_2124,N_1934,N_1931);
xnor U2125 (N_2125,N_1859,N_1983);
nand U2126 (N_2126,N_1926,N_1854);
and U2127 (N_2127,N_1842,N_1943);
nand U2128 (N_2128,N_1975,N_1825);
nand U2129 (N_2129,N_1829,N_1901);
nor U2130 (N_2130,N_1811,N_1950);
and U2131 (N_2131,N_1909,N_1809);
xor U2132 (N_2132,N_1815,N_1849);
nor U2133 (N_2133,N_1816,N_1904);
nor U2134 (N_2134,N_1805,N_1896);
or U2135 (N_2135,N_1910,N_1873);
nand U2136 (N_2136,N_1872,N_1832);
nor U2137 (N_2137,N_1896,N_1953);
nand U2138 (N_2138,N_1831,N_1983);
or U2139 (N_2139,N_1834,N_1837);
or U2140 (N_2140,N_1913,N_1905);
and U2141 (N_2141,N_1890,N_1801);
or U2142 (N_2142,N_1984,N_1938);
or U2143 (N_2143,N_1989,N_1806);
or U2144 (N_2144,N_1887,N_1801);
nor U2145 (N_2145,N_1975,N_1965);
or U2146 (N_2146,N_1811,N_1812);
nor U2147 (N_2147,N_1977,N_1915);
or U2148 (N_2148,N_1837,N_1891);
nand U2149 (N_2149,N_1987,N_1838);
nand U2150 (N_2150,N_1917,N_1834);
nor U2151 (N_2151,N_1960,N_1873);
and U2152 (N_2152,N_1951,N_1842);
nand U2153 (N_2153,N_1893,N_1835);
nor U2154 (N_2154,N_1933,N_1809);
nor U2155 (N_2155,N_1805,N_1984);
or U2156 (N_2156,N_1811,N_1891);
or U2157 (N_2157,N_1992,N_1808);
or U2158 (N_2158,N_1822,N_1886);
and U2159 (N_2159,N_1896,N_1804);
nand U2160 (N_2160,N_1900,N_1896);
nand U2161 (N_2161,N_1820,N_1907);
nor U2162 (N_2162,N_1932,N_1941);
or U2163 (N_2163,N_1900,N_1970);
nor U2164 (N_2164,N_1995,N_1806);
and U2165 (N_2165,N_1844,N_1908);
or U2166 (N_2166,N_1953,N_1943);
nor U2167 (N_2167,N_1924,N_1818);
xor U2168 (N_2168,N_1864,N_1847);
nand U2169 (N_2169,N_1921,N_1981);
nand U2170 (N_2170,N_1821,N_1928);
or U2171 (N_2171,N_1964,N_1945);
and U2172 (N_2172,N_1967,N_1836);
nand U2173 (N_2173,N_1871,N_1957);
nor U2174 (N_2174,N_1930,N_1844);
nor U2175 (N_2175,N_1983,N_1903);
and U2176 (N_2176,N_1889,N_1893);
and U2177 (N_2177,N_1824,N_1892);
nor U2178 (N_2178,N_1951,N_1868);
nand U2179 (N_2179,N_1877,N_1813);
nor U2180 (N_2180,N_1898,N_1933);
or U2181 (N_2181,N_1974,N_1804);
nor U2182 (N_2182,N_1822,N_1948);
nor U2183 (N_2183,N_1805,N_1835);
and U2184 (N_2184,N_1997,N_1967);
nand U2185 (N_2185,N_1918,N_1858);
nand U2186 (N_2186,N_1870,N_1932);
xnor U2187 (N_2187,N_1928,N_1976);
xor U2188 (N_2188,N_1982,N_1805);
nand U2189 (N_2189,N_1803,N_1956);
and U2190 (N_2190,N_1834,N_1848);
and U2191 (N_2191,N_1833,N_1906);
and U2192 (N_2192,N_1827,N_1841);
nand U2193 (N_2193,N_1907,N_1928);
or U2194 (N_2194,N_1938,N_1995);
xnor U2195 (N_2195,N_1819,N_1950);
and U2196 (N_2196,N_1915,N_1913);
nand U2197 (N_2197,N_1921,N_1875);
or U2198 (N_2198,N_1859,N_1865);
nand U2199 (N_2199,N_1822,N_1880);
nand U2200 (N_2200,N_2177,N_2046);
and U2201 (N_2201,N_2172,N_2060);
and U2202 (N_2202,N_2113,N_2003);
nor U2203 (N_2203,N_2057,N_2047);
and U2204 (N_2204,N_2085,N_2009);
and U2205 (N_2205,N_2173,N_2011);
xnor U2206 (N_2206,N_2073,N_2038);
or U2207 (N_2207,N_2028,N_2114);
or U2208 (N_2208,N_2170,N_2098);
nand U2209 (N_2209,N_2184,N_2005);
or U2210 (N_2210,N_2029,N_2145);
and U2211 (N_2211,N_2023,N_2040);
nor U2212 (N_2212,N_2193,N_2151);
nor U2213 (N_2213,N_2002,N_2055);
or U2214 (N_2214,N_2006,N_2137);
or U2215 (N_2215,N_2075,N_2014);
nand U2216 (N_2216,N_2051,N_2026);
nor U2217 (N_2217,N_2016,N_2128);
nand U2218 (N_2218,N_2167,N_2076);
nand U2219 (N_2219,N_2130,N_2069);
or U2220 (N_2220,N_2061,N_2065);
xnor U2221 (N_2221,N_2082,N_2067);
or U2222 (N_2222,N_2086,N_2070);
and U2223 (N_2223,N_2135,N_2168);
nand U2224 (N_2224,N_2106,N_2150);
nand U2225 (N_2225,N_2125,N_2102);
nand U2226 (N_2226,N_2068,N_2066);
or U2227 (N_2227,N_2189,N_2183);
and U2228 (N_2228,N_2131,N_2089);
xor U2229 (N_2229,N_2115,N_2105);
and U2230 (N_2230,N_2097,N_2000);
nand U2231 (N_2231,N_2101,N_2186);
xnor U2232 (N_2232,N_2136,N_2163);
or U2233 (N_2233,N_2013,N_2141);
and U2234 (N_2234,N_2071,N_2160);
nand U2235 (N_2235,N_2117,N_2034);
and U2236 (N_2236,N_2093,N_2024);
nor U2237 (N_2237,N_2153,N_2157);
nand U2238 (N_2238,N_2036,N_2008);
nor U2239 (N_2239,N_2081,N_2165);
or U2240 (N_2240,N_2156,N_2022);
or U2241 (N_2241,N_2030,N_2010);
nand U2242 (N_2242,N_2012,N_2110);
and U2243 (N_2243,N_2142,N_2017);
nor U2244 (N_2244,N_2092,N_2166);
nor U2245 (N_2245,N_2180,N_2133);
nor U2246 (N_2246,N_2127,N_2149);
nand U2247 (N_2247,N_2095,N_2094);
nand U2248 (N_2248,N_2155,N_2045);
nand U2249 (N_2249,N_2041,N_2143);
xor U2250 (N_2250,N_2072,N_2198);
nand U2251 (N_2251,N_2112,N_2126);
or U2252 (N_2252,N_2171,N_2139);
nor U2253 (N_2253,N_2091,N_2132);
xnor U2254 (N_2254,N_2162,N_2096);
and U2255 (N_2255,N_2129,N_2004);
nor U2256 (N_2256,N_2104,N_2083);
and U2257 (N_2257,N_2182,N_2074);
or U2258 (N_2258,N_2175,N_2174);
nor U2259 (N_2259,N_2032,N_2191);
and U2260 (N_2260,N_2107,N_2148);
nand U2261 (N_2261,N_2018,N_2048);
and U2262 (N_2262,N_2176,N_2144);
or U2263 (N_2263,N_2140,N_2181);
and U2264 (N_2264,N_2001,N_2059);
nand U2265 (N_2265,N_2120,N_2108);
nand U2266 (N_2266,N_2161,N_2037);
or U2267 (N_2267,N_2197,N_2195);
and U2268 (N_2268,N_2042,N_2146);
or U2269 (N_2269,N_2015,N_2169);
nor U2270 (N_2270,N_2134,N_2053);
nor U2271 (N_2271,N_2088,N_2190);
nand U2272 (N_2272,N_2147,N_2178);
nor U2273 (N_2273,N_2077,N_2056);
or U2274 (N_2274,N_2138,N_2121);
and U2275 (N_2275,N_2019,N_2062);
and U2276 (N_2276,N_2099,N_2063);
and U2277 (N_2277,N_2090,N_2192);
and U2278 (N_2278,N_2084,N_2111);
nand U2279 (N_2279,N_2100,N_2025);
and U2280 (N_2280,N_2109,N_2199);
and U2281 (N_2281,N_2007,N_2158);
and U2282 (N_2282,N_2103,N_2124);
nand U2283 (N_2283,N_2123,N_2064);
and U2284 (N_2284,N_2122,N_2043);
or U2285 (N_2285,N_2050,N_2049);
and U2286 (N_2286,N_2159,N_2033);
nand U2287 (N_2287,N_2179,N_2196);
nor U2288 (N_2288,N_2058,N_2044);
nand U2289 (N_2289,N_2027,N_2039);
xnor U2290 (N_2290,N_2116,N_2052);
nor U2291 (N_2291,N_2188,N_2194);
nor U2292 (N_2292,N_2187,N_2079);
or U2293 (N_2293,N_2035,N_2118);
nand U2294 (N_2294,N_2087,N_2021);
nor U2295 (N_2295,N_2164,N_2152);
and U2296 (N_2296,N_2185,N_2078);
or U2297 (N_2297,N_2119,N_2020);
and U2298 (N_2298,N_2080,N_2154);
or U2299 (N_2299,N_2031,N_2054);
and U2300 (N_2300,N_2138,N_2194);
nand U2301 (N_2301,N_2009,N_2103);
and U2302 (N_2302,N_2030,N_2095);
nor U2303 (N_2303,N_2146,N_2155);
or U2304 (N_2304,N_2009,N_2049);
nand U2305 (N_2305,N_2084,N_2133);
and U2306 (N_2306,N_2064,N_2063);
nand U2307 (N_2307,N_2194,N_2095);
xor U2308 (N_2308,N_2103,N_2104);
xnor U2309 (N_2309,N_2139,N_2046);
nor U2310 (N_2310,N_2124,N_2036);
and U2311 (N_2311,N_2033,N_2154);
and U2312 (N_2312,N_2099,N_2082);
xor U2313 (N_2313,N_2070,N_2183);
nor U2314 (N_2314,N_2117,N_2049);
nand U2315 (N_2315,N_2170,N_2011);
nand U2316 (N_2316,N_2015,N_2070);
and U2317 (N_2317,N_2151,N_2098);
and U2318 (N_2318,N_2109,N_2104);
nor U2319 (N_2319,N_2055,N_2172);
and U2320 (N_2320,N_2177,N_2151);
nor U2321 (N_2321,N_2079,N_2134);
nor U2322 (N_2322,N_2065,N_2127);
and U2323 (N_2323,N_2059,N_2073);
xor U2324 (N_2324,N_2045,N_2124);
nand U2325 (N_2325,N_2005,N_2085);
and U2326 (N_2326,N_2075,N_2125);
and U2327 (N_2327,N_2060,N_2190);
nor U2328 (N_2328,N_2116,N_2037);
nand U2329 (N_2329,N_2142,N_2089);
xnor U2330 (N_2330,N_2017,N_2081);
nand U2331 (N_2331,N_2115,N_2005);
nor U2332 (N_2332,N_2142,N_2100);
nor U2333 (N_2333,N_2114,N_2131);
nand U2334 (N_2334,N_2097,N_2100);
nand U2335 (N_2335,N_2148,N_2179);
nor U2336 (N_2336,N_2147,N_2065);
nand U2337 (N_2337,N_2032,N_2093);
or U2338 (N_2338,N_2170,N_2032);
or U2339 (N_2339,N_2036,N_2105);
nand U2340 (N_2340,N_2159,N_2009);
xor U2341 (N_2341,N_2111,N_2132);
xor U2342 (N_2342,N_2169,N_2050);
nand U2343 (N_2343,N_2057,N_2191);
and U2344 (N_2344,N_2136,N_2085);
xor U2345 (N_2345,N_2092,N_2169);
and U2346 (N_2346,N_2081,N_2167);
nand U2347 (N_2347,N_2100,N_2076);
or U2348 (N_2348,N_2111,N_2115);
and U2349 (N_2349,N_2169,N_2091);
or U2350 (N_2350,N_2067,N_2135);
xor U2351 (N_2351,N_2060,N_2184);
nor U2352 (N_2352,N_2100,N_2050);
nand U2353 (N_2353,N_2134,N_2108);
and U2354 (N_2354,N_2094,N_2020);
nand U2355 (N_2355,N_2126,N_2098);
or U2356 (N_2356,N_2044,N_2163);
or U2357 (N_2357,N_2129,N_2012);
or U2358 (N_2358,N_2066,N_2196);
nand U2359 (N_2359,N_2124,N_2052);
xor U2360 (N_2360,N_2151,N_2165);
and U2361 (N_2361,N_2071,N_2054);
or U2362 (N_2362,N_2163,N_2042);
nand U2363 (N_2363,N_2191,N_2148);
and U2364 (N_2364,N_2152,N_2157);
nor U2365 (N_2365,N_2035,N_2092);
nand U2366 (N_2366,N_2041,N_2023);
nor U2367 (N_2367,N_2015,N_2180);
nand U2368 (N_2368,N_2159,N_2028);
or U2369 (N_2369,N_2161,N_2090);
nor U2370 (N_2370,N_2053,N_2049);
and U2371 (N_2371,N_2110,N_2093);
nor U2372 (N_2372,N_2042,N_2034);
xor U2373 (N_2373,N_2012,N_2024);
or U2374 (N_2374,N_2081,N_2179);
nand U2375 (N_2375,N_2057,N_2190);
nor U2376 (N_2376,N_2110,N_2030);
or U2377 (N_2377,N_2177,N_2069);
nand U2378 (N_2378,N_2170,N_2145);
nand U2379 (N_2379,N_2190,N_2005);
or U2380 (N_2380,N_2168,N_2125);
or U2381 (N_2381,N_2191,N_2042);
and U2382 (N_2382,N_2044,N_2013);
nor U2383 (N_2383,N_2136,N_2078);
nor U2384 (N_2384,N_2014,N_2052);
or U2385 (N_2385,N_2011,N_2167);
and U2386 (N_2386,N_2189,N_2193);
nor U2387 (N_2387,N_2084,N_2015);
and U2388 (N_2388,N_2188,N_2161);
nor U2389 (N_2389,N_2055,N_2199);
nand U2390 (N_2390,N_2041,N_2058);
or U2391 (N_2391,N_2179,N_2067);
nor U2392 (N_2392,N_2140,N_2125);
xnor U2393 (N_2393,N_2028,N_2061);
and U2394 (N_2394,N_2082,N_2024);
and U2395 (N_2395,N_2163,N_2132);
or U2396 (N_2396,N_2085,N_2051);
nand U2397 (N_2397,N_2163,N_2009);
nor U2398 (N_2398,N_2021,N_2003);
and U2399 (N_2399,N_2094,N_2136);
nor U2400 (N_2400,N_2253,N_2255);
nor U2401 (N_2401,N_2284,N_2261);
nand U2402 (N_2402,N_2297,N_2285);
and U2403 (N_2403,N_2264,N_2306);
nor U2404 (N_2404,N_2397,N_2211);
and U2405 (N_2405,N_2218,N_2357);
and U2406 (N_2406,N_2250,N_2200);
nor U2407 (N_2407,N_2299,N_2335);
nor U2408 (N_2408,N_2302,N_2392);
and U2409 (N_2409,N_2203,N_2311);
or U2410 (N_2410,N_2230,N_2280);
and U2411 (N_2411,N_2377,N_2294);
nand U2412 (N_2412,N_2269,N_2224);
nand U2413 (N_2413,N_2214,N_2365);
or U2414 (N_2414,N_2229,N_2221);
or U2415 (N_2415,N_2304,N_2216);
nor U2416 (N_2416,N_2205,N_2395);
nand U2417 (N_2417,N_2346,N_2271);
xor U2418 (N_2418,N_2345,N_2359);
xor U2419 (N_2419,N_2265,N_2301);
nor U2420 (N_2420,N_2233,N_2303);
nor U2421 (N_2421,N_2333,N_2223);
nand U2422 (N_2422,N_2393,N_2246);
nor U2423 (N_2423,N_2351,N_2226);
and U2424 (N_2424,N_2344,N_2360);
nor U2425 (N_2425,N_2252,N_2307);
xnor U2426 (N_2426,N_2249,N_2212);
xnor U2427 (N_2427,N_2352,N_2355);
nand U2428 (N_2428,N_2277,N_2368);
or U2429 (N_2429,N_2347,N_2381);
or U2430 (N_2430,N_2309,N_2283);
nand U2431 (N_2431,N_2362,N_2275);
nor U2432 (N_2432,N_2279,N_2206);
nand U2433 (N_2433,N_2259,N_2262);
or U2434 (N_2434,N_2213,N_2263);
nand U2435 (N_2435,N_2353,N_2322);
or U2436 (N_2436,N_2289,N_2228);
nand U2437 (N_2437,N_2243,N_2260);
nor U2438 (N_2438,N_2256,N_2308);
nor U2439 (N_2439,N_2232,N_2274);
nand U2440 (N_2440,N_2323,N_2376);
nor U2441 (N_2441,N_2325,N_2340);
or U2442 (N_2442,N_2241,N_2286);
nand U2443 (N_2443,N_2349,N_2358);
nor U2444 (N_2444,N_2379,N_2296);
nand U2445 (N_2445,N_2372,N_2219);
nand U2446 (N_2446,N_2231,N_2394);
xor U2447 (N_2447,N_2399,N_2317);
or U2448 (N_2448,N_2316,N_2375);
and U2449 (N_2449,N_2204,N_2338);
and U2450 (N_2450,N_2348,N_2278);
nand U2451 (N_2451,N_2290,N_2273);
or U2452 (N_2452,N_2398,N_2364);
nor U2453 (N_2453,N_2383,N_2324);
nand U2454 (N_2454,N_2371,N_2209);
nor U2455 (N_2455,N_2374,N_2287);
nor U2456 (N_2456,N_2390,N_2272);
or U2457 (N_2457,N_2326,N_2356);
nor U2458 (N_2458,N_2339,N_2334);
nor U2459 (N_2459,N_2244,N_2282);
xor U2460 (N_2460,N_2288,N_2373);
nand U2461 (N_2461,N_2267,N_2291);
nor U2462 (N_2462,N_2292,N_2378);
nand U2463 (N_2463,N_2266,N_2336);
and U2464 (N_2464,N_2391,N_2328);
nor U2465 (N_2465,N_2254,N_2210);
and U2466 (N_2466,N_2202,N_2320);
nand U2467 (N_2467,N_2248,N_2208);
nor U2468 (N_2468,N_2350,N_2367);
nand U2469 (N_2469,N_2319,N_2315);
nor U2470 (N_2470,N_2380,N_2235);
nor U2471 (N_2471,N_2295,N_2268);
nor U2472 (N_2472,N_2215,N_2329);
or U2473 (N_2473,N_2236,N_2201);
and U2474 (N_2474,N_2220,N_2369);
nand U2475 (N_2475,N_2207,N_2388);
nor U2476 (N_2476,N_2363,N_2217);
or U2477 (N_2477,N_2354,N_2240);
xor U2478 (N_2478,N_2396,N_2343);
and U2479 (N_2479,N_2258,N_2242);
nand U2480 (N_2480,N_2298,N_2222);
and U2481 (N_2481,N_2300,N_2321);
and U2482 (N_2482,N_2239,N_2389);
nand U2483 (N_2483,N_2245,N_2247);
and U2484 (N_2484,N_2342,N_2225);
or U2485 (N_2485,N_2387,N_2330);
nand U2486 (N_2486,N_2234,N_2331);
and U2487 (N_2487,N_2293,N_2337);
nor U2488 (N_2488,N_2251,N_2327);
and U2489 (N_2489,N_2237,N_2238);
or U2490 (N_2490,N_2270,N_2382);
xnor U2491 (N_2491,N_2305,N_2227);
nand U2492 (N_2492,N_2281,N_2386);
nand U2493 (N_2493,N_2366,N_2385);
and U2494 (N_2494,N_2384,N_2341);
or U2495 (N_2495,N_2310,N_2314);
nor U2496 (N_2496,N_2276,N_2257);
nor U2497 (N_2497,N_2318,N_2312);
nand U2498 (N_2498,N_2361,N_2313);
or U2499 (N_2499,N_2332,N_2370);
and U2500 (N_2500,N_2364,N_2279);
xnor U2501 (N_2501,N_2209,N_2375);
nor U2502 (N_2502,N_2276,N_2308);
and U2503 (N_2503,N_2234,N_2307);
nand U2504 (N_2504,N_2261,N_2294);
or U2505 (N_2505,N_2278,N_2286);
xor U2506 (N_2506,N_2305,N_2385);
nand U2507 (N_2507,N_2396,N_2232);
nor U2508 (N_2508,N_2224,N_2344);
and U2509 (N_2509,N_2335,N_2230);
nor U2510 (N_2510,N_2215,N_2292);
or U2511 (N_2511,N_2297,N_2374);
nand U2512 (N_2512,N_2289,N_2214);
xor U2513 (N_2513,N_2364,N_2349);
and U2514 (N_2514,N_2221,N_2344);
or U2515 (N_2515,N_2297,N_2223);
nand U2516 (N_2516,N_2363,N_2232);
and U2517 (N_2517,N_2284,N_2210);
nor U2518 (N_2518,N_2363,N_2242);
xor U2519 (N_2519,N_2259,N_2337);
nand U2520 (N_2520,N_2232,N_2203);
nand U2521 (N_2521,N_2378,N_2231);
nand U2522 (N_2522,N_2221,N_2366);
nand U2523 (N_2523,N_2220,N_2293);
xnor U2524 (N_2524,N_2319,N_2357);
xor U2525 (N_2525,N_2299,N_2249);
and U2526 (N_2526,N_2395,N_2240);
and U2527 (N_2527,N_2378,N_2204);
nand U2528 (N_2528,N_2333,N_2377);
or U2529 (N_2529,N_2354,N_2217);
and U2530 (N_2530,N_2220,N_2392);
nand U2531 (N_2531,N_2288,N_2349);
nor U2532 (N_2532,N_2270,N_2301);
nor U2533 (N_2533,N_2298,N_2380);
nand U2534 (N_2534,N_2358,N_2210);
or U2535 (N_2535,N_2223,N_2248);
and U2536 (N_2536,N_2321,N_2350);
nor U2537 (N_2537,N_2351,N_2306);
and U2538 (N_2538,N_2308,N_2200);
or U2539 (N_2539,N_2356,N_2395);
nand U2540 (N_2540,N_2272,N_2378);
or U2541 (N_2541,N_2305,N_2201);
and U2542 (N_2542,N_2263,N_2278);
and U2543 (N_2543,N_2299,N_2393);
nand U2544 (N_2544,N_2327,N_2254);
nand U2545 (N_2545,N_2263,N_2297);
nor U2546 (N_2546,N_2319,N_2327);
or U2547 (N_2547,N_2218,N_2332);
or U2548 (N_2548,N_2304,N_2366);
and U2549 (N_2549,N_2328,N_2269);
nor U2550 (N_2550,N_2338,N_2247);
and U2551 (N_2551,N_2347,N_2264);
and U2552 (N_2552,N_2283,N_2319);
nand U2553 (N_2553,N_2322,N_2236);
nor U2554 (N_2554,N_2205,N_2211);
nand U2555 (N_2555,N_2292,N_2357);
xor U2556 (N_2556,N_2223,N_2219);
nor U2557 (N_2557,N_2300,N_2222);
nor U2558 (N_2558,N_2320,N_2251);
and U2559 (N_2559,N_2224,N_2270);
xnor U2560 (N_2560,N_2349,N_2313);
or U2561 (N_2561,N_2283,N_2313);
or U2562 (N_2562,N_2254,N_2332);
or U2563 (N_2563,N_2380,N_2319);
or U2564 (N_2564,N_2325,N_2269);
and U2565 (N_2565,N_2280,N_2274);
nor U2566 (N_2566,N_2354,N_2256);
or U2567 (N_2567,N_2294,N_2306);
and U2568 (N_2568,N_2391,N_2320);
and U2569 (N_2569,N_2220,N_2274);
nor U2570 (N_2570,N_2297,N_2392);
and U2571 (N_2571,N_2220,N_2216);
or U2572 (N_2572,N_2331,N_2397);
or U2573 (N_2573,N_2324,N_2202);
or U2574 (N_2574,N_2236,N_2356);
nand U2575 (N_2575,N_2348,N_2205);
nor U2576 (N_2576,N_2325,N_2332);
nor U2577 (N_2577,N_2225,N_2363);
xor U2578 (N_2578,N_2343,N_2212);
and U2579 (N_2579,N_2336,N_2243);
nand U2580 (N_2580,N_2350,N_2392);
and U2581 (N_2581,N_2247,N_2241);
or U2582 (N_2582,N_2397,N_2275);
and U2583 (N_2583,N_2214,N_2357);
nor U2584 (N_2584,N_2234,N_2384);
nand U2585 (N_2585,N_2350,N_2270);
and U2586 (N_2586,N_2341,N_2213);
nor U2587 (N_2587,N_2278,N_2200);
nor U2588 (N_2588,N_2230,N_2265);
or U2589 (N_2589,N_2347,N_2353);
or U2590 (N_2590,N_2235,N_2243);
and U2591 (N_2591,N_2236,N_2376);
nor U2592 (N_2592,N_2338,N_2283);
or U2593 (N_2593,N_2220,N_2384);
nor U2594 (N_2594,N_2392,N_2253);
or U2595 (N_2595,N_2230,N_2296);
and U2596 (N_2596,N_2235,N_2314);
nand U2597 (N_2597,N_2346,N_2334);
or U2598 (N_2598,N_2208,N_2300);
nand U2599 (N_2599,N_2380,N_2255);
xor U2600 (N_2600,N_2515,N_2486);
xnor U2601 (N_2601,N_2428,N_2512);
nand U2602 (N_2602,N_2415,N_2470);
or U2603 (N_2603,N_2524,N_2536);
or U2604 (N_2604,N_2432,N_2410);
and U2605 (N_2605,N_2584,N_2566);
and U2606 (N_2606,N_2438,N_2561);
xnor U2607 (N_2607,N_2416,N_2436);
xor U2608 (N_2608,N_2586,N_2429);
nor U2609 (N_2609,N_2417,N_2533);
xor U2610 (N_2610,N_2419,N_2479);
and U2611 (N_2611,N_2402,N_2505);
and U2612 (N_2612,N_2459,N_2591);
nand U2613 (N_2613,N_2472,N_2597);
nor U2614 (N_2614,N_2446,N_2593);
and U2615 (N_2615,N_2458,N_2526);
nand U2616 (N_2616,N_2480,N_2498);
and U2617 (N_2617,N_2504,N_2590);
or U2618 (N_2618,N_2453,N_2581);
xnor U2619 (N_2619,N_2406,N_2457);
nand U2620 (N_2620,N_2563,N_2440);
and U2621 (N_2621,N_2476,N_2535);
xnor U2622 (N_2622,N_2468,N_2525);
nor U2623 (N_2623,N_2587,N_2595);
nor U2624 (N_2624,N_2585,N_2451);
and U2625 (N_2625,N_2541,N_2449);
nand U2626 (N_2626,N_2576,N_2464);
or U2627 (N_2627,N_2471,N_2484);
nand U2628 (N_2628,N_2510,N_2425);
xor U2629 (N_2629,N_2599,N_2488);
nand U2630 (N_2630,N_2475,N_2528);
or U2631 (N_2631,N_2434,N_2569);
xnor U2632 (N_2632,N_2575,N_2435);
and U2633 (N_2633,N_2550,N_2572);
nand U2634 (N_2634,N_2592,N_2431);
and U2635 (N_2635,N_2496,N_2534);
and U2636 (N_2636,N_2495,N_2404);
and U2637 (N_2637,N_2422,N_2439);
or U2638 (N_2638,N_2571,N_2527);
or U2639 (N_2639,N_2430,N_2529);
nor U2640 (N_2640,N_2433,N_2481);
and U2641 (N_2641,N_2461,N_2570);
nor U2642 (N_2642,N_2426,N_2447);
or U2643 (N_2643,N_2483,N_2482);
xnor U2644 (N_2644,N_2588,N_2560);
nand U2645 (N_2645,N_2567,N_2448);
nor U2646 (N_2646,N_2474,N_2409);
or U2647 (N_2647,N_2580,N_2582);
nand U2648 (N_2648,N_2564,N_2478);
nor U2649 (N_2649,N_2543,N_2418);
xnor U2650 (N_2650,N_2531,N_2462);
nand U2651 (N_2651,N_2513,N_2443);
or U2652 (N_2652,N_2518,N_2562);
nand U2653 (N_2653,N_2509,N_2424);
xor U2654 (N_2654,N_2460,N_2540);
nor U2655 (N_2655,N_2491,N_2530);
and U2656 (N_2656,N_2423,N_2452);
nand U2657 (N_2657,N_2493,N_2594);
nor U2658 (N_2658,N_2412,N_2532);
nand U2659 (N_2659,N_2538,N_2455);
or U2660 (N_2660,N_2552,N_2517);
or U2661 (N_2661,N_2401,N_2573);
nand U2662 (N_2662,N_2492,N_2554);
nor U2663 (N_2663,N_2542,N_2544);
nor U2664 (N_2664,N_2500,N_2467);
xor U2665 (N_2665,N_2520,N_2477);
nand U2666 (N_2666,N_2523,N_2579);
or U2667 (N_2667,N_2485,N_2403);
nor U2668 (N_2668,N_2547,N_2441);
or U2669 (N_2669,N_2568,N_2413);
nor U2670 (N_2670,N_2508,N_2420);
and U2671 (N_2671,N_2549,N_2589);
or U2672 (N_2672,N_2414,N_2450);
xor U2673 (N_2673,N_2522,N_2565);
nand U2674 (N_2674,N_2521,N_2411);
or U2675 (N_2675,N_2465,N_2499);
nor U2676 (N_2676,N_2489,N_2559);
and U2677 (N_2677,N_2407,N_2514);
or U2678 (N_2678,N_2545,N_2553);
and U2679 (N_2679,N_2574,N_2506);
or U2680 (N_2680,N_2405,N_2583);
xor U2681 (N_2681,N_2557,N_2442);
nand U2682 (N_2682,N_2511,N_2539);
nand U2683 (N_2683,N_2445,N_2537);
or U2684 (N_2684,N_2494,N_2558);
nor U2685 (N_2685,N_2556,N_2487);
nor U2686 (N_2686,N_2497,N_2473);
nor U2687 (N_2687,N_2503,N_2437);
nand U2688 (N_2688,N_2466,N_2501);
or U2689 (N_2689,N_2519,N_2555);
xnor U2690 (N_2690,N_2516,N_2546);
nand U2691 (N_2691,N_2507,N_2548);
nor U2692 (N_2692,N_2502,N_2400);
and U2693 (N_2693,N_2463,N_2454);
and U2694 (N_2694,N_2578,N_2456);
nand U2695 (N_2695,N_2444,N_2421);
nor U2696 (N_2696,N_2408,N_2577);
or U2697 (N_2697,N_2596,N_2490);
nand U2698 (N_2698,N_2427,N_2551);
nand U2699 (N_2699,N_2469,N_2598);
and U2700 (N_2700,N_2449,N_2533);
nor U2701 (N_2701,N_2583,N_2584);
nor U2702 (N_2702,N_2562,N_2461);
or U2703 (N_2703,N_2566,N_2491);
or U2704 (N_2704,N_2556,N_2563);
nor U2705 (N_2705,N_2566,N_2423);
nor U2706 (N_2706,N_2506,N_2434);
xnor U2707 (N_2707,N_2426,N_2527);
nand U2708 (N_2708,N_2433,N_2536);
nand U2709 (N_2709,N_2474,N_2587);
and U2710 (N_2710,N_2581,N_2459);
and U2711 (N_2711,N_2564,N_2593);
nor U2712 (N_2712,N_2502,N_2497);
nor U2713 (N_2713,N_2510,N_2537);
xor U2714 (N_2714,N_2408,N_2483);
xor U2715 (N_2715,N_2520,N_2470);
nor U2716 (N_2716,N_2432,N_2428);
and U2717 (N_2717,N_2595,N_2506);
nor U2718 (N_2718,N_2517,N_2576);
or U2719 (N_2719,N_2496,N_2527);
and U2720 (N_2720,N_2501,N_2441);
nor U2721 (N_2721,N_2408,N_2511);
xnor U2722 (N_2722,N_2479,N_2548);
xnor U2723 (N_2723,N_2513,N_2560);
and U2724 (N_2724,N_2507,N_2429);
nor U2725 (N_2725,N_2538,N_2596);
nand U2726 (N_2726,N_2576,N_2527);
or U2727 (N_2727,N_2573,N_2415);
nor U2728 (N_2728,N_2598,N_2468);
nand U2729 (N_2729,N_2495,N_2430);
nand U2730 (N_2730,N_2420,N_2569);
and U2731 (N_2731,N_2488,N_2573);
nand U2732 (N_2732,N_2428,N_2537);
and U2733 (N_2733,N_2556,N_2525);
nor U2734 (N_2734,N_2421,N_2522);
xor U2735 (N_2735,N_2478,N_2544);
nand U2736 (N_2736,N_2454,N_2573);
nor U2737 (N_2737,N_2453,N_2480);
and U2738 (N_2738,N_2524,N_2558);
nand U2739 (N_2739,N_2439,N_2468);
nor U2740 (N_2740,N_2588,N_2407);
nor U2741 (N_2741,N_2475,N_2510);
nand U2742 (N_2742,N_2527,N_2588);
nor U2743 (N_2743,N_2583,N_2449);
and U2744 (N_2744,N_2550,N_2548);
nand U2745 (N_2745,N_2454,N_2583);
or U2746 (N_2746,N_2500,N_2579);
nor U2747 (N_2747,N_2510,N_2428);
nand U2748 (N_2748,N_2566,N_2430);
nand U2749 (N_2749,N_2496,N_2521);
nand U2750 (N_2750,N_2541,N_2585);
or U2751 (N_2751,N_2580,N_2424);
nand U2752 (N_2752,N_2440,N_2503);
or U2753 (N_2753,N_2575,N_2440);
nand U2754 (N_2754,N_2513,N_2561);
nand U2755 (N_2755,N_2560,N_2494);
nor U2756 (N_2756,N_2548,N_2411);
nor U2757 (N_2757,N_2460,N_2532);
or U2758 (N_2758,N_2485,N_2529);
or U2759 (N_2759,N_2423,N_2425);
nand U2760 (N_2760,N_2550,N_2405);
and U2761 (N_2761,N_2536,N_2489);
nand U2762 (N_2762,N_2535,N_2589);
and U2763 (N_2763,N_2493,N_2410);
nand U2764 (N_2764,N_2570,N_2470);
or U2765 (N_2765,N_2514,N_2438);
nor U2766 (N_2766,N_2533,N_2494);
and U2767 (N_2767,N_2440,N_2407);
nand U2768 (N_2768,N_2573,N_2570);
and U2769 (N_2769,N_2522,N_2404);
nor U2770 (N_2770,N_2503,N_2571);
nand U2771 (N_2771,N_2529,N_2535);
xnor U2772 (N_2772,N_2447,N_2559);
and U2773 (N_2773,N_2414,N_2580);
or U2774 (N_2774,N_2528,N_2510);
nand U2775 (N_2775,N_2576,N_2450);
nand U2776 (N_2776,N_2539,N_2559);
nor U2777 (N_2777,N_2568,N_2444);
or U2778 (N_2778,N_2570,N_2511);
xnor U2779 (N_2779,N_2411,N_2559);
or U2780 (N_2780,N_2597,N_2557);
or U2781 (N_2781,N_2523,N_2402);
nor U2782 (N_2782,N_2496,N_2573);
nor U2783 (N_2783,N_2573,N_2472);
nor U2784 (N_2784,N_2497,N_2525);
nor U2785 (N_2785,N_2555,N_2459);
nor U2786 (N_2786,N_2412,N_2451);
xor U2787 (N_2787,N_2576,N_2547);
nand U2788 (N_2788,N_2553,N_2527);
or U2789 (N_2789,N_2455,N_2451);
and U2790 (N_2790,N_2501,N_2563);
nor U2791 (N_2791,N_2464,N_2487);
and U2792 (N_2792,N_2527,N_2506);
nand U2793 (N_2793,N_2448,N_2495);
and U2794 (N_2794,N_2520,N_2435);
and U2795 (N_2795,N_2533,N_2570);
nor U2796 (N_2796,N_2573,N_2563);
and U2797 (N_2797,N_2458,N_2482);
xor U2798 (N_2798,N_2407,N_2592);
and U2799 (N_2799,N_2434,N_2448);
or U2800 (N_2800,N_2732,N_2757);
xor U2801 (N_2801,N_2781,N_2796);
and U2802 (N_2802,N_2655,N_2669);
nor U2803 (N_2803,N_2638,N_2612);
xnor U2804 (N_2804,N_2738,N_2728);
or U2805 (N_2805,N_2798,N_2767);
and U2806 (N_2806,N_2793,N_2659);
and U2807 (N_2807,N_2689,N_2666);
or U2808 (N_2808,N_2733,N_2622);
and U2809 (N_2809,N_2663,N_2606);
nor U2810 (N_2810,N_2644,N_2610);
or U2811 (N_2811,N_2681,N_2656);
or U2812 (N_2812,N_2660,N_2640);
nor U2813 (N_2813,N_2672,N_2706);
nor U2814 (N_2814,N_2772,N_2770);
nand U2815 (N_2815,N_2671,N_2741);
nor U2816 (N_2816,N_2698,N_2619);
and U2817 (N_2817,N_2694,N_2712);
and U2818 (N_2818,N_2608,N_2740);
nor U2819 (N_2819,N_2686,N_2683);
and U2820 (N_2820,N_2613,N_2784);
xnor U2821 (N_2821,N_2618,N_2667);
and U2822 (N_2822,N_2773,N_2760);
or U2823 (N_2823,N_2725,N_2739);
xor U2824 (N_2824,N_2790,N_2684);
nand U2825 (N_2825,N_2752,N_2748);
nor U2826 (N_2826,N_2641,N_2720);
nor U2827 (N_2827,N_2670,N_2652);
nor U2828 (N_2828,N_2701,N_2677);
xor U2829 (N_2829,N_2727,N_2674);
or U2830 (N_2830,N_2782,N_2629);
or U2831 (N_2831,N_2620,N_2768);
nand U2832 (N_2832,N_2799,N_2704);
or U2833 (N_2833,N_2700,N_2614);
nor U2834 (N_2834,N_2717,N_2697);
or U2835 (N_2835,N_2662,N_2688);
nand U2836 (N_2836,N_2664,N_2765);
and U2837 (N_2837,N_2616,N_2621);
or U2838 (N_2838,N_2676,N_2635);
nand U2839 (N_2839,N_2682,N_2795);
nor U2840 (N_2840,N_2630,N_2731);
and U2841 (N_2841,N_2719,N_2746);
and U2842 (N_2842,N_2705,N_2699);
and U2843 (N_2843,N_2787,N_2771);
nor U2844 (N_2844,N_2714,N_2661);
nor U2845 (N_2845,N_2753,N_2749);
or U2846 (N_2846,N_2665,N_2774);
nand U2847 (N_2847,N_2736,N_2775);
nor U2848 (N_2848,N_2791,N_2650);
xor U2849 (N_2849,N_2716,N_2611);
or U2850 (N_2850,N_2709,N_2762);
nand U2851 (N_2851,N_2668,N_2600);
xnor U2852 (N_2852,N_2657,N_2678);
or U2853 (N_2853,N_2624,N_2627);
and U2854 (N_2854,N_2761,N_2722);
nor U2855 (N_2855,N_2754,N_2715);
xor U2856 (N_2856,N_2785,N_2637);
and U2857 (N_2857,N_2713,N_2744);
nor U2858 (N_2858,N_2797,N_2685);
nand U2859 (N_2859,N_2696,N_2605);
nand U2860 (N_2860,N_2609,N_2632);
nand U2861 (N_2861,N_2648,N_2778);
xor U2862 (N_2862,N_2623,N_2690);
or U2863 (N_2863,N_2658,N_2747);
and U2864 (N_2864,N_2711,N_2737);
and U2865 (N_2865,N_2708,N_2607);
xnor U2866 (N_2866,N_2789,N_2634);
nor U2867 (N_2867,N_2691,N_2631);
nor U2868 (N_2868,N_2653,N_2729);
nand U2869 (N_2869,N_2603,N_2675);
nand U2870 (N_2870,N_2724,N_2792);
xor U2871 (N_2871,N_2602,N_2764);
nor U2872 (N_2872,N_2750,N_2766);
and U2873 (N_2873,N_2643,N_2654);
xnor U2874 (N_2874,N_2751,N_2794);
nand U2875 (N_2875,N_2625,N_2687);
nand U2876 (N_2876,N_2642,N_2718);
nand U2877 (N_2877,N_2645,N_2601);
nor U2878 (N_2878,N_2692,N_2626);
xor U2879 (N_2879,N_2759,N_2649);
xnor U2880 (N_2880,N_2723,N_2769);
nand U2881 (N_2881,N_2779,N_2758);
nor U2882 (N_2882,N_2745,N_2628);
nor U2883 (N_2883,N_2673,N_2763);
xnor U2884 (N_2884,N_2617,N_2735);
nand U2885 (N_2885,N_2703,N_2647);
and U2886 (N_2886,N_2646,N_2604);
and U2887 (N_2887,N_2783,N_2742);
and U2888 (N_2888,N_2780,N_2743);
and U2889 (N_2889,N_2786,N_2695);
and U2890 (N_2890,N_2730,N_2777);
or U2891 (N_2891,N_2636,N_2755);
and U2892 (N_2892,N_2721,N_2756);
and U2893 (N_2893,N_2639,N_2788);
nor U2894 (N_2894,N_2615,N_2651);
and U2895 (N_2895,N_2702,N_2680);
and U2896 (N_2896,N_2693,N_2679);
nor U2897 (N_2897,N_2707,N_2776);
or U2898 (N_2898,N_2633,N_2734);
nand U2899 (N_2899,N_2710,N_2726);
nand U2900 (N_2900,N_2722,N_2686);
and U2901 (N_2901,N_2614,N_2770);
or U2902 (N_2902,N_2739,N_2699);
or U2903 (N_2903,N_2684,N_2616);
xor U2904 (N_2904,N_2659,N_2611);
or U2905 (N_2905,N_2757,N_2717);
and U2906 (N_2906,N_2673,N_2771);
or U2907 (N_2907,N_2658,N_2644);
and U2908 (N_2908,N_2650,N_2753);
xnor U2909 (N_2909,N_2795,N_2654);
nand U2910 (N_2910,N_2645,N_2797);
nand U2911 (N_2911,N_2660,N_2618);
nor U2912 (N_2912,N_2652,N_2762);
nand U2913 (N_2913,N_2722,N_2663);
nor U2914 (N_2914,N_2761,N_2684);
nand U2915 (N_2915,N_2784,N_2799);
nand U2916 (N_2916,N_2664,N_2689);
xnor U2917 (N_2917,N_2748,N_2664);
or U2918 (N_2918,N_2686,N_2633);
or U2919 (N_2919,N_2776,N_2642);
or U2920 (N_2920,N_2604,N_2703);
nor U2921 (N_2921,N_2775,N_2711);
or U2922 (N_2922,N_2675,N_2798);
or U2923 (N_2923,N_2789,N_2786);
or U2924 (N_2924,N_2714,N_2664);
and U2925 (N_2925,N_2708,N_2608);
nand U2926 (N_2926,N_2601,N_2712);
nand U2927 (N_2927,N_2691,N_2633);
and U2928 (N_2928,N_2602,N_2666);
xor U2929 (N_2929,N_2673,N_2622);
and U2930 (N_2930,N_2676,N_2619);
nand U2931 (N_2931,N_2751,N_2739);
nand U2932 (N_2932,N_2722,N_2756);
and U2933 (N_2933,N_2765,N_2796);
and U2934 (N_2934,N_2674,N_2675);
nor U2935 (N_2935,N_2762,N_2732);
xor U2936 (N_2936,N_2650,N_2609);
nand U2937 (N_2937,N_2741,N_2676);
nor U2938 (N_2938,N_2656,N_2708);
and U2939 (N_2939,N_2756,N_2696);
and U2940 (N_2940,N_2661,N_2625);
nand U2941 (N_2941,N_2711,N_2688);
nor U2942 (N_2942,N_2727,N_2626);
or U2943 (N_2943,N_2666,N_2670);
and U2944 (N_2944,N_2765,N_2607);
and U2945 (N_2945,N_2735,N_2680);
nand U2946 (N_2946,N_2702,N_2717);
xnor U2947 (N_2947,N_2759,N_2730);
and U2948 (N_2948,N_2620,N_2794);
or U2949 (N_2949,N_2743,N_2765);
nor U2950 (N_2950,N_2685,N_2693);
and U2951 (N_2951,N_2752,N_2638);
and U2952 (N_2952,N_2745,N_2600);
nor U2953 (N_2953,N_2616,N_2754);
nor U2954 (N_2954,N_2696,N_2705);
nor U2955 (N_2955,N_2673,N_2736);
and U2956 (N_2956,N_2717,N_2737);
nand U2957 (N_2957,N_2799,N_2677);
nor U2958 (N_2958,N_2643,N_2689);
and U2959 (N_2959,N_2698,N_2743);
nand U2960 (N_2960,N_2696,N_2627);
nand U2961 (N_2961,N_2650,N_2621);
nor U2962 (N_2962,N_2682,N_2654);
nor U2963 (N_2963,N_2633,N_2775);
and U2964 (N_2964,N_2734,N_2765);
or U2965 (N_2965,N_2740,N_2706);
and U2966 (N_2966,N_2783,N_2692);
and U2967 (N_2967,N_2699,N_2731);
and U2968 (N_2968,N_2765,N_2676);
nand U2969 (N_2969,N_2698,N_2664);
xnor U2970 (N_2970,N_2613,N_2797);
and U2971 (N_2971,N_2760,N_2611);
nor U2972 (N_2972,N_2744,N_2786);
and U2973 (N_2973,N_2692,N_2696);
and U2974 (N_2974,N_2748,N_2709);
nand U2975 (N_2975,N_2699,N_2646);
nor U2976 (N_2976,N_2685,N_2790);
nand U2977 (N_2977,N_2689,N_2732);
and U2978 (N_2978,N_2620,N_2796);
nand U2979 (N_2979,N_2764,N_2737);
or U2980 (N_2980,N_2752,N_2701);
or U2981 (N_2981,N_2713,N_2730);
or U2982 (N_2982,N_2706,N_2622);
nor U2983 (N_2983,N_2722,N_2633);
and U2984 (N_2984,N_2690,N_2784);
and U2985 (N_2985,N_2760,N_2618);
nor U2986 (N_2986,N_2653,N_2667);
nor U2987 (N_2987,N_2660,N_2764);
and U2988 (N_2988,N_2731,N_2684);
and U2989 (N_2989,N_2757,N_2704);
or U2990 (N_2990,N_2746,N_2685);
nand U2991 (N_2991,N_2718,N_2721);
and U2992 (N_2992,N_2655,N_2651);
nor U2993 (N_2993,N_2646,N_2686);
nand U2994 (N_2994,N_2768,N_2799);
or U2995 (N_2995,N_2670,N_2752);
or U2996 (N_2996,N_2621,N_2637);
nand U2997 (N_2997,N_2728,N_2600);
xor U2998 (N_2998,N_2744,N_2649);
nand U2999 (N_2999,N_2644,N_2616);
xnor UO_0 (O_0,N_2942,N_2933);
and UO_1 (O_1,N_2856,N_2915);
nor UO_2 (O_2,N_2886,N_2957);
and UO_3 (O_3,N_2894,N_2917);
nand UO_4 (O_4,N_2919,N_2809);
nand UO_5 (O_5,N_2861,N_2891);
and UO_6 (O_6,N_2881,N_2863);
nand UO_7 (O_7,N_2975,N_2979);
nand UO_8 (O_8,N_2811,N_2876);
and UO_9 (O_9,N_2832,N_2938);
nand UO_10 (O_10,N_2946,N_2966);
nor UO_11 (O_11,N_2888,N_2914);
nand UO_12 (O_12,N_2995,N_2828);
nor UO_13 (O_13,N_2805,N_2867);
nand UO_14 (O_14,N_2997,N_2889);
or UO_15 (O_15,N_2978,N_2880);
nand UO_16 (O_16,N_2952,N_2922);
or UO_17 (O_17,N_2980,N_2926);
and UO_18 (O_18,N_2987,N_2836);
nand UO_19 (O_19,N_2847,N_2884);
xor UO_20 (O_20,N_2996,N_2857);
nor UO_21 (O_21,N_2815,N_2989);
and UO_22 (O_22,N_2974,N_2941);
nor UO_23 (O_23,N_2951,N_2993);
and UO_24 (O_24,N_2906,N_2920);
nand UO_25 (O_25,N_2913,N_2887);
and UO_26 (O_26,N_2969,N_2905);
nand UO_27 (O_27,N_2898,N_2877);
nor UO_28 (O_28,N_2949,N_2862);
nand UO_29 (O_29,N_2858,N_2967);
or UO_30 (O_30,N_2814,N_2934);
nand UO_31 (O_31,N_2936,N_2959);
and UO_32 (O_32,N_2945,N_2838);
nand UO_33 (O_33,N_2883,N_2866);
xnor UO_34 (O_34,N_2854,N_2879);
xor UO_35 (O_35,N_2924,N_2850);
nand UO_36 (O_36,N_2897,N_2970);
or UO_37 (O_37,N_2841,N_2872);
nand UO_38 (O_38,N_2901,N_2823);
and UO_39 (O_39,N_2868,N_2939);
nor UO_40 (O_40,N_2944,N_2827);
nor UO_41 (O_41,N_2929,N_2902);
nor UO_42 (O_42,N_2831,N_2983);
or UO_43 (O_43,N_2813,N_2981);
or UO_44 (O_44,N_2992,N_2928);
xor UO_45 (O_45,N_2892,N_2954);
and UO_46 (O_46,N_2882,N_2918);
and UO_47 (O_47,N_2953,N_2925);
or UO_48 (O_48,N_2912,N_2991);
nor UO_49 (O_49,N_2962,N_2986);
or UO_50 (O_50,N_2998,N_2835);
or UO_51 (O_51,N_2931,N_2916);
or UO_52 (O_52,N_2911,N_2808);
nand UO_53 (O_53,N_2890,N_2895);
and UO_54 (O_54,N_2830,N_2972);
nor UO_55 (O_55,N_2842,N_2825);
and UO_56 (O_56,N_2829,N_2803);
nand UO_57 (O_57,N_2904,N_2816);
xnor UO_58 (O_58,N_2955,N_2848);
and UO_59 (O_59,N_2930,N_2927);
nand UO_60 (O_60,N_2900,N_2818);
nand UO_61 (O_61,N_2982,N_2859);
xor UO_62 (O_62,N_2860,N_2965);
nand UO_63 (O_63,N_2864,N_2963);
or UO_64 (O_64,N_2851,N_2961);
xor UO_65 (O_65,N_2804,N_2819);
nand UO_66 (O_66,N_2923,N_2843);
nand UO_67 (O_67,N_2824,N_2869);
nor UO_68 (O_68,N_2806,N_2855);
or UO_69 (O_69,N_2846,N_2940);
and UO_70 (O_70,N_2849,N_2870);
and UO_71 (O_71,N_2985,N_2839);
nand UO_72 (O_72,N_2908,N_2874);
and UO_73 (O_73,N_2840,N_2935);
or UO_74 (O_74,N_2844,N_2826);
nand UO_75 (O_75,N_2921,N_2817);
xor UO_76 (O_76,N_2910,N_2976);
nor UO_77 (O_77,N_2833,N_2802);
or UO_78 (O_78,N_2973,N_2820);
nand UO_79 (O_79,N_2937,N_2812);
or UO_80 (O_80,N_2907,N_2834);
xnor UO_81 (O_81,N_2853,N_2932);
and UO_82 (O_82,N_2943,N_2971);
xor UO_83 (O_83,N_2873,N_2822);
and UO_84 (O_84,N_2960,N_2865);
and UO_85 (O_85,N_2990,N_2988);
and UO_86 (O_86,N_2999,N_2909);
xnor UO_87 (O_87,N_2837,N_2950);
or UO_88 (O_88,N_2968,N_2885);
nand UO_89 (O_89,N_2899,N_2807);
or UO_90 (O_90,N_2801,N_2903);
or UO_91 (O_91,N_2893,N_2994);
nand UO_92 (O_92,N_2896,N_2948);
nand UO_93 (O_93,N_2800,N_2977);
and UO_94 (O_94,N_2964,N_2956);
nand UO_95 (O_95,N_2878,N_2810);
nand UO_96 (O_96,N_2852,N_2871);
nand UO_97 (O_97,N_2821,N_2845);
nand UO_98 (O_98,N_2947,N_2875);
nor UO_99 (O_99,N_2984,N_2958);
nand UO_100 (O_100,N_2900,N_2909);
and UO_101 (O_101,N_2915,N_2983);
xnor UO_102 (O_102,N_2835,N_2975);
nand UO_103 (O_103,N_2892,N_2882);
and UO_104 (O_104,N_2801,N_2994);
xor UO_105 (O_105,N_2883,N_2916);
or UO_106 (O_106,N_2846,N_2814);
and UO_107 (O_107,N_2918,N_2810);
or UO_108 (O_108,N_2844,N_2934);
nand UO_109 (O_109,N_2833,N_2821);
nand UO_110 (O_110,N_2836,N_2880);
and UO_111 (O_111,N_2827,N_2817);
nor UO_112 (O_112,N_2889,N_2862);
and UO_113 (O_113,N_2976,N_2909);
nand UO_114 (O_114,N_2968,N_2848);
xor UO_115 (O_115,N_2944,N_2865);
xnor UO_116 (O_116,N_2811,N_2884);
and UO_117 (O_117,N_2971,N_2904);
or UO_118 (O_118,N_2897,N_2985);
nor UO_119 (O_119,N_2999,N_2885);
xnor UO_120 (O_120,N_2890,N_2894);
nand UO_121 (O_121,N_2953,N_2800);
nor UO_122 (O_122,N_2915,N_2961);
nand UO_123 (O_123,N_2960,N_2964);
or UO_124 (O_124,N_2816,N_2938);
nor UO_125 (O_125,N_2938,N_2927);
xor UO_126 (O_126,N_2865,N_2855);
nand UO_127 (O_127,N_2956,N_2950);
and UO_128 (O_128,N_2969,N_2966);
nand UO_129 (O_129,N_2952,N_2902);
or UO_130 (O_130,N_2810,N_2832);
or UO_131 (O_131,N_2813,N_2840);
nand UO_132 (O_132,N_2909,N_2807);
and UO_133 (O_133,N_2973,N_2919);
nand UO_134 (O_134,N_2812,N_2824);
xnor UO_135 (O_135,N_2965,N_2818);
nand UO_136 (O_136,N_2927,N_2849);
and UO_137 (O_137,N_2873,N_2858);
nand UO_138 (O_138,N_2954,N_2863);
xnor UO_139 (O_139,N_2932,N_2861);
xnor UO_140 (O_140,N_2920,N_2882);
nand UO_141 (O_141,N_2804,N_2956);
and UO_142 (O_142,N_2910,N_2833);
nand UO_143 (O_143,N_2975,N_2934);
xnor UO_144 (O_144,N_2917,N_2803);
and UO_145 (O_145,N_2838,N_2946);
and UO_146 (O_146,N_2863,N_2978);
nor UO_147 (O_147,N_2822,N_2811);
nor UO_148 (O_148,N_2866,N_2856);
nand UO_149 (O_149,N_2940,N_2976);
nand UO_150 (O_150,N_2880,N_2865);
or UO_151 (O_151,N_2968,N_2907);
nor UO_152 (O_152,N_2875,N_2953);
nor UO_153 (O_153,N_2828,N_2826);
nand UO_154 (O_154,N_2909,N_2942);
and UO_155 (O_155,N_2900,N_2843);
nor UO_156 (O_156,N_2960,N_2985);
and UO_157 (O_157,N_2998,N_2902);
xor UO_158 (O_158,N_2804,N_2875);
xnor UO_159 (O_159,N_2837,N_2947);
xor UO_160 (O_160,N_2815,N_2878);
nor UO_161 (O_161,N_2947,N_2857);
nand UO_162 (O_162,N_2957,N_2965);
nor UO_163 (O_163,N_2801,N_2982);
nand UO_164 (O_164,N_2999,N_2935);
or UO_165 (O_165,N_2984,N_2857);
nor UO_166 (O_166,N_2926,N_2832);
and UO_167 (O_167,N_2866,N_2877);
and UO_168 (O_168,N_2874,N_2937);
nand UO_169 (O_169,N_2838,N_2947);
or UO_170 (O_170,N_2901,N_2999);
or UO_171 (O_171,N_2815,N_2816);
and UO_172 (O_172,N_2992,N_2851);
nor UO_173 (O_173,N_2918,N_2821);
and UO_174 (O_174,N_2828,N_2923);
and UO_175 (O_175,N_2915,N_2889);
nor UO_176 (O_176,N_2996,N_2999);
nand UO_177 (O_177,N_2950,N_2924);
and UO_178 (O_178,N_2972,N_2896);
and UO_179 (O_179,N_2895,N_2806);
nor UO_180 (O_180,N_2941,N_2856);
xnor UO_181 (O_181,N_2927,N_2884);
or UO_182 (O_182,N_2937,N_2893);
or UO_183 (O_183,N_2877,N_2809);
nor UO_184 (O_184,N_2808,N_2994);
nor UO_185 (O_185,N_2818,N_2930);
and UO_186 (O_186,N_2962,N_2934);
nand UO_187 (O_187,N_2986,N_2841);
and UO_188 (O_188,N_2966,N_2843);
or UO_189 (O_189,N_2930,N_2951);
nor UO_190 (O_190,N_2850,N_2953);
and UO_191 (O_191,N_2991,N_2917);
and UO_192 (O_192,N_2924,N_2975);
nor UO_193 (O_193,N_2997,N_2841);
nand UO_194 (O_194,N_2948,N_2991);
nor UO_195 (O_195,N_2816,N_2834);
and UO_196 (O_196,N_2850,N_2819);
or UO_197 (O_197,N_2967,N_2943);
nor UO_198 (O_198,N_2828,N_2990);
nand UO_199 (O_199,N_2837,N_2971);
nand UO_200 (O_200,N_2873,N_2984);
nor UO_201 (O_201,N_2953,N_2993);
and UO_202 (O_202,N_2948,N_2980);
and UO_203 (O_203,N_2864,N_2941);
xor UO_204 (O_204,N_2885,N_2870);
and UO_205 (O_205,N_2844,N_2995);
or UO_206 (O_206,N_2925,N_2890);
nand UO_207 (O_207,N_2805,N_2865);
nor UO_208 (O_208,N_2964,N_2856);
and UO_209 (O_209,N_2948,N_2858);
nor UO_210 (O_210,N_2960,N_2892);
nand UO_211 (O_211,N_2940,N_2824);
and UO_212 (O_212,N_2915,N_2867);
xor UO_213 (O_213,N_2843,N_2868);
xor UO_214 (O_214,N_2853,N_2866);
xor UO_215 (O_215,N_2955,N_2972);
nor UO_216 (O_216,N_2937,N_2931);
and UO_217 (O_217,N_2996,N_2874);
nand UO_218 (O_218,N_2906,N_2977);
or UO_219 (O_219,N_2848,N_2967);
nor UO_220 (O_220,N_2850,N_2949);
and UO_221 (O_221,N_2917,N_2943);
or UO_222 (O_222,N_2957,N_2992);
nand UO_223 (O_223,N_2895,N_2802);
or UO_224 (O_224,N_2849,N_2824);
and UO_225 (O_225,N_2904,N_2837);
or UO_226 (O_226,N_2832,N_2878);
nor UO_227 (O_227,N_2970,N_2998);
or UO_228 (O_228,N_2998,N_2900);
nand UO_229 (O_229,N_2985,N_2801);
nor UO_230 (O_230,N_2810,N_2923);
nor UO_231 (O_231,N_2840,N_2812);
or UO_232 (O_232,N_2889,N_2933);
nand UO_233 (O_233,N_2933,N_2999);
and UO_234 (O_234,N_2890,N_2853);
and UO_235 (O_235,N_2904,N_2996);
and UO_236 (O_236,N_2812,N_2850);
and UO_237 (O_237,N_2979,N_2810);
nand UO_238 (O_238,N_2976,N_2854);
or UO_239 (O_239,N_2928,N_2934);
nor UO_240 (O_240,N_2852,N_2934);
and UO_241 (O_241,N_2985,N_2963);
nand UO_242 (O_242,N_2804,N_2910);
and UO_243 (O_243,N_2885,N_2912);
nand UO_244 (O_244,N_2971,N_2856);
and UO_245 (O_245,N_2861,N_2828);
nor UO_246 (O_246,N_2947,N_2940);
or UO_247 (O_247,N_2817,N_2911);
xnor UO_248 (O_248,N_2818,N_2814);
and UO_249 (O_249,N_2879,N_2958);
nor UO_250 (O_250,N_2982,N_2967);
or UO_251 (O_251,N_2843,N_2846);
nor UO_252 (O_252,N_2926,N_2995);
nand UO_253 (O_253,N_2948,N_2974);
nor UO_254 (O_254,N_2825,N_2953);
or UO_255 (O_255,N_2813,N_2873);
and UO_256 (O_256,N_2946,N_2924);
nor UO_257 (O_257,N_2802,N_2960);
nor UO_258 (O_258,N_2956,N_2851);
and UO_259 (O_259,N_2807,N_2824);
and UO_260 (O_260,N_2949,N_2829);
xor UO_261 (O_261,N_2909,N_2861);
xor UO_262 (O_262,N_2800,N_2814);
or UO_263 (O_263,N_2949,N_2803);
nor UO_264 (O_264,N_2845,N_2850);
xor UO_265 (O_265,N_2965,N_2855);
nor UO_266 (O_266,N_2843,N_2907);
xnor UO_267 (O_267,N_2844,N_2933);
or UO_268 (O_268,N_2916,N_2982);
and UO_269 (O_269,N_2984,N_2832);
or UO_270 (O_270,N_2883,N_2836);
or UO_271 (O_271,N_2874,N_2809);
nor UO_272 (O_272,N_2981,N_2926);
nor UO_273 (O_273,N_2819,N_2864);
nor UO_274 (O_274,N_2859,N_2987);
and UO_275 (O_275,N_2968,N_2864);
and UO_276 (O_276,N_2931,N_2820);
nor UO_277 (O_277,N_2841,N_2832);
nand UO_278 (O_278,N_2957,N_2858);
xor UO_279 (O_279,N_2832,N_2918);
nor UO_280 (O_280,N_2957,N_2802);
or UO_281 (O_281,N_2804,N_2995);
or UO_282 (O_282,N_2808,N_2918);
and UO_283 (O_283,N_2862,N_2882);
or UO_284 (O_284,N_2934,N_2988);
or UO_285 (O_285,N_2924,N_2897);
nand UO_286 (O_286,N_2947,N_2850);
or UO_287 (O_287,N_2965,N_2886);
and UO_288 (O_288,N_2879,N_2830);
xnor UO_289 (O_289,N_2938,N_2923);
or UO_290 (O_290,N_2913,N_2842);
and UO_291 (O_291,N_2999,N_2965);
nand UO_292 (O_292,N_2846,N_2904);
and UO_293 (O_293,N_2994,N_2957);
and UO_294 (O_294,N_2962,N_2928);
nor UO_295 (O_295,N_2852,N_2928);
or UO_296 (O_296,N_2824,N_2882);
nand UO_297 (O_297,N_2955,N_2999);
or UO_298 (O_298,N_2833,N_2806);
nand UO_299 (O_299,N_2916,N_2997);
and UO_300 (O_300,N_2986,N_2965);
nor UO_301 (O_301,N_2846,N_2942);
nand UO_302 (O_302,N_2961,N_2920);
xor UO_303 (O_303,N_2832,N_2968);
or UO_304 (O_304,N_2891,N_2855);
nor UO_305 (O_305,N_2920,N_2927);
nor UO_306 (O_306,N_2999,N_2840);
nand UO_307 (O_307,N_2904,N_2997);
or UO_308 (O_308,N_2826,N_2848);
and UO_309 (O_309,N_2815,N_2994);
nand UO_310 (O_310,N_2917,N_2845);
and UO_311 (O_311,N_2847,N_2874);
or UO_312 (O_312,N_2952,N_2914);
or UO_313 (O_313,N_2914,N_2921);
nand UO_314 (O_314,N_2870,N_2905);
nand UO_315 (O_315,N_2995,N_2881);
xor UO_316 (O_316,N_2971,N_2980);
xor UO_317 (O_317,N_2805,N_2888);
nand UO_318 (O_318,N_2916,N_2970);
and UO_319 (O_319,N_2889,N_2827);
xor UO_320 (O_320,N_2838,N_2902);
or UO_321 (O_321,N_2914,N_2989);
and UO_322 (O_322,N_2823,N_2845);
xnor UO_323 (O_323,N_2970,N_2892);
and UO_324 (O_324,N_2965,N_2951);
nor UO_325 (O_325,N_2920,N_2990);
nand UO_326 (O_326,N_2831,N_2869);
xor UO_327 (O_327,N_2920,N_2841);
or UO_328 (O_328,N_2836,N_2852);
nand UO_329 (O_329,N_2935,N_2866);
xnor UO_330 (O_330,N_2929,N_2832);
nand UO_331 (O_331,N_2941,N_2996);
nor UO_332 (O_332,N_2994,N_2852);
nor UO_333 (O_333,N_2966,N_2882);
nand UO_334 (O_334,N_2985,N_2970);
nor UO_335 (O_335,N_2996,N_2960);
nor UO_336 (O_336,N_2867,N_2973);
nand UO_337 (O_337,N_2930,N_2937);
or UO_338 (O_338,N_2899,N_2822);
nand UO_339 (O_339,N_2934,N_2973);
nand UO_340 (O_340,N_2892,N_2957);
nor UO_341 (O_341,N_2818,N_2858);
and UO_342 (O_342,N_2903,N_2982);
or UO_343 (O_343,N_2849,N_2839);
nor UO_344 (O_344,N_2832,N_2976);
nor UO_345 (O_345,N_2874,N_2976);
or UO_346 (O_346,N_2824,N_2821);
xor UO_347 (O_347,N_2985,N_2976);
nand UO_348 (O_348,N_2831,N_2957);
or UO_349 (O_349,N_2958,N_2954);
nand UO_350 (O_350,N_2834,N_2936);
or UO_351 (O_351,N_2810,N_2870);
and UO_352 (O_352,N_2901,N_2926);
and UO_353 (O_353,N_2893,N_2844);
or UO_354 (O_354,N_2857,N_2892);
or UO_355 (O_355,N_2801,N_2943);
and UO_356 (O_356,N_2851,N_2966);
or UO_357 (O_357,N_2931,N_2823);
nor UO_358 (O_358,N_2821,N_2890);
or UO_359 (O_359,N_2913,N_2936);
and UO_360 (O_360,N_2991,N_2953);
nor UO_361 (O_361,N_2997,N_2985);
or UO_362 (O_362,N_2876,N_2891);
xnor UO_363 (O_363,N_2881,N_2915);
or UO_364 (O_364,N_2863,N_2807);
nand UO_365 (O_365,N_2813,N_2886);
nor UO_366 (O_366,N_2873,N_2925);
nor UO_367 (O_367,N_2806,N_2807);
nor UO_368 (O_368,N_2814,N_2887);
nor UO_369 (O_369,N_2948,N_2806);
and UO_370 (O_370,N_2839,N_2853);
nand UO_371 (O_371,N_2808,N_2842);
and UO_372 (O_372,N_2894,N_2812);
and UO_373 (O_373,N_2910,N_2918);
nand UO_374 (O_374,N_2827,N_2840);
nor UO_375 (O_375,N_2954,N_2906);
and UO_376 (O_376,N_2909,N_2848);
xnor UO_377 (O_377,N_2948,N_2802);
or UO_378 (O_378,N_2890,N_2878);
nand UO_379 (O_379,N_2991,N_2980);
xnor UO_380 (O_380,N_2899,N_2987);
nor UO_381 (O_381,N_2824,N_2903);
or UO_382 (O_382,N_2872,N_2914);
nand UO_383 (O_383,N_2997,N_2821);
nor UO_384 (O_384,N_2965,N_2800);
nand UO_385 (O_385,N_2943,N_2855);
nand UO_386 (O_386,N_2900,N_2921);
or UO_387 (O_387,N_2819,N_2940);
and UO_388 (O_388,N_2829,N_2999);
nor UO_389 (O_389,N_2810,N_2967);
and UO_390 (O_390,N_2913,N_2984);
or UO_391 (O_391,N_2952,N_2970);
and UO_392 (O_392,N_2944,N_2962);
nor UO_393 (O_393,N_2829,N_2951);
or UO_394 (O_394,N_2830,N_2979);
nor UO_395 (O_395,N_2878,N_2876);
xnor UO_396 (O_396,N_2897,N_2899);
and UO_397 (O_397,N_2848,N_2953);
nand UO_398 (O_398,N_2849,N_2897);
nor UO_399 (O_399,N_2975,N_2806);
and UO_400 (O_400,N_2853,N_2984);
nand UO_401 (O_401,N_2899,N_2990);
or UO_402 (O_402,N_2817,N_2986);
or UO_403 (O_403,N_2929,N_2849);
nor UO_404 (O_404,N_2891,N_2805);
and UO_405 (O_405,N_2989,N_2816);
nor UO_406 (O_406,N_2996,N_2835);
nand UO_407 (O_407,N_2869,N_2807);
or UO_408 (O_408,N_2896,N_2939);
xor UO_409 (O_409,N_2992,N_2881);
xnor UO_410 (O_410,N_2937,N_2984);
nor UO_411 (O_411,N_2913,N_2879);
nor UO_412 (O_412,N_2820,N_2921);
nand UO_413 (O_413,N_2833,N_2954);
or UO_414 (O_414,N_2889,N_2942);
nor UO_415 (O_415,N_2913,N_2970);
nand UO_416 (O_416,N_2928,N_2940);
nand UO_417 (O_417,N_2879,N_2971);
nor UO_418 (O_418,N_2951,N_2944);
nor UO_419 (O_419,N_2815,N_2830);
nand UO_420 (O_420,N_2830,N_2814);
nor UO_421 (O_421,N_2827,N_2870);
nor UO_422 (O_422,N_2962,N_2923);
nand UO_423 (O_423,N_2917,N_2864);
and UO_424 (O_424,N_2933,N_2851);
or UO_425 (O_425,N_2874,N_2872);
nand UO_426 (O_426,N_2913,N_2954);
xnor UO_427 (O_427,N_2942,N_2924);
and UO_428 (O_428,N_2880,N_2804);
or UO_429 (O_429,N_2912,N_2959);
and UO_430 (O_430,N_2954,N_2800);
nand UO_431 (O_431,N_2816,N_2987);
or UO_432 (O_432,N_2927,N_2933);
nand UO_433 (O_433,N_2950,N_2902);
nor UO_434 (O_434,N_2815,N_2931);
nand UO_435 (O_435,N_2972,N_2934);
xnor UO_436 (O_436,N_2962,N_2893);
nand UO_437 (O_437,N_2871,N_2921);
xnor UO_438 (O_438,N_2898,N_2861);
and UO_439 (O_439,N_2961,N_2869);
or UO_440 (O_440,N_2859,N_2978);
nand UO_441 (O_441,N_2905,N_2834);
and UO_442 (O_442,N_2994,N_2929);
and UO_443 (O_443,N_2911,N_2961);
nand UO_444 (O_444,N_2817,N_2904);
or UO_445 (O_445,N_2922,N_2967);
or UO_446 (O_446,N_2806,N_2899);
and UO_447 (O_447,N_2954,N_2979);
and UO_448 (O_448,N_2933,N_2923);
nand UO_449 (O_449,N_2966,N_2979);
or UO_450 (O_450,N_2892,N_2864);
nand UO_451 (O_451,N_2922,N_2930);
and UO_452 (O_452,N_2988,N_2853);
or UO_453 (O_453,N_2924,N_2847);
or UO_454 (O_454,N_2871,N_2821);
nor UO_455 (O_455,N_2928,N_2893);
or UO_456 (O_456,N_2929,N_2891);
nand UO_457 (O_457,N_2817,N_2980);
nor UO_458 (O_458,N_2931,N_2803);
and UO_459 (O_459,N_2891,N_2863);
xnor UO_460 (O_460,N_2907,N_2800);
nand UO_461 (O_461,N_2897,N_2896);
and UO_462 (O_462,N_2837,N_2961);
and UO_463 (O_463,N_2978,N_2801);
or UO_464 (O_464,N_2866,N_2900);
nand UO_465 (O_465,N_2979,N_2984);
nand UO_466 (O_466,N_2904,N_2947);
nand UO_467 (O_467,N_2854,N_2955);
nor UO_468 (O_468,N_2805,N_2871);
and UO_469 (O_469,N_2805,N_2967);
nand UO_470 (O_470,N_2994,N_2997);
or UO_471 (O_471,N_2834,N_2918);
and UO_472 (O_472,N_2810,N_2899);
nor UO_473 (O_473,N_2885,N_2871);
xnor UO_474 (O_474,N_2870,N_2806);
or UO_475 (O_475,N_2918,N_2973);
nor UO_476 (O_476,N_2905,N_2846);
or UO_477 (O_477,N_2907,N_2851);
nor UO_478 (O_478,N_2812,N_2897);
nor UO_479 (O_479,N_2868,N_2848);
and UO_480 (O_480,N_2868,N_2876);
or UO_481 (O_481,N_2823,N_2937);
nand UO_482 (O_482,N_2852,N_2900);
xnor UO_483 (O_483,N_2856,N_2907);
or UO_484 (O_484,N_2979,N_2832);
nor UO_485 (O_485,N_2993,N_2885);
or UO_486 (O_486,N_2879,N_2933);
nor UO_487 (O_487,N_2969,N_2885);
nor UO_488 (O_488,N_2971,N_2948);
nand UO_489 (O_489,N_2987,N_2939);
or UO_490 (O_490,N_2963,N_2921);
nor UO_491 (O_491,N_2992,N_2927);
or UO_492 (O_492,N_2914,N_2820);
and UO_493 (O_493,N_2812,N_2839);
nor UO_494 (O_494,N_2882,N_2905);
or UO_495 (O_495,N_2876,N_2927);
nand UO_496 (O_496,N_2807,N_2916);
nor UO_497 (O_497,N_2849,N_2938);
nand UO_498 (O_498,N_2886,N_2944);
and UO_499 (O_499,N_2994,N_2841);
endmodule